magic
tech ihp-sg13g2
magscale 1 2
timestamp 1747537721
<< nwell >>
rect -48 350 432 834
<< pwell >>
rect 5 56 386 288
rect -26 -56 410 56
<< nmos >>
rect 150 152 176 262
rect 266 114 292 262
<< pmos >>
rect 153 468 179 636
rect 259 412 285 636
<< ndiff >>
rect 31 247 150 262
rect 31 215 92 247
rect 124 215 150 247
rect 31 201 150 215
rect 96 152 150 201
rect 176 195 266 262
rect 176 163 204 195
rect 236 163 266 195
rect 176 152 266 163
rect 191 114 266 152
rect 292 245 360 262
rect 292 213 314 245
rect 346 213 360 245
rect 292 162 360 213
rect 292 130 314 162
rect 346 130 360 162
rect 292 114 360 130
<< pdiff >>
rect 81 620 153 636
rect 81 588 95 620
rect 127 588 153 620
rect 81 550 153 588
rect 81 518 95 550
rect 127 518 153 550
rect 81 468 153 518
rect 179 620 259 636
rect 179 588 203 620
rect 235 588 259 620
rect 179 468 259 588
rect 206 412 259 468
rect 285 620 357 636
rect 285 588 311 620
rect 343 588 357 620
rect 285 540 357 588
rect 285 508 311 540
rect 343 508 357 540
rect 285 464 357 508
rect 285 432 311 464
rect 343 432 357 464
rect 285 412 357 432
<< ndiffc >>
rect 92 215 124 247
rect 204 163 236 195
rect 314 213 346 245
rect 314 130 346 162
<< pdiffc >>
rect 95 588 127 620
rect 95 518 127 550
rect 203 588 235 620
rect 311 588 343 620
rect 311 508 343 540
rect 311 432 343 464
<< psubdiff >>
rect 0 16 384 30
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 384 16
rect 0 -30 384 -16
<< nsubdiff >>
rect 0 772 384 786
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 384 772
rect 0 726 384 740
<< psubdiffcont >>
rect 32 -16 64 16
rect 128 -16 160 16
rect 224 -16 256 16
rect 320 -16 352 16
<< nsubdiffcont >>
rect 32 740 64 772
rect 128 740 160 772
rect 224 740 256 772
rect 320 740 352 772
<< poly >>
rect 153 636 179 672
rect 259 636 285 672
rect 153 449 179 468
rect 146 414 182 449
rect 146 396 176 414
rect 40 379 176 396
rect 259 393 285 412
rect 40 347 57 379
rect 89 347 125 379
rect 157 347 176 379
rect 256 366 292 393
rect 40 330 176 347
rect 150 262 176 330
rect 224 349 292 366
rect 224 317 241 349
rect 273 317 292 349
rect 224 300 292 317
rect 266 262 292 300
rect 150 116 176 152
rect 266 78 292 114
<< polycont >>
rect 57 347 89 379
rect 125 347 157 379
rect 241 317 273 349
<< metal1 >>
rect 0 772 384 800
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 384 772
rect 0 712 384 740
rect 86 620 140 636
rect 86 588 95 620
rect 127 588 140 620
rect 86 550 140 588
rect 189 620 249 712
rect 189 588 203 620
rect 235 588 249 620
rect 189 568 249 588
rect 298 620 358 636
rect 298 588 311 620
rect 343 588 358 620
rect 86 518 95 550
rect 127 524 140 550
rect 298 540 358 588
rect 127 518 252 524
rect 86 488 252 518
rect 20 379 174 423
rect 20 347 57 379
rect 89 347 125 379
rect 157 347 174 379
rect 20 330 174 347
rect 218 366 252 488
rect 298 508 311 540
rect 343 508 358 540
rect 298 464 358 508
rect 298 432 311 464
rect 343 432 358 464
rect 298 404 358 432
rect 218 349 283 366
rect 218 317 241 349
rect 273 317 283 349
rect 218 300 283 317
rect 218 293 252 300
rect 63 258 252 293
rect 320 258 358 404
rect 63 247 141 258
rect 63 215 92 247
rect 124 215 141 247
rect 63 200 141 215
rect 300 245 358 258
rect 300 213 314 245
rect 346 213 358 245
rect 187 195 253 205
rect 187 163 204 195
rect 236 163 253 195
rect 187 44 253 163
rect 300 162 358 213
rect 300 130 314 162
rect 346 130 358 162
rect 300 110 358 130
rect 0 16 384 44
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 384 16
rect 0 -44 384 -16
<< labels >>
flabel metal1 s 0 -44 384 44 0 FreeSans 400 0 0 0 VSS
port 3 nsew
flabel metal1 s 0 712 384 800 0 FreeSans 400 0 0 0 VDD
port 2 nsew
<< properties >>
string FIXED_BBOX 0 0 384 756
string GDS_END 186940
string GDS_FILE ../gds/controller.gds
string GDS_START 183652
<< end >>
