magic
tech ihp-sg13g2
magscale 1 2
timestamp 1747056038
<< nwell >>
rect -48 350 1200 834
<< pwell >>
rect 19 56 1152 314
rect -26 -56 1178 56
<< nmos >>
rect 114 140 140 288
rect 216 140 242 288
rect 420 140 446 288
rect 522 140 548 288
rect 624 140 650 288
rect 726 140 752 288
rect 930 140 956 288
rect 1032 140 1058 288
<< pmos >>
rect 114 412 140 636
rect 216 412 242 636
rect 420 412 446 636
rect 522 412 548 636
rect 624 412 650 636
rect 726 412 752 636
rect 930 412 956 636
rect 1032 412 1058 636
<< ndiff >>
rect 45 274 114 288
rect 45 242 60 274
rect 92 242 114 274
rect 45 186 114 242
rect 45 154 60 186
rect 92 154 114 186
rect 45 140 114 154
rect 140 274 216 288
rect 140 242 162 274
rect 194 242 216 274
rect 140 186 216 242
rect 140 154 162 186
rect 194 154 216 186
rect 140 140 216 154
rect 242 186 420 288
rect 242 154 264 186
rect 296 154 366 186
rect 398 154 420 186
rect 242 140 420 154
rect 446 274 522 288
rect 446 242 468 274
rect 500 242 522 274
rect 446 186 522 242
rect 446 154 468 186
rect 500 154 522 186
rect 446 140 522 154
rect 548 186 624 288
rect 548 154 570 186
rect 602 154 624 186
rect 548 140 624 154
rect 650 274 726 288
rect 650 242 672 274
rect 704 242 726 274
rect 650 186 726 242
rect 650 154 672 186
rect 704 154 726 186
rect 650 140 726 154
rect 752 186 930 288
rect 752 154 774 186
rect 806 154 876 186
rect 908 154 930 186
rect 752 140 930 154
rect 956 274 1032 288
rect 956 242 978 274
rect 1010 242 1032 274
rect 956 186 1032 242
rect 956 154 978 186
rect 1010 154 1032 186
rect 956 140 1032 154
rect 1058 274 1126 288
rect 1058 242 1080 274
rect 1112 242 1126 274
rect 1058 186 1126 242
rect 1058 154 1080 186
rect 1112 154 1126 186
rect 1058 140 1126 154
<< pdiff >>
rect 45 622 114 636
rect 45 590 60 622
rect 92 590 114 622
rect 45 543 114 590
rect 45 511 60 543
rect 92 511 114 543
rect 45 458 114 511
rect 45 426 60 458
rect 92 426 114 458
rect 45 412 114 426
rect 140 622 216 636
rect 140 590 162 622
rect 194 590 216 622
rect 140 543 216 590
rect 140 511 162 543
rect 194 511 216 543
rect 140 458 216 511
rect 140 426 162 458
rect 194 426 216 458
rect 140 412 216 426
rect 242 622 310 636
rect 242 590 264 622
rect 296 590 310 622
rect 242 543 310 590
rect 242 511 264 543
rect 296 511 310 543
rect 242 412 310 511
rect 352 622 420 636
rect 352 590 366 622
rect 398 590 420 622
rect 352 543 420 590
rect 352 511 366 543
rect 398 511 420 543
rect 352 412 420 511
rect 446 543 522 636
rect 446 511 468 543
rect 500 511 522 543
rect 446 458 522 511
rect 446 426 468 458
rect 500 426 522 458
rect 446 412 522 426
rect 548 622 624 636
rect 548 590 570 622
rect 602 590 624 622
rect 548 543 624 590
rect 548 511 570 543
rect 602 511 624 543
rect 548 458 624 511
rect 548 426 570 458
rect 602 426 624 458
rect 548 412 624 426
rect 650 543 726 636
rect 650 511 672 543
rect 704 511 726 543
rect 650 458 726 511
rect 650 426 672 458
rect 704 426 726 458
rect 650 412 726 426
rect 752 622 820 636
rect 752 590 774 622
rect 806 590 820 622
rect 752 543 820 590
rect 752 511 774 543
rect 806 511 820 543
rect 752 412 820 511
rect 862 622 930 636
rect 862 590 876 622
rect 908 590 930 622
rect 862 543 930 590
rect 862 511 876 543
rect 908 511 930 543
rect 862 458 930 511
rect 862 426 876 458
rect 908 426 930 458
rect 862 412 930 426
rect 956 543 1032 636
rect 956 511 978 543
rect 1010 511 1032 543
rect 956 458 1032 511
rect 956 426 978 458
rect 1010 426 1032 458
rect 956 412 1032 426
rect 1058 622 1126 636
rect 1058 590 1080 622
rect 1112 590 1126 622
rect 1058 543 1126 590
rect 1058 511 1080 543
rect 1112 511 1126 543
rect 1058 458 1126 511
rect 1058 426 1080 458
rect 1112 426 1126 458
rect 1058 412 1126 426
<< ndiffc >>
rect 60 242 92 274
rect 60 154 92 186
rect 162 242 194 274
rect 162 154 194 186
rect 264 154 296 186
rect 366 154 398 186
rect 468 242 500 274
rect 468 154 500 186
rect 570 154 602 186
rect 672 242 704 274
rect 672 154 704 186
rect 774 154 806 186
rect 876 154 908 186
rect 978 242 1010 274
rect 978 154 1010 186
rect 1080 242 1112 274
rect 1080 154 1112 186
<< pdiffc >>
rect 60 590 92 622
rect 60 511 92 543
rect 60 426 92 458
rect 162 590 194 622
rect 162 511 194 543
rect 162 426 194 458
rect 264 590 296 622
rect 264 511 296 543
rect 366 590 398 622
rect 366 511 398 543
rect 468 511 500 543
rect 468 426 500 458
rect 570 590 602 622
rect 570 511 602 543
rect 570 426 602 458
rect 672 511 704 543
rect 672 426 704 458
rect 774 590 806 622
rect 774 511 806 543
rect 876 590 908 622
rect 876 511 908 543
rect 876 426 908 458
rect 978 511 1010 543
rect 978 426 1010 458
rect 1080 590 1112 622
rect 1080 511 1112 543
rect 1080 426 1112 458
<< psubdiff >>
rect 0 16 1152 30
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 608 16
rect 640 -16 704 16
rect 736 -16 800 16
rect 832 -16 896 16
rect 928 -16 992 16
rect 1024 -16 1088 16
rect 1120 -16 1152 16
rect 0 -30 1152 -16
<< nsubdiff >>
rect 0 772 1152 786
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 608 772
rect 640 740 704 772
rect 736 740 800 772
rect 832 740 896 772
rect 928 740 992 772
rect 1024 740 1088 772
rect 1120 740 1152 772
rect 0 726 1152 740
<< psubdiffcont >>
rect 32 -16 64 16
rect 128 -16 160 16
rect 224 -16 256 16
rect 320 -16 352 16
rect 416 -16 448 16
rect 512 -16 544 16
rect 608 -16 640 16
rect 704 -16 736 16
rect 800 -16 832 16
rect 896 -16 928 16
rect 992 -16 1024 16
rect 1088 -16 1120 16
<< nsubdiffcont >>
rect 32 740 64 772
rect 128 740 160 772
rect 224 740 256 772
rect 320 740 352 772
rect 416 740 448 772
rect 512 740 544 772
rect 608 740 640 772
rect 704 740 736 772
rect 800 740 832 772
rect 896 740 928 772
rect 992 740 1024 772
rect 1088 740 1120 772
<< poly >>
rect 114 636 140 672
rect 216 636 242 672
rect 420 636 446 672
rect 522 636 548 672
rect 624 636 650 672
rect 726 636 752 672
rect 930 636 956 672
rect 1032 636 1058 672
rect 114 380 140 412
rect 216 380 242 412
rect 420 380 446 412
rect 522 380 548 412
rect 624 380 650 412
rect 726 380 752 412
rect 930 380 956 412
rect 1032 380 1058 412
rect 97 366 259 380
rect 97 334 111 366
rect 143 334 213 366
rect 245 334 259 366
rect 97 320 259 334
rect 403 366 565 380
rect 403 334 417 366
rect 449 334 519 366
rect 551 334 565 366
rect 403 320 565 334
rect 607 366 769 380
rect 607 334 621 366
rect 653 334 723 366
rect 755 334 769 366
rect 607 320 769 334
rect 872 366 1075 380
rect 872 334 886 366
rect 918 334 1075 366
rect 872 320 1075 334
rect 114 288 140 320
rect 216 288 242 320
rect 420 288 446 320
rect 522 288 548 320
rect 624 288 650 320
rect 726 288 752 320
rect 930 288 956 320
rect 1032 288 1058 320
rect 114 104 140 140
rect 216 104 242 140
rect 420 104 446 140
rect 522 104 548 140
rect 624 104 650 140
rect 726 104 752 140
rect 930 104 956 140
rect 1032 104 1058 140
<< polycont >>
rect 111 334 143 366
rect 213 334 245 366
rect 417 334 449 366
rect 519 334 551 366
rect 621 334 653 366
rect 723 334 755 366
rect 886 334 918 366
<< metal1 >>
rect 0 772 1152 800
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 608 772
rect 640 740 704 772
rect 736 740 800 772
rect 832 740 896 772
rect 928 740 992 772
rect 1024 740 1088 772
rect 1120 740 1152 772
rect 0 712 1152 740
rect 50 622 102 712
rect 50 590 60 622
rect 92 590 102 622
rect 50 543 102 590
rect 50 511 60 543
rect 92 511 102 543
rect 50 458 102 511
rect 50 426 60 458
rect 92 426 102 458
rect 50 416 102 426
rect 152 622 204 632
rect 152 590 162 622
rect 194 590 204 622
rect 152 543 204 590
rect 152 511 162 543
rect 194 511 204 543
rect 152 468 204 511
rect 254 622 306 712
rect 254 590 264 622
rect 296 590 306 622
rect 254 543 306 590
rect 254 511 264 543
rect 296 511 306 543
rect 254 504 306 511
rect 356 622 816 641
rect 356 590 366 622
rect 398 590 570 622
rect 602 590 774 622
rect 806 590 816 622
rect 356 589 816 590
rect 356 543 408 589
rect 356 511 366 543
rect 398 511 408 543
rect 356 504 408 511
rect 458 543 510 553
rect 458 511 468 543
rect 500 511 510 543
rect 458 468 510 511
rect 152 458 510 468
rect 152 426 162 458
rect 194 426 468 458
rect 500 426 510 458
rect 152 425 510 426
rect 560 543 612 589
rect 560 511 570 543
rect 602 511 612 543
rect 560 458 612 511
rect 560 426 570 458
rect 602 426 612 458
rect 560 416 612 426
rect 662 543 714 553
rect 662 511 672 543
rect 704 511 714 543
rect 662 461 714 511
rect 764 543 816 589
rect 764 511 774 543
rect 806 511 816 543
rect 764 501 816 511
rect 866 622 1122 641
rect 866 590 876 622
rect 908 590 1080 622
rect 1112 590 1122 622
rect 866 589 1122 590
rect 866 543 918 589
rect 866 511 876 543
rect 908 511 918 543
rect 866 461 918 511
rect 662 458 918 461
rect 662 426 672 458
rect 704 426 876 458
rect 908 426 918 458
rect 662 425 918 426
rect 968 543 1020 553
rect 968 511 978 543
rect 1010 511 1020 543
rect 968 458 1020 511
rect 968 426 978 458
rect 1010 426 1020 458
rect 97 366 259 380
rect 97 334 111 366
rect 143 334 213 366
rect 245 334 259 366
rect 97 315 259 334
rect 403 366 565 380
rect 403 334 417 366
rect 449 334 519 366
rect 551 334 565 366
rect 403 315 565 334
rect 607 366 769 380
rect 607 334 621 366
rect 653 334 723 366
rect 755 334 769 366
rect 607 315 769 334
rect 805 366 932 380
rect 805 334 886 366
rect 918 334 932 366
rect 805 315 932 334
rect 968 275 1020 426
rect 1070 543 1122 589
rect 1070 511 1080 543
rect 1112 511 1122 543
rect 1070 458 1122 511
rect 1070 426 1080 458
rect 1112 426 1122 458
rect 1070 416 1122 426
rect 50 274 102 275
rect 50 242 60 274
rect 92 242 102 274
rect 50 186 102 242
rect 50 154 60 186
rect 92 154 102 186
rect 50 44 102 154
rect 152 274 1020 275
rect 152 242 162 274
rect 194 242 468 274
rect 500 242 672 274
rect 704 242 978 274
rect 1010 242 1020 274
rect 152 235 1020 242
rect 152 186 204 235
rect 152 154 162 186
rect 194 154 204 186
rect 152 144 204 154
rect 254 186 408 196
rect 254 154 264 186
rect 296 154 366 186
rect 398 154 408 186
rect 254 44 408 154
rect 458 186 510 235
rect 458 154 468 186
rect 500 154 510 186
rect 458 144 510 154
rect 560 186 612 196
rect 560 154 570 186
rect 602 154 612 186
rect 560 44 612 154
rect 662 186 714 235
rect 662 154 672 186
rect 704 154 714 186
rect 662 144 714 154
rect 764 186 918 196
rect 764 154 774 186
rect 806 154 876 186
rect 908 154 918 186
rect 764 44 918 154
rect 968 186 1020 235
rect 968 154 978 186
rect 1010 154 1020 186
rect 968 144 1020 154
rect 1070 274 1122 284
rect 1070 242 1080 274
rect 1112 242 1122 274
rect 1070 186 1122 242
rect 1070 154 1080 186
rect 1112 154 1122 186
rect 1070 44 1122 154
rect 0 16 1152 44
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 608 16
rect 640 -16 704 16
rect 736 -16 800 16
rect 832 -16 896 16
rect 928 -16 992 16
rect 1024 -16 1088 16
rect 1120 -16 1152 16
rect 0 -44 1152 -16
<< labels >>
flabel metal1 s 968 144 1020 553 0 FreeSans 500 0 0 0 Y
port 4 nsew
flabel metal1 s 805 316 932 380 0 FreeSans 500 0 0 0 D
port 1 nsew
flabel metal1 s 0 712 1152 800 0 FreeSans 500 0 0 0 VDD
port 5 nsew
flabel metal1 s 403 316 565 380 0 FreeSans 500 0 0 0 B
port 2 nsew
flabel metal1 s 97 316 259 380 0 FreeSans 500 0 0 0 A
port 7 nsew
flabel metal1 s 0 -44 1152 44 0 FreeSans 500 0 0 0 VSS
port 6 nsew
flabel metal1 s 607 316 769 380 0 FreeSans 500 0 0 0 C
port 3 nsew
<< properties >>
string FIXED_BBOX 0 0 1152 756
string GDS_END 248748
string GDS_FILE ../gds/controller.gds
string GDS_START 240490
<< end >>
