magic
tech ihp-sg13g2
magscale 1 2
timestamp 1747537721
<< nwell >>
rect -48 350 624 834
<< pwell >>
rect 30 56 550 292
rect -26 -56 602 56
<< nmos >>
rect 124 118 150 266
rect 226 118 252 266
rect 328 118 354 266
rect 430 118 456 266
<< pmos >>
rect 124 412 150 636
rect 226 412 252 636
rect 328 412 354 636
rect 430 412 456 636
<< ndiff >>
rect 56 252 124 266
rect 56 220 70 252
rect 102 220 124 252
rect 56 164 124 220
rect 56 132 70 164
rect 102 132 124 164
rect 56 118 124 132
rect 150 252 226 266
rect 150 220 172 252
rect 204 220 226 252
rect 150 164 226 220
rect 150 132 172 164
rect 204 132 226 164
rect 150 118 226 132
rect 252 164 328 266
rect 252 132 274 164
rect 306 132 328 164
rect 252 118 328 132
rect 354 252 430 266
rect 354 220 376 252
rect 408 220 430 252
rect 354 164 430 220
rect 354 132 376 164
rect 408 132 430 164
rect 354 118 430 132
rect 456 164 524 266
rect 456 132 478 164
rect 510 132 524 164
rect 456 118 524 132
<< pdiff >>
rect 52 622 124 636
rect 52 590 70 622
rect 102 590 124 622
rect 52 551 124 590
rect 52 519 70 551
rect 102 519 124 551
rect 52 458 124 519
rect 52 426 70 458
rect 102 426 124 458
rect 52 412 124 426
rect 150 622 226 636
rect 150 590 172 622
rect 204 590 226 622
rect 150 551 226 590
rect 150 519 172 551
rect 204 519 226 551
rect 150 412 226 519
rect 252 622 328 636
rect 252 590 274 622
rect 306 590 328 622
rect 252 551 328 590
rect 252 519 274 551
rect 306 519 328 551
rect 252 458 328 519
rect 252 426 274 458
rect 306 426 328 458
rect 252 412 328 426
rect 354 458 430 636
rect 354 426 376 458
rect 408 426 430 458
rect 354 412 430 426
rect 456 622 524 636
rect 456 590 478 622
rect 510 590 524 622
rect 456 551 524 590
rect 456 519 478 551
rect 510 519 524 551
rect 456 412 524 519
<< ndiffc >>
rect 70 220 102 252
rect 70 132 102 164
rect 172 220 204 252
rect 172 132 204 164
rect 274 132 306 164
rect 376 220 408 252
rect 376 132 408 164
rect 478 132 510 164
<< pdiffc >>
rect 70 590 102 622
rect 70 519 102 551
rect 70 426 102 458
rect 172 590 204 622
rect 172 519 204 551
rect 274 590 306 622
rect 274 519 306 551
rect 274 426 306 458
rect 376 426 408 458
rect 478 590 510 622
rect 478 519 510 551
<< psubdiff >>
rect 0 16 576 30
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 576 16
rect 0 -30 576 -16
<< nsubdiff >>
rect 0 772 576 786
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 576 772
rect 0 726 576 740
<< psubdiffcont >>
rect 32 -16 64 16
rect 128 -16 160 16
rect 224 -16 256 16
rect 320 -16 352 16
rect 416 -16 448 16
rect 512 -16 544 16
<< nsubdiffcont >>
rect 32 740 64 772
rect 128 740 160 772
rect 224 740 256 772
rect 320 740 352 772
rect 416 740 448 772
rect 512 740 544 772
<< poly >>
rect 124 636 150 672
rect 226 636 252 672
rect 328 636 354 672
rect 430 636 456 672
rect 124 368 150 412
rect 226 368 252 412
rect 124 353 252 368
rect 124 321 172 353
rect 204 321 252 353
rect 124 306 252 321
rect 124 266 150 306
rect 226 266 252 306
rect 328 368 354 412
rect 430 368 456 412
rect 328 353 456 368
rect 328 321 376 353
rect 408 321 456 353
rect 328 306 456 321
rect 328 266 354 306
rect 430 266 456 306
rect 124 82 150 118
rect 226 82 252 118
rect 328 82 354 118
rect 430 82 456 118
<< polycont >>
rect 172 321 204 353
rect 376 321 408 353
<< metal1 >>
rect 0 772 576 800
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 576 772
rect 0 712 576 740
rect 60 622 112 635
rect 60 590 70 622
rect 102 590 112 622
rect 60 551 112 590
rect 60 519 70 551
rect 102 519 112 551
rect 60 473 112 519
rect 162 622 214 712
rect 162 590 172 622
rect 204 590 214 622
rect 162 551 214 590
rect 162 519 172 551
rect 204 519 214 551
rect 162 509 214 519
rect 264 622 520 640
rect 264 590 274 622
rect 306 590 478 622
rect 510 590 520 622
rect 264 573 520 590
rect 264 551 316 573
rect 264 519 274 551
rect 306 519 316 551
rect 468 551 520 573
rect 264 473 316 519
rect 60 458 316 473
rect 60 426 70 458
rect 102 426 274 458
rect 306 426 316 458
rect 60 411 316 426
rect 356 472 426 528
rect 468 519 478 551
rect 510 519 520 551
rect 468 509 520 519
rect 356 458 520 472
rect 356 426 376 458
rect 408 426 520 458
rect 356 411 520 426
rect 155 353 221 365
rect 155 321 172 353
rect 204 321 221 353
rect 155 304 221 321
rect 361 353 425 365
rect 361 321 376 353
rect 408 321 425 353
rect 361 304 425 321
rect 60 252 112 264
rect 469 263 520 411
rect 60 220 70 252
rect 102 220 112 252
rect 60 164 112 220
rect 60 132 70 164
rect 102 132 112 164
rect 60 44 112 132
rect 162 252 520 263
rect 162 220 172 252
rect 204 220 376 252
rect 408 220 520 252
rect 162 215 520 220
rect 162 164 213 215
rect 162 132 172 164
rect 204 132 213 164
rect 162 118 213 132
rect 264 164 316 173
rect 264 132 274 164
rect 306 132 316 164
rect 264 44 316 132
rect 366 164 417 215
rect 366 132 376 164
rect 408 132 417 164
rect 366 118 417 132
rect 468 164 520 173
rect 468 132 478 164
rect 510 132 520 164
rect 468 44 520 132
rect 0 16 576 44
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 576 16
rect 0 -44 576 -16
<< labels >>
flabel metal1 s 155 304 221 365 0 FreeSans 400 0 0 0 A
port 2 nsew
flabel metal1 s 0 712 576 800 0 FreeSans 400 0 0 0 VDD
port 3 nsew
flabel metal1 s 356 411 426 528 0 FreeSans 400 0 0 0 Y
port 4 nsew
flabel metal1 s 0 -44 576 44 0 FreeSans 400 0 0 0 VSS
port 5 nsew
flabel metal1 s 361 304 425 365 0 FreeSans 400 0 0 0 B
port 6 nsew
<< properties >>
string FIXED_BBOX 0 0 576 756
string GDS_END 153712
string GDS_FILE ../gds/controller.gds
string GDS_START 144890
<< end >>
