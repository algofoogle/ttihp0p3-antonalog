magic
tech ihp-sg13g2
magscale 1 2
timestamp 1747492089
<< metal1 >>
rect 288 25724 2304 25748
rect 288 25684 1544 25724
rect 1912 25684 2304 25724
rect 288 25660 2304 25684
rect 268 24968 2304 24992
rect 268 24928 304 24968
rect 672 24928 2304 24968
rect 268 24904 2304 24928
rect 288 24212 2304 24236
rect 288 24172 1544 24212
rect 1912 24172 2304 24212
rect 288 24148 2304 24172
rect 268 23456 2304 23480
rect 268 23416 304 23456
rect 672 23416 2304 23456
rect 268 23392 2304 23416
rect 1515 23036 1557 23045
rect 1515 22996 1516 23036
rect 1556 22996 1557 23036
rect 1515 22987 1557 22996
rect 730 22868 788 22869
rect 730 22828 739 22868
rect 779 22828 788 22868
rect 730 22827 788 22828
rect 288 22700 2304 22724
rect 288 22660 1544 22700
rect 1912 22660 2304 22700
rect 288 22636 2304 22660
rect 1611 22364 1653 22373
rect 1611 22324 1612 22364
rect 1652 22324 1653 22364
rect 1611 22315 1653 22324
rect 826 22112 884 22113
rect 826 22072 835 22112
rect 875 22072 884 22112
rect 826 22071 884 22072
rect 268 21944 2304 21968
rect 268 21904 304 21944
rect 672 21904 2304 21944
rect 268 21880 2304 21904
rect 2091 21524 2133 21533
rect 2091 21484 2092 21524
rect 2132 21484 2133 21524
rect 2091 21475 2133 21484
rect 1306 21356 1364 21357
rect 1306 21316 1315 21356
rect 1355 21316 1364 21356
rect 1306 21315 1364 21316
rect 288 21188 2304 21212
rect 288 21148 1544 21188
rect 1912 21148 2304 21188
rect 288 21124 2304 21148
rect 2091 20852 2133 20861
rect 2091 20812 2092 20852
rect 2132 20812 2133 20852
rect 2091 20803 2133 20812
rect 1306 20600 1364 20601
rect 1306 20560 1315 20600
rect 1355 20560 1364 20600
rect 1306 20559 1364 20560
rect 268 20432 2304 20456
rect 268 20392 304 20432
rect 672 20392 2304 20432
rect 268 20368 2304 20392
rect 1515 20012 1557 20021
rect 1515 19972 1516 20012
rect 1556 19972 1557 20012
rect 1515 19963 1557 19972
rect 730 19844 788 19845
rect 730 19804 739 19844
rect 779 19804 788 19844
rect 730 19803 788 19804
rect 288 19676 2304 19700
rect 288 19636 1544 19676
rect 1912 19636 2304 19676
rect 288 19612 2304 19636
rect 1515 19340 1557 19349
rect 1515 19300 1516 19340
rect 1556 19300 1557 19340
rect 1515 19291 1557 19300
rect 730 19088 788 19089
rect 730 19048 739 19088
rect 779 19048 788 19088
rect 730 19047 788 19048
rect 268 18920 2304 18944
rect 268 18880 304 18920
rect 672 18880 2304 18920
rect 268 18856 2304 18880
rect 2091 18500 2133 18509
rect 2091 18460 2092 18500
rect 2132 18460 2133 18500
rect 2091 18451 2133 18460
rect 1306 18332 1364 18333
rect 1306 18292 1315 18332
rect 1355 18292 1364 18332
rect 1306 18291 1364 18292
rect 288 18164 2304 18188
rect 288 18124 1544 18164
rect 1912 18124 2304 18164
rect 288 18100 2304 18124
rect 1515 17828 1557 17837
rect 1515 17788 1516 17828
rect 1556 17788 1557 17828
rect 1515 17779 1557 17788
rect 730 17576 788 17577
rect 730 17536 739 17576
rect 779 17536 788 17576
rect 730 17535 788 17536
rect 268 17408 2304 17432
rect 268 17368 304 17408
rect 672 17368 2304 17408
rect 268 17344 2304 17368
rect 288 16652 2304 16676
rect 288 16612 1544 16652
rect 1912 16612 2304 16652
rect 288 16588 2304 16612
rect 268 15896 2304 15920
rect 268 15856 304 15896
rect 672 15856 2304 15896
rect 268 15832 2304 15856
rect 2091 15476 2133 15485
rect 2091 15436 2092 15476
rect 2132 15436 2133 15476
rect 2091 15427 2133 15436
rect 1306 15308 1364 15309
rect 1306 15268 1315 15308
rect 1355 15268 1364 15308
rect 1306 15267 1364 15268
rect 288 15140 2304 15164
rect 288 15100 1544 15140
rect 1912 15100 2304 15140
rect 288 15076 2304 15100
rect 1515 14804 1557 14813
rect 1515 14764 1516 14804
rect 1556 14764 1557 14804
rect 1515 14755 1557 14764
rect 730 14552 788 14553
rect 730 14512 739 14552
rect 779 14512 788 14552
rect 730 14511 788 14512
rect 268 14384 2304 14408
rect 268 14344 304 14384
rect 672 14344 2304 14384
rect 268 14320 2304 14344
rect 1515 13964 1557 13973
rect 1515 13924 1516 13964
rect 1556 13924 1557 13964
rect 1515 13915 1557 13924
rect 730 13796 788 13797
rect 730 13756 739 13796
rect 779 13756 788 13796
rect 730 13755 788 13756
rect 288 13628 2304 13652
rect 288 13588 1544 13628
rect 1912 13588 2304 13628
rect 288 13564 2304 13588
rect 2091 13292 2133 13301
rect 2091 13252 2092 13292
rect 2132 13252 2133 13292
rect 2091 13243 2133 13252
rect 1306 13040 1364 13041
rect 1306 13000 1315 13040
rect 1355 13000 1364 13040
rect 1306 12999 1364 13000
rect 268 12872 2304 12896
rect 268 12832 304 12872
rect 672 12832 2304 12872
rect 268 12808 2304 12832
rect 2091 12452 2133 12461
rect 2091 12412 2092 12452
rect 2132 12412 2133 12452
rect 2091 12403 2133 12412
rect 1306 12284 1364 12285
rect 1306 12244 1315 12284
rect 1355 12244 1364 12284
rect 1306 12243 1364 12244
rect 288 12116 2304 12140
rect 288 12076 1544 12116
rect 1912 12076 2304 12116
rect 288 12052 2304 12076
rect 1515 11780 1557 11789
rect 1515 11740 1516 11780
rect 1556 11740 1557 11780
rect 1515 11731 1557 11740
rect 730 11528 788 11529
rect 730 11488 739 11528
rect 779 11488 788 11528
rect 730 11487 788 11488
rect 268 11360 2304 11384
rect 268 11320 304 11360
rect 672 11320 2304 11360
rect 268 11296 2304 11320
rect 1515 10940 1557 10949
rect 1515 10900 1516 10940
rect 1556 10900 1557 10940
rect 1515 10891 1557 10900
rect 730 10772 788 10773
rect 730 10732 739 10772
rect 779 10732 788 10772
rect 730 10731 788 10732
rect 288 10604 2304 10628
rect 288 10564 1544 10604
rect 1912 10564 2304 10604
rect 288 10540 2304 10564
rect 2091 10268 2133 10277
rect 2091 10228 2092 10268
rect 2132 10228 2133 10268
rect 2091 10219 2133 10228
rect 1306 10016 1364 10017
rect 1306 9976 1315 10016
rect 1355 9976 1364 10016
rect 1306 9975 1364 9976
rect 268 9848 2304 9872
rect 268 9808 304 9848
rect 672 9808 2304 9848
rect 268 9784 2304 9808
rect 288 9092 2304 9116
rect 288 9052 1544 9092
rect 1912 9052 2304 9092
rect 288 9028 2304 9052
rect 268 8336 2304 8360
rect 268 8296 304 8336
rect 672 8296 2304 8336
rect 268 8272 2304 8296
rect 1515 7916 1557 7925
rect 1515 7876 1516 7916
rect 1556 7876 1557 7916
rect 1515 7867 1557 7876
rect 730 7748 788 7749
rect 730 7708 739 7748
rect 779 7708 788 7748
rect 730 7707 788 7708
rect 288 7580 2304 7604
rect 288 7540 1544 7580
rect 1912 7540 2304 7580
rect 288 7516 2304 7540
rect 1803 7244 1845 7253
rect 1803 7204 1804 7244
rect 1844 7204 1845 7244
rect 1803 7195 1845 7204
rect 1018 6992 1076 6993
rect 1018 6952 1027 6992
rect 1067 6952 1076 6992
rect 1018 6951 1076 6952
rect 268 6824 2304 6848
rect 268 6784 304 6824
rect 672 6784 2304 6824
rect 268 6760 2304 6784
rect 1515 6404 1557 6413
rect 1515 6364 1516 6404
rect 1556 6364 1557 6404
rect 1515 6355 1557 6364
rect 730 6236 788 6237
rect 730 6196 739 6236
rect 779 6196 788 6236
rect 730 6195 788 6196
rect 288 6068 2304 6092
rect 288 6028 1544 6068
rect 1912 6028 2304 6068
rect 288 6004 2304 6028
rect 2091 5732 2133 5741
rect 2091 5692 2092 5732
rect 2132 5692 2133 5732
rect 2091 5683 2133 5692
rect 1306 5480 1364 5481
rect 1306 5440 1315 5480
rect 1355 5440 1364 5480
rect 1306 5439 1364 5440
rect 268 5312 2304 5336
rect 268 5272 304 5312
rect 672 5272 2304 5312
rect 268 5248 2304 5272
rect 2091 4892 2133 4901
rect 2091 4852 2092 4892
rect 2132 4852 2133 4892
rect 2091 4843 2133 4852
rect 1306 4724 1364 4725
rect 1306 4684 1315 4724
rect 1355 4684 1364 4724
rect 1306 4683 1364 4684
rect 288 4556 2304 4580
rect 288 4516 1544 4556
rect 1912 4516 2304 4556
rect 288 4492 2304 4516
rect 1515 4220 1557 4229
rect 1515 4180 1516 4220
rect 1556 4180 1557 4220
rect 1515 4171 1557 4180
rect 730 3968 788 3969
rect 730 3928 739 3968
rect 779 3928 788 3968
rect 730 3927 788 3928
rect 268 3800 2304 3824
rect 268 3760 304 3800
rect 672 3760 2304 3800
rect 268 3736 2304 3760
rect 2091 3380 2133 3389
rect 2091 3340 2092 3380
rect 2132 3340 2133 3380
rect 2091 3331 2133 3340
rect 1306 3212 1364 3213
rect 1306 3172 1315 3212
rect 1355 3172 1364 3212
rect 1306 3171 1364 3172
rect 288 3044 2304 3068
rect 288 3004 1544 3044
rect 1912 3004 2304 3044
rect 288 2980 2304 3004
rect 1515 2708 1557 2717
rect 1515 2668 1516 2708
rect 1556 2668 1557 2708
rect 1515 2659 1557 2668
rect 730 2456 788 2457
rect 730 2416 739 2456
rect 779 2416 788 2456
rect 730 2415 788 2416
rect 268 2288 2304 2312
rect 268 2248 304 2288
rect 672 2248 2304 2288
rect 268 2224 2304 2248
rect 288 1532 2304 1556
rect 288 1492 1544 1532
rect 1912 1492 2304 1532
rect 288 1468 2304 1492
rect 268 776 2304 800
rect 268 736 304 776
rect 672 736 2304 776
rect 268 712 2304 736
rect 288 20 2304 44
rect 288 -20 1544 20
rect 1912 -20 2304 20
rect 288 -44 2304 -20
<< via1 >>
rect 1544 25684 1912 25724
rect 304 24928 672 24968
rect 1544 24172 1912 24212
rect 304 23416 672 23456
rect 1516 22996 1556 23036
rect 739 22828 779 22868
rect 1544 22660 1912 22700
rect 1612 22324 1652 22364
rect 835 22072 875 22112
rect 304 21904 672 21944
rect 2092 21484 2132 21524
rect 1315 21316 1355 21356
rect 1544 21148 1912 21188
rect 2092 20812 2132 20852
rect 1315 20560 1355 20600
rect 304 20392 672 20432
rect 1516 19972 1556 20012
rect 739 19804 779 19844
rect 1544 19636 1912 19676
rect 1516 19300 1556 19340
rect 739 19048 779 19088
rect 304 18880 672 18920
rect 2092 18460 2132 18500
rect 1315 18292 1355 18332
rect 1544 18124 1912 18164
rect 1516 17788 1556 17828
rect 739 17536 779 17576
rect 304 17368 672 17408
rect 1544 16612 1912 16652
rect 304 15856 672 15896
rect 2092 15436 2132 15476
rect 1315 15268 1355 15308
rect 1544 15100 1912 15140
rect 1516 14764 1556 14804
rect 739 14512 779 14552
rect 304 14344 672 14384
rect 1516 13924 1556 13964
rect 739 13756 779 13796
rect 1544 13588 1912 13628
rect 2092 13252 2132 13292
rect 1315 13000 1355 13040
rect 304 12832 672 12872
rect 2092 12412 2132 12452
rect 1315 12244 1355 12284
rect 1544 12076 1912 12116
rect 1516 11740 1556 11780
rect 739 11488 779 11528
rect 304 11320 672 11360
rect 1516 10900 1556 10940
rect 739 10732 779 10772
rect 1544 10564 1912 10604
rect 2092 10228 2132 10268
rect 1315 9976 1355 10016
rect 304 9808 672 9848
rect 1544 9052 1912 9092
rect 304 8296 672 8336
rect 1516 7876 1556 7916
rect 739 7708 779 7748
rect 1544 7540 1912 7580
rect 1804 7204 1844 7244
rect 1027 6952 1067 6992
rect 304 6784 672 6824
rect 1516 6364 1556 6404
rect 739 6196 779 6236
rect 1544 6028 1912 6068
rect 2092 5692 2132 5732
rect 1315 5440 1355 5480
rect 304 5272 672 5312
rect 2092 4852 2132 4892
rect 1315 4684 1355 4724
rect 1544 4516 1912 4556
rect 1516 4180 1556 4220
rect 739 3928 779 3968
rect 304 3760 672 3800
rect 2092 3340 2132 3380
rect 1315 3172 1355 3212
rect 1544 3004 1912 3044
rect 1516 2668 1556 2708
rect 739 2416 779 2456
rect 304 2248 672 2288
rect 1544 1492 1912 1532
rect 304 736 672 776
rect 1544 -20 1912 20
<< metal2 >>
rect 1535 25684 1544 25724
rect 1912 25684 1921 25724
rect 295 24928 304 24968
rect 672 24928 681 24968
rect 1535 24172 1544 24212
rect 1912 24172 1921 24212
rect 295 23416 304 23456
rect 672 23416 681 23456
rect 1507 22996 1516 23036
rect 1556 22996 1996 23036
rect 2036 22996 2045 23036
rect 730 22828 739 22868
rect 779 22828 788 22868
rect 0 22784 100 22804
rect 748 22784 788 22828
rect 0 22744 788 22784
rect 0 22724 100 22744
rect 1535 22660 1544 22700
rect 1912 22660 1921 22700
rect 1603 22324 1612 22364
rect 1652 22324 2188 22364
rect 2228 22324 2237 22364
rect 826 22072 835 22112
rect 875 22072 884 22112
rect 0 22028 100 22048
rect 844 22028 884 22072
rect 0 21988 884 22028
rect 0 21968 100 21988
rect 295 21904 304 21944
rect 672 21904 681 21944
rect 2083 21484 2092 21524
rect 2132 21484 2284 21524
rect 2324 21484 2333 21524
rect 1306 21316 1315 21356
rect 1355 21316 1364 21356
rect 0 21272 100 21292
rect 1324 21272 1364 21316
rect 0 21232 1364 21272
rect 0 21212 100 21232
rect 1535 21148 1544 21188
rect 1912 21148 1921 21188
rect 2500 21104 2600 21124
rect 1987 21064 1996 21104
rect 2036 21064 2600 21104
rect 2500 21044 2600 21064
rect 1961 20812 2092 20852
rect 2132 20812 2141 20852
rect 2500 20684 2600 20704
rect 2179 20644 2188 20684
rect 2228 20644 2600 20684
rect 2500 20624 2600 20644
rect 1306 20560 1315 20600
rect 1355 20560 1364 20600
rect 0 20516 100 20536
rect 1324 20516 1364 20560
rect 0 20476 1364 20516
rect 0 20456 100 20476
rect 295 20392 304 20432
rect 672 20392 681 20432
rect 2500 20264 2600 20284
rect 2275 20224 2284 20264
rect 2324 20224 2600 20264
rect 2500 20204 2600 20224
rect 1507 19972 1516 20012
rect 1556 19972 1996 20012
rect 2036 19972 2045 20012
rect 2500 19844 2600 19864
rect 730 19804 739 19844
rect 779 19804 788 19844
rect 2083 19804 2092 19844
rect 2132 19804 2600 19844
rect 0 19760 100 19780
rect 748 19760 788 19804
rect 2500 19784 2600 19804
rect 0 19720 788 19760
rect 0 19700 100 19720
rect 1535 19636 1544 19676
rect 1912 19636 1921 19676
rect 2500 19424 2600 19444
rect 1987 19384 1996 19424
rect 2036 19384 2600 19424
rect 2500 19364 2600 19384
rect 1507 19300 1516 19340
rect 1556 19300 1940 19340
rect 730 19048 739 19088
rect 779 19048 788 19088
rect 0 19004 100 19024
rect 748 19004 788 19048
rect 0 18964 788 19004
rect 1900 19004 1940 19300
rect 2500 19004 2600 19024
rect 1900 18964 2600 19004
rect 0 18944 100 18964
rect 2500 18944 2600 18964
rect 295 18880 304 18920
rect 672 18880 681 18920
rect 2500 18584 2600 18604
rect 2092 18544 2600 18584
rect 2092 18500 2132 18544
rect 2500 18524 2600 18544
rect 2083 18460 2092 18500
rect 2132 18460 2141 18500
rect 1306 18292 1315 18332
rect 1355 18292 1364 18332
rect 0 18248 100 18268
rect 1324 18248 1364 18292
rect 0 18208 1364 18248
rect 0 18188 100 18208
rect 2500 18164 2600 18184
rect 1535 18124 1544 18164
rect 1912 18124 1921 18164
rect 1996 18124 2600 18164
rect 1996 17828 2036 18124
rect 2500 18104 2600 18124
rect 1507 17788 1516 17828
rect 1556 17788 2036 17828
rect 730 17536 739 17576
rect 779 17536 788 17576
rect 0 17492 100 17512
rect 748 17492 788 17536
rect 0 17452 788 17492
rect 0 17432 100 17452
rect 295 17368 304 17408
rect 672 17368 681 17408
rect 1535 16612 1544 16652
rect 1912 16612 1921 16652
rect 295 15856 304 15896
rect 672 15856 681 15896
rect 1961 15436 2092 15476
rect 2132 15436 2141 15476
rect 1306 15268 1315 15308
rect 1355 15268 1364 15308
rect 0 15224 100 15244
rect 1324 15224 1364 15268
rect 0 15184 1364 15224
rect 0 15164 100 15184
rect 1535 15100 1544 15140
rect 1912 15100 1921 15140
rect 1507 14764 1516 14804
rect 1556 14764 1708 14804
rect 1748 14764 1757 14804
rect 730 14512 739 14552
rect 779 14512 788 14552
rect 0 14468 100 14488
rect 748 14468 788 14512
rect 0 14428 788 14468
rect 0 14408 100 14428
rect 2500 14384 2600 14404
rect 295 14344 304 14384
rect 672 14344 681 14384
rect 2083 14344 2092 14384
rect 2132 14344 2600 14384
rect 2500 14324 2600 14344
rect 2500 13964 2600 13984
rect 1507 13924 1516 13964
rect 1556 13924 1565 13964
rect 1699 13924 1708 13964
rect 1748 13924 2600 13964
rect 1516 13880 1556 13924
rect 2500 13904 2600 13924
rect 1516 13840 2036 13880
rect 730 13756 739 13796
rect 779 13756 788 13796
rect 0 13712 100 13732
rect 748 13712 788 13756
rect 0 13672 788 13712
rect 0 13652 100 13672
rect 1535 13588 1544 13628
rect 1912 13588 1921 13628
rect 1996 13544 2036 13840
rect 2500 13544 2600 13564
rect 1996 13504 2600 13544
rect 2500 13484 2600 13504
rect 2083 13252 2092 13292
rect 2132 13252 2141 13292
rect 2092 13124 2132 13252
rect 2500 13124 2600 13144
rect 2092 13084 2600 13124
rect 2500 13064 2600 13084
rect 1306 13000 1315 13040
rect 1355 13000 1364 13040
rect 0 12956 100 12976
rect 1324 12956 1364 13000
rect 0 12916 1364 12956
rect 0 12896 100 12916
rect 295 12832 304 12872
rect 672 12832 681 12872
rect 2500 12704 2600 12724
rect 2092 12664 2600 12704
rect 2092 12452 2132 12664
rect 2500 12644 2600 12664
rect 2083 12412 2092 12452
rect 2132 12412 2141 12452
rect 2500 12284 2600 12304
rect 1306 12244 1315 12284
rect 1355 12244 1364 12284
rect 1987 12244 1996 12284
rect 2036 12244 2600 12284
rect 0 12200 100 12220
rect 1324 12200 1364 12244
rect 2500 12224 2600 12244
rect 0 12160 1364 12200
rect 0 12140 100 12160
rect 1535 12076 1544 12116
rect 1912 12076 1921 12116
rect 2500 11864 2600 11884
rect 1507 11824 1516 11864
rect 1556 11824 2600 11864
rect 2500 11804 2600 11824
rect 1507 11740 1516 11780
rect 1556 11740 1996 11780
rect 2036 11740 2045 11780
rect 730 11488 739 11528
rect 779 11488 788 11528
rect 0 11444 100 11464
rect 748 11444 788 11488
rect 2500 11444 2600 11464
rect 0 11404 788 11444
rect 2083 11404 2092 11444
rect 2132 11404 2600 11444
rect 0 11384 100 11404
rect 2500 11384 2600 11404
rect 295 11320 304 11360
rect 672 11320 681 11360
rect 1385 10900 1516 10940
rect 1556 10900 1565 10940
rect 730 10732 739 10772
rect 779 10732 788 10772
rect 0 10688 100 10708
rect 748 10688 788 10732
rect 0 10648 788 10688
rect 0 10628 100 10648
rect 1535 10564 1544 10604
rect 1912 10564 1921 10604
rect 1961 10228 2092 10268
rect 2132 10228 2141 10268
rect 1306 9976 1315 10016
rect 1355 9976 1364 10016
rect 0 9932 100 9952
rect 1324 9932 1364 9976
rect 0 9892 1364 9932
rect 0 9872 100 9892
rect 295 9808 304 9848
rect 672 9808 681 9848
rect 1535 9052 1544 9092
rect 1912 9052 1921 9092
rect 295 8296 304 8336
rect 672 8296 681 8336
rect 1507 7876 1516 7916
rect 1556 7876 1565 7916
rect 730 7708 739 7748
rect 779 7708 788 7748
rect 0 7664 100 7684
rect 748 7664 788 7708
rect 0 7624 788 7664
rect 1516 7664 1556 7876
rect 2500 7664 2600 7684
rect 1516 7624 2600 7664
rect 0 7604 100 7624
rect 2500 7604 2600 7624
rect 1535 7540 1544 7580
rect 1912 7540 1921 7580
rect 2500 7244 2600 7264
rect 1795 7204 1804 7244
rect 1844 7204 2600 7244
rect 2500 7184 2600 7204
rect 1018 6952 1027 6992
rect 1067 6952 1076 6992
rect 0 6908 100 6928
rect 1036 6908 1076 6952
rect 0 6868 1076 6908
rect 0 6848 100 6868
rect 2500 6824 2600 6844
rect 295 6784 304 6824
rect 672 6784 681 6824
rect 1507 6784 1516 6824
rect 1556 6784 2600 6824
rect 2500 6764 2600 6784
rect 2500 6404 2600 6424
rect 1385 6364 1516 6404
rect 1556 6364 1565 6404
rect 2083 6364 2092 6404
rect 2132 6364 2600 6404
rect 2500 6344 2600 6364
rect 730 6196 739 6236
rect 779 6196 788 6236
rect 0 6152 100 6172
rect 748 6152 788 6196
rect 0 6112 788 6152
rect 0 6092 100 6112
rect 1535 6028 1544 6068
rect 1912 6028 1921 6068
rect 2500 5984 2600 6004
rect 2275 5944 2284 5984
rect 2324 5944 2600 5984
rect 2500 5924 2600 5944
rect 1961 5692 2092 5732
rect 2132 5692 2141 5732
rect 2500 5564 2600 5584
rect 2179 5524 2188 5564
rect 2228 5524 2600 5564
rect 2500 5504 2600 5524
rect 1306 5440 1315 5480
rect 1355 5440 1364 5480
rect 0 5396 100 5416
rect 1324 5396 1364 5440
rect 0 5356 1364 5396
rect 0 5336 100 5356
rect 295 5272 304 5312
rect 672 5272 681 5312
rect 2500 5144 2600 5164
rect 2083 5104 2092 5144
rect 2132 5104 2600 5144
rect 2500 5084 2600 5104
rect 2083 4852 2092 4892
rect 2132 4852 2284 4892
rect 2324 4852 2333 4892
rect 2500 4724 2600 4744
rect 1306 4684 1315 4724
rect 1355 4684 1364 4724
rect 1987 4684 1996 4724
rect 2036 4684 2600 4724
rect 0 4640 100 4660
rect 1324 4640 1364 4684
rect 2500 4664 2600 4684
rect 0 4600 1364 4640
rect 0 4580 100 4600
rect 1535 4516 1544 4556
rect 1912 4516 1921 4556
rect 1507 4180 1516 4220
rect 1556 4180 2188 4220
rect 2228 4180 2237 4220
rect 730 3928 739 3968
rect 779 3928 788 3968
rect 0 3884 100 3904
rect 748 3884 788 3928
rect 0 3844 788 3884
rect 0 3824 100 3844
rect 295 3760 304 3800
rect 672 3760 681 3800
rect 1961 3340 2092 3380
rect 2132 3340 2141 3380
rect 1306 3172 1315 3212
rect 1355 3172 1364 3212
rect 0 3128 100 3148
rect 1324 3128 1364 3172
rect 0 3088 1364 3128
rect 0 3068 100 3088
rect 1535 3004 1544 3044
rect 1912 3004 1921 3044
rect 1507 2668 1516 2708
rect 1556 2668 1996 2708
rect 2036 2668 2045 2708
rect 730 2416 739 2456
rect 779 2416 788 2456
rect 0 2372 100 2392
rect 748 2372 788 2416
rect 0 2332 788 2372
rect 0 2312 100 2332
rect 295 2248 304 2288
rect 672 2248 681 2288
rect 1535 1492 1544 1532
rect 1912 1492 1921 1532
rect 295 736 304 776
rect 672 736 681 776
rect 1535 -20 1544 20
rect 1912 -20 1921 20
<< via2 >>
rect 1544 25684 1912 25724
rect 304 24928 672 24968
rect 1544 24172 1912 24212
rect 304 23416 672 23456
rect 1996 22996 2036 23036
rect 1544 22660 1912 22700
rect 2188 22324 2228 22364
rect 304 21904 672 21944
rect 2284 21484 2324 21524
rect 1544 21148 1912 21188
rect 1996 21064 2036 21104
rect 2092 20812 2132 20852
rect 2188 20644 2228 20684
rect 304 20392 672 20432
rect 2284 20224 2324 20264
rect 1996 19972 2036 20012
rect 2092 19804 2132 19844
rect 1544 19636 1912 19676
rect 1996 19384 2036 19424
rect 304 18880 672 18920
rect 1544 18124 1912 18164
rect 304 17368 672 17408
rect 1544 16612 1912 16652
rect 304 15856 672 15896
rect 2092 15436 2132 15476
rect 1544 15100 1912 15140
rect 1708 14764 1748 14804
rect 304 14344 672 14384
rect 2092 14344 2132 14384
rect 1708 13924 1748 13964
rect 1544 13588 1912 13628
rect 304 12832 672 12872
rect 1996 12244 2036 12284
rect 1544 12076 1912 12116
rect 1516 11824 1556 11864
rect 1996 11740 2036 11780
rect 2092 11404 2132 11444
rect 304 11320 672 11360
rect 1516 10900 1556 10940
rect 1544 10564 1912 10604
rect 2092 10228 2132 10268
rect 304 9808 672 9848
rect 1544 9052 1912 9092
rect 304 8296 672 8336
rect 1544 7540 1912 7580
rect 304 6784 672 6824
rect 1516 6784 1556 6824
rect 1516 6364 1556 6404
rect 2092 6364 2132 6404
rect 1544 6028 1912 6068
rect 2284 5944 2324 5984
rect 2092 5692 2132 5732
rect 2188 5524 2228 5564
rect 304 5272 672 5312
rect 2092 5104 2132 5144
rect 2284 4852 2324 4892
rect 1996 4684 2036 4724
rect 1544 4516 1912 4556
rect 2188 4180 2228 4220
rect 304 3760 672 3800
rect 2092 3340 2132 3380
rect 1544 3004 1912 3044
rect 1996 2668 2036 2708
rect 304 2248 672 2288
rect 1544 1492 1912 1532
rect 304 736 672 776
rect 1544 -20 1912 20
<< metal3 >>
rect 1544 25724 1912 25733
rect 1544 25675 1912 25684
rect 304 24968 672 24977
rect 304 24919 672 24928
rect 1544 24212 1912 24221
rect 1544 24163 1912 24172
rect 304 23456 672 23465
rect 304 23407 672 23416
rect 1996 23036 2036 23045
rect 1544 22700 1912 22709
rect 1544 22651 1912 22660
rect 304 21944 672 21953
rect 304 21895 672 21904
rect 1544 21188 1912 21197
rect 1544 21139 1912 21148
rect 1996 21104 2036 22996
rect 1996 21055 2036 21064
rect 2188 22364 2228 22373
rect 2092 20852 2132 20861
rect 304 20432 672 20441
rect 304 20383 672 20392
rect 1996 20012 2036 20021
rect 1544 19676 1912 19685
rect 1544 19627 1912 19636
rect 1996 19424 2036 19972
rect 2092 19844 2132 20812
rect 2188 20684 2228 22324
rect 2188 20635 2228 20644
rect 2284 21524 2324 21533
rect 2284 20264 2324 21484
rect 2284 20215 2324 20224
rect 2092 19795 2132 19804
rect 1996 19375 2036 19384
rect 304 18920 672 18929
rect 304 18871 672 18880
rect 1544 18164 1912 18173
rect 1544 18115 1912 18124
rect 304 17408 672 17417
rect 304 17359 672 17368
rect 1544 16652 1912 16661
rect 1544 16603 1912 16612
rect 304 15896 672 15905
rect 304 15847 672 15856
rect 2092 15476 2132 15485
rect 1544 15140 1912 15149
rect 1544 15091 1912 15100
rect 1708 14804 1748 14813
rect 304 14384 672 14393
rect 304 14335 672 14344
rect 1708 13964 1748 14764
rect 2092 14384 2132 15436
rect 2092 14335 2132 14344
rect 1708 13915 1748 13924
rect 1544 13628 1912 13637
rect 1544 13579 1912 13588
rect 304 12872 672 12881
rect 304 12823 672 12832
rect 1996 12284 2036 12293
rect 1544 12116 1912 12125
rect 1544 12067 1912 12076
rect 1516 11864 1556 11873
rect 304 11360 672 11369
rect 304 11311 672 11320
rect 1516 10940 1556 11824
rect 1996 11780 2036 12244
rect 1996 11731 2036 11740
rect 1516 10891 1556 10900
rect 2092 11444 2132 11453
rect 1544 10604 1912 10613
rect 1544 10555 1912 10564
rect 2092 10268 2132 11404
rect 2092 10219 2132 10228
rect 304 9848 672 9857
rect 304 9799 672 9808
rect 1544 9092 1912 9101
rect 1544 9043 1912 9052
rect 304 8336 672 8345
rect 304 8287 672 8296
rect 1544 7580 1912 7589
rect 1544 7531 1912 7540
rect 304 6824 672 6833
rect 304 6775 672 6784
rect 1516 6824 1556 6833
rect 1516 6404 1556 6784
rect 1516 6355 1556 6364
rect 2092 6404 2132 6413
rect 1544 6068 1912 6077
rect 1544 6019 1912 6028
rect 2092 5732 2132 6364
rect 2092 5683 2132 5692
rect 2284 5984 2324 5993
rect 2188 5564 2228 5573
rect 304 5312 672 5321
rect 304 5263 672 5272
rect 2092 5144 2132 5153
rect 1996 4724 2036 4733
rect 1544 4556 1912 4565
rect 1544 4507 1912 4516
rect 304 3800 672 3809
rect 304 3751 672 3760
rect 1544 3044 1912 3053
rect 1544 2995 1912 3004
rect 1996 2708 2036 4684
rect 2092 3380 2132 5104
rect 2188 4220 2228 5524
rect 2284 4892 2324 5944
rect 2284 4843 2324 4852
rect 2188 4171 2228 4180
rect 2092 3331 2132 3340
rect 1996 2659 2036 2668
rect 304 2288 672 2297
rect 304 2239 672 2248
rect 1544 1532 1912 1541
rect 1544 1483 1912 1492
rect 304 776 672 785
rect 304 727 672 736
rect 1544 20 1912 29
rect 1544 -29 1912 -20
<< via3 >>
rect 1544 25684 1912 25724
rect 304 24928 672 24968
rect 1544 24172 1912 24212
rect 304 23416 672 23456
rect 1544 22660 1912 22700
rect 304 21904 672 21944
rect 1544 21148 1912 21188
rect 304 20392 672 20432
rect 1544 19636 1912 19676
rect 304 18880 672 18920
rect 1544 18124 1912 18164
rect 304 17368 672 17408
rect 1544 16612 1912 16652
rect 304 15856 672 15896
rect 1544 15100 1912 15140
rect 304 14344 672 14384
rect 1544 13588 1912 13628
rect 304 12832 672 12872
rect 1544 12076 1912 12116
rect 304 11320 672 11360
rect 1544 10564 1912 10604
rect 304 9808 672 9848
rect 1544 9052 1912 9092
rect 304 8296 672 8336
rect 1544 7540 1912 7580
rect 304 6784 672 6824
rect 1544 6028 1912 6068
rect 304 5272 672 5312
rect 1544 4516 1912 4556
rect 304 3760 672 3800
rect 1544 3004 1912 3044
rect 304 2248 672 2288
rect 1544 1492 1912 1532
rect 304 736 672 776
rect 1544 -20 1912 20
<< metal4 >>
rect 1535 25684 1544 25724
rect 1912 25684 1921 25724
rect 295 24928 304 24968
rect 672 24928 681 24968
rect 1535 24172 1544 24212
rect 1912 24172 1921 24212
rect 295 23416 304 23456
rect 672 23416 681 23456
rect 1535 22660 1544 22700
rect 1912 22660 1921 22700
rect 295 21904 304 21944
rect 672 21904 681 21944
rect 1535 21148 1544 21188
rect 1912 21148 1921 21188
rect 295 20392 304 20432
rect 672 20392 681 20432
rect 1535 19636 1544 19676
rect 1912 19636 1921 19676
rect 295 18880 304 18920
rect 672 18880 681 18920
rect 1535 18124 1544 18164
rect 1912 18124 1921 18164
rect 295 17368 304 17408
rect 672 17368 681 17408
rect 1535 16612 1544 16652
rect 1912 16612 1921 16652
rect 295 15856 304 15896
rect 672 15856 681 15896
rect 1535 15100 1544 15140
rect 1912 15100 1921 15140
rect 295 14344 304 14384
rect 672 14344 681 14384
rect 1535 13588 1544 13628
rect 1912 13588 1921 13628
rect 295 12832 304 12872
rect 672 12832 681 12872
rect 1535 12076 1544 12116
rect 1912 12076 1921 12116
rect 295 11320 304 11360
rect 672 11320 681 11360
rect 1535 10564 1544 10604
rect 1912 10564 1921 10604
rect 295 9808 304 9848
rect 672 9808 681 9848
rect 1535 9052 1544 9092
rect 1912 9052 1921 9092
rect 295 8296 304 8336
rect 672 8296 681 8336
rect 1535 7540 1544 7580
rect 1912 7540 1921 7580
rect 295 6784 304 6824
rect 672 6784 681 6824
rect 1535 6028 1544 6068
rect 1912 6028 1921 6068
rect 295 5272 304 5312
rect 672 5272 681 5312
rect 1535 4516 1544 4556
rect 1912 4516 1921 4556
rect 295 3760 304 3800
rect 672 3760 681 3800
rect 1535 3004 1544 3044
rect 1912 3004 1921 3044
rect 295 2248 304 2288
rect 672 2248 681 2288
rect 1535 1492 1544 1532
rect 1912 1492 1921 1532
rect 295 736 304 776
rect 672 736 681 776
rect 1535 -20 1544 20
rect 1912 -20 1921 20
<< via4 >>
rect 1544 25684 1912 25724
rect 304 24928 672 24968
rect 1544 24172 1912 24212
rect 304 23416 672 23456
rect 1544 22660 1912 22700
rect 304 21904 672 21944
rect 1544 21148 1912 21188
rect 304 20392 672 20432
rect 1544 19636 1912 19676
rect 304 18880 672 18920
rect 1544 18124 1912 18164
rect 304 17368 672 17408
rect 1544 16612 1912 16652
rect 304 15856 672 15896
rect 1544 15100 1912 15140
rect 304 14344 672 14384
rect 1544 13588 1912 13628
rect 304 12832 672 12872
rect 1544 12076 1912 12116
rect 304 11320 672 11360
rect 1544 10564 1912 10604
rect 304 9808 672 9848
rect 1544 9052 1912 9092
rect 304 8296 672 8336
rect 1544 7540 1912 7580
rect 304 6784 672 6824
rect 1544 6028 1912 6068
rect 304 5272 672 5312
rect 1544 4516 1912 4556
rect 304 3760 672 3800
rect 1544 3004 1912 3044
rect 304 2248 672 2288
rect 1544 1492 1912 1532
rect 304 736 672 776
rect 1544 -20 1912 20
<< metal5 >>
rect 268 24968 708 25748
rect 268 24928 304 24968
rect 672 24928 708 24968
rect 268 23456 708 24928
rect 268 23416 304 23456
rect 672 23416 708 23456
rect 268 21944 708 23416
rect 268 21904 304 21944
rect 672 21904 708 21944
rect 268 20432 708 21904
rect 268 20392 304 20432
rect 672 20392 708 20432
rect 268 18920 708 20392
rect 268 18880 304 18920
rect 672 18880 708 18920
rect 268 17408 708 18880
rect 268 17368 304 17408
rect 672 17368 708 17408
rect 268 15896 708 17368
rect 268 15856 304 15896
rect 672 15856 708 15896
rect 268 14384 708 15856
rect 268 14344 304 14384
rect 672 14344 708 14384
rect 268 12872 708 14344
rect 268 12832 304 12872
rect 672 12832 708 12872
rect 268 11360 708 12832
rect 268 11320 304 11360
rect 672 11320 708 11360
rect 268 9848 708 11320
rect 268 9808 304 9848
rect 672 9808 708 9848
rect 268 8336 708 9808
rect 268 8296 304 8336
rect 672 8296 708 8336
rect 268 6824 708 8296
rect 268 6784 304 6824
rect 672 6784 708 6824
rect 268 5312 708 6784
rect 268 5272 304 5312
rect 672 5272 708 5312
rect 268 3800 708 5272
rect 268 3760 304 3800
rect 672 3760 708 3800
rect 268 2288 708 3760
rect 268 2248 304 2288
rect 672 2248 708 2288
rect 268 776 708 2248
rect 268 736 304 776
rect 672 736 708 776
rect 268 -44 708 736
rect 1508 25724 1948 25748
rect 1508 25684 1544 25724
rect 1912 25684 1948 25724
rect 1508 24212 1948 25684
rect 1508 24172 1544 24212
rect 1912 24172 1948 24212
rect 1508 22700 1948 24172
rect 1508 22660 1544 22700
rect 1912 22660 1948 22700
rect 1508 21188 1948 22660
rect 1508 21148 1544 21188
rect 1912 21148 1948 21188
rect 1508 19676 1948 21148
rect 1508 19636 1544 19676
rect 1912 19636 1948 19676
rect 1508 18164 1948 19636
rect 1508 18124 1544 18164
rect 1912 18124 1948 18164
rect 1508 16652 1948 18124
rect 1508 16612 1544 16652
rect 1912 16612 1948 16652
rect 1508 15140 1948 16612
rect 1508 15100 1544 15140
rect 1912 15100 1948 15140
rect 1508 13628 1948 15100
rect 1508 13588 1544 13628
rect 1912 13588 1948 13628
rect 1508 12116 1948 13588
rect 1508 12076 1544 12116
rect 1912 12076 1948 12116
rect 1508 10604 1948 12076
rect 1508 10564 1544 10604
rect 1912 10564 1948 10604
rect 1508 9092 1948 10564
rect 1508 9052 1544 9092
rect 1912 9052 1948 9092
rect 1508 7580 1948 9052
rect 1508 7540 1544 7580
rect 1912 7540 1948 7580
rect 1508 6068 1948 7540
rect 1508 6028 1544 6068
rect 1912 6028 1948 6068
rect 1508 4556 1948 6028
rect 1508 4516 1544 4556
rect 1912 4516 1948 4556
rect 1508 3044 1948 4516
rect 1508 3004 1544 3044
rect 1912 3004 1948 3044
rect 1508 1532 1948 3004
rect 1508 1492 1544 1532
rect 1912 1492 1948 1532
rect 1508 20 1948 1492
rect 1508 -20 1544 20
rect 1912 -20 1948 20
rect 1508 -44 1948 -20
use sg13g2_decap_8  FILLER_0_0
timestamp 1747491194
transform 1 0 288 0 1 0
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_7
timestamp 1747491194
transform 1 0 960 0 1 0
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_14
timestamp 1747491194
transform 1 0 1632 0 1 0
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_0
timestamp 1747491194
transform 1 0 288 0 -1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_7
timestamp 1747491194
transform 1 0 960 0 -1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_14
timestamp 1747491194
transform 1 0 1632 0 -1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_0
timestamp 1747491194
transform 1 0 288 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_7
timestamp 1747491194
transform 1 0 960 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_14
timestamp 1747491194
transform 1 0 1632 0 1 1512
box -48 -56 720 834
use sg13g2_fill_1  FILLER_3_0
timestamp 1747491194
transform 1 0 288 0 -1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_14
timestamp 1747491194
transform 1 0 1632 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_0
timestamp 1747491194
transform 1 0 288 0 1 3024
box -48 -56 720 834
use sg13g2_fill_1  FILLER_4_20
timestamp 1747491194
transform 1 0 2208 0 1 3024
box -48 -56 144 834
use sg13g2_fill_1  FILLER_5_0
timestamp 1747491194
transform 1 0 288 0 -1 4536
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_14
timestamp 1747491194
transform 1 0 1632 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_0
timestamp 1747491194
transform 1 0 288 0 1 4536
box -48 -56 720 834
use sg13g2_fill_1  FILLER_6_20
timestamp 1747491194
transform 1 0 2208 0 1 4536
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_0
timestamp 1747491194
transform 1 0 288 0 -1 6048
box -48 -56 720 834
use sg13g2_fill_1  FILLER_7_20
timestamp 1747491194
transform 1 0 2208 0 -1 6048
box -48 -56 144 834
use sg13g2_fill_1  FILLER_8_0
timestamp 1747491194
transform 1 0 288 0 1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_14
timestamp 1747491194
transform 1 0 1632 0 1 6048
box -48 -56 720 834
use sg13g2_decap_4  FILLER_9_0
timestamp 1747491194
transform 1 0 288 0 -1 7560
box -48 -56 432 834
use sg13g2_decap_4  FILLER_9_17
timestamp 1747491194
transform 1 0 1920 0 -1 7560
box -48 -56 432 834
use sg13g2_fill_1  FILLER_10_0
timestamp 1747491194
transform 1 0 288 0 1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_14
timestamp 1747491194
transform 1 0 1632 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_0
timestamp 1747491194
transform 1 0 288 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_7
timestamp 1747491194
transform 1 0 960 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_14
timestamp 1747491194
transform 1 0 1632 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_0
timestamp 1747491194
transform 1 0 288 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_7
timestamp 1747491194
transform 1 0 960 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_14
timestamp 1747491194
transform 1 0 1632 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_0
timestamp 1747491194
transform 1 0 288 0 -1 10584
box -48 -56 720 834
use sg13g2_fill_1  FILLER_13_20
timestamp 1747491194
transform 1 0 2208 0 -1 10584
box -48 -56 144 834
use sg13g2_fill_1  FILLER_14_0
timestamp 1747491194
transform 1 0 288 0 1 10584
box -48 -56 144 834
use sg13g2_decap_8  FILLER_14_14
timestamp 1747491194
transform 1 0 1632 0 1 10584
box -48 -56 720 834
use sg13g2_fill_1  FILLER_15_0
timestamp 1747491194
transform 1 0 288 0 -1 12096
box -48 -56 144 834
use sg13g2_decap_8  FILLER_15_14
timestamp 1747491194
transform 1 0 1632 0 -1 12096
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_0
timestamp 1747491194
transform 1 0 288 0 1 12096
box -48 -56 720 834
use sg13g2_fill_1  FILLER_16_20
timestamp 1747491194
transform 1 0 2208 0 1 12096
box -48 -56 144 834
use sg13g2_decap_8  FILLER_17_0
timestamp 1747491194
transform 1 0 288 0 -1 13608
box -48 -56 720 834
use sg13g2_fill_1  FILLER_17_20
timestamp 1747491194
transform 1 0 2208 0 -1 13608
box -48 -56 144 834
use sg13g2_fill_1  FILLER_18_0
timestamp 1747491194
transform 1 0 288 0 1 13608
box -48 -56 144 834
use sg13g2_decap_8  FILLER_18_14
timestamp 1747491194
transform 1 0 1632 0 1 13608
box -48 -56 720 834
use sg13g2_fill_1  FILLER_19_0
timestamp 1747491194
transform 1 0 288 0 -1 15120
box -48 -56 144 834
use sg13g2_decap_8  FILLER_19_14
timestamp 1747491194
transform 1 0 1632 0 -1 15120
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_0
timestamp 1747491194
transform 1 0 288 0 1 15120
box -48 -56 720 834
use sg13g2_fill_1  FILLER_20_20
timestamp 1747491194
transform 1 0 2208 0 1 15120
box -48 -56 144 834
use sg13g2_decap_8  FILLER_21_0
timestamp 1747491194
transform 1 0 288 0 -1 16632
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_7
timestamp 1747491194
transform 1 0 960 0 -1 16632
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_14
timestamp 1747491194
transform 1 0 1632 0 -1 16632
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_0
timestamp 1747491194
transform 1 0 288 0 1 16632
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_7
timestamp 1747491194
transform 1 0 960 0 1 16632
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_14
timestamp 1747491194
transform 1 0 1632 0 1 16632
box -48 -56 720 834
use sg13g2_fill_1  FILLER_23_0
timestamp 1747491194
transform 1 0 288 0 -1 18144
box -48 -56 144 834
use sg13g2_decap_8  FILLER_23_14
timestamp 1747491194
transform 1 0 1632 0 -1 18144
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_0
timestamp 1747491194
transform 1 0 288 0 1 18144
box -48 -56 720 834
use sg13g2_fill_1  FILLER_24_20
timestamp 1747491194
transform 1 0 2208 0 1 18144
box -48 -56 144 834
use sg13g2_fill_1  FILLER_25_0
timestamp 1747491194
transform 1 0 288 0 -1 19656
box -48 -56 144 834
use sg13g2_decap_8  FILLER_25_14
timestamp 1747491194
transform 1 0 1632 0 -1 19656
box -48 -56 720 834
use sg13g2_fill_1  FILLER_26_0
timestamp 1747491194
transform 1 0 288 0 1 19656
box -48 -56 144 834
use sg13g2_decap_8  FILLER_26_14
timestamp 1747491194
transform 1 0 1632 0 1 19656
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_0
timestamp 1747491194
transform 1 0 288 0 -1 21168
box -48 -56 720 834
use sg13g2_fill_1  FILLER_27_20
timestamp 1747491194
transform 1 0 2208 0 -1 21168
box -48 -56 144 834
use sg13g2_decap_8  FILLER_28_0
timestamp 1747491194
transform 1 0 288 0 1 21168
box -48 -56 720 834
use sg13g2_fill_1  FILLER_28_20
timestamp 1747491194
transform 1 0 2208 0 1 21168
box -48 -56 144 834
use sg13g2_fill_2  FILLER_29_0
timestamp 1747491194
transform 1 0 288 0 -1 22680
box -48 -56 240 834
use sg13g2_decap_4  FILLER_29_15
timestamp 1747491194
transform 1 0 1728 0 -1 22680
box -48 -56 432 834
use sg13g2_fill_2  FILLER_29_19
timestamp 1747491194
transform 1 0 2112 0 -1 22680
box -48 -56 240 834
use sg13g2_fill_1  FILLER_30_0
timestamp 1747491194
transform 1 0 288 0 1 22680
box -48 -56 144 834
use sg13g2_decap_8  FILLER_30_14
timestamp 1747491194
transform 1 0 1632 0 1 22680
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_0
timestamp 1747491194
transform 1 0 288 0 -1 24192
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_7
timestamp 1747491194
transform 1 0 960 0 -1 24192
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_14
timestamp 1747491194
transform 1 0 1632 0 -1 24192
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_0
timestamp 1747491194
transform 1 0 288 0 1 24192
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_7
timestamp 1747491194
transform 1 0 960 0 1 24192
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_14
timestamp 1747491194
transform 1 0 1632 0 1 24192
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_0
timestamp 1747491194
transform 1 0 288 0 -1 25704
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_7
timestamp 1747491194
transform 1 0 960 0 -1 25704
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_14
timestamp 1747491194
transform 1 0 1632 0 -1 25704
box -48 -56 720 834
use sg13g2_buf_8  rgb_buffer_cell\[0\]
timestamp 1747491194
transform -1 0 1632 0 1 7560
box -48 -56 1296 834
use sg13g2_buf_8  rgb_buffer_cell\[1\]
timestamp 1747491194
transform -1 0 1920 0 -1 7560
box -48 -56 1296 834
use sg13g2_buf_8  rgb_buffer_cell\[2\]
timestamp 1747491194
transform -1 0 1632 0 1 6048
box -48 -56 1296 834
use sg13g2_buf_8  rgb_buffer_cell\[3\]
timestamp 1747491194
transform -1 0 2208 0 -1 6048
box -48 -56 1296 834
use sg13g2_buf_8  rgb_buffer_cell\[4\]
timestamp 1747491194
transform -1 0 2208 0 1 4536
box -48 -56 1296 834
use sg13g2_buf_8  rgb_buffer_cell\[5\]
timestamp 1747491194
transform -1 0 1632 0 -1 4536
box -48 -56 1296 834
use sg13g2_buf_8  rgb_buffer_cell\[6\]
timestamp 1747491194
transform -1 0 2208 0 1 3024
box -48 -56 1296 834
use sg13g2_buf_8  rgb_buffer_cell\[7\]
timestamp 1747491194
transform -1 0 1632 0 -1 3024
box -48 -56 1296 834
use sg13g2_buf_8  rgb_buffer_cell\[8\]
timestamp 1747491194
transform -1 0 2208 0 1 15120
box -48 -56 1296 834
use sg13g2_buf_8  rgb_buffer_cell\[9\]
timestamp 1747491194
transform -1 0 1632 0 -1 15120
box -48 -56 1296 834
use sg13g2_buf_8  rgb_buffer_cell\[10\]
timestamp 1747491194
transform -1 0 1632 0 1 13608
box -48 -56 1296 834
use sg13g2_buf_8  rgb_buffer_cell\[11\]
timestamp 1747491194
transform -1 0 2208 0 -1 13608
box -48 -56 1296 834
use sg13g2_buf_8  rgb_buffer_cell\[12\]
timestamp 1747491194
transform -1 0 2208 0 1 12096
box -48 -56 1296 834
use sg13g2_buf_8  rgb_buffer_cell\[13\]
timestamp 1747491194
transform -1 0 1632 0 -1 12096
box -48 -56 1296 834
use sg13g2_buf_8  rgb_buffer_cell\[14\]
timestamp 1747491194
transform -1 0 1632 0 1 10584
box -48 -56 1296 834
use sg13g2_buf_8  rgb_buffer_cell\[15\]
timestamp 1747491194
transform -1 0 2208 0 -1 10584
box -48 -56 1296 834
use sg13g2_buf_8  rgb_buffer_cell\[16\]
timestamp 1747491194
transform -1 0 1632 0 1 22680
box -48 -56 1296 834
use sg13g2_buf_8  rgb_buffer_cell\[17\]
timestamp 1747491194
transform -1 0 1728 0 -1 22680
box -48 -56 1296 834
use sg13g2_buf_8  rgb_buffer_cell\[18\]
timestamp 1747491194
transform -1 0 2208 0 1 21168
box -48 -56 1296 834
use sg13g2_buf_8  rgb_buffer_cell\[19\]
timestamp 1747491194
transform -1 0 2208 0 -1 21168
box -48 -56 1296 834
use sg13g2_buf_8  rgb_buffer_cell\[20\]
timestamp 1747491194
transform -1 0 1632 0 1 19656
box -48 -56 1296 834
use sg13g2_buf_8  rgb_buffer_cell\[21\]
timestamp 1747491194
transform -1 0 1632 0 -1 19656
box -48 -56 1296 834
use sg13g2_buf_8  rgb_buffer_cell\[22\]
timestamp 1747491194
transform -1 0 2208 0 1 18144
box -48 -56 1296 834
use sg13g2_buf_8  rgb_buffer_cell\[23\]
timestamp 1747491194
transform -1 0 1632 0 -1 18144
box -48 -56 1296 834
<< labels >>
flabel metal5 s 1508 -44 1948 25748 0 FreeSans 3200 90 0 0 VGND
port 1 nsew
flabel metal5 s 268 -44 708 25748 0 FreeSans 3200 90 0 0 VPWR
port 2 nsew
flabel metal2 s 0 7604 100 7684 0 FreeSans 400 0 0 0 b[0]
port 3 nsew
flabel metal2 s 0 6848 100 6928 0 FreeSans 400 0 0 0 b[1]
port 4 nsew
flabel metal2 s 0 6092 100 6172 0 FreeSans 400 0 0 0 b[2]
port 5 nsew
flabel metal2 s 0 5336 100 5416 0 FreeSans 400 0 0 0 b[3]
port 6 nsew
flabel metal2 s 0 4580 100 4660 0 FreeSans 400 0 0 0 b[4]
port 7 nsew
flabel metal2 s 0 3824 100 3904 0 FreeSans 400 0 0 0 b[5]
port 8 nsew
flabel metal2 s 0 3068 100 3148 0 FreeSans 400 0 0 0 b[6]
port 9 nsew
flabel metal2 s 0 2312 100 2392 0 FreeSans 400 0 0 0 b[7]
port 10 nsew
flabel metal2 s 2500 7604 2600 7684 0 FreeSans 400 0 0 0 db[0]
port 11 nsew
flabel metal2 s 2500 7184 2600 7264 0 FreeSans 400 0 0 0 db[1]
port 12 nsew
flabel metal2 s 2500 6764 2600 6844 0 FreeSans 400 0 0 0 db[2]
port 13 nsew
flabel metal2 s 2500 6344 2600 6424 0 FreeSans 400 0 0 0 db[3]
port 14 nsew
flabel metal2 s 2500 5924 2600 6004 0 FreeSans 400 0 0 0 db[4]
port 15 nsew
flabel metal2 s 2500 5504 2600 5584 0 FreeSans 400 0 0 0 db[5]
port 16 nsew
flabel metal2 s 2500 5084 2600 5164 0 FreeSans 400 0 0 0 db[6]
port 17 nsew
flabel metal2 s 2500 4664 2600 4744 0 FreeSans 400 0 0 0 db[7]
port 18 nsew
flabel metal2 s 2500 14324 2600 14404 0 FreeSans 400 0 0 0 dg[0]
port 19 nsew
flabel metal2 s 2500 13904 2600 13984 0 FreeSans 400 0 0 0 dg[1]
port 20 nsew
flabel metal2 s 2500 13484 2600 13564 0 FreeSans 400 0 0 0 dg[2]
port 21 nsew
flabel metal2 s 2500 13064 2600 13144 0 FreeSans 400 0 0 0 dg[3]
port 22 nsew
flabel metal2 s 2500 12644 2600 12724 0 FreeSans 400 0 0 0 dg[4]
port 23 nsew
flabel metal2 s 2500 12224 2600 12304 0 FreeSans 400 0 0 0 dg[5]
port 24 nsew
flabel metal2 s 2500 11804 2600 11884 0 FreeSans 400 0 0 0 dg[6]
port 25 nsew
flabel metal2 s 2500 11384 2600 11464 0 FreeSans 400 0 0 0 dg[7]
port 26 nsew
flabel metal2 s 2500 21044 2600 21124 0 FreeSans 400 0 0 0 dr[0]
port 27 nsew
flabel metal2 s 2500 20624 2600 20704 0 FreeSans 400 0 0 0 dr[1]
port 28 nsew
flabel metal2 s 2500 20204 2600 20284 0 FreeSans 400 0 0 0 dr[2]
port 29 nsew
flabel metal2 s 2500 19784 2600 19864 0 FreeSans 400 0 0 0 dr[3]
port 30 nsew
flabel metal2 s 2500 19364 2600 19444 0 FreeSans 400 0 0 0 dr[4]
port 31 nsew
flabel metal2 s 2500 18944 2600 19024 0 FreeSans 400 0 0 0 dr[5]
port 32 nsew
flabel metal2 s 2500 18524 2600 18604 0 FreeSans 400 0 0 0 dr[6]
port 33 nsew
flabel metal2 s 2500 18104 2600 18184 0 FreeSans 400 0 0 0 dr[7]
port 34 nsew
flabel metal2 s 0 15164 100 15244 0 FreeSans 400 0 0 0 g[0]
port 35 nsew
flabel metal2 s 0 14408 100 14488 0 FreeSans 400 0 0 0 g[1]
port 36 nsew
flabel metal2 s 0 13652 100 13732 0 FreeSans 400 0 0 0 g[2]
port 37 nsew
flabel metal2 s 0 12896 100 12976 0 FreeSans 400 0 0 0 g[3]
port 38 nsew
flabel metal2 s 0 12140 100 12220 0 FreeSans 400 0 0 0 g[4]
port 39 nsew
flabel metal2 s 0 11384 100 11464 0 FreeSans 400 0 0 0 g[5]
port 40 nsew
flabel metal2 s 0 10628 100 10708 0 FreeSans 400 0 0 0 g[6]
port 41 nsew
flabel metal2 s 0 9872 100 9952 0 FreeSans 400 0 0 0 g[7]
port 42 nsew
flabel metal2 s 0 22724 100 22804 0 FreeSans 400 0 0 0 r[0]
port 43 nsew
flabel metal2 s 0 21968 100 22048 0 FreeSans 400 0 0 0 r[1]
port 44 nsew
flabel metal2 s 0 21212 100 21292 0 FreeSans 400 0 0 0 r[2]
port 45 nsew
flabel metal2 s 0 20456 100 20536 0 FreeSans 400 0 0 0 r[3]
port 46 nsew
flabel metal2 s 0 19700 100 19780 0 FreeSans 400 0 0 0 r[4]
port 47 nsew
flabel metal2 s 0 18944 100 19024 0 FreeSans 400 0 0 0 r[5]
port 48 nsew
flabel metal2 s 0 18188 100 18268 0 FreeSans 400 0 0 0 r[6]
port 49 nsew
flabel metal2 s 0 17432 100 17512 0 FreeSans 400 0 0 0 r[7]
port 50 nsew
<< properties >>
string FIXED_BBOX 0 0 2600 26000
string GDS_END 109962
string GDS_FILE ../gds/rgb_buffers.gds
string GDS_START 18750
<< end >>
