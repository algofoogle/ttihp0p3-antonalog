magic
tech ihp-sg13g2
magscale 1 2
timestamp 1746816402
<< nwell >>
rect -48 350 912 834
<< pwell >>
rect 19 56 846 314
rect -26 -56 890 56
<< nmos >>
rect 114 140 140 288
rect 216 140 242 288
rect 420 140 446 288
rect 522 140 548 288
rect 624 140 650 288
rect 726 140 752 288
<< pmos >>
rect 114 412 140 636
rect 216 412 242 636
rect 420 412 446 636
rect 522 412 548 636
rect 624 412 650 636
rect 726 412 752 636
<< ndiff >>
rect 45 274 114 288
rect 45 242 60 274
rect 92 242 114 274
rect 45 186 114 242
rect 45 154 60 186
rect 92 154 114 186
rect 45 140 114 154
rect 140 274 216 288
rect 140 242 162 274
rect 194 242 216 274
rect 140 186 216 242
rect 140 154 162 186
rect 194 154 216 186
rect 140 140 216 154
rect 242 186 420 288
rect 242 154 264 186
rect 296 154 366 186
rect 398 154 420 186
rect 242 140 420 154
rect 446 274 522 288
rect 446 242 468 274
rect 500 242 522 274
rect 446 186 522 242
rect 446 154 468 186
rect 500 154 522 186
rect 446 140 522 154
rect 548 274 624 288
rect 548 242 570 274
rect 602 242 624 274
rect 548 186 624 242
rect 548 154 570 186
rect 602 154 624 186
rect 548 140 624 154
rect 650 274 726 288
rect 650 242 672 274
rect 704 242 726 274
rect 650 186 726 242
rect 650 154 672 186
rect 704 154 726 186
rect 650 140 726 154
rect 752 274 820 288
rect 752 242 774 274
rect 806 242 820 274
rect 752 186 820 242
rect 752 154 774 186
rect 806 154 820 186
rect 752 140 820 154
<< pdiff >>
rect 45 622 114 636
rect 45 590 60 622
rect 92 590 114 622
rect 45 543 114 590
rect 45 511 60 543
rect 92 511 114 543
rect 45 458 114 511
rect 45 426 60 458
rect 92 426 114 458
rect 45 412 114 426
rect 140 622 216 636
rect 140 590 162 622
rect 194 590 216 622
rect 140 543 216 590
rect 140 511 162 543
rect 194 511 216 543
rect 140 458 216 511
rect 140 426 162 458
rect 194 426 216 458
rect 140 412 216 426
rect 242 622 310 636
rect 242 590 264 622
rect 296 590 310 622
rect 242 543 310 590
rect 242 511 264 543
rect 296 511 310 543
rect 242 412 310 511
rect 352 622 420 636
rect 352 590 366 622
rect 398 590 420 622
rect 352 543 420 590
rect 352 511 366 543
rect 398 511 420 543
rect 352 412 420 511
rect 446 543 522 636
rect 446 511 468 543
rect 500 511 522 543
rect 446 458 522 511
rect 446 426 468 458
rect 500 426 522 458
rect 446 412 522 426
rect 548 622 624 636
rect 548 590 570 622
rect 602 590 624 622
rect 548 543 624 590
rect 548 511 570 543
rect 602 511 624 543
rect 548 458 624 511
rect 548 426 570 458
rect 602 426 624 458
rect 548 412 624 426
rect 650 543 726 636
rect 650 511 672 543
rect 704 511 726 543
rect 650 458 726 511
rect 650 426 672 458
rect 704 426 726 458
rect 650 412 726 426
rect 752 622 820 636
rect 752 590 774 622
rect 806 590 820 622
rect 752 543 820 590
rect 752 511 774 543
rect 806 511 820 543
rect 752 458 820 511
rect 752 426 774 458
rect 806 426 820 458
rect 752 412 820 426
<< ndiffc >>
rect 60 242 92 274
rect 60 154 92 186
rect 162 242 194 274
rect 162 154 194 186
rect 264 154 296 186
rect 366 154 398 186
rect 468 242 500 274
rect 468 154 500 186
rect 570 242 602 274
rect 570 154 602 186
rect 672 242 704 274
rect 672 154 704 186
rect 774 242 806 274
rect 774 154 806 186
<< pdiffc >>
rect 60 590 92 622
rect 60 511 92 543
rect 60 426 92 458
rect 162 590 194 622
rect 162 511 194 543
rect 162 426 194 458
rect 264 590 296 622
rect 264 511 296 543
rect 366 590 398 622
rect 366 511 398 543
rect 468 511 500 543
rect 468 426 500 458
rect 570 590 602 622
rect 570 511 602 543
rect 570 426 602 458
rect 672 511 704 543
rect 672 426 704 458
rect 774 590 806 622
rect 774 511 806 543
rect 774 426 806 458
<< psubdiff >>
rect 0 16 864 30
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 608 16
rect 640 -16 704 16
rect 736 -16 800 16
rect 832 -16 864 16
rect 0 -30 864 -16
<< nsubdiff >>
rect 0 772 864 786
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 608 772
rect 640 740 704 772
rect 736 740 800 772
rect 832 740 864 772
rect 0 726 864 740
<< psubdiffcont >>
rect 32 -16 64 16
rect 128 -16 160 16
rect 224 -16 256 16
rect 320 -16 352 16
rect 416 -16 448 16
rect 512 -16 544 16
rect 608 -16 640 16
rect 704 -16 736 16
rect 800 -16 832 16
<< nsubdiffcont >>
rect 32 740 64 772
rect 128 740 160 772
rect 224 740 256 772
rect 320 740 352 772
rect 416 740 448 772
rect 512 740 544 772
rect 608 740 640 772
rect 704 740 736 772
rect 800 740 832 772
<< poly >>
rect 114 636 140 672
rect 216 636 242 672
rect 420 636 446 672
rect 522 636 548 672
rect 624 636 650 672
rect 726 636 752 672
rect 114 380 140 412
rect 216 380 242 412
rect 420 380 446 412
rect 522 380 548 412
rect 624 380 650 412
rect 726 380 752 412
rect 97 366 259 380
rect 97 334 163 366
rect 195 334 259 366
rect 97 320 259 334
rect 351 366 565 380
rect 351 334 369 366
rect 401 334 565 366
rect 351 320 565 334
rect 607 366 817 380
rect 607 334 770 366
rect 802 334 817 366
rect 607 320 817 334
rect 114 288 140 320
rect 216 288 242 320
rect 420 288 446 320
rect 522 288 548 320
rect 624 288 650 320
rect 726 288 752 320
rect 114 104 140 140
rect 216 104 242 140
rect 420 104 446 140
rect 522 104 548 140
rect 624 104 650 140
rect 726 104 752 140
<< polycont >>
rect 163 334 195 366
rect 369 334 401 366
rect 770 334 802 366
<< metal1 >>
rect 0 772 864 800
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 608 772
rect 640 740 704 772
rect 736 740 800 772
rect 832 740 864 772
rect 0 712 864 740
rect 50 622 102 712
rect 50 590 60 622
rect 92 590 102 622
rect 50 543 102 590
rect 50 511 60 543
rect 92 511 102 543
rect 50 458 102 511
rect 50 426 60 458
rect 92 426 102 458
rect 50 416 102 426
rect 152 622 204 632
rect 152 590 162 622
rect 194 590 204 622
rect 152 543 204 590
rect 152 511 162 543
rect 194 511 204 543
rect 152 468 204 511
rect 254 622 306 712
rect 254 590 264 622
rect 296 590 306 622
rect 254 543 306 590
rect 254 511 264 543
rect 296 511 306 543
rect 254 504 306 511
rect 356 622 816 641
rect 356 590 366 622
rect 398 590 570 622
rect 602 590 774 622
rect 806 590 816 622
rect 356 589 816 590
rect 356 543 408 589
rect 356 511 366 543
rect 398 511 408 543
rect 356 504 408 511
rect 458 543 510 553
rect 458 511 468 543
rect 500 511 510 543
rect 458 468 510 511
rect 152 458 510 468
rect 152 426 162 458
rect 194 426 468 458
rect 500 426 510 458
rect 152 425 510 426
rect 560 543 612 589
rect 560 511 570 543
rect 602 511 612 543
rect 560 458 612 511
rect 560 426 570 458
rect 602 426 612 458
rect 560 416 612 426
rect 662 543 714 553
rect 662 511 672 543
rect 704 511 714 543
rect 662 458 714 511
rect 662 426 672 458
rect 704 426 714 458
rect 97 366 259 380
rect 97 334 163 366
rect 195 334 259 366
rect 97 315 259 334
rect 319 366 415 380
rect 662 372 714 426
rect 764 543 816 589
rect 764 511 774 543
rect 806 511 816 543
rect 764 458 816 511
rect 764 426 774 458
rect 806 426 816 458
rect 764 416 816 426
rect 319 334 369 366
rect 401 334 415 366
rect 319 315 415 334
rect 458 320 714 372
rect 458 275 510 320
rect 50 274 102 275
rect 50 242 60 274
rect 92 242 102 274
rect 50 186 102 242
rect 50 154 60 186
rect 92 154 102 186
rect 50 44 102 154
rect 152 274 510 275
rect 152 242 162 274
rect 194 242 468 274
rect 500 242 510 274
rect 152 235 510 242
rect 152 186 204 235
rect 152 154 162 186
rect 194 154 204 186
rect 152 144 204 154
rect 254 186 408 196
rect 254 154 264 186
rect 296 154 366 186
rect 398 154 408 186
rect 254 44 408 154
rect 458 186 510 235
rect 458 154 468 186
rect 500 154 510 186
rect 458 144 510 154
rect 560 274 612 284
rect 560 242 570 274
rect 602 242 612 274
rect 560 186 612 242
rect 560 154 570 186
rect 602 154 612 186
rect 560 44 612 154
rect 662 274 714 320
rect 764 366 833 380
rect 764 334 770 366
rect 802 334 833 366
rect 764 315 833 334
rect 662 242 672 274
rect 704 242 714 274
rect 662 186 714 242
rect 662 154 672 186
rect 704 154 714 186
rect 662 144 714 154
rect 764 274 816 275
rect 764 242 774 274
rect 806 242 816 274
rect 764 186 816 242
rect 764 154 774 186
rect 806 154 816 186
rect 764 44 816 154
rect 0 16 865 44
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 608 16
rect 640 -16 704 16
rect 736 -16 800 16
rect 832 -16 865 16
rect 0 -44 865 -16
<< labels >>
flabel metal1 s 0 712 864 800 0 FreeSans 500 0 0 0 VDD
port 4 nsew
flabel metal1 s 662 144 714 553 0 FreeSans 500 0 0 0 Y
port 3 nsew
flabel metal1 s 319 315 415 380 0 FreeSans 500 0 0 0 B
port 1 nsew
flabel metal1 s 97 315 259 380 0 FreeSans 500 0 0 0 A
port 6 nsew
flabel metal1 s 0 -44 864 44 0 FreeSans 500 0 0 0 VSS
port 5 nsew
flabel metal1 s 764 315 833 380 0 FreeSans 500 0 0 0 C
port 2 nsew
<< properties >>
string FIXED_BBOX 0 0 864 756
string GDS_END 237652
string GDS_FILE ../gds/controller.gds
string GDS_START 231296
<< end >>
