magic
tech ihp-sg13g2
timestamp 1747537721
<< nwell >>
rect -24 175 264 417
<< pwell >>
rect 0 28 223 146
rect -13 -28 253 28
<< nmos >>
rect 47 78 60 133
rect 132 59 145 133
rect 163 59 176 133
<< pmos >>
rect 47 206 60 290
rect 101 206 114 318
rect 152 206 165 318
<< ndiff >>
rect 13 113 47 133
rect 13 97 20 113
rect 36 97 47 113
rect 13 78 47 97
rect 60 100 132 133
rect 60 84 71 100
rect 87 99 132 100
rect 87 84 105 99
rect 60 83 105 84
rect 121 83 132 99
rect 60 78 132 83
rect 67 59 132 78
rect 145 59 163 133
rect 176 126 210 133
rect 176 110 187 126
rect 203 110 210 126
rect 176 82 210 110
rect 176 66 187 82
rect 203 66 210 82
rect 176 59 210 66
<< pdiff >>
rect 67 309 101 318
rect 67 293 74 309
rect 90 293 101 309
rect 67 290 101 293
rect 13 283 47 290
rect 13 267 20 283
rect 36 267 47 283
rect 13 241 47 267
rect 13 225 20 241
rect 36 225 47 241
rect 13 206 47 225
rect 60 275 101 290
rect 60 259 74 275
rect 90 259 101 275
rect 60 206 101 259
rect 114 311 152 318
rect 114 295 125 311
rect 141 295 152 311
rect 114 275 152 295
rect 114 259 125 275
rect 141 259 152 275
rect 114 206 152 259
rect 165 311 199 318
rect 165 295 176 311
rect 192 295 199 311
rect 165 206 199 295
<< ndiffc >>
rect 20 97 36 113
rect 71 84 87 100
rect 105 83 121 99
rect 187 110 203 126
rect 187 66 203 82
<< pdiffc >>
rect 74 293 90 309
rect 20 267 36 283
rect 20 225 36 241
rect 74 259 90 275
rect 125 295 141 311
rect 125 259 141 275
rect 176 295 192 311
<< psubdiff >>
rect 0 8 240 15
rect 0 -8 16 8
rect 32 -8 64 8
rect 80 -8 112 8
rect 128 -8 160 8
rect 176 -8 208 8
rect 224 -8 240 8
rect 0 -15 240 -8
<< nsubdiff >>
rect 0 386 240 393
rect 0 370 16 386
rect 32 370 64 386
rect 80 370 112 386
rect 128 370 160 386
rect 176 370 208 386
rect 224 370 240 386
rect 0 363 240 370
<< psubdiffcont >>
rect 16 -8 32 8
rect 64 -8 80 8
rect 112 -8 128 8
rect 160 -8 176 8
rect 208 -8 224 8
<< nsubdiffcont >>
rect 16 370 32 386
rect 64 370 80 386
rect 112 370 128 386
rect 160 370 176 386
rect 208 370 224 386
<< poly >>
rect 101 318 114 336
rect 152 318 165 336
rect 47 290 60 308
rect 47 185 60 206
rect 10 176 77 185
rect 10 160 18 176
rect 34 160 52 176
rect 68 160 77 176
rect 10 152 77 160
rect 101 183 114 206
rect 152 192 165 206
rect 101 176 131 183
rect 152 177 193 192
rect 101 160 108 176
rect 124 160 131 176
rect 101 154 131 160
rect 163 176 193 177
rect 163 160 170 176
rect 186 160 193 176
rect 47 133 60 152
rect 101 140 145 154
rect 132 133 145 140
rect 163 152 193 160
rect 163 133 176 152
rect 47 60 60 78
rect 132 41 145 59
rect 163 41 176 59
<< polycont >>
rect 18 160 34 176
rect 52 160 68 176
rect 108 160 124 176
rect 170 160 186 176
<< metal1 >>
rect 0 386 240 400
rect 0 370 16 386
rect 32 370 64 386
rect 80 370 112 386
rect 128 370 160 386
rect 176 370 208 386
rect 224 370 240 386
rect 0 356 240 370
rect 73 309 91 356
rect 73 293 74 309
rect 90 293 91 309
rect 19 283 38 290
rect 19 267 20 283
rect 36 267 38 283
rect 19 241 38 267
rect 73 275 91 293
rect 73 259 74 275
rect 90 259 91 275
rect 73 254 91 259
rect 120 311 146 312
rect 120 295 125 311
rect 141 295 146 311
rect 120 275 146 295
rect 171 311 197 356
rect 171 295 176 311
rect 192 295 197 311
rect 171 293 197 295
rect 120 259 125 275
rect 141 268 146 275
rect 141 259 225 268
rect 120 251 225 259
rect 19 225 20 241
rect 36 233 38 241
rect 36 225 189 233
rect 19 217 189 225
rect 10 176 77 189
rect 10 160 18 176
rect 34 160 52 176
rect 68 160 77 176
rect 10 153 77 160
rect 101 176 133 194
rect 101 160 108 176
rect 124 160 133 176
rect 162 176 189 217
rect 162 170 170 176
rect 101 155 133 160
rect 151 160 170 170
rect 186 160 189 176
rect 151 152 189 160
rect 151 135 168 152
rect 15 119 168 135
rect 208 131 225 251
rect 186 126 225 131
rect 15 113 41 119
rect 15 97 20 113
rect 36 97 41 113
rect 186 110 187 126
rect 203 110 225 126
rect 15 92 41 97
rect 66 84 71 100
rect 87 99 126 100
rect 87 84 105 99
rect 66 83 105 84
rect 121 83 126 99
rect 66 22 126 83
rect 186 82 225 110
rect 186 66 187 82
rect 203 66 225 82
rect 186 61 225 66
rect 0 8 240 22
rect 0 -8 16 8
rect 32 -8 64 8
rect 80 -8 112 8
rect 128 -8 160 8
rect 176 -8 208 8
rect 224 -8 240 8
rect 0 -22 240 -8
<< labels >>
flabel metal1 s 0 -22 240 22 0 FreeSans 200 0 0 0 VSS
port 2 nsew
flabel metal1 s 10 153 77 189 0 FreeSans 200 0 0 0 A_N
port 3 nsew
flabel metal1 s 186 61 225 131 0 FreeSans 200 0 0 0 Y
port 4 nsew
flabel metal1 s 101 155 133 194 0 FreeSans 200 0 0 0 B
port 5 nsew
flabel metal1 s 0 356 240 400 0 FreeSans 200 0 0 0 VDD
port 6 nsew
<< properties >>
string FIXED_BBOX 0 0 240 378
string GDS_END 118104
string GDS_FILE ../gds/controller.gds
string GDS_START 113616
<< end >>
