magic
tech ihp-sg13g2
magscale 1 2
timestamp 1747537721
<< nwell >>
rect -48 350 432 834
<< pwell >>
rect 49 56 325 292
rect -26 -56 410 56
<< nmos >>
rect 143 118 169 266
rect 205 118 231 266
<< pmos >>
rect 128 412 154 636
rect 230 412 256 636
<< ndiff >>
rect 75 245 143 266
rect 75 213 89 245
rect 121 213 143 245
rect 75 166 143 213
rect 75 134 89 166
rect 121 134 143 166
rect 75 118 143 134
rect 169 118 205 266
rect 231 245 299 266
rect 231 213 253 245
rect 285 213 299 245
rect 231 166 299 213
rect 231 134 253 166
rect 285 134 299 166
rect 231 118 299 134
<< pdiff >>
rect 60 622 128 636
rect 60 590 74 622
rect 106 590 128 622
rect 60 540 128 590
rect 60 508 74 540
rect 106 508 128 540
rect 60 460 128 508
rect 60 428 74 460
rect 106 428 128 460
rect 60 412 128 428
rect 154 622 230 636
rect 154 590 176 622
rect 208 590 230 622
rect 154 540 230 590
rect 154 508 176 540
rect 208 508 230 540
rect 154 460 230 508
rect 154 428 176 460
rect 208 428 230 460
rect 154 412 230 428
rect 256 622 324 636
rect 256 590 278 622
rect 310 590 324 622
rect 256 540 324 590
rect 256 508 278 540
rect 310 508 324 540
rect 256 460 324 508
rect 256 428 278 460
rect 310 428 324 460
rect 256 412 324 428
<< ndiffc >>
rect 89 213 121 245
rect 89 134 121 166
rect 253 213 285 245
rect 253 134 285 166
<< pdiffc >>
rect 74 590 106 622
rect 74 508 106 540
rect 74 428 106 460
rect 176 590 208 622
rect 176 508 208 540
rect 176 428 208 460
rect 278 590 310 622
rect 278 508 310 540
rect 278 428 310 460
<< psubdiff >>
rect 0 16 384 30
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 384 16
rect 0 -30 384 -16
<< nsubdiff >>
rect 0 772 384 786
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 384 772
rect 0 726 384 740
<< psubdiffcont >>
rect 32 -16 64 16
rect 128 -16 160 16
rect 224 -16 256 16
rect 320 -16 352 16
<< nsubdiffcont >>
rect 32 740 64 772
rect 128 740 160 772
rect 224 740 256 772
rect 320 740 352 772
<< poly >>
rect 128 636 154 672
rect 230 636 256 672
rect 128 354 154 412
rect 230 354 256 412
rect 66 337 169 354
rect 66 305 80 337
rect 112 305 169 337
rect 66 288 169 305
rect 143 266 169 288
rect 205 334 312 354
rect 205 302 266 334
rect 298 302 312 334
rect 205 288 312 302
rect 205 266 231 288
rect 143 82 169 118
rect 205 82 231 118
<< polycont >>
rect 80 305 112 337
rect 266 302 298 334
<< metal1 >>
rect 0 772 384 800
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 384 772
rect 0 712 384 740
rect 64 622 116 712
rect 64 590 74 622
rect 106 590 116 622
rect 64 540 116 590
rect 64 508 74 540
rect 106 508 116 540
rect 64 460 116 508
rect 64 428 74 460
rect 106 428 116 460
rect 64 425 116 428
rect 166 622 218 625
rect 166 590 176 622
rect 208 590 218 622
rect 166 540 218 590
rect 166 508 176 540
rect 208 508 218 540
rect 166 460 218 508
rect 166 428 176 460
rect 208 428 218 460
rect 58 337 124 362
rect 58 305 80 337
rect 112 305 124 337
rect 58 288 124 305
rect 166 273 218 428
rect 268 622 320 712
rect 268 590 278 622
rect 310 590 320 622
rect 268 540 320 590
rect 268 508 278 540
rect 310 508 320 540
rect 268 460 320 508
rect 268 428 278 460
rect 310 428 320 460
rect 268 425 320 428
rect 254 334 320 362
rect 254 302 266 334
rect 298 302 320 334
rect 254 288 320 302
rect 172 249 218 273
rect 79 245 131 249
rect 79 213 89 245
rect 121 213 131 245
rect 79 166 131 213
rect 172 245 295 249
rect 172 213 253 245
rect 285 213 295 245
rect 172 212 295 213
rect 79 134 89 166
rect 121 134 131 166
rect 79 44 131 134
rect 243 166 295 212
rect 243 134 253 166
rect 285 134 295 166
rect 243 131 295 134
rect 0 16 384 44
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 384 16
rect 0 -44 384 -16
<< labels >>
flabel metal1 s 166 273 218 625 0 FreeSans 400 0 0 0 Y
port 2 nsew
flabel metal1 s 0 712 384 800 0 FreeSans 400 0 0 0 VDD
port 3 nsew
flabel metal1 s 254 288 320 362 0 FreeSans 400 0 0 0 A
port 4 nsew
flabel metal1 s 0 -44 384 44 0 FreeSans 400 0 0 0 VSS
port 5 nsew
flabel metal1 s 58 288 124 362 0 FreeSans 400 0 0 0 B
port 6 nsew
<< properties >>
string FIXED_BBOX 0 0 384 756
string GDS_END 73720
string GDS_FILE ../gds/controller.gds
string GDS_START 69874
<< end >>
