magic
tech ihp-sg13g2
timestamp 1746839677
<< pwell >>
rect -1401 -512 2631 528
<< psubdiff >>
rect -1370 490 2600 497
rect -1370 474 -1324 490
rect 2554 474 2600 490
rect -1370 467 2600 474
rect -1370 451 -1340 467
rect -1370 -435 -1363 451
rect -1347 -435 -1340 451
rect -1370 -451 -1340 -435
rect 2570 451 2600 467
rect 2570 -435 2577 451
rect 2593 -435 2600 451
rect 2570 -451 2600 -435
rect -1370 -458 2600 -451
rect -1370 -474 -1324 -458
rect 2554 -474 2600 -458
rect -1370 -481 2600 -474
<< psubdiffcont >>
rect -1324 474 2554 490
rect -1363 -435 -1347 451
rect 2577 -435 2593 451
rect -1324 -474 2554 -458
<< metal1 >>
rect -1363 474 -1324 490
rect 2554 474 2593 490
rect -1363 451 -1347 474
rect -1363 -458 -1347 -435
rect 2577 451 2593 474
rect 2577 -458 2593 -435
rect -1363 -474 -1324 -458
rect 2554 -474 2593 -458
use rhigh  rhigh_0
array 0 24 148 0 0 686
timestamp 1746838591
transform 1 0 -1208 0 1 -284
box 0 -43 100 643
<< labels >>
rlabel psubdiffcont 0 -466 0 -466 0 B
port 1 nsew
<< end >>
