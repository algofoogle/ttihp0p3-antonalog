magic
tech ihp-sg13g2
magscale 1 2
timestamp 1747056179
<< metal1 >>
rect 2026 30244 3192 30322
rect 2026 30118 2268 30244
rect 2936 30118 3192 30244
rect 2026 29124 2148 30118
rect 3040 30040 3192 30118
rect 4340 30118 4950 30256
rect 4340 30040 4496 30118
rect 2420 29730 2768 30014
rect 3040 29910 4496 30040
rect 3040 29750 3276 29910
rect 3484 29834 3630 29910
rect 3944 29882 4496 29910
rect 4768 30040 4950 30118
rect 4768 29916 7132 30040
rect 4768 29882 6184 29916
rect 3944 29750 4314 29882
rect 2420 29124 2768 29500
rect 3040 29124 3262 29750
rect 3652 29596 3846 29680
rect 3534 29124 3846 29596
rect 4118 29652 4314 29750
rect 4982 29876 6184 29882
rect 4982 29756 5250 29876
rect 5918 29756 6184 29876
rect 6392 29840 6538 29916
rect 6852 29756 7132 29916
rect 4982 29652 5174 29756
rect 4118 29124 4496 29652
rect 4768 29262 5174 29652
rect 5446 29354 5724 29646
rect 5996 29262 6170 29756
rect 6560 29602 6754 29686
rect 4768 29124 5258 29262
rect 5926 29130 6170 29262
rect 6442 29130 6754 29602
rect 7026 29130 7132 29756
rect 5926 29124 7132 29130
rect 2026 29012 7132 29124
rect 2420 28876 2770 28888
rect 2226 28846 2770 28876
rect 2226 27664 2252 28846
rect 2556 28154 2770 28846
rect 2556 27664 2576 28154
rect 2226 27634 2576 27664
rect 2512 27419 2644 27420
rect 2512 27307 2521 27419
rect 2635 27307 2644 27419
rect 2512 27306 2644 27307
rect 4069 26514 4187 26515
rect 4069 26416 4078 26514
rect 4178 26416 4187 26514
rect 4069 26415 4187 26416
rect 2504 25711 2629 25712
rect 2504 25606 2513 25711
rect 2620 25606 2629 25711
rect 2504 25605 2629 25606
rect 4062 24811 4194 24812
rect 4062 24699 4071 24811
rect 4185 24699 4194 24811
rect 4062 24698 4194 24699
rect 2496 23915 2637 23916
rect 2496 23794 2505 23915
rect 2628 23794 2637 23915
rect 2496 23793 2637 23794
rect 4070 23025 4202 23026
rect 4070 22913 4079 23025
rect 4193 22913 4202 23025
rect 4070 22912 4202 22913
rect 2511 22118 2627 22127
rect 2511 22002 2512 22118
rect 2626 22002 2627 22118
rect 2511 21993 2627 22002
rect 4047 21696 4227 21705
rect 4047 21516 4048 21696
rect 4226 21516 4227 21696
rect 4047 21507 4227 21516
rect 4062 21253 4203 21254
rect 4062 21132 4071 21253
rect 4194 21132 4203 21253
rect 4062 21131 4203 21132
rect 2162 20634 4374 20992
rect 2162 19794 2734 20634
rect 2162 19774 4374 19794
rect 2114 19568 4374 19774
rect 2114 18988 2320 19568
rect 2656 19414 4374 19568
rect 2830 19312 4374 19414
rect 2114 18944 2656 18988
rect 4051 12464 4231 12473
rect 4051 12284 4052 12464
rect 4230 12284 4231 12464
rect 4051 12275 4231 12284
rect 2162 11394 4374 11752
rect 2162 10554 2734 11394
rect 2162 10366 4374 10554
rect 2162 10072 2252 10366
rect 2226 9184 2252 10072
rect 2556 10072 4374 10366
rect 2556 9674 2770 10072
rect 2556 9184 2576 9674
rect 2226 9154 2576 9184
rect 4047 3204 4227 3213
rect 4047 3024 4048 3204
rect 4226 3024 4227 3204
rect 4047 3015 4227 3024
rect 2276 2314 4398 2494
rect 2276 2012 2316 2314
rect 4358 2012 4398 2314
rect 2276 1972 4398 2012
<< via1 >>
rect 2252 27664 2556 28846
rect 2521 27307 2635 27419
rect 4078 26416 4178 26514
rect 2513 25606 2620 25711
rect 4071 24699 4185 24811
rect 2505 23794 2628 23915
rect 4079 22913 4193 23025
rect 2512 22002 2626 22118
rect 4048 21516 4226 21696
rect 4071 21132 4194 21253
rect 2320 18988 2656 19568
rect 2521 18067 2635 18179
rect 4078 17176 4178 17274
rect 2513 16366 2620 16471
rect 4071 15459 4185 15571
rect 2505 14554 2628 14675
rect 4079 13673 4193 13785
rect 2512 12762 2626 12878
rect 4052 12284 4230 12464
rect 4071 11892 4194 12013
rect 2252 9184 2556 10366
rect 2521 8827 2635 8939
rect 4078 7936 4178 8034
rect 2513 7126 2620 7231
rect 4071 6219 4185 6331
rect 2505 5314 2628 5435
rect 4079 4433 4193 4545
rect 2512 3522 2626 3638
rect 4048 3024 4226 3204
rect 4071 2652 4194 2773
rect 2316 2012 4358 2314
<< metal2 >>
rect 2026 30244 3192 30322
rect 2026 30118 2268 30244
rect 2936 30118 3192 30244
rect 2026 29124 2148 30118
rect 3040 30040 3192 30118
rect 4340 30118 4950 30256
rect 4340 30040 4496 30118
rect 2420 29730 2768 30014
rect 3040 29910 4496 30040
rect 3040 29750 3276 29910
rect 3484 29834 3630 29910
rect 3944 29882 4496 29910
rect 4768 30040 4950 30118
rect 4768 29916 7132 30040
rect 4768 29882 6184 29916
rect 3944 29750 4314 29882
rect 2420 29124 2768 29500
rect 3040 29124 3262 29750
rect 3652 29596 3846 29680
rect 3534 29124 3846 29596
rect 4118 29652 4314 29750
rect 4982 29876 6184 29882
rect 4982 29756 5250 29876
rect 5918 29756 6184 29876
rect 6392 29840 6538 29916
rect 6852 29756 7132 29916
rect 4982 29652 5174 29756
rect 4118 29124 4496 29652
rect 4768 29262 5174 29652
rect 5446 29354 5724 29646
rect 5996 29262 6170 29756
rect 6560 29602 6754 29686
rect 4768 29124 5258 29262
rect 5926 29130 6170 29262
rect 6442 29130 6754 29602
rect 7026 29130 7132 29756
rect 5926 29124 7132 29130
rect 2026 29012 7132 29124
rect 2216 28846 2596 28880
rect 2216 27664 2252 28846
rect 2556 27664 2596 28846
rect 2216 27624 2596 27664
rect 2521 27488 2635 27505
rect 2521 27419 4732 27488
rect 2635 27408 4732 27419
rect 2521 27298 2635 27307
rect 4078 26564 4178 26574
rect 4078 26514 4732 26564
rect 4178 26484 4732 26514
rect 4078 26407 4178 26416
rect 2513 25711 2620 25720
rect 2620 25606 4732 25640
rect 2513 25560 4732 25606
rect 2513 25547 2620 25560
rect 4071 24811 4185 24820
rect 4185 24699 4732 24716
rect 4071 24636 4732 24699
rect 4071 24619 4185 24636
rect 2505 23915 2628 23924
rect 2505 23792 2628 23794
rect 2505 23712 4732 23792
rect 2505 23691 2628 23712
rect 7176 23460 7458 23540
rect 7176 23040 7458 23120
rect 4079 23025 4193 23034
rect 4079 22868 4193 22913
rect 4079 22788 4732 22868
rect 4079 22771 4193 22788
rect 7176 22620 7458 22700
rect 7176 22200 7458 22280
rect 2500 22002 2512 22118
rect 2626 22100 2780 22118
rect 2626 22020 4732 22100
rect 2626 22002 2780 22020
rect 1960 21976 2140 21985
rect 4652 21864 4732 22020
rect 1960 21696 2140 21796
rect 7176 21780 7458 21860
rect 1960 21516 4048 21696
rect 4226 21516 4235 21696
rect 7176 21360 7458 21440
rect 4071 21253 4194 21262
rect 4071 21020 4194 21132
rect 4071 20940 4732 21020
rect 7176 20940 7458 21020
rect 4071 20919 4194 20940
rect 7176 20520 7458 20600
rect 2240 19606 2736 19646
rect 1955 18628 1964 18808
rect 2144 18628 2153 18808
rect 1964 12464 2144 18628
rect 2240 18424 2280 19606
rect 2696 18424 2736 19606
rect 2240 18384 2736 18424
rect 2521 18248 2635 18265
rect 2521 18179 4732 18248
rect 2635 18168 4732 18179
rect 2521 18058 2635 18067
rect 4078 17324 4178 17334
rect 4078 17274 4732 17324
rect 4178 17244 4732 17274
rect 4078 17167 4178 17176
rect 7176 16740 7458 16820
rect 2513 16471 2620 16480
rect 2620 16366 4732 16400
rect 2513 16320 4732 16366
rect 7176 16320 7458 16400
rect 2513 16307 2620 16320
rect 7176 15900 7458 15980
rect 4071 15571 4185 15580
rect 7176 15480 7458 15560
rect 4185 15459 4732 15476
rect 4071 15396 4732 15459
rect 4071 15379 4185 15396
rect 7176 15060 7458 15140
rect 2505 14675 2628 14684
rect 7176 14640 7458 14720
rect 2505 14552 2628 14554
rect 2505 14472 4732 14552
rect 2505 14451 2628 14472
rect 7176 14220 7458 14300
rect 7176 13800 7458 13880
rect 4079 13785 4193 13794
rect 4079 13628 4193 13673
rect 4079 13548 4732 13628
rect 4079 13531 4193 13548
rect 2500 12762 2512 12878
rect 2626 12860 2780 12878
rect 2626 12780 4732 12860
rect 2626 12762 2780 12780
rect 4652 12624 4732 12780
rect 1964 12284 4052 12464
rect 4230 12284 4239 12464
rect 4071 12013 4194 12022
rect 4071 11780 4194 11892
rect 4071 11700 4732 11780
rect 4071 11679 4194 11700
rect 2216 10366 2596 10400
rect 2216 9184 2252 10366
rect 2556 9184 2596 10366
rect 7176 10020 7458 10100
rect 7176 9600 7458 9680
rect 2216 9144 2596 9184
rect 7176 9180 7458 9260
rect 2521 9008 2635 9025
rect 2521 8939 4732 9008
rect 2635 8928 4732 8939
rect 2521 8818 2635 8827
rect 7176 8760 7458 8840
rect 7176 8340 7458 8420
rect 4078 8084 4178 8094
rect 4078 8034 4732 8084
rect 4178 8004 4732 8034
rect 4078 7927 4178 7936
rect 7176 7920 7458 8000
rect 7176 7500 7458 7580
rect 2513 7231 2620 7240
rect 2620 7126 4732 7160
rect 2513 7080 4732 7126
rect 7176 7080 7458 7160
rect 2513 7067 2620 7080
rect 4071 6331 4185 6340
rect 4185 6219 4732 6236
rect 4071 6156 4732 6219
rect 4071 6139 4185 6156
rect 2505 5435 2628 5444
rect 2505 5312 2628 5314
rect 2505 5232 4732 5312
rect 2505 5211 2628 5232
rect 4079 4545 4193 4554
rect 4079 4388 4193 4433
rect 4079 4308 4732 4388
rect 4079 4291 4193 4308
rect 2500 3522 2512 3638
rect 2626 3620 2780 3638
rect 2626 3540 4732 3620
rect 2626 3522 2780 3540
rect 4652 3384 4732 3540
rect 1660 3204 1840 3213
rect 1840 3024 4048 3204
rect 4226 3024 4235 3204
rect 1660 3015 1840 3024
rect 4071 2773 4194 2782
rect 4071 2540 4194 2652
rect 4071 2460 4732 2540
rect 4071 2439 4194 2460
rect 2276 2314 4398 2354
rect 2276 2012 2316 2314
rect 4358 2012 4398 2314
rect 2276 1972 4398 2012
<< via2 >>
rect 2252 27664 2556 28846
rect 1960 21796 2140 21976
rect 1964 18628 2144 18808
rect 2280 19568 2696 19606
rect 2280 18988 2320 19568
rect 2320 18988 2656 19568
rect 2656 18988 2696 19568
rect 2280 18424 2696 18988
rect 2252 9184 2556 10366
rect 1660 3024 1840 3204
rect 2316 2012 4358 2314
<< metal3 >>
rect 10502 30465 10621 30479
rect 10502 30373 10515 30465
rect 10607 30373 10621 30465
rect 2026 30244 3192 30322
rect 2026 30118 2268 30244
rect 2936 30118 3192 30244
rect 2026 29124 2148 30118
rect 3040 30040 3192 30118
rect 4340 30118 4950 30256
rect 4340 30040 4496 30118
rect 2420 29730 2768 30014
rect 3040 29910 4496 30040
rect 3040 29750 3276 29910
rect 3484 29834 3630 29910
rect 3944 29882 4496 29910
rect 4768 30040 4950 30118
rect 4768 29916 7132 30040
rect 10502 30019 10621 30373
rect 11270 30465 11389 30479
rect 11270 30373 11283 30465
rect 11375 30373 11389 30465
rect 11270 30019 11389 30373
rect 12038 30465 12157 30479
rect 12038 30373 12051 30465
rect 12143 30373 12157 30465
rect 12038 30019 12157 30373
rect 12806 30465 12925 30479
rect 12806 30373 12819 30465
rect 12911 30373 12925 30465
rect 12806 30019 12925 30373
rect 13574 30465 13693 30479
rect 13574 30373 13587 30465
rect 13679 30373 13693 30465
rect 13574 30019 13693 30373
rect 14342 30465 14461 30479
rect 14342 30373 14355 30465
rect 14447 30373 14461 30465
rect 14342 30019 14461 30373
rect 15110 30465 15229 30479
rect 15110 30373 15123 30465
rect 15215 30373 15229 30465
rect 15110 30019 15229 30373
rect 15878 30465 15997 30479
rect 15878 30373 15891 30465
rect 15983 30373 15997 30465
rect 15878 30019 15997 30373
rect 16646 30465 16765 30479
rect 16646 30373 16659 30465
rect 16751 30373 16765 30465
rect 16646 30019 16765 30373
rect 17414 30465 17533 30479
rect 17414 30373 17427 30465
rect 17519 30373 17533 30465
rect 17414 30019 17533 30373
rect 18182 30465 18301 30479
rect 18182 30373 18195 30465
rect 18287 30373 18301 30465
rect 18182 30019 18301 30373
rect 18950 30465 19069 30479
rect 18950 30373 18963 30465
rect 19055 30373 19069 30465
rect 18950 30019 19069 30373
rect 19718 30465 19837 30479
rect 19718 30373 19731 30465
rect 19823 30373 19837 30465
rect 19718 30019 19837 30373
rect 20486 30465 20605 30479
rect 20486 30373 20499 30465
rect 20591 30373 20605 30465
rect 20486 30019 20605 30373
rect 21254 30465 21373 30479
rect 21254 30373 21267 30465
rect 21359 30373 21373 30465
rect 21254 30019 21373 30373
rect 22022 30465 22141 30479
rect 22022 30373 22035 30465
rect 22127 30373 22141 30465
rect 22022 30019 22141 30373
rect 22790 30465 22909 30479
rect 22790 30373 22803 30465
rect 22895 30373 22909 30465
rect 22790 30019 22909 30373
rect 23558 30465 23677 30479
rect 23558 30373 23571 30465
rect 23663 30373 23677 30465
rect 23558 30019 23677 30373
rect 30471 30362 30480 30458
rect 30576 30362 30585 30458
rect 31239 30362 31248 30458
rect 31344 30362 31353 30458
rect 32007 30362 32016 30458
rect 32112 30362 32121 30458
rect 32775 30362 32784 30458
rect 32880 30362 32889 30458
rect 33543 30362 33552 30458
rect 33648 30362 33657 30458
rect 34311 30362 34320 30458
rect 34416 30362 34425 30458
rect 35079 30362 35088 30458
rect 35184 30362 35193 30458
rect 35847 30362 35856 30458
rect 35952 30362 35961 30458
rect 36615 30362 36624 30458
rect 36720 30362 36729 30458
rect 37383 30362 37392 30458
rect 37488 30362 37497 30458
rect 38151 30362 38160 30458
rect 38256 30362 38265 30458
rect 30480 30010 30576 30362
rect 31248 30010 31344 30362
rect 32016 30010 32112 30362
rect 32784 30010 32880 30362
rect 33552 30010 33648 30362
rect 34320 30010 34416 30362
rect 35088 30010 35184 30362
rect 35856 30010 35952 30362
rect 36624 30010 36720 30362
rect 37392 30010 37488 30362
rect 38160 30010 38256 30362
rect 4768 29882 6184 29916
rect 3944 29750 4314 29882
rect 2420 29124 2768 29500
rect 3040 29124 3262 29750
rect 3652 29596 3846 29680
rect 3534 29124 3846 29596
rect 4118 29652 4314 29750
rect 4982 29876 6184 29882
rect 4982 29756 5250 29876
rect 5918 29756 6184 29876
rect 6392 29840 6538 29916
rect 6852 29756 7132 29916
rect 4982 29652 5174 29756
rect 4118 29124 4496 29652
rect 4768 29262 5174 29652
rect 5446 29354 5724 29646
rect 5996 29262 6170 29756
rect 6560 29602 6754 29686
rect 4768 29124 5258 29262
rect 5926 29130 6170 29262
rect 6442 29130 6754 29602
rect 7026 29130 7132 29756
rect 5926 29124 7132 29130
rect 2026 29012 7132 29124
rect 2212 28846 2596 28886
rect 2212 27664 2252 28846
rect 2556 27664 2596 28846
rect 2212 27624 2596 27664
rect 425 21976 605 21985
rect 605 21796 1960 21976
rect 2140 21796 2149 21976
rect 425 21787 605 21796
rect 2240 19606 2736 19646
rect 1964 18808 2144 18817
rect 418 18628 427 18808
rect 607 18628 1964 18808
rect 1964 18619 2144 18628
rect 2240 18424 2280 19606
rect 2696 18424 2736 19606
rect 2240 18384 2736 18424
rect 2212 10366 2596 10406
rect 2212 9184 2252 10366
rect 2556 9184 2596 10366
rect 2212 9144 2596 9184
rect 401 3204 581 3213
rect 581 3024 1660 3204
rect 1840 3024 1849 3204
rect 401 3015 581 3024
rect 2276 2314 4398 2354
rect 2276 2012 2316 2314
rect 4358 2012 4398 2314
rect 2276 1972 4398 2012
<< via3 >>
rect 10515 30373 10607 30465
rect 11283 30373 11375 30465
rect 12051 30373 12143 30465
rect 12819 30373 12911 30465
rect 13587 30373 13679 30465
rect 14355 30373 14447 30465
rect 15123 30373 15215 30465
rect 15891 30373 15983 30465
rect 16659 30373 16751 30465
rect 17427 30373 17519 30465
rect 18195 30373 18287 30465
rect 18963 30373 19055 30465
rect 19731 30373 19823 30465
rect 20499 30373 20591 30465
rect 21267 30373 21359 30465
rect 22035 30373 22127 30465
rect 22803 30373 22895 30465
rect 23571 30373 23663 30465
rect 30480 30362 30576 30458
rect 31248 30362 31344 30458
rect 32016 30362 32112 30458
rect 32784 30362 32880 30458
rect 33552 30362 33648 30458
rect 34320 30362 34416 30458
rect 35088 30362 35184 30458
rect 35856 30362 35952 30458
rect 36624 30362 36720 30458
rect 37392 30362 37488 30458
rect 38160 30362 38256 30458
rect 2252 27664 2556 28846
rect 425 21796 605 21976
rect 427 18628 607 18808
rect 2280 18424 2696 19606
rect 2252 9184 2556 10366
rect 401 3024 581 3204
rect 2316 2012 4358 2314
<< metal4 >>
rect 10515 30465 10607 30474
rect 11283 30465 11375 30474
rect 12051 30465 12143 30474
rect 12819 30465 12911 30474
rect 13587 30465 13679 30474
rect 14355 30465 14447 30474
rect 15123 30465 15215 30474
rect 15891 30465 15983 30474
rect 16659 30465 16751 30474
rect 17427 30465 17519 30474
rect 18195 30465 18287 30474
rect 18963 30465 19055 30474
rect 19731 30465 19823 30474
rect 20499 30465 20591 30474
rect 21267 30465 21359 30474
rect 22035 30465 22127 30474
rect 22803 30465 22895 30474
rect 23571 30465 23663 30474
rect 10508 30375 10515 30462
rect 10607 30375 10613 30462
rect 11276 30375 11283 30462
rect 11375 30375 11381 30462
rect 12044 30375 12051 30462
rect 12143 30375 12149 30462
rect 12812 30375 12819 30462
rect 12911 30375 12917 30462
rect 13580 30375 13587 30462
rect 13679 30375 13685 30462
rect 14348 30375 14355 30462
rect 14447 30375 14453 30462
rect 15116 30375 15123 30462
rect 15215 30375 15221 30462
rect 15884 30375 15891 30462
rect 15983 30375 15989 30462
rect 16652 30375 16659 30462
rect 16751 30375 16757 30462
rect 17420 30375 17427 30462
rect 17519 30375 17525 30462
rect 18188 30375 18195 30462
rect 18287 30375 18293 30462
rect 18956 30375 18963 30462
rect 19055 30375 19061 30462
rect 19724 30375 19731 30462
rect 19823 30375 19829 30462
rect 20492 30375 20499 30462
rect 20591 30375 20597 30462
rect 21260 30375 21267 30462
rect 21359 30375 21365 30462
rect 22028 30375 22035 30462
rect 22127 30375 22133 30462
rect 22796 30375 22803 30462
rect 22895 30375 22901 30462
rect 23564 30375 23571 30462
rect 23663 30375 23669 30462
rect 30480 30458 30576 30467
rect 31248 30458 31344 30467
rect 32016 30458 32112 30467
rect 32784 30458 32880 30467
rect 33552 30458 33648 30467
rect 34320 30458 34416 30467
rect 35088 30458 35184 30467
rect 35856 30458 35952 30467
rect 36624 30458 36720 30467
rect 37392 30458 37488 30467
rect 38160 30458 38256 30467
rect 10515 30364 10607 30373
rect 11283 30364 11375 30373
rect 12051 30364 12143 30373
rect 12819 30364 12911 30373
rect 13587 30364 13679 30373
rect 14355 30364 14447 30373
rect 15123 30364 15215 30373
rect 15891 30364 15983 30373
rect 16659 30364 16751 30373
rect 17427 30364 17519 30373
rect 18195 30364 18287 30373
rect 18963 30364 19055 30373
rect 19731 30364 19823 30373
rect 20499 30364 20591 30373
rect 21267 30364 21359 30373
rect 22035 30364 22127 30373
rect 22803 30364 22895 30373
rect 23571 30364 23663 30373
rect 30471 30362 30480 30458
rect 30576 30362 30585 30458
rect 31239 30362 31248 30458
rect 31344 30362 31353 30458
rect 32007 30362 32016 30458
rect 32112 30362 32121 30458
rect 32775 30362 32784 30458
rect 32880 30362 32889 30458
rect 33543 30362 33552 30458
rect 33648 30362 33657 30458
rect 34311 30362 34320 30458
rect 34416 30362 34425 30458
rect 35079 30362 35088 30458
rect 35184 30362 35193 30458
rect 35847 30362 35856 30458
rect 35952 30362 35961 30458
rect 36615 30362 36624 30458
rect 36720 30362 36729 30458
rect 37383 30362 37392 30458
rect 37488 30362 37497 30458
rect 38151 30362 38160 30458
rect 38256 30362 38265 30458
rect 30480 30353 30576 30362
rect 31248 30353 31344 30362
rect 32016 30353 32112 30362
rect 32784 30353 32880 30362
rect 33552 30353 33648 30362
rect 34320 30353 34416 30362
rect 35088 30353 35184 30362
rect 35856 30353 35952 30362
rect 36624 30353 36720 30362
rect 37392 30353 37488 30362
rect 38160 30353 38256 30362
rect 2026 30244 3192 30322
rect 2026 30118 2268 30244
rect 2936 30118 3192 30244
rect 2026 29124 2148 30118
rect 3040 30040 3192 30118
rect 4340 30118 4950 30256
rect 4340 30040 4496 30118
rect 2420 29730 2768 30014
rect 3040 29910 4496 30040
rect 3040 29750 3276 29910
rect 3484 29834 3630 29910
rect 3944 29882 4496 29910
rect 4768 30040 4950 30118
rect 4768 29916 7132 30040
rect 10528 29917 10841 29926
rect 18296 29917 18609 29926
rect 26055 29917 26368 29926
rect 33840 29917 34153 29926
rect 38530 29917 38924 29930
rect 4768 29882 6184 29916
rect 3944 29750 4314 29882
rect 2420 29124 2768 29500
rect 3040 29124 3262 29750
rect 3652 29596 3846 29680
rect 3534 29124 3846 29596
rect 4118 29652 4314 29750
rect 4982 29876 6184 29882
rect 4982 29756 5250 29876
rect 5918 29756 6184 29876
rect 6392 29840 6538 29916
rect 6852 29756 7132 29916
rect 4982 29652 5174 29756
rect 4118 29124 4496 29652
rect 4768 29262 5174 29652
rect 5446 29354 5724 29646
rect 5996 29262 6170 29756
rect 6560 29602 6754 29686
rect 4768 29124 5258 29262
rect 5926 29130 6170 29262
rect 6442 29130 6754 29602
rect 7026 29130 7132 29756
rect 9984 29612 10528 29917
rect 10841 29612 18296 29917
rect 18609 29612 26055 29917
rect 26368 29612 33840 29917
rect 34153 29884 38924 29917
rect 39102 29884 39542 29893
rect 34153 29612 39102 29884
rect 10528 29603 10841 29612
rect 18296 29603 18609 29612
rect 26055 29603 26368 29612
rect 33840 29603 34153 29612
rect 38530 29474 39102 29612
rect 38844 29444 39102 29474
rect 39102 29435 39542 29444
rect 5926 29124 7132 29130
rect 2026 29012 7132 29124
rect 2212 28846 2596 28886
rect 2212 27664 2252 28846
rect 2556 27664 2596 28846
rect 2212 27624 2596 27664
rect 416 24596 425 24776
rect 605 24596 614 24776
rect 425 21976 605 24596
rect 416 21796 425 21976
rect 605 21796 614 21976
rect 427 21576 607 21585
rect 427 18808 607 21396
rect 427 18619 607 18628
rect 2240 19606 2736 19646
rect 2240 18424 2280 19606
rect 2696 18424 2736 19606
rect 2240 18384 2736 18424
rect 392 18196 401 18376
rect 581 18196 590 18376
rect 401 3204 581 18196
rect 2212 10366 2596 10406
rect 2212 9184 2252 10366
rect 2556 9184 2596 10366
rect 2212 9144 2596 9184
rect 392 3024 401 3204
rect 581 3024 590 3204
rect 2276 2314 4398 2354
rect 2276 2012 2316 2314
rect 4358 2012 4398 2314
rect 2276 1972 4398 2012
rect 3894 1628 38332 1659
rect 3894 1576 6140 1628
rect 3894 1136 4060 1576
rect 4500 1136 6140 1576
rect 3894 1100 6140 1136
rect 6668 1584 38332 1628
rect 6668 1144 11718 1584
rect 12158 1144 19492 1584
rect 19932 1578 38332 1584
rect 19932 1144 27266 1578
rect 6668 1138 27266 1144
rect 27706 1570 38332 1578
rect 27706 1138 35040 1570
rect 6668 1130 35040 1138
rect 35480 1130 38332 1570
rect 6668 1100 38332 1130
rect 3894 1054 38332 1100
<< via4 >>
rect 10517 30375 10604 30462
rect 11285 30375 11372 30462
rect 12053 30375 12140 30462
rect 12821 30375 12908 30462
rect 13589 30375 13676 30462
rect 14357 30375 14444 30462
rect 15125 30375 15212 30462
rect 15893 30375 15980 30462
rect 16661 30375 16748 30462
rect 17429 30375 17516 30462
rect 18197 30375 18284 30462
rect 18965 30375 19052 30462
rect 19733 30375 19820 30462
rect 20501 30375 20588 30462
rect 21269 30375 21356 30462
rect 22037 30375 22124 30462
rect 22805 30375 22892 30462
rect 23573 30375 23660 30462
rect 30480 30362 30576 30458
rect 31248 30362 31344 30458
rect 32016 30362 32112 30458
rect 32784 30362 32880 30458
rect 33552 30362 33648 30458
rect 34320 30362 34416 30458
rect 35088 30362 35184 30458
rect 35856 30362 35952 30458
rect 36624 30362 36720 30458
rect 37392 30362 37488 30458
rect 38160 30362 38256 30458
rect 10528 29612 10841 29917
rect 18296 29612 18609 29917
rect 26055 29612 26368 29917
rect 33840 29612 34153 29917
rect 39102 29444 39542 29884
rect 2252 27664 2556 28846
rect 425 24596 605 24776
rect 427 21396 607 21576
rect 2280 18424 2696 19606
rect 401 18196 581 18376
rect 2252 9184 2556 10366
rect 2316 2012 4358 2314
rect 4060 1136 4500 1576
rect 6140 1100 6668 1628
rect 11718 1144 12158 1584
rect 19492 1144 19932 1584
rect 27266 1138 27706 1578
rect 35040 1130 35480 1570
<< metal5 >>
rect 958 30596 1732 30678
rect 791 30592 1732 30596
rect 5922 30592 5982 30996
rect 6690 30592 6750 30996
rect 7458 30592 7518 30996
rect 8226 30592 8286 30996
rect 8994 30592 9054 30996
rect 9762 30592 9822 30996
rect 791 30532 9822 30592
rect 791 30456 1732 30532
rect 10530 30522 10590 30996
rect 11298 30522 11358 30996
rect 12066 30522 12126 30996
rect 12834 30522 12894 30996
rect 13602 30522 13662 30996
rect 14370 30522 14430 30996
rect 15138 30522 15198 30996
rect 15906 30522 15966 30996
rect 16674 30522 16734 30996
rect 17442 30522 17502 30996
rect 18210 30522 18270 30996
rect 18978 30522 19038 30996
rect 19746 30522 19806 30996
rect 20514 30522 20574 30996
rect 21282 30522 21342 30996
rect 22050 30522 22110 30996
rect 22818 30522 22878 30996
rect 23586 30522 23646 30996
rect 24354 30796 24414 30996
rect 25122 30796 25182 30996
rect 25890 30796 25950 30996
rect 26658 30796 26718 30996
rect 27426 30796 27486 30996
rect 28194 30796 28254 30996
rect 28962 30796 29022 30996
rect 29730 30796 29790 30996
rect 30498 30522 30558 30996
rect 31266 30522 31326 30996
rect 32034 30522 32094 30996
rect 32802 30522 32862 30996
rect 33570 30522 33630 30996
rect 34338 30522 34398 30996
rect 35106 30522 35166 30996
rect 35874 30522 35934 30996
rect 36642 30522 36702 30996
rect 37410 30522 37470 30996
rect 38178 30522 38238 30996
rect 800 30446 1732 30456
rect 10517 30462 10604 30522
rect 800 28886 1240 30446
rect 10517 30366 10604 30375
rect 11285 30462 11372 30522
rect 11285 30366 11372 30375
rect 12053 30462 12140 30522
rect 12053 30366 12140 30375
rect 12821 30462 12908 30522
rect 12821 30366 12908 30375
rect 13589 30462 13676 30522
rect 13589 30366 13676 30375
rect 14357 30462 14444 30522
rect 14357 30366 14444 30375
rect 15125 30462 15212 30522
rect 15125 30366 15212 30375
rect 15893 30462 15980 30522
rect 15893 30366 15980 30375
rect 16661 30462 16748 30522
rect 16661 30366 16748 30375
rect 17429 30462 17516 30522
rect 17429 30366 17516 30375
rect 18197 30462 18284 30522
rect 18197 30366 18284 30375
rect 18965 30462 19052 30522
rect 18965 30366 19052 30375
rect 19733 30462 19820 30522
rect 19733 30366 19820 30375
rect 20501 30462 20588 30522
rect 20501 30366 20588 30375
rect 21269 30462 21356 30522
rect 21269 30366 21356 30375
rect 22037 30462 22124 30522
rect 22037 30366 22124 30375
rect 22805 30462 22892 30522
rect 22805 30366 22892 30375
rect 23573 30462 23660 30522
rect 23573 30366 23660 30375
rect 30480 30458 30576 30522
rect 30480 30353 30576 30362
rect 31248 30458 31344 30522
rect 31248 30353 31344 30362
rect 32016 30458 32112 30522
rect 32016 30353 32112 30362
rect 32784 30458 32880 30522
rect 32784 30353 32880 30362
rect 33552 30458 33648 30522
rect 33552 30353 33648 30362
rect 34320 30458 34416 30522
rect 34320 30353 34416 30362
rect 35088 30458 35184 30522
rect 35088 30353 35184 30362
rect 35856 30458 35952 30522
rect 35856 30353 35952 30362
rect 36624 30458 36720 30522
rect 36624 30353 36720 30362
rect 37392 30458 37488 30522
rect 37392 30353 37488 30362
rect 38160 30458 38256 30522
rect 38160 30353 38256 30362
rect 2268 30118 2936 30244
rect 2148 30014 3040 30118
rect 2148 29730 2420 30014
rect 2768 29730 3040 30014
rect 3276 29834 3484 29910
rect 3630 29834 3944 29910
rect 4496 29882 4768 30118
rect 7482 30000 38626 30276
rect 3276 29750 3944 29834
rect 2148 29500 3040 29730
rect 2148 29124 2420 29500
rect 2768 29124 3040 29500
rect 3262 29680 4118 29750
rect 3262 29596 3652 29680
rect 3262 29124 3534 29596
rect 3846 29124 4118 29680
rect 4314 29652 4982 29882
rect 5250 29756 5918 29876
rect 6184 29840 6392 29916
rect 6538 29840 6852 29916
rect 6184 29756 6852 29840
rect 4496 29124 4768 29652
rect 5174 29646 5996 29756
rect 5174 29354 5446 29646
rect 5724 29354 5996 29646
rect 5174 29262 5996 29354
rect 6170 29686 7026 29756
rect 6170 29602 6560 29686
rect 5258 29124 5926 29262
rect 6170 29130 6442 29602
rect 6754 29130 7026 29686
rect 800 28846 2596 28886
rect 800 27664 2252 28846
rect 2556 28722 2596 28846
rect 7482 28722 7758 30000
rect 10519 29612 10528 29917
rect 10841 29612 10850 29917
rect 10532 28760 10837 29612
rect 11792 28740 12068 30000
rect 18287 29612 18296 29917
rect 18609 29612 18618 29917
rect 18300 28812 18605 29612
rect 19562 28740 19838 30000
rect 26046 29612 26055 29917
rect 26368 29612 26377 29917
rect 26059 28838 26364 29612
rect 27348 28844 27624 30000
rect 33831 29612 33840 29917
rect 34153 29612 34162 29917
rect 33844 28812 34149 29612
rect 35100 28810 35376 30000
rect 39800 29884 40240 30596
rect 39093 29444 39102 29884
rect 39542 29444 40240 29884
rect 2556 28446 7758 28722
rect 2556 27664 2596 28446
rect 800 27624 2596 27664
rect 425 24776 605 24785
rect 0 24596 425 24776
rect 425 24587 605 24596
rect 0 21396 427 21576
rect 607 21396 616 21576
rect 800 19646 1240 27624
rect 6240 27602 6516 28446
rect 800 19606 2736 19646
rect 800 18424 2280 19606
rect 2696 18424 2736 19606
rect 401 18376 581 18385
rect 0 18196 401 18376
rect 401 18187 581 18196
rect 800 18384 2736 18424
rect 0 14996 200 15176
rect 800 10406 1240 18384
rect 800 10366 2596 10406
rect 800 9184 2252 10366
rect 2556 9184 2596 10366
rect 800 9144 2596 9184
rect 800 1576 1240 9144
rect 2188 2354 3514 2406
rect 2188 2314 4398 2354
rect 2188 2012 2316 2314
rect 4358 2012 4398 2314
rect 2188 1972 4398 2012
rect 2188 1576 3514 1972
rect 800 1136 4060 1576
rect 4500 1136 4509 1576
rect 800 0 1240 1136
rect 4890 792 5406 3116
rect 6102 1628 6707 3082
rect 6102 1100 6140 1628
rect 6668 1100 6707 1628
rect 6102 1040 6707 1100
rect 10448 796 10968 2534
rect 11718 1584 12158 2488
rect 11718 1135 12158 1144
rect 18214 796 18734 2540
rect 19492 1584 19932 2372
rect 19492 1135 19932 1144
rect 25998 796 26518 2556
rect 27266 1578 27706 2372
rect 27266 1129 27706 1138
rect 33750 796 34270 2482
rect 35040 1570 35480 2372
rect 35040 1121 35480 1130
rect 39800 796 40240 29444
rect 7828 792 40240 796
rect 4890 276 40240 792
rect 39800 0 40240 276
use r2r_dac  blue_dac
timestamp 1746839692
transform 0 1 2318 -1 0 10142
box -142 -18 7922 2062
use controller  controller_0
timestamp 1747056179
transform 1 0 7402 0 1 1156
box 0 700 31440 29000
use r2r_dac  green_dac
timestamp 1746839692
transform 0 1 2318 -1 0 19382
box -142 -18 7922 2062
use r2r_dac  red_dac
timestamp 1746839692
transform 0 1 2318 -1 0 28622
box -142 -18 7922 2062
use rgb_buffers  rgb_buffers_0
timestamp 1747056179
transform 1 0 4652 0 1 2416
box 0 -56 2600 25760
<< labels >>
flabel metal5 s 37410 30796 37470 30996 4 FreeSans 320 0 0 0 clk
port 2 nsew
flabel metal5 s 38178 30796 38238 30996 4 FreeSans 320 0 0 0 ena
port 3 nsew
flabel metal5 s 36642 30796 36702 30996 4 FreeSans 320 0 0 0 rst_n
port 4 nsew
flabel metal5 s 35874 30796 35934 30996 4 FreeSans 320 0 0 0 ui_in[0]
port 5 nsew
flabel metal5 s 35106 30796 35166 30996 4 FreeSans 320 0 0 0 ui_in[1]
port 6 nsew
flabel metal5 s 34338 30796 34398 30996 4 FreeSans 320 0 0 0 ui_in[2]
port 7 nsew
flabel metal5 s 33570 30796 33630 30996 4 FreeSans 320 0 0 0 ui_in[3]
port 8 nsew
flabel metal5 s 32802 30796 32862 30996 4 FreeSans 320 0 0 0 ui_in[4]
port 9 nsew
flabel metal5 s 32034 30796 32094 30996 4 FreeSans 320 0 0 0 ui_in[5]
port 10 nsew
flabel metal5 s 31266 30796 31326 30996 4 FreeSans 320 0 0 0 ui_in[6]
port 11 nsew
flabel metal5 s 30498 30796 30558 30996 4 FreeSans 320 0 0 0 ui_in[7]
port 12 nsew
flabel metal5 s 29730 30796 29790 30996 4 FreeSans 320 0 0 0 uio_in[0]
port 13 nsew
flabel metal5 s 28962 30796 29022 30996 4 FreeSans 320 0 0 0 uio_in[1]
port 14 nsew
flabel metal5 s 28194 30796 28254 30996 4 FreeSans 320 0 0 0 uio_in[2]
port 15 nsew
flabel metal5 s 27426 30796 27486 30996 4 FreeSans 320 0 0 0 uio_in[3]
port 16 nsew
flabel metal5 s 26658 30796 26718 30996 4 FreeSans 320 0 0 0 uio_in[4]
port 17 nsew
flabel metal5 s 25890 30796 25950 30996 4 FreeSans 320 0 0 0 uio_in[5]
port 18 nsew
flabel metal5 s 25122 30796 25182 30996 4 FreeSans 320 0 0 0 uio_in[6]
port 19 nsew
flabel metal5 s 24354 30796 24414 30996 4 FreeSans 320 0 0 0 uio_in[7]
port 20 nsew
flabel metal5 s 11298 30796 11358 30996 4 FreeSans 320 0 0 0 uio_oe[0]
port 21 nsew
flabel metal5 s 10530 30796 10590 30996 4 FreeSans 320 0 0 0 uio_oe[1]
port 22 nsew
flabel metal5 s 9762 30796 9822 30996 4 FreeSans 320 0 0 0 uio_oe[2]
port 23 nsew
flabel metal5 s 8994 30796 9054 30996 4 FreeSans 320 0 0 0 uio_oe[3]
port 24 nsew
flabel metal5 s 8226 30796 8286 30996 4 FreeSans 320 0 0 0 uio_oe[4]
port 25 nsew
flabel metal5 s 7458 30796 7518 30996 4 FreeSans 320 0 0 0 uio_oe[5]
port 26 nsew
flabel metal5 s 6690 30796 6750 30996 4 FreeSans 320 0 0 0 uio_oe[6]
port 27 nsew
flabel metal5 s 5922 30796 5982 30996 4 FreeSans 320 0 0 0 uio_oe[7]
port 28 nsew
flabel metal5 s 17442 30796 17502 30996 4 FreeSans 320 0 0 0 uio_out[0]
port 29 nsew
flabel metal5 s 16674 30796 16734 30996 4 FreeSans 320 0 0 0 uio_out[1]
port 30 nsew
flabel metal5 s 15906 30796 15966 30996 4 FreeSans 320 0 0 0 uio_out[2]
port 31 nsew
flabel metal5 s 15138 30796 15198 30996 4 FreeSans 320 0 0 0 uio_out[3]
port 32 nsew
flabel metal5 s 14370 30796 14430 30996 4 FreeSans 320 0 0 0 uio_out[4]
port 33 nsew
flabel metal5 s 13602 30796 13662 30996 4 FreeSans 320 0 0 0 uio_out[5]
port 34 nsew
flabel metal5 s 12834 30796 12894 30996 4 FreeSans 320 0 0 0 uio_out[6]
port 35 nsew
flabel metal5 s 12066 30796 12126 30996 4 FreeSans 320 0 0 0 uio_out[7]
port 36 nsew
flabel metal5 s 23586 30796 23646 30996 4 FreeSans 320 0 0 0 uo_out[0]
port 37 nsew
flabel metal5 s 22818 30796 22878 30996 4 FreeSans 320 0 0 0 uo_out[1]
port 38 nsew
flabel metal5 s 22050 30796 22110 30996 4 FreeSans 320 0 0 0 uo_out[2]
port 39 nsew
flabel metal5 s 21282 30796 21342 30996 4 FreeSans 320 0 0 0 uo_out[3]
port 40 nsew
flabel metal5 s 20514 30796 20574 30996 4 FreeSans 320 0 0 0 uo_out[4]
port 41 nsew
flabel metal5 s 19746 30796 19806 30996 4 FreeSans 320 0 0 0 uo_out[5]
port 42 nsew
flabel metal5 s 18978 30796 19038 30996 4 FreeSans 320 0 0 0 uo_out[6]
port 43 nsew
flabel metal5 s 18210 30796 18270 30996 4 FreeSans 320 0 0 0 uo_out[7]
port 44 nsew
flabel metal5 s 0 24596 200 24776 0 FreeSans 320 0 0 0 ua[0]
port 45 nsew
flabel metal5 s 0 21396 200 21576 0 FreeSans 320 0 0 0 ua[1]
port 46 nsew
flabel metal5 s 0 18196 200 18376 0 FreeSans 320 0 0 0 ua[2]
port 47 nsew
flabel metal5 s 0 14996 200 15176 0 FreeSans 320 0 0 0 ua[3]
port 48 nsew
flabel metal5 s 800 0 1240 30596 0 FreeSans 320 0 0 0 VGND
port 49 nsew
flabel metal5 s 39800 0 40240 30596 0 FreeSans 320 0 0 0 VPWR
port 50 nsew
<< properties >>
string FIXED_BBOX 0 0 40416 30996
<< end >>
