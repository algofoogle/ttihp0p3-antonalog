magic
tech ihp-sg13g2
timestamp 1747537721
<< nwell >>
rect -24 175 312 417
<< pwell >>
rect 8 28 273 148
rect -13 -28 301 28
<< nmos >>
rect 60 61 73 135
rect 110 61 123 135
rect 162 61 175 135
rect 213 61 226 135
<< pmos >>
rect 60 213 73 325
rect 111 213 124 325
rect 162 213 175 325
rect 213 213 226 325
<< ndiff >>
rect 21 128 60 135
rect 21 112 28 128
rect 44 112 60 128
rect 21 84 60 112
rect 21 68 28 84
rect 44 68 60 84
rect 21 61 60 68
rect 73 61 110 135
rect 123 61 162 135
rect 175 61 213 135
rect 226 128 260 135
rect 226 112 237 128
rect 253 112 260 128
rect 226 84 260 112
rect 226 68 237 84
rect 253 68 260 84
rect 226 61 260 68
<< pdiff >>
rect 26 317 60 325
rect 26 301 33 317
rect 49 301 60 317
rect 26 278 60 301
rect 26 262 33 278
rect 49 262 60 278
rect 26 236 60 262
rect 26 220 33 236
rect 49 220 60 236
rect 26 213 60 220
rect 73 317 111 325
rect 73 301 84 317
rect 100 301 111 317
rect 73 278 111 301
rect 73 262 84 278
rect 100 262 111 278
rect 73 236 111 262
rect 73 220 84 236
rect 100 220 111 236
rect 73 213 111 220
rect 124 317 162 325
rect 124 301 135 317
rect 151 301 162 317
rect 124 278 162 301
rect 124 262 135 278
rect 151 262 162 278
rect 124 213 162 262
rect 175 317 213 325
rect 175 301 186 317
rect 202 301 213 317
rect 175 278 213 301
rect 175 262 186 278
rect 202 262 213 278
rect 175 236 213 262
rect 175 220 186 236
rect 202 220 213 236
rect 175 213 213 220
rect 226 317 260 325
rect 226 301 237 317
rect 253 301 260 317
rect 226 278 260 301
rect 226 262 237 278
rect 253 262 260 278
rect 226 213 260 262
<< ndiffc >>
rect 28 112 44 128
rect 28 68 44 84
rect 237 112 253 128
rect 237 68 253 84
<< pdiffc >>
rect 33 301 49 317
rect 33 262 49 278
rect 33 220 49 236
rect 84 301 100 317
rect 84 262 100 278
rect 84 220 100 236
rect 135 301 151 317
rect 135 262 151 278
rect 186 301 202 317
rect 186 262 202 278
rect 186 220 202 236
rect 237 301 253 317
rect 237 262 253 278
<< psubdiff >>
rect 0 8 288 15
rect 0 -8 16 8
rect 32 -8 64 8
rect 80 -8 112 8
rect 128 -8 160 8
rect 176 -8 208 8
rect 224 -8 256 8
rect 272 -8 288 8
rect 0 -15 288 -8
<< nsubdiff >>
rect 0 386 288 393
rect 0 370 16 386
rect 32 370 64 386
rect 80 370 112 386
rect 128 370 160 386
rect 176 370 208 386
rect 224 370 256 386
rect 272 370 288 386
rect 0 363 288 370
<< psubdiffcont >>
rect 16 -8 32 8
rect 64 -8 80 8
rect 112 -8 128 8
rect 160 -8 176 8
rect 208 -8 224 8
rect 256 -8 272 8
<< nsubdiffcont >>
rect 16 370 32 386
rect 64 370 80 386
rect 112 370 128 386
rect 160 370 176 386
rect 208 370 224 386
rect 256 370 272 386
<< poly >>
rect 60 325 73 343
rect 111 325 124 343
rect 162 325 175 343
rect 213 325 226 343
rect 60 187 73 213
rect 111 190 124 213
rect 36 180 73 187
rect 36 164 43 180
rect 59 164 73 180
rect 36 157 73 164
rect 102 181 132 190
rect 162 185 175 213
rect 213 196 226 213
rect 204 189 234 196
rect 102 165 109 181
rect 125 165 132 181
rect 102 158 132 165
rect 153 178 183 185
rect 153 162 160 178
rect 176 162 183 178
rect 204 173 211 189
rect 227 173 234 189
rect 204 166 234 173
rect 60 135 73 157
rect 110 135 123 158
rect 153 155 183 162
rect 162 135 175 155
rect 213 135 226 166
rect 60 43 73 61
rect 110 43 123 61
rect 162 43 175 61
rect 213 43 226 61
<< polycont >>
rect 43 164 59 180
rect 109 165 125 181
rect 160 162 176 178
rect 211 173 227 189
<< metal1 >>
rect 0 386 288 400
rect 0 370 16 386
rect 32 370 64 386
rect 80 370 112 386
rect 128 370 160 386
rect 176 370 208 386
rect 224 370 256 386
rect 272 370 288 386
rect 0 356 288 370
rect 28 317 54 356
rect 28 301 33 317
rect 49 301 54 317
rect 28 278 54 301
rect 28 262 33 278
rect 49 262 54 278
rect 28 236 54 262
rect 28 220 33 236
rect 49 220 54 236
rect 28 218 54 220
rect 79 317 105 322
rect 79 301 84 317
rect 100 301 105 317
rect 79 278 105 301
rect 79 262 84 278
rect 100 262 105 278
rect 79 239 105 262
rect 130 317 156 356
rect 130 301 135 317
rect 151 301 156 317
rect 130 278 156 301
rect 130 262 135 278
rect 151 262 156 278
rect 130 257 156 262
rect 181 317 207 322
rect 181 301 186 317
rect 202 301 207 317
rect 181 278 207 301
rect 181 262 186 278
rect 202 262 207 278
rect 181 239 207 262
rect 232 317 258 356
rect 232 301 237 317
rect 253 301 258 317
rect 232 278 258 301
rect 232 262 237 278
rect 253 262 258 278
rect 232 257 258 262
rect 79 236 270 239
rect 79 220 84 236
rect 100 220 186 236
rect 202 220 270 236
rect 79 218 270 220
rect 36 180 69 200
rect 36 164 43 180
rect 59 164 69 180
rect 36 155 69 164
rect 95 181 132 200
rect 95 165 109 181
rect 125 165 132 181
rect 95 155 132 165
rect 150 178 183 200
rect 150 162 160 178
rect 176 162 183 178
rect 150 155 183 162
rect 201 189 228 200
rect 201 173 211 189
rect 227 173 228 189
rect 201 155 228 173
rect 246 133 270 218
rect 22 128 49 133
rect 22 112 28 128
rect 44 112 49 128
rect 22 84 49 112
rect 22 68 28 84
rect 44 68 49 84
rect 22 22 49 68
rect 232 128 270 133
rect 232 112 237 128
rect 253 112 270 128
rect 232 84 270 112
rect 232 68 237 84
rect 253 68 270 84
rect 232 63 270 68
rect 0 8 288 22
rect 0 -8 16 8
rect 32 -8 64 8
rect 80 -8 112 8
rect 128 -8 160 8
rect 176 -8 208 8
rect 224 -8 256 8
rect 272 -8 288 8
rect 0 -22 288 -8
<< labels >>
flabel metal1 s 0 356 288 400 0 FreeSans 200 0 0 0 VDD
port 2 nsew
flabel metal1 s 246 63 270 239 0 FreeSans 200 0 0 0 Y
port 3 nsew
flabel metal1 s 150 155 183 200 0 FreeSans 200 0 0 0 B
port 4 nsew
flabel metal1 s 95 155 132 200 0 FreeSans 200 0 0 0 C
port 5 nsew
flabel metal1 s 0 -22 288 22 0 FreeSans 200 0 0 0 VSS
port 6 nsew
flabel metal1 s 201 155 228 200 0 FreeSans 200 0 0 0 A
port 7 nsew
flabel metal1 s 36 155 69 200 0 FreeSans 250 0 0 0 D
port 8 nsew
<< properties >>
string FIXED_BBOX 0 0 288 378
string GDS_END 191660
string GDS_FILE ../gds/controller.gds
string GDS_START 186986
<< end >>
