magic
tech ihp-sg13g2
magscale 1 2
timestamp 1747056038
<< nwell >>
rect -54 350 528 834
<< pwell >>
rect 20 56 464 292
rect -26 -56 506 56
<< nmos >>
rect 114 156 140 266
rect 242 118 268 266
rect 344 118 370 266
<< pmos >>
rect 114 412 140 580
rect 242 412 268 636
rect 310 412 336 636
<< ndiff >>
rect 46 252 114 266
rect 46 220 60 252
rect 92 220 114 252
rect 46 156 114 220
rect 140 164 242 266
rect 140 156 188 164
rect 174 132 188 156
rect 220 132 242 164
rect 174 118 242 132
rect 268 252 344 266
rect 268 220 290 252
rect 322 220 344 252
rect 268 164 344 220
rect 268 132 290 164
rect 322 132 344 164
rect 268 118 344 132
rect 370 252 438 266
rect 370 220 392 252
rect 424 220 438 252
rect 370 164 438 220
rect 370 132 392 164
rect 424 132 438 164
rect 370 118 438 132
<< pdiff >>
rect 174 622 242 636
rect 174 590 188 622
rect 220 590 242 622
rect 174 580 242 590
rect 46 566 114 580
rect 46 534 60 566
rect 92 534 114 566
rect 46 458 114 534
rect 46 426 60 458
rect 92 426 114 458
rect 46 412 114 426
rect 140 553 242 580
rect 140 521 188 553
rect 220 521 242 553
rect 140 412 242 521
rect 268 412 310 636
rect 336 622 404 636
rect 336 590 358 622
rect 390 590 404 622
rect 336 553 404 590
rect 336 521 358 553
rect 390 521 404 553
rect 336 483 404 521
rect 336 451 358 483
rect 390 451 404 483
rect 336 412 404 451
<< ndiffc >>
rect 60 220 92 252
rect 188 132 220 164
rect 290 220 322 252
rect 290 132 322 164
rect 392 220 424 252
rect 392 132 424 164
<< pdiffc >>
rect 188 590 220 622
rect 60 534 92 566
rect 60 426 92 458
rect 188 521 220 553
rect 358 590 390 622
rect 358 521 390 553
rect 358 451 390 483
<< psubdiff >>
rect 0 16 480 30
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 480 16
rect 0 -30 480 -16
<< nsubdiff >>
rect 0 772 480 786
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 480 772
rect 0 726 480 740
<< psubdiffcont >>
rect 32 -16 64 16
rect 128 -16 160 16
rect 224 -16 256 16
rect 320 -16 352 16
rect 416 -16 448 16
<< nsubdiffcont >>
rect 32 740 64 772
rect 128 740 160 772
rect 224 740 256 772
rect 320 740 352 772
rect 416 740 448 772
<< poly >>
rect 242 636 268 672
rect 310 636 336 672
rect 114 580 140 616
rect 114 356 140 412
rect 54 342 140 356
rect 242 354 268 412
rect 54 310 68 342
rect 100 310 140 342
rect 54 296 140 310
rect 114 266 140 296
rect 176 340 268 354
rect 176 308 190 340
rect 222 308 268 340
rect 176 294 268 308
rect 310 397 336 412
rect 310 370 346 397
rect 310 353 406 370
rect 310 321 357 353
rect 389 321 406 353
rect 310 304 406 321
rect 242 266 268 294
rect 344 266 370 304
rect 114 120 140 156
rect 242 82 268 118
rect 344 82 370 118
<< polycont >>
rect 68 310 100 342
rect 190 308 222 340
rect 357 321 389 353
<< metal1 >>
rect 0 772 480 800
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 480 772
rect 0 712 480 740
rect 178 622 230 712
rect 178 590 188 622
rect 220 590 230 622
rect 50 566 102 576
rect 50 534 60 566
rect 92 534 102 566
rect 50 458 102 534
rect 178 553 230 590
rect 178 521 188 553
rect 220 521 230 553
rect 178 511 230 521
rect 346 622 406 625
rect 346 590 358 622
rect 390 590 406 622
rect 346 553 406 590
rect 346 521 358 553
rect 390 521 406 553
rect 346 487 406 521
rect 50 426 60 458
rect 92 452 102 458
rect 272 483 406 487
rect 92 426 230 452
rect 50 416 230 426
rect 54 342 114 374
rect 54 310 68 342
rect 100 310 114 342
rect 54 300 114 310
rect 178 340 230 416
rect 178 308 190 340
rect 222 308 230 340
rect 178 262 230 308
rect 50 252 230 262
rect 50 220 60 252
rect 92 220 230 252
rect 50 210 230 220
rect 272 451 358 483
rect 390 451 406 483
rect 272 447 406 451
rect 272 270 306 447
rect 342 353 406 400
rect 342 321 357 353
rect 389 321 406 353
rect 342 304 406 321
rect 272 252 325 270
rect 272 220 290 252
rect 322 220 325 252
rect 178 164 230 174
rect 178 132 188 164
rect 220 132 230 164
rect 178 44 230 132
rect 272 164 325 220
rect 272 132 290 164
rect 322 132 325 164
rect 272 121 325 132
rect 382 252 434 257
rect 382 220 392 252
rect 424 220 434 252
rect 382 164 434 220
rect 382 132 392 164
rect 424 132 434 164
rect 382 44 434 132
rect 0 16 480 44
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 480 16
rect 0 -44 480 -16
<< labels >>
flabel metal1 s 342 304 406 400 0 FreeSans 400 0 0 0 A
port 2 nsew
flabel metal1 s 54 300 114 374 0 FreeSans 400 0 0 0 B_N
port 3 nsew
flabel metal1 s 0 712 480 800 0 FreeSans 400 0 0 0 VDD
port 4 nsew
flabel metal1 s 346 447 406 625 0 FreeSans 400 0 0 0 Y
port 5 nsew
flabel metal1 s 0 -44 480 44 0 FreeSans 400 0 0 0 VSS
port 6 nsew
<< properties >>
string FIXED_BBOX 0 0 480 756
string GDS_END 112448
string GDS_FILE ../gds/controller.gds
string GDS_START 108680
<< end >>
