magic
tech ihp-sg13g2
magscale 1 2
timestamp 1747056038
<< nwell >>
rect -48 350 816 834
<< pwell >>
rect 17 56 731 292
rect -26 -56 794 56
<< nmos >>
rect 111 118 137 266
rect 213 118 239 266
rect 315 118 341 266
rect 417 118 443 266
rect 607 118 633 266
<< pmos >>
rect 111 412 137 636
rect 213 412 239 636
rect 315 412 341 636
rect 417 412 443 636
rect 519 412 545 580
rect 621 412 647 580
<< ndiff >>
rect 43 196 111 266
rect 43 164 57 196
rect 89 164 111 196
rect 43 118 111 164
rect 137 252 213 266
rect 137 220 159 252
rect 191 220 213 252
rect 137 164 213 220
rect 137 132 159 164
rect 191 132 213 164
rect 137 118 213 132
rect 239 174 315 266
rect 239 142 261 174
rect 293 142 315 174
rect 239 118 315 142
rect 341 252 417 266
rect 341 220 363 252
rect 395 220 417 252
rect 341 164 417 220
rect 341 132 363 164
rect 395 132 417 164
rect 341 118 417 132
rect 443 164 607 266
rect 443 132 485 164
rect 517 132 553 164
rect 585 132 607 164
rect 443 118 607 132
rect 633 252 705 266
rect 633 220 659 252
rect 691 220 705 252
rect 633 164 705 220
rect 633 132 659 164
rect 691 132 705 164
rect 633 118 705 132
<< pdiff >>
rect 43 622 111 636
rect 43 590 57 622
rect 89 590 111 622
rect 43 540 111 590
rect 43 508 57 540
rect 89 508 111 540
rect 43 458 111 508
rect 43 426 57 458
rect 89 426 111 458
rect 43 412 111 426
rect 137 622 213 636
rect 137 590 159 622
rect 191 590 213 622
rect 137 540 213 590
rect 137 508 159 540
rect 191 508 213 540
rect 137 458 213 508
rect 137 426 159 458
rect 191 426 213 458
rect 137 412 213 426
rect 239 622 315 636
rect 239 590 261 622
rect 293 590 315 622
rect 239 505 315 590
rect 239 473 261 505
rect 293 473 315 505
rect 239 412 315 473
rect 341 622 417 636
rect 341 590 363 622
rect 395 590 417 622
rect 341 540 417 590
rect 341 508 363 540
rect 395 508 417 540
rect 341 458 417 508
rect 341 426 363 458
rect 395 426 417 458
rect 341 412 417 426
rect 443 580 505 636
rect 443 565 519 580
rect 443 533 465 565
rect 497 533 519 565
rect 443 494 519 533
rect 443 462 465 494
rect 497 462 519 494
rect 443 412 519 462
rect 545 551 621 580
rect 545 519 567 551
rect 599 519 621 551
rect 545 483 621 519
rect 545 451 567 483
rect 599 451 621 483
rect 545 412 621 451
rect 647 566 715 580
rect 647 534 669 566
rect 701 534 715 566
rect 647 412 715 534
<< ndiffc >>
rect 57 164 89 196
rect 159 220 191 252
rect 159 132 191 164
rect 261 142 293 174
rect 363 220 395 252
rect 363 132 395 164
rect 485 132 517 164
rect 553 132 585 164
rect 659 220 691 252
rect 659 132 691 164
<< pdiffc >>
rect 57 590 89 622
rect 57 508 89 540
rect 57 426 89 458
rect 159 590 191 622
rect 159 508 191 540
rect 159 426 191 458
rect 261 590 293 622
rect 261 473 293 505
rect 363 590 395 622
rect 363 508 395 540
rect 363 426 395 458
rect 465 533 497 565
rect 465 462 497 494
rect 567 519 599 551
rect 567 451 599 483
rect 669 534 701 566
<< psubdiff >>
rect 0 16 768 30
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 608 16
rect 640 -16 704 16
rect 736 -16 768 16
rect 0 -30 768 -16
<< nsubdiff >>
rect 0 772 768 786
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 608 772
rect 640 740 704 772
rect 736 740 768 772
rect 0 726 768 740
<< psubdiffcont >>
rect 32 -16 64 16
rect 128 -16 160 16
rect 224 -16 256 16
rect 320 -16 352 16
rect 416 -16 448 16
rect 512 -16 544 16
rect 608 -16 640 16
rect 704 -16 736 16
<< nsubdiffcont >>
rect 32 740 64 772
rect 128 740 160 772
rect 224 740 256 772
rect 320 740 352 772
rect 416 740 448 772
rect 512 740 544 772
rect 608 740 640 772
rect 704 740 736 772
<< poly >>
rect 111 636 137 672
rect 213 636 239 672
rect 315 636 341 672
rect 417 636 443 672
rect 519 580 545 616
rect 621 580 647 616
rect 111 334 137 412
rect 213 370 239 412
rect 315 370 341 412
rect 417 370 443 412
rect 519 380 545 412
rect 621 380 647 412
rect 213 353 464 370
rect 213 334 278 353
rect 111 321 278 334
rect 310 321 346 353
rect 378 321 414 353
rect 446 321 464 353
rect 519 363 647 380
rect 519 350 581 363
rect 111 304 464 321
rect 564 331 581 350
rect 613 331 647 363
rect 564 314 647 331
rect 111 266 137 304
rect 213 266 239 304
rect 315 266 341 304
rect 417 266 443 304
rect 607 266 633 314
rect 111 82 137 118
rect 213 82 239 118
rect 315 82 341 118
rect 417 82 443 118
rect 607 82 633 118
<< polycont >>
rect 278 321 310 353
rect 346 321 378 353
rect 414 321 446 353
rect 581 331 613 363
<< metal1 >>
rect 0 772 768 800
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 608 772
rect 640 740 704 772
rect 736 740 768 772
rect 0 712 768 740
rect 47 622 99 712
rect 47 590 57 622
rect 89 590 99 622
rect 47 540 99 590
rect 47 508 57 540
rect 89 508 99 540
rect 47 458 99 508
rect 47 426 57 458
rect 89 426 99 458
rect 47 423 99 426
rect 149 622 201 626
rect 149 590 159 622
rect 191 590 201 622
rect 149 540 201 590
rect 149 508 159 540
rect 191 508 201 540
rect 149 458 201 508
rect 251 622 303 712
rect 251 590 261 622
rect 293 590 303 622
rect 251 505 303 590
rect 251 473 261 505
rect 293 473 303 505
rect 251 469 303 473
rect 353 622 405 626
rect 353 590 363 622
rect 395 590 405 622
rect 353 540 405 590
rect 353 508 363 540
rect 395 508 405 540
rect 149 426 159 458
rect 191 433 201 458
rect 353 458 405 508
rect 353 433 363 458
rect 191 426 363 433
rect 395 426 405 458
rect 455 565 507 712
rect 455 533 465 565
rect 497 533 507 565
rect 659 566 711 712
rect 455 494 507 533
rect 455 462 465 494
rect 497 462 507 494
rect 455 457 507 462
rect 557 551 609 554
rect 557 519 567 551
rect 599 519 609 551
rect 659 534 669 566
rect 701 534 711 566
rect 659 528 711 534
rect 557 484 609 519
rect 557 483 718 484
rect 557 451 567 483
rect 599 451 718 483
rect 557 441 718 451
rect 149 399 405 426
rect 149 257 201 399
rect 554 363 630 400
rect 261 353 506 363
rect 261 321 278 353
rect 310 321 346 353
rect 378 321 414 353
rect 446 321 506 353
rect 261 311 506 321
rect 554 331 581 363
rect 613 331 630 363
rect 554 314 630 331
rect 472 270 506 311
rect 680 270 718 441
rect 149 252 405 257
rect 149 220 159 252
rect 191 220 363 252
rect 395 220 405 252
rect 472 252 718 270
rect 472 236 659 252
rect 149 213 405 220
rect 47 196 99 200
rect 47 164 57 196
rect 89 164 99 196
rect 47 44 99 164
rect 149 164 201 213
rect 149 132 159 164
rect 191 132 201 164
rect 149 126 201 132
rect 251 174 303 176
rect 251 142 261 174
rect 293 142 303 174
rect 251 44 303 142
rect 353 164 405 213
rect 649 220 659 236
rect 691 220 718 252
rect 353 132 363 164
rect 395 132 405 164
rect 353 129 405 132
rect 482 164 588 174
rect 482 132 485 164
rect 517 132 553 164
rect 585 132 588 164
rect 482 119 588 132
rect 649 164 718 220
rect 649 132 659 164
rect 691 132 718 164
rect 649 128 718 132
rect 509 44 561 119
rect 0 16 768 44
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 608 16
rect 640 -16 704 16
rect 736 -16 768 16
rect 0 -44 768 -16
<< labels >>
flabel metal1 s 149 126 201 626 0 FreeSans 400 0 0 0 X
port 2 nsew
flabel metal1 s 0 -44 768 44 0 FreeSans 400 0 0 0 VSS
port 3 nsew
flabel metal1 s 554 314 630 400 0 FreeSans 400 0 0 0 A
port 4 nsew
flabel metal1 s 0 712 768 800 0 FreeSans 400 0 0 0 VDD
port 5 nsew
<< properties >>
string FIXED_BBOX 0 0 768 756
string GDS_END 61080
string GDS_FILE ../gds/controller.gds
string GDS_START 54848
<< end >>
