* NGSPICE file created from rgb_buffers_parax.ext - technology: ihp-sg13g2

.subckt rgb_buffers_parax VGND VPWR b[0] b[1] b[2] b[3] b[4] b[5] b[6] b[7] db[0]
+ db[1] db[2] db[3] db[4] db[5] db[6] db[7] dg[0] dg[1] dg[2] dg[3] dg[4] dg[5] dg[6]
+ dg[7] dr[0] dr[1] dr[2] dr[3] dr[4] dr[5] dr[6] dr[7] g[0] g[1] g[2] g[3] g[4] g[5]
+ g[6] g[7] r[0] r[1] r[2] r[3] r[4] r[5] r[6] r[7]
X0 b[5].t4 a_490_3864# VGND.t446 VGND.t456 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X1 VGND.t372 VPWR.t443 VGND.t372 VGND.t169 sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
X2 VGND.t378 VPWR.t444 VGND.t376 VGND.t377 sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
X3 VPWR.t301 VGND.t600 VPWR.t194 VPWR.t79 sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
X4 a_586_22008# dr[1].t0 VGND.t497 VGND.t559 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X5 a_1066_5376# db[3].t0 VGND.t368 VGND.t371 sg13_lv_nmos ad=0.2553p pd=2.17u as=0.1406p ps=1.12u w=0.74u l=0.13u
X6 VPWR.t235 VGND.t601 VPWR.t235 VPWR.t26 sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
X7 VGND.t380 VPWR.t445 VGND.t380 VGND.t382 sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
X8 VPWR.t205 VGND.t602 VPWR.t205 VPWR.t180 sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
X9 VGND.t586 dr[4].t0 a_490_19738# VGND.t154 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X10 a_490_3864# db[5].t0 VPWR.t126 VPWR.t123 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X11 VPWR.t297 VGND.t603 VPWR.t296 VPWR.t35 sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
X12 VGND.t289 dr[6].t0 a_1066_18226# VGND.t290 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X13 b[5].t3 a_490_3864# VGND.t455 VGND.t454 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.2516p ps=2.16u w=0.74u l=0.13u
X14 VGND.t385 VPWR.t446 VGND.t383 VGND.t260 sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
X15 VGND.t386 VPWR.t447 VGND.t386 VGND.t193 sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
X16 VGND.t31 a_1066_18226# r[6].t1 VGND.t35 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X17 VPWR.t349 a_1066_5376# b[3].t6 VPWR.t61 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X18 VPWR.t290 VGND.t604 VPWR.t290 VPWR.t26 sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
X19 VGND.t426 VPWR.t448 VGND.t424 VGND.t425 sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
X20 VGND.t240 a_490_18984# r[5].t1 VGND.t242 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X21 VPWR.t386 a_586_22008# r[1].t5 VPWR.t13 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X22 VGND.t33 a_1066_18226# r[6].t0 VGND.t34 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X23 b[3].t7 a_1066_5376# VPWR.t355 VPWR.t61 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X24 VPWR.t316 a_778_6888# b[1].t6 VPWR.t35 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X25 VPWR.t356 a_1066_5376# b[3].t4 VPWR.t61 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X26 VGND.t430 VPWR.t449 VGND.t428 VGND.t429 sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
X27 VPWR.t278 VGND.t605 VPWR.t278 VPWR.t61 sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
X28 VGND.t69 a_490_10666# g[6].t1 VGND.t73 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X29 VGND.t432 VPWR.t450 VGND.t432 VGND.t434 sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
X30 g[1].t3 a_490_14448# VGND.t79 VGND.t86 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X31 VPWR.t219 VGND.t606 VPWR.t219 VPWR.t9 sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
X32 VPWR.t217 VGND.t607 VPWR.t217 VPWR.t79 sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
X33 VPWR.t48 a_490_10666# g[6].t5 VPWR.t9 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X34 VGND.t437 VPWR.t451 VGND.t435 VGND.t164 sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
X35 a_490_19738# dr[4].t0 VPWR.t392 VPWR.t0 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X36 b[5].t6 a_490_3864# VPWR.t362 VPWR.t123 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X37 VGND.t570 a_490_13690# g[2].t2 VGND.t572 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X38 b[2].t3 a_490_6130# VGND.t52 VGND.t61 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X39 VPWR.t291 VGND.t608 VPWR.t290 VPWR.t26 sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
X40 VPWR.t85 a_490_22762# r[0].t5 VPWR.t79 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X41 VPWR.t289 VGND.t609 VPWR.t204 VPWR.t9 sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
X42 r[7].t3 a_490_17472# VGND.t323 VGND.t332 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X43 a_490_18984# dr[5].t0 VPWR.t90 VPWR.t17 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X44 VGND.t204 db[7].t0 a_490_2352# VGND.t205 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X45 b[5].t7 a_490_3864# VPWR.t368 VPWR.t123 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3864p ps=2.93u w=1.12u l=0.13u
X46 a_490_19738# dr[4].t0 VGND.t586 VGND.t152 sg13_lv_nmos ad=0.2553p pd=2.17u as=0.1406p ps=1.12u w=0.74u l=0.13u
X47 VPWR.t57 a_490_14448# g[1].t5 VPWR.t52 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X48 VGND.t306 a_1066_3106# b[6].t2 VGND.t305 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X49 VGND.t440 VPWR.t452 VGND.t438 VGND.t256 sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
X50 r[4].t3 a_490_19738# VGND.t509 VGND.t239 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X51 VGND.t590 dg[0].t0 a_1066_15202# VGND.t591 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X52 b[6].t3 a_1066_3106# VGND.t297 VGND.t304 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X53 VGND.t444 VPWR.t453 VGND.t442 VGND.t443 sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
X54 VGND.t299 a_1066_3106# b[6].t0 VGND.t303 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X55 VGND.t582 a_490_2352# b[7].t1 VGND.t584 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X56 a_1066_3106# db[6].t0 VPWR.t304 VPWR.t123 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X57 a_490_7642# db[0].t0 VGND.t265 VGND.t267 sg13_lv_nmos ad=0.2553p pd=2.17u as=0.1406p ps=1.12u w=0.74u l=0.13u
X58 VGND.t108 a_1066_15202# g[0].t1 VGND.t112 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X59 VPWR.t287 VGND.t610 VPWR.t286 VPWR.t13 sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
X60 r[6].t2 a_1066_18226# VGND.t33 VGND.t32 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X61 b[2].t2 a_490_6130# VGND.t50 VGND.t60 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X62 VGND.t471 VPWR.t454 VGND.t469 VGND.t379 sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
X63 VPWR.t308 a_1066_3106# b[6].t5 VPWR.t123 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X64 VGND.t48 a_490_7642# b[0].t1 VGND.t47 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X65 VGND.t362 a_490_11424# g[5].t1 VGND.t366 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X66 VGND.t475 VPWR.t455 VGND.t473 VGND.t474 sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
X67 VGND.t477 VPWR.t456 VGND.t477 VGND.t479 sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
X68 VGND.t110 a_1066_15202# g[0].t0 VGND.t111 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X69 VGND.t480 VPWR.t457 VGND.t480 VGND.t375 sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
X70 r[6].t7 a_1066_18226# VPWR.t20 VPWR.t17 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X71 g[2].t7 a_490_13690# VPWR.t417 VPWR.t52 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X72 a_1066_5376# db[3].t0 VPWR.t348 VPWR.t61 sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
X73 VPWR.t273 VGND.t611 VPWR.t273 VPWR.t91 sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
X74 VGND.t373 VPWR.t443 VGND.t372 VGND.t166 sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
X75 g[6].t3 a_490_10666# VGND.t72 VGND.t71 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.2516p ps=2.16u w=0.74u l=0.13u
X76 g[3].t7 a_1066_12936# VPWR.t328 VPWR.t180 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X77 r[0].t3 a_490_22762# VGND.t116 VGND.t125 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X78 VGND.t83 a_490_14448# g[1].t1 VGND.t85 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X79 g[6].t7 a_490_10666# VPWR.t50 VPWR.t9 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3864p ps=2.93u w=1.12u l=0.13u
X80 a_1066_4618# db[4].t0 VGND.t92 VGND.t464 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X81 b[2].t7 a_490_6130# VPWR.t37 VPWR.t35 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X82 VPWR.t395 a_490_19738# r[4].t5 VPWR.t0 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X83 VGND.t98 a_1066_4618# b[4].t1 VGND.t99 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X84 VGND.t580 a_490_2352# b[7].t0 VGND.t583 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X85 g[5].t7 a_490_11424# VPWR.t341 VPWR.t9 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X86 VPWR.t284 VGND.t612 VPWR.t179 VPWR.t91 sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
X87 VPWR.t374 db[4].t0 a_1066_4618# VPWR.t61 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X88 a_490_13690# dg[2].t0 VGND.t563 VGND.t595 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X89 VGND.t45 a_490_7642# b[0].t0 VGND.t46 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X90 VPWR.t120 a_490_18984# r[5].t5 VPWR.t17 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X91 VGND.t598 dr[7].t0 a_490_17472# VGND.t599 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X92 VPWR.t282 VGND.t613 VPWR.t193 VPWR.t52 sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
X93 b[4].t6 a_1066_4618# VPWR.t62 VPWR.t61 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X94 a_1066_12178# dg[4].t0 VGND.t507 VGND.t506 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X95 VGND.t486 VPWR.t458 VGND.t484 VGND.t485 sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
X96 VGND.t487 VPWR.t459 VGND.t487 VGND.t422 sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
X97 VGND.t519 VPWR.t460 VGND.t517 VGND.t518 sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
X98 VPWR.t260 VGND.t614 VPWR.t260 VPWR.t106 sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
X99 g[4].t3 a_1066_12178# VGND.t545 VGND.t555 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X100 g[1].t7 a_490_14448# VPWR.t59 VPWR.t52 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3864p ps=2.93u w=1.12u l=0.13u
X101 VPWR.t279 VGND.t615 VPWR.t278 VPWR.t61 sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
X102 VPWR.t435 dg[0].t0 a_1066_15202# VPWR.t70 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X103 g[4].t2 a_1066_12178# VGND.t554 VGND.t553 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.2516p ps=2.16u w=0.74u l=0.13u
X104 a_1066_3106# db[6].t0 VGND.t347 VGND.t349 sg13_lv_nmos ad=0.2553p pd=2.17u as=0.1406p ps=1.12u w=0.74u l=0.13u
X105 b[4].t7 a_1066_4618# VPWR.t63 VPWR.t61 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X106 VPWR.t181 VGND.t616 VPWR.t181 VPWR.t180 sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
X107 a_490_7642# db[0].t0 VPWR.t127 VPWR.t26 sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
X108 VPWR.t75 a_1066_15202# g[0].t5 VPWR.t70 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X109 b[2].t6 a_490_6130# VPWR.t36 VPWR.t35 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X110 g[0].t2 a_1066_15202# VGND.t110 VGND.t109 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X111 VPWR.t34 a_490_7642# b[0].t5 VPWR.t26 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X112 VGND.t292 dr[3].t0 a_1066_20496# VGND.t22 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X113 r[7].t7 a_490_17472# VPWR.t319 VPWR.t147 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X114 VPWR.t24 a_1066_18226# r[6].t7 VPWR.t17 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X115 VPWR.t76 a_1066_15202# g[0].t4 VPWR.t70 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X116 a_490_2352# db[7].t0 VPWR.t94 VPWR.t91 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X117 g[5].t3 a_490_11424# VGND.t365 VGND.t364 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.2516p ps=2.16u w=0.74u l=0.13u
X118 VGND.t521 VPWR.t461 VGND.t521 VGND.t523 sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
X119 VGND.t8 a_1066_20496# r[3].t1 VGND.t12 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X120 VPWR.t22 a_1066_18226# r[6].t4 VPWR.t17 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X121 VPWR.t419 a_490_13690# g[2].t5 VPWR.t52 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X122 VPWR.t332 a_1066_12936# g[3].t7 VPWR.t180 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X123 a_1066_5376# db[3].t0 VGND.t370 VGND.t369 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X124 VGND.t403 a_1066_5376# b[3].t1 VGND.t404 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X125 VGND.t10 a_1066_20496# r[3].t0 VGND.t11 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X126 VPWR.t330 a_1066_12936# g[3].t4 VPWR.t180 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X127 VGND.t501 a_586_22008# r[1].t1 VGND.t502 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X128 VGND.t391 db[1].t0 a_778_6888# VGND.t392 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X129 VGND.t17 a_490_10666# g[6].t0 VGND.t70 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X130 VGND.t538 dr[0].t0 a_490_22762# VGND.t539 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X131 a_490_14448# dg[1].t0 VGND.t75 VGND.t209 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X132 VPWR.t198 VGND.t617 VPWR.t198 VPWR.t79 sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
X133 VGND.t21 dr[2].t0 a_1066_21250# VGND.t22 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X134 VPWR.t12 a_490_10666# g[6].t4 VPWR.t9 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X135 a_1066_12936# dg[3].t0 VGND.t336 VGND.t460 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X136 a_1066_20496# dr[3].t0 VPWR.t2 VPWR.t0 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X137 a_490_17472# dr[7].t0 VGND.t598 VGND.t597 sg13_lv_nmos ad=0.2553p pd=2.17u as=0.1406p ps=1.12u w=0.74u l=0.13u
X138 VPWR.t32 a_490_7642# b[0].t4 VPWR.t26 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X139 VGND.t214 a_1066_21250# r[2].t1 VGND.t12 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X140 VGND.t568 a_490_13690# g[2].t0 VGND.t571 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X141 g[3].t3 a_1066_12936# VGND.t334 VGND.t345 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X142 r[3].t7 a_1066_20496# VPWR.t1 VPWR.t0 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X143 VGND.t524 VPWR.t462 VGND.t524 VGND.t197 sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
X144 VPWR.t338 dg[5].t0 a_490_11424# VPWR.t9 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X145 r[1].t7 a_586_22008# VPWR.t379 VPWR.t13 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X146 r[5].t3 a_490_18984# VGND.t232 VGND.t241 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X147 r[7].t2 a_490_17472# VGND.t321 VGND.t331 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X148 b[7].t7 a_490_2352# VPWR.t423 VPWR.t91 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X149 VPWR.t166 VGND.t618 VPWR.t166 VPWR.t140 sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
X150 VGND.t215 a_1066_21250# r[2].t0 VGND.t11 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X151 g[3].t2 a_1066_12936# VGND.t344 VGND.t343 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.2516p ps=2.16u w=0.74u l=0.13u
X152 VGND.t529 VPWR.t463 VGND.t528 VGND.t527 sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
X153 r[1].t6 a_586_22008# VPWR.t384 VPWR.t13 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3864p ps=2.93u w=1.12u l=0.13u
X154 r[3].t6 a_1066_20496# VPWR.t7 VPWR.t0 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3864p ps=2.93u w=1.12u l=0.13u
X155 VPWR.t274 VGND.t619 VPWR.t273 VPWR.t91 sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
X156 VGND.t246 db[5].t0 a_490_3864# VGND.t247 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X157 VPWR.t388 dg[4].t0 a_1066_12178# VPWR.t180 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X158 a_1066_18226# dr[6].t0 VGND.t289 VGND.t288 sg13_lv_nmos ad=0.2553p pd=2.17u as=0.1406p ps=1.12u w=0.74u l=0.13u
X159 VPWR.t58 a_490_14448# g[1].t4 VPWR.t52 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X160 b[7].t6 a_490_2352# VPWR.t429 VPWR.t91 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3864p ps=2.93u w=1.12u l=0.13u
X161 VPWR.t111 a_1066_9912# g[7].t4 VPWR.t106 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X162 VPWR.t408 a_1066_12178# g[4].t5 VPWR.t180 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X163 VPWR.t272 VGND.t620 VPWR.t201 VPWR.t147 sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
X164 g[0].t6 a_1066_15202# VPWR.t76 VPWR.t70 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X165 g[7].t7 a_1066_9912# VPWR.t113 VPWR.t106 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3864p ps=2.93u w=1.12u l=0.13u
X166 r[0].t7 a_490_22762# VPWR.t80 VPWR.t79 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X167 VGND.t451 a_490_3864# b[5].t4 VGND.t453 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X168 VPWR.t409 a_1066_12178# g[4].t4 VPWR.t180 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X169 VPWR.t352 db[1].t0 a_778_6888# VPWR.t35 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X170 b[1].t3 a_778_6888# VGND.t308 VGND.t319 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X171 VPWR.t270 VGND.t621 VPWR.t173 VPWR.t17 sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
X172 VGND.t532 VPWR.t464 VGND.t531 VGND.t530 sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
X173 VPWR.t441 dr[7].t0 a_490_17472# VPWR.t147 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X174 r[3].t2 a_1066_20496# VGND.t10 VGND.t9 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X175 VGND.t354 a_490_11424# g[5].t0 VGND.t363 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X176 VGND.t535 VPWR.t465 VGND.t533 VGND.t476 sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
X177 r[1].t3 a_586_22008# VGND.t501 VGND.t500 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X178 VPWR.t268 VGND.t622 VPWR.t197 VPWR.t70 sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
X179 VPWR.t266 VGND.t623 VPWR.t169 VPWR.t0 sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
X180 VGND.t178 VPWR.t466 VGND.t178 VGND.t180 sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
X181 a_490_13690# dg[2].t0 VPWR.t415 VPWR.t52 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X182 VGND.t488 VPWR.t459 VGND.t487 VGND.t419 sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
X183 a_490_22762# dr[0].t0 VGND.t538 VGND.t537 sg13_lv_nmos ad=0.2553p pd=2.17u as=0.1406p ps=1.12u w=0.74u l=0.13u
X184 VPWR.t239 VGND.t624 VPWR.t239 VPWR.t123 sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
X185 VPWR.t263 VGND.t625 VPWR.t196 VPWR.t13 sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
X186 VPWR.t261 VGND.t626 VPWR.t260 VPWR.t106 sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
X187 VGND.t511 a_490_19738# r[4].t0 VGND.t238 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X188 VGND.t182 VPWR.t467 VGND.t182 VGND.t184 sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
X189 VPWR.t259 VGND.t627 VPWR.t258 VPWR.t35 sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
X190 r[0].t2 a_490_22762# VGND.t114 VGND.t124 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X191 VGND.t81 a_490_14448# g[1].t3 VGND.t84 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X192 VGND.t186 VPWR.t468 VGND.t186 VGND.t188 sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
X193 VPWR.t15 dr[2].t0 a_1066_21250# VPWR.t13 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X194 a_1066_9912# dg[7].t0 VGND.t221 VGND.t543 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X195 a_490_11424# dg[5].t0 VPWR.t338 VPWR.t9 sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
X196 VPWR.t124 db[5].t0 a_490_3864# VPWR.t123 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X197 VPWR.t102 a_1066_21250# r[2].t5 VPWR.t13 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X198 g[7].t3 a_1066_9912# VGND.t219 VGND.t230 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X199 r[2].t2 a_1066_21250# VGND.t215 VGND.t9 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X200 VGND.t449 a_490_3864# b[5].t3 VGND.t452 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X201 VGND.t192 VPWR.t469 VGND.t190 VGND.t191 sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
X202 g[5].t6 a_490_11424# VPWR.t340 VPWR.t9 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X203 VPWR.t103 a_1066_21250# r[2].t4 VPWR.t13 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X204 g[7].t2 a_1066_9912# VGND.t229 VGND.t228 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.2516p ps=2.16u w=0.74u l=0.13u
X205 VGND.t196 VPWR.t470 VGND.t194 VGND.t195 sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
X206 a_1066_5376# db[3].t0 VPWR.t349 VPWR.t61 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X207 VGND.t153 dr[5].t0 a_490_18984# VGND.t154 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X208 VPWR.t257 VGND.t628 VPWR.t148 VPWR.t147 sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
X209 VPWR.t365 a_490_3864# b[5].t6 VPWR.t123 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X210 VGND.t183 VPWR.t467 VGND.t182 VGND.t181 sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
X211 VPWR.t357 a_1066_5376# b[3].t7 VPWR.t61 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X212 a_1066_15202# dg[0].t0 VGND.t590 VGND.t589 sg13_lv_nmos ad=0.2553p pd=2.17u as=0.1406p ps=1.12u w=0.74u l=0.13u
X213 VPWR.t229 VGND.t629 VPWR.t229 VPWR.t106 sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
X214 b[1].t7 a_778_6888# VPWR.t316 VPWR.t35 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X215 g[4].t6 a_1066_12178# VPWR.t409 VPWR.t180 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X216 r[4].t7 a_490_19738# VPWR.t390 VPWR.t0 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X217 VGND.t200 VPWR.t471 VGND.t198 VGND.t199 sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
X218 VPWR.t254 VGND.t630 VPWR.t143 VPWR.t70 sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
X219 VPWR.t153 VGND.t631 VPWR.t153 VPWR.t140 sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
X220 r[1].t2 a_586_22008# VGND.t491 VGND.t499 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X221 a_490_17472# dr[7].t0 VPWR.t441 VPWR.t147 sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
X222 a_490_6130# db[2].t0 VGND.t466 VGND.t468 sg13_lv_nmos ad=0.2553p pd=2.17u as=0.1406p ps=1.12u w=0.74u l=0.13u
X223 VPWR.t399 dr[0].t0 a_490_22762# VPWR.t79 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X224 VGND.t156 VPWR.t472 VGND.t156 VGND.t158 sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
X225 VGND.t59 a_490_6130# b[2].t3 VGND.t58 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X226 r[5].t7 a_490_18984# VPWR.t115 VPWR.t17 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X227 r[7].t6 a_490_17472# VPWR.t318 VPWR.t147 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X228 VPWR.t251 VGND.t632 VPWR.t146 VPWR.t106 sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
X229 VGND.t161 VPWR.t473 VGND.t159 VGND.t142 sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
X230 VGND.t165 VPWR.t474 VGND.t163 VGND.t164 sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
X231 VPWR.t249 VGND.t633 VPWR.t188 VPWR.t0 sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
X232 VPWR.t418 a_490_13690# g[2].t7 VPWR.t52 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X233 VGND.t557 dr[1].t0 a_586_22008# VGND.t558 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X234 VGND.t167 VPWR.t475 VGND.t167 VGND.t169 sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
X235 VPWR.t247 VGND.t634 VPWR.t185 VPWR.t17 sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
X236 r[4].t2 a_490_19738# VGND.t513 VGND.t236 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.2516p ps=2.16u w=0.74u l=0.13u
X237 VPWR.t364 a_490_3864# b[5].t7 VPWR.t123 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X238 VPWR.t175 VGND.t635 VPWR.t175 VPWR.t147 sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
X239 VPWR.t380 a_586_22008# r[1].t7 VPWR.t13 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X240 a_1066_3106# db[6].t0 VGND.t306 VGND.t348 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X241 VGND.t301 a_1066_3106# b[6].t3 VGND.t302 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X242 VGND.t157 VPWR.t472 VGND.t156 VGND.t155 sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
X243 r[2].t6 a_1066_21250# VPWR.t103 VPWR.t13 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X244 b[7].t3 a_490_2352# VGND.t582 VGND.t581 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X245 a_490_18984# dr[5].t0 VGND.t153 VGND.t152 sg13_lv_nmos ad=0.2553p pd=2.17u as=0.1406p ps=1.12u w=0.74u l=0.13u
X246 VPWR.t171 VGND.t636 VPWR.t171 VPWR.t70 sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
X247 VPWR.t334 db[6].t0 a_1066_3106# VPWR.t123 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X248 r[6].t3 a_1066_18226# VGND.t31 VGND.t30 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X249 VGND.t172 VPWR.t476 VGND.t170 VGND.t130 sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
X250 VGND.t56 a_490_6130# b[2].t2 VGND.t57 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X251 b[6].t6 a_1066_3106# VPWR.t308 VPWR.t123 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X252 a_490_7642# db[0].t0 VGND.t48 VGND.t266 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X253 VPWR.t243 VGND.t637 VPWR.t152 VPWR.t140 sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
X254 r[5].t2 a_490_18984# VGND.t240 VGND.t239 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X255 a_586_22008# dr[1].t0 VPWR.t386 VPWR.t13 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X256 a_1066_15202# dg[0].t0 VPWR.t435 VPWR.t70 sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
X257 VPWR.t222 VGND.t638 VPWR.t222 VPWR.t26 sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
X258 g[6].t2 a_490_10666# VGND.t69 VGND.t68 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X259 VPWR.t240 VGND.t639 VPWR.t239 VPWR.t123 sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
X260 g[6].t6 a_490_10666# VPWR.t48 VPWR.t9 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X261 a_1066_20496# dr[3].t0 VGND.t292 VGND.t20 sg13_lv_nmos ad=0.2553p pd=2.17u as=0.1406p ps=1.12u w=0.74u l=0.13u
X262 b[6].t7 a_1066_3106# VPWR.t302 VPWR.t123 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X263 VPWR.t231 VGND.t640 VPWR.t231 VPWR.t26 sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
X264 VPWR.t144 VGND.t641 VPWR.t144 VPWR.t79 sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
X265 a_490_22762# dr[0].t0 VPWR.t399 VPWR.t79 sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
X266 a_490_6130# db[2].t0 VPWR.t376 VPWR.t35 sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
X267 VGND.t462 db[4].t0 a_1066_4618# VGND.t463 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X268 VGND.t174 VPWR.t477 VGND.t174 VGND.t176 sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
X269 VPWR.t431 dr[4].t0 a_490_19738# VPWR.t0 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X270 VPWR.t41 a_490_6130# b[2].t7 VPWR.t35 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X271 g[2].t3 a_490_13690# VGND.t570 VGND.t569 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X272 b[4].t2 a_1066_4618# VGND.t98 VGND.t97 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X273 r[0].t6 a_490_22762# VPWR.t85 VPWR.t79 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X274 VGND.t325 a_490_17472# r[7].t3 VGND.t330 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X275 b[7].t2 a_490_2352# VGND.t580 VGND.t579 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X276 VPWR.t236 VGND.t642 VPWR.t235 VPWR.t26 sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
X277 VPWR.t88 dr[5].t0 a_490_18984# VPWR.t17 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X278 b[0].t3 a_490_7642# VGND.t45 VGND.t44 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X279 VGND.t129 VPWR.t478 VGND.t127 VGND.t128 sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
X280 VPWR.t234 VGND.t643 VPWR.t168 VPWR.t70 sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
X281 g[1].t6 a_490_14448# VPWR.t57 VPWR.t52 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X282 b[4].t3 a_1066_4618# VGND.t88 VGND.t96 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X283 VPWR.t232 VGND.t644 VPWR.t231 VPWR.t26 sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
X284 a_1066_21250# dr[2].t0 VGND.t21 VGND.t20 sg13_lv_nmos ad=0.2553p pd=2.17u as=0.1406p ps=1.12u w=0.74u l=0.13u
X285 VGND.t131 VPWR.t479 VGND.t131 VGND.t133 sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
X286 VPWR.t230 VGND.t645 VPWR.t229 VPWR.t106 sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
X287 VPWR.t228 VGND.t646 VPWR.t149 VPWR.t147 sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
X288 VGND.t512 a_490_19738# r[4].t3 VGND.t235 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X289 VGND.t137 VPWR.t480 VGND.t135 VGND.t136 sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
X290 VGND.t139 VPWR.t481 VGND.t139 VGND.t141 sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
X291 VGND.t29 a_1066_18226# r[6].t3 VGND.t28 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X292 b[0].t2 a_490_7642# VGND.t43 VGND.t42 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.2516p ps=2.16u w=0.74u l=0.13u
X293 VPWR.t64 a_1066_4618# b[4].t7 VPWR.t61 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X294 g[0].t3 a_1066_15202# VGND.t108 VGND.t107 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X295 b[4].t5 a_1066_4618# VPWR.t66 VPWR.t61 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3864p ps=2.93u w=1.12u l=0.13u
X296 VPWR.t39 a_490_6130# b[2].t6 VPWR.t35 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X297 a_490_7642# db[0].t0 VPWR.t34 VPWR.t26 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X298 VGND.t143 VPWR.t482 VGND.t143 VGND.t145 sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
X299 VGND.t26 a_1066_18226# r[6].t2 VGND.t27 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X300 g[5].t2 a_490_11424# VGND.t362 VGND.t361 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X301 VGND.t147 VPWR.t483 VGND.t147 VGND.t149 sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
X302 VPWR.t92 db[7].t0 a_490_2352# VPWR.t91 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X303 a_1066_12178# dg[4].t0 VPWR.t388 VPWR.t180 sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
X304 VGND.t376 VPWR.t444 VGND.t376 VGND.t375 sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
X305 VPWR.t183 VGND.t647 VPWR.t183 VPWR.t155 sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
X306 VGND.t368 db[3].t0 a_1066_5376# VGND.t367 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X307 VGND.t140 VPWR.t481 VGND.t139 VGND.t138 sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
X308 VGND.t65 a_490_10666# g[6].t3 VGND.t67 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X309 VGND.t168 VPWR.t475 VGND.t167 VGND.t166 sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
X310 VGND.t118 a_490_22762# r[0].t3 VGND.t123 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X311 g[1].t2 a_490_14448# VGND.t83 VGND.t82 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X312 b[3].t2 a_1066_5376# VGND.t403 VGND.t402 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X313 a_490_19738# dr[4].t0 VPWR.t431 VPWR.t0 sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
X314 a_778_6888# db[1].t0 VGND.t391 VGND.t390 sg13_lv_nmos ad=0.2553p pd=2.17u as=0.1406p ps=1.12u w=0.74u l=0.13u
X315 VPWR.t45 a_490_10666# g[6].t7 VPWR.t9 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X316 VGND.t271 VPWR.t484 VGND.t269 VGND.t270 sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
X317 VPWR.t426 a_490_2352# b[7].t7 VPWR.t91 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X318 VPWR.t225 VGND.t648 VPWR.t141 VPWR.t140 sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
X319 r[4].t6 a_490_19738# VPWR.t395 VPWR.t0 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X320 VGND.t148 VPWR.t483 VGND.t147 VGND.t146 sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
X321 a_490_18984# dr[5].t0 VPWR.t88 VPWR.t17 sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
X322 VPWR.t342 a_490_11424# g[5].t7 VPWR.t9 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X323 r[7].t1 a_490_17472# VGND.t329 VGND.t328 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.2516p ps=2.16u w=0.74u l=0.13u
X324 VGND.t593 dg[2].t0 a_490_13690# VGND.t594 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X325 b[3].t3 a_1066_5376# VGND.t394 VGND.t401 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X326 b[0].t7 a_490_7642# VPWR.t32 VPWR.t26 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X327 r[5].t6 a_490_18984# VPWR.t120 VPWR.t17 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X328 b[1].t2 a_778_6888# VGND.t310 VGND.t318 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X329 VGND.t274 VPWR.t485 VGND.t273 VGND.t272 sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
X330 VGND.t504 dg[4].t0 a_1066_12178# VGND.t505 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X331 VGND.t312 a_778_6888# b[1].t3 VGND.t317 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X332 a_1066_21250# dr[2].t0 VPWR.t15 VPWR.t13 sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
X333 VGND.t276 VPWR.t486 VGND.t276 VGND.t278 sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
X334 VGND.t548 a_1066_12178# g[4].t3 VGND.t552 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X335 VPWR.t54 a_490_14448# g[1].t7 VPWR.t52 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X336 VPWR.t223 VGND.t649 VPWR.t222 VPWR.t26 sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
X337 VGND.t106 a_1066_15202# g[0].t3 VGND.t105 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X338 b[0].t6 a_490_7642# VPWR.t31 VPWR.t26 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3864p ps=2.93u w=1.12u l=0.13u
X339 VPWR.t112 a_1066_9912# g[7].t5 VPWR.t106 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X340 VGND.t550 a_1066_12178# g[4].t2 VGND.t551 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X341 VGND.t435 VPWR.t451 VGND.t435 VGND.t162 sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
X342 g[0].t7 a_1066_15202# VPWR.t75 VPWR.t70 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X343 VPWR.t425 a_490_2352# b[7].t6 VPWR.t91 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X344 g[7].t6 a_1066_9912# VPWR.t111 VPWR.t106 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X345 VGND.t103 a_1066_15202# g[0].t2 VGND.t104 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X346 VGND.t175 VPWR.t477 VGND.t174 VGND.t173 sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
X347 VPWR.t107 a_1066_9912# g[7].t7 VPWR.t106 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X348 VPWR.t320 a_490_17472# r[7].t7 VPWR.t147 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X349 a_1066_18226# dr[6].t0 VPWR.t24 VPWR.t17 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X350 b[5].t2 a_490_3864# VGND.t451 VGND.t450 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X351 VGND.t358 a_490_11424# g[5].t3 VGND.t360 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X352 a_778_6888# db[1].t0 VPWR.t352 VPWR.t35 sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
X353 VGND.t387 VPWR.t447 VGND.t386 VGND.t195 sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
X354 r[3].t3 a_1066_20496# VGND.t8 VGND.t7 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X355 r[6].t6 a_1066_18226# VPWR.t22 VPWR.t17 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X356 g[2].t6 a_490_13690# VPWR.t419 VPWR.t52 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X357 b[1].t0 a_778_6888# VGND.t316 VGND.t315 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.2516p ps=2.16u w=0.74u l=0.13u
X358 a_1066_12936# dg[3].t0 VPWR.t332 VPWR.t180 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X359 VPWR.t214 VGND.t650 VPWR.t214 VPWR.t123 sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
X360 g[3].t6 a_1066_12936# VPWR.t330 VPWR.t180 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X361 r[0].t1 a_490_22762# VGND.t122 VGND.t121 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.2516p ps=2.16u w=0.74u l=0.13u
X362 r[6].t5 a_1066_18226# VPWR.t21 VPWR.t17 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3864p ps=2.93u w=1.12u l=0.13u
X363 a_490_10666# dg[6].t0 VGND.t17 VGND.t16 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X364 VGND.t433 VPWR.t450 VGND.t432 VGND.t431 sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
X365 b[1].t5 a_778_6888# VPWR.t310 VPWR.t35 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X366 VPWR.t220 VGND.t651 VPWR.t219 VPWR.t9 sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
X367 VPWR.t218 VGND.t652 VPWR.t217 VPWR.t79 sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
X368 VGND.t207 dg[1].t0 a_490_14448# VGND.t208 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X369 g[3].t5 a_1066_12936# VPWR.t329 VPWR.t180 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3864p ps=2.93u w=1.12u l=0.13u
X370 VGND.t282 VPWR.t487 VGND.t280 VGND.t281 sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
X371 a_490_13690# dg[2].t0 VGND.t593 VGND.t592 sg13_lv_nmos ad=0.2553p pd=2.17u as=0.1406p ps=1.12u w=0.74u l=0.13u
X372 a_490_10666# dg[6].t0 VPWR.t12 VPWR.t9 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X373 VGND.t458 dg[3].t0 a_1066_12936# VGND.t459 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X374 VPWR.t311 a_778_6888# b[1].t7 VPWR.t35 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X375 VPWR.t133 dr[3].t0 a_1066_20496# VPWR.t0 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X376 VGND.t469 VPWR.t454 VGND.t469 VGND.t382 sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
X377 g[5].t5 a_490_11424# VPWR.t344 VPWR.t9 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3864p ps=2.93u w=1.12u l=0.13u
X378 VPWR.t158 VGND.t653 VPWR.t158 VPWR.t140 sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
X379 r[2].t3 a_1066_21250# VGND.t214 VGND.t7 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X380 g[2].t1 a_490_13690# VGND.t568 VGND.t567 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X381 VGND.t338 a_1066_12936# g[3].t3 VGND.t342 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X382 VPWR.t3 a_1066_20496# r[3].t7 VPWR.t0 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X383 b[5].t1 a_490_3864# VGND.t449 VGND.t448 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X384 VGND.t234 a_490_18984# r[5].t3 VGND.t238 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X385 VGND.t327 a_490_17472# r[7].t2 VGND.t326 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X386 VGND.t340 a_1066_12936# g[3].t2 VGND.t341 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X387 VPWR.t215 VGND.t654 VPWR.t214 VPWR.t123 sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
X388 VPWR.t348 db[3].t0 a_1066_5376# VPWR.t61 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X389 VPWR.t4 a_1066_20496# r[3].t6 VPWR.t0 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X390 VPWR.t202 VGND.t655 VPWR.t202 VPWR.t155 sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
X391 g[4].t0 a_1066_12178# VGND.t550 VGND.t549 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X392 VPWR.t381 a_586_22008# r[1].t6 VPWR.t13 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X393 VPWR.t74 a_1066_15202# g[0].t7 VPWR.t70 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X394 b[5].t0 a_490_3864# VPWR.t365 VPWR.t123 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X395 b[3].t6 a_1066_5376# VPWR.t357 VPWR.t61 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X396 a_490_14448# dg[1].t0 VPWR.t58 VPWR.t52 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X397 g[4].t7 a_1066_12178# VPWR.t408 VPWR.t180 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X398 VGND.t284 VPWR.t488 VGND.t284 VGND.t286 sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
X399 b[1].t6 a_778_6888# VPWR.t313 VPWR.t35 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3864p ps=2.93u w=1.12u l=0.13u
X400 VPWR.t72 a_1066_15202# g[0].t6 VPWR.t70 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X401 a_1066_9912# dg[7].t0 VPWR.t401 VPWR.t106 sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
X402 VPWR.t81 a_490_22762# r[0].t7 VPWR.t79 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X403 VGND.t6 a_1066_20496# r[3].t3 VGND.t5 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X404 r[7].t5 a_490_17472# VPWR.t322 VPWR.t147 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3864p ps=2.93u w=1.12u l=0.13u
X405 VPWR.t136 VGND.t656 VPWR.t136 VPWR.t52 sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
X406 b[3].t5 a_1066_5376# VPWR.t356 VPWR.t61 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X407 VGND.t484 VPWR.t458 VGND.t484 VGND.t483 sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
X408 a_490_6130# db[2].t0 VGND.t59 VGND.t467 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X409 VGND.t517 VPWR.t460 VGND.t517 VGND.t516 sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
X410 VGND.t3 a_1066_20496# r[3].t2 VGND.t4 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X411 a_490_11424# dg[5].t0 VGND.t354 VGND.t353 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X412 VGND.t495 a_586_22008# r[1].t3 VGND.t498 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X413 VGND.t478 VPWR.t456 VGND.t477 VGND.t476 sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
X414 VPWR.t437 dg[2].t0 a_490_13690# VPWR.t52 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X415 VPWR.t156 VGND.t657 VPWR.t156 VPWR.t155 sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
X416 a_490_14448# dg[1].t0 VGND.t207 VGND.t206 sg13_lv_nmos ad=0.2553p pd=2.17u as=0.1406p ps=1.12u w=0.74u l=0.13u
X417 VGND.t249 VPWR.t489 VGND.t249 VGND.t251 sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
X418 VGND.t63 a_490_10666# g[6].t2 VGND.t66 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X419 r[4].t1 a_490_19738# VGND.t511 VGND.t233 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X420 b[5].t5 a_490_3864# VPWR.t364 VPWR.t123 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X421 VGND.t120 a_490_22762# r[0].t2 VGND.t119 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X422 g[1].t0 a_490_14448# VGND.t81 VGND.t80 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X423 VGND.t255 VPWR.t490 VGND.t253 VGND.t254 sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
X424 VPWR.t208 VGND.t658 VPWR.t208 VPWR.t35 sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
X425 VGND.t541 dg[7].t0 a_1066_9912# VGND.t542 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X426 VGND.t19 a_1066_21250# r[2].t3 VGND.t5 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X427 VGND.t347 db[6].t0 a_1066_3106# VGND.t346 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X428 VPWR.t44 a_490_10666# g[6].t6 VPWR.t9 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X429 a_490_2352# db[7].t0 VGND.t204 VGND.t203 sg13_lv_nmos ad=0.2553p pd=2.17u as=0.1406p ps=1.12u w=0.74u l=0.13u
X430 r[2].t7 a_1066_21250# VPWR.t102 VPWR.t13 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X431 b[6].t2 a_1066_3106# VGND.t301 VGND.t300 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X432 VGND.t223 a_1066_9912# g[7].t3 VGND.t227 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X433 VGND.t211 a_1066_21250# r[2].t2 VGND.t4 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X434 g[3].t0 a_1066_12936# VGND.t340 VGND.t339 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X435 VGND.t202 a_490_2352# b[7].t3 VGND.t578 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X436 r[3].t4 a_1066_20496# VPWR.t4 VPWR.t0 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X437 VPWR.t337 a_490_11424# g[5].t6 VPWR.t9 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X438 r[1].t4 a_586_22008# VPWR.t381 VPWR.t13 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X439 r[5].t0 a_490_18984# VGND.t237 VGND.t236 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.2516p ps=2.16u w=0.74u l=0.13u
X440 VGND.t225 a_1066_9912# g[7].t2 VGND.t226 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X441 VGND.t250 VPWR.t489 VGND.t249 VGND.t248 sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
X442 b[2].t1 a_490_6130# VGND.t56 VGND.t55 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X443 VGND.t265 db[0].t0 a_490_7642# VGND.t264 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X444 b[6].t1 a_1066_3106# VGND.t299 VGND.t298 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X445 VPWR.t387 a_1066_12178# g[4].t7 VPWR.t180 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X446 VPWR.t209 VGND.t659 VPWR.t208 VPWR.t35 sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
X447 VPWR.t53 a_490_14448# g[1].t6 VPWR.t52 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X448 VGND.t381 VPWR.t445 VGND.t380 VGND.t379 sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
X449 VPWR.t150 VGND.t660 VPWR.t150 VPWR.t140 sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
X450 VPWR.t405 a_1066_12178# g[4].t6 VPWR.t180 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X451 VPWR.t206 VGND.t661 VPWR.t205 VPWR.t180 sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
X452 VPWR.t391 a_490_19738# r[4].t7 VPWR.t0 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X453 b[2].t0 a_490_6130# VGND.t54 VGND.t53 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.2516p ps=2.16u w=0.74u l=0.13u
X454 VGND.t39 a_490_7642# b[0].t3 VGND.t41 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X455 r[0].t4 a_490_22762# VPWR.t83 VPWR.t79 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3864p ps=2.93u w=1.12u l=0.13u
X456 VPWR.t303 a_1066_3106# b[6].t7 VPWR.t123 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X457 VPWR.t204 VGND.t662 VPWR.t204 VPWR.t9 sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
X458 b[6].t4 a_1066_3106# VPWR.t305 VPWR.t123 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3864p ps=2.93u w=1.12u l=0.13u
X459 a_490_6130# db[2].t0 VPWR.t41 VPWR.t35 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X460 VPWR.t116 a_490_18984# r[5].t7 VPWR.t17 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X461 VPWR.t321 a_490_17472# r[7].t6 VPWR.t147 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X462 a_490_13690# dg[2].t0 VPWR.t437 VPWR.t52 sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
X463 VGND.t576 a_490_2352# b[7].t2 VGND.t577 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X464 VGND.t356 a_490_11424# g[5].t2 VGND.t359 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X465 VPWR.t203 VGND.t663 VPWR.t202 VPWR.t155 sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
X466 g[2].t4 a_490_13690# VPWR.t418 VPWR.t52 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X467 a_586_22008# dr[1].t0 VGND.t557 VGND.t556 sg13_lv_nmos ad=0.2553p pd=2.17u as=0.1406p ps=1.12u w=0.74u l=0.13u
X468 VGND.t508 a_490_19738# r[4].t2 VGND.t231 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X469 VGND.t90 a_1066_4618# b[4].t3 VGND.t95 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X470 VPWR.t14 a_1066_21250# r[2].t7 VPWR.t13 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X471 VPWR.t201 VGND.t664 VPWR.t201 VPWR.t147 sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
X472 r[1].t5 a_586_22008# VPWR.t380 VPWR.t13 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X473 VPWR.t190 VGND.t665 VPWR.t190 VPWR.t155 sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
X474 b[4].t0 a_1066_4618# VGND.t94 VGND.t93 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.2516p ps=2.16u w=0.74u l=0.13u
X475 VPWR.t199 VGND.t666 VPWR.t198 VPWR.t79 sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
X476 VPWR.t65 a_1066_4618# b[4].t6 VPWR.t61 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X477 VGND.t285 VPWR.t488 VGND.t284 VGND.t283 sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
X478 VPWR.t99 a_1066_21250# r[2].t6 VPWR.t13 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X479 VGND.t37 a_490_7642# b[0].t2 VGND.t40 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X480 g[7].t0 a_1066_9912# VGND.t225 VGND.t224 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X481 a_1066_12178# dg[4].t0 VGND.t504 VGND.t503 sg13_lv_nmos ad=0.2553p pd=2.17u as=0.1406p ps=1.12u w=0.74u l=0.13u
X482 b[4].t4 a_1066_4618# VPWR.t64 VPWR.t61 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X483 VGND.t473 VPWR.t455 VGND.t473 VGND.t472 sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
X484 VPWR.t197 VGND.t667 VPWR.t197 VPWR.t70 sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
X485 VPWR.t63 a_1066_4618# b[4].t5 VPWR.t61 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X486 b[2].t5 a_490_6130# VPWR.t39 VPWR.t35 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X487 VPWR.t127 db[0].t0 a_490_7642# VPWR.t26 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X488 VGND.t151 a_490_18984# r[5].t2 VGND.t235 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X489 VPWR.t412 dr[1].t0 a_586_22008# VPWR.t13 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X490 VPWR.t196 VGND.t668 VPWR.t196 VPWR.t13 sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
X491 VGND.t257 VPWR.t491 VGND.t257 VGND.t259 sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
X492 VPWR.t177 VGND.t669 VPWR.t177 VPWR.t155 sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
X493 VPWR.t194 VGND.t670 VPWR.t194 VPWR.t79 sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
X494 b[2].t4 a_490_6130# VPWR.t38 VPWR.t35 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3864p ps=2.93u w=1.12u l=0.13u
X495 r[4].t4 a_490_19738# VPWR.t393 VPWR.t0 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3864p ps=2.93u w=1.12u l=0.13u
X496 VPWR.t28 a_490_7642# b[0].t7 VPWR.t26 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X497 b[7].t5 a_490_2352# VPWR.t426 VPWR.t91 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X498 VGND.t561 a_490_13690# g[2].t3 VGND.t566 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X499 VPWR.t82 a_490_22762# r[0].t6 VPWR.t79 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X500 VPWR.t193 VGND.t671 VPWR.t193 VPWR.t52 sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
X501 r[5].t4 a_490_18984# VPWR.t118 VPWR.t17 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3864p ps=2.93u w=1.12u l=0.13u
X502 r[7].t0 a_490_17472# VGND.t325 VGND.t324 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X503 VGND.t261 VPWR.t492 VGND.t261 VGND.t263 sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
X504 VGND.t396 a_1066_5376# b[3].t3 VGND.t400 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X505 VGND.t314 a_778_6888# b[1].t2 VGND.t313 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X506 VGND.t481 VPWR.t457 VGND.t480 VGND.t377 sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
X507 VGND.t497 a_586_22008# r[1].t2 VGND.t496 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X508 b[3].t0 a_1066_5376# VGND.t399 VGND.t398 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.2516p ps=2.16u w=0.74u l=0.13u
X509 VPWR.t186 VGND.t672 VPWR.t186 VPWR.t91 sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
X510 VPWR.t191 VGND.t673 VPWR.t190 VPWR.t155 sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
X511 b[1].t1 a_778_6888# VGND.t312 VGND.t311 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X512 a_1066_12936# dg[3].t0 VGND.t458 VGND.t457 sg13_lv_nmos ad=0.2553p pd=2.17u as=0.1406p ps=1.12u w=0.74u l=0.13u
X513 a_1066_20496# dr[3].t0 VPWR.t133 VPWR.t0 sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
X514 a_490_19738# dr[4].t0 VGND.t512 VGND.t150 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X515 VGND.t198 VPWR.t471 VGND.t198 VGND.t197 sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
X516 a_1066_18226# dr[6].t0 VGND.t29 VGND.t287 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X517 VPWR.t27 a_490_7642# b[0].t6 VPWR.t26 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X518 a_1066_9912# dg[7].t0 VPWR.t112 VPWR.t106 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X519 VGND.t187 VPWR.t468 VGND.t186 VGND.t185 sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
X520 VPWR.t162 VGND.t674 VPWR.t162 VPWR.t61 sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
X521 b[7].t4 a_490_2352# VPWR.t425 VPWR.t91 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X522 VGND.t262 VPWR.t492 VGND.t261 VGND.t260 sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
X523 VPWR.t108 a_1066_9912# g[7].t6 VPWR.t106 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X524 a_490_3864# db[5].t0 VGND.t246 VGND.t245 sg13_lv_nmos ad=0.2553p pd=2.17u as=0.1406p ps=1.12u w=0.74u l=0.13u
X525 a_1066_4618# db[4].t0 VPWR.t374 VPWR.t61 sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
X526 r[6].t1 a_1066_18226# VGND.t26 VGND.t25 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X527 VGND.t159 VPWR.t473 VGND.t159 VGND.t145 sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
X528 VGND.t163 VPWR.t474 VGND.t163 VGND.t162 sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
X529 VGND.t244 a_490_3864# b[5].t2 VGND.t447 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X530 VGND.t424 VPWR.t448 VGND.t424 VGND.t423 sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
X531 VPWR.t188 VGND.t675 VPWR.t188 VPWR.t0 sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
X532 VPWR.t187 VGND.t676 VPWR.t186 VPWR.t91 sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
X533 VPWR.t185 VGND.t677 VPWR.t185 VPWR.t17 sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
X534 r[6].t0 a_1066_18226# VGND.t24 VGND.t23 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.2516p ps=2.16u w=0.74u l=0.13u
X535 VPWR.t184 VGND.t678 VPWR.t183 VPWR.t155 sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
X536 g[6].t1 a_490_10666# VGND.t65 VGND.t64 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X537 r[0].t0 a_490_22762# VGND.t118 VGND.t117 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X538 VGND.t79 a_490_14448# g[1].t2 VGND.t78 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X539 g[6].t5 a_490_10666# VPWR.t45 VPWR.t9 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X540 VPWR.t312 a_778_6888# b[1].t5 VPWR.t35 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X541 VPWR.t182 VGND.t679 VPWR.t181 VPWR.t180 sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
X542 VPWR.t392 a_490_19738# r[4].t6 VPWR.t0 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X543 g[2].t2 a_490_13690# VGND.t565 VGND.t564 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.2516p ps=2.16u w=0.74u l=0.13u
X544 b[1].t4 a_778_6888# VPWR.t311 VPWR.t35 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X545 g[5].t4 a_490_11424# VPWR.t342 VPWR.t9 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X546 VGND.t323 a_490_17472# r[7].t1 VGND.t322 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X547 VPWR.t90 a_490_18984# r[5].t6 VPWR.t17 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X548 VGND.t522 VPWR.t461 VGND.t521 VGND.t520 sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
X549 VGND.t446 a_490_3864# b[5].t1 VGND.t445 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X550 VPWR.t179 VGND.t680 VPWR.t179 VPWR.t91 sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
X551 VPWR.t178 VGND.t681 VPWR.t177 VPWR.t155 sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
X552 a_1066_9912# dg[7].t0 VGND.t541 VGND.t540 sg13_lv_nmos ad=0.2553p pd=2.17u as=0.1406p ps=1.12u w=0.74u l=0.13u
X553 g[4].t1 a_1066_12178# VGND.t548 VGND.t547 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X554 g[1].t5 a_490_14448# VPWR.t54 VPWR.t52 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X555 a_490_3864# db[5].t0 VPWR.t124 VPWR.t123 sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
X556 VGND.t258 VPWR.t491 VGND.t257 VGND.t256 sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
X557 VGND.t509 a_490_19738# r[4].t1 VGND.t242 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X558 VPWR.t176 VGND.t682 VPWR.t175 VPWR.t147 sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
X559 a_1066_15202# dg[0].t0 VGND.t106 VGND.t588 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X560 VPWR.t126 a_490_3864# b[5].t0 VPWR.t123 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X561 VGND.t406 VPWR.t493 VGND.t406 VGND.t408 sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
X562 VPWR.t160 VGND.t683 VPWR.t160 VPWR.t155 sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
X563 g[0].t1 a_1066_15202# VGND.t103 VGND.t102 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X564 VPWR.t173 VGND.t684 VPWR.t173 VPWR.t17 sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
X565 r[7].t4 a_490_17472# VPWR.t320 VPWR.t147 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X566 VPWR.t130 dr[6].t0 a_1066_18226# VPWR.t17 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X567 g[5].t1 a_490_11424# VGND.t358 VGND.t357 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X568 VGND.t533 VPWR.t465 VGND.t533 VGND.t479 sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
X569 VPWR.t172 VGND.t685 VPWR.t171 VPWR.t70 sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
X570 VPWR.t164 VGND.t686 VPWR.t164 VPWR.t91 sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
X571 VPWR.t169 VGND.t687 VPWR.t169 VPWR.t0 sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
X572 VPWR.t168 VGND.t688 VPWR.t168 VPWR.t70 sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
X573 g[0].t0 a_1066_15202# VGND.t101 VGND.t100 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.2516p ps=2.16u w=0.74u l=0.13u
X574 VPWR.t355 a_1066_5376# b[3].t5 VPWR.t61 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X575 VGND.t525 VPWR.t462 VGND.t524 VGND.t199 sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
X576 VGND.t466 db[2].t0 a_490_6130# VGND.t465 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X577 VPWR.t20 a_1066_18226# r[6].t6 VPWR.t17 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X578 VPWR.t417 a_490_13690# g[2].t6 VPWR.t52 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X579 b[3].t4 a_1066_5376# VPWR.t354 VPWR.t61 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3864p ps=2.93u w=1.12u l=0.13u
X580 VPWR.t370 dg[3].t0 a_1066_12936# VPWR.t180 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X581 VPWR.t167 VGND.t689 VPWR.t166 VPWR.t140 sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
X582 VGND.t409 VPWR.t494 VGND.t409 VGND.t286 sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
X583 VPWR.t328 a_1066_12936# g[3].t6 VPWR.t180 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X584 VGND.t116 a_490_22762# r[0].t1 VGND.t115 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X585 VPWR.t18 a_1066_18226# r[6].t5 VPWR.t17 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X586 g[1].t1 a_490_14448# VGND.t77 VGND.t76 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.2516p ps=2.16u w=0.74u l=0.13u
X587 VGND.t135 VPWR.t480 VGND.t135 VGND.t134 sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
X588 VGND.t14 dg[6].t0 a_490_10666# VGND.t15 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X589 VPWR.t362 a_490_3864# b[5].t5 VPWR.t123 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X590 VGND.t52 a_490_6130# b[2].t1 VGND.t51 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X591 VPWR.t10 dg[6].t0 a_490_10666# VPWR.t9 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X592 VPWR.t326 a_1066_12936# g[3].t5 VPWR.t180 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X593 VPWR.t165 VGND.t690 VPWR.t164 VPWR.t91 sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
X594 VPWR.t163 VGND.t691 VPWR.t162 VPWR.t61 sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
X595 VGND.t190 VPWR.t469 VGND.t190 VGND.t189 sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
X596 VPWR.t341 a_490_11424# g[5].t5 VPWR.t9 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X597 VGND.t412 VPWR.t495 VGND.t412 VGND.t251 sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
X598 VGND.t563 a_490_13690# g[2].t1 VGND.t562 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X599 g[3].t1 a_1066_12936# VGND.t338 VGND.t337 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X600 r[3].t5 a_1066_20496# VPWR.t3 VPWR.t0 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X601 VGND.t194 VPWR.t470 VGND.t194 VGND.t193 sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
X602 r[5].t1 a_490_18984# VGND.t234 VGND.t233 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X603 a_490_17472# dr[7].t0 VGND.t327 VGND.t596 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X604 a_490_2352# db[7].t0 VGND.t202 VGND.t201 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X605 VGND.t507 a_1066_12178# g[4].t1 VGND.t546 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X606 VGND.t416 VPWR.t496 VGND.t416 VGND.t418 sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
X607 VGND.t545 a_1066_12178# g[4].t0 VGND.t544 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X608 VGND.t179 VPWR.t466 VGND.t178 VGND.t177 sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
X609 a_1066_15202# dg[0].t0 VPWR.t74 VPWR.t70 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X610 VPWR.t161 VGND.t692 VPWR.t160 VPWR.t155 sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
X611 VPWR.t95 dg[1].t0 a_490_14448# VPWR.t52 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X612 VGND.t297 a_1066_3106# b[6].t1 VGND.t296 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X613 VGND.t132 VPWR.t479 VGND.t131 VGND.t130 sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
X614 b[6].t0 a_1066_3106# VGND.t295 VGND.t294 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.2516p ps=2.16u w=0.74u l=0.13u
X615 g[0].t5 a_1066_15202# VPWR.t72 VPWR.t70 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X616 VPWR.t304 a_1066_3106# b[6].t6 VPWR.t123 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X617 VPWR.t159 VGND.t693 VPWR.t158 VPWR.t140 sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
X618 VGND.t413 VPWR.t495 VGND.t412 VGND.t248 sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
X619 VGND.t50 a_490_6130# b[2].t0 VGND.t49 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X620 r[0].t5 a_490_22762# VPWR.t81 VPWR.t79 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X621 b[6].t5 a_1066_3106# VPWR.t303 VPWR.t123 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X622 b[0].t1 a_490_7642# VGND.t39 VGND.t38 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X623 a_1066_20496# dr[3].t0 VGND.t6 VGND.t18 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X624 VPWR.t319 a_490_17472# r[7].t5 VPWR.t147 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X625 g[0].t4 a_1066_15202# VPWR.t71 VPWR.t70 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3864p ps=2.93u w=1.12u l=0.13u
X626 VPWR.t302 a_1066_3106# b[6].t4 VPWR.t123 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X627 VPWR.t376 db[2].t0 a_490_6130# VPWR.t35 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X628 r[3].t1 a_1066_20496# VGND.t3 VGND.t2 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X629 VGND.t351 dg[5].t0 a_490_11424# VGND.t352 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X630 r[1].t0 a_586_22008# VGND.t495 VGND.t494 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X631 r[6].t4 a_1066_18226# VPWR.t18 VPWR.t17 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X632 g[2].t5 a_490_13690# VPWR.t416 VPWR.t52 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3864p ps=2.93u w=1.12u l=0.13u
X633 b[7].t1 a_490_2352# VGND.t576 VGND.t575 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X634 a_490_10666# dg[6].t0 VGND.t14 VGND.t13 sg13_lv_nmos ad=0.2553p pd=2.17u as=0.1406p ps=1.12u w=0.74u l=0.13u
X635 VPWR.t157 VGND.t694 VPWR.t156 VPWR.t155 sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
X636 r[3].t0 a_1066_20496# VGND.t1 VGND.t0 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.2516p ps=2.16u w=0.74u l=0.13u
X637 a_490_10666# dg[6].t0 VPWR.t10 VPWR.t9 sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
X638 g[3].t4 a_1066_12936# VPWR.t326 VPWR.t180 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X639 r[1].t1 a_586_22008# VGND.t493 VGND.t492 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.2516p ps=2.16u w=0.74u l=0.13u
X640 VGND.t92 a_1066_4618# b[4].t2 VGND.t91 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X641 g[6].t0 a_490_10666# VGND.t63 VGND.t62 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X642 a_490_22762# dr[0].t0 VGND.t120 VGND.t536 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X643 VGND.t75 a_490_14448# g[1].t0 VGND.t74 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X644 VGND.t420 VPWR.t497 VGND.t420 VGND.t422 sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
X645 VPWR.t37 a_490_6130# b[2].t5 VPWR.t35 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X646 b[4].t1 a_1066_4618# VGND.t90 VGND.t89 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X647 a_1066_21250# dr[2].t0 VGND.t19 VGND.t18 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X648 b[7].t0 a_490_2352# VGND.t574 VGND.t573 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.2516p ps=2.16u w=0.74u l=0.13u
X649 g[6].t4 a_490_10666# VPWR.t44 VPWR.t9 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X650 VGND.t336 a_1066_12936# g[3].t1 VGND.t335 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X651 VGND.t88 a_1066_4618# b[4].t0 VGND.t87 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X652 VPWR.t2 a_1066_20496# r[3].t5 VPWR.t0 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X653 VGND.t407 VPWR.t493 VGND.t406 VGND.t405 sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
X654 VPWR.t154 VGND.t695 VPWR.t153 VPWR.t140 sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
X655 a_1066_4618# db[4].t0 VPWR.t65 VPWR.t61 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X656 g[7].t1 a_1066_9912# VGND.t223 VGND.t222 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X657 VGND.t170 VPWR.t476 VGND.t170 VGND.t133 sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
X658 b[0].t0 a_490_7642# VGND.t37 VGND.t36 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X659 r[2].t1 a_1066_21250# VGND.t211 VGND.t2 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X660 VGND.t334 a_1066_12936# g[3].t0 VGND.t333 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X661 VPWR.t62 a_1066_4618# b[4].t4 VPWR.t61 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X662 VPWR.t152 VGND.t696 VPWR.t152 VPWR.t140 sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
X663 VPWR.t1 a_1066_20496# r[3].t4 VPWR.t0 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X664 a_490_11424# dg[5].t0 VPWR.t337 VPWR.t9 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X665 VPWR.t379 a_586_22008# r[1].t4 VPWR.t13 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X666 VGND.t232 a_490_18984# r[5].t0 VGND.t231 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X667 VGND.t321 a_490_17472# r[7].t0 VGND.t320 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X668 r[2].t0 a_1066_21250# VGND.t210 VGND.t0 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.2516p ps=2.16u w=0.74u l=0.13u
X669 a_490_14448# dg[1].t0 VPWR.t95 VPWR.t52 sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
X670 VGND.t410 VPWR.t494 VGND.t409 VGND.t283 sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
X671 a_1066_12178# dg[4].t0 VPWR.t387 VPWR.t180 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X672 g[1].t4 a_490_14448# VPWR.t53 VPWR.t52 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X673 VGND.t277 VPWR.t486 VGND.t276 VGND.t275 sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
X674 VGND.t280 VPWR.t487 VGND.t280 VGND.t279 sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
X675 g[4].t5 a_1066_12178# VPWR.t405 VPWR.t180 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X676 VPWR.t36 a_490_6130# b[2].t4 VPWR.t35 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X677 r[4].t5 a_490_19738# VPWR.t391 VPWR.t0 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X678 a_490_2352# db[7].t0 VPWR.t92 VPWR.t91 sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
X679 b[0].t5 a_490_7642# VPWR.t28 VPWR.t26 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X680 VPWR.t80 a_490_22762# r[0].t4 VPWR.t79 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X681 g[4].t4 a_1066_12178# VPWR.t404 VPWR.t180 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3864p ps=2.93u w=1.12u l=0.13u
X682 a_1066_3106# db[6].t0 VPWR.t334 VPWR.t123 sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
X683 VPWR.t94 a_490_2352# b[7].t5 VPWR.t91 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X684 a_490_11424# dg[5].t0 VGND.t351 VGND.t350 sg13_lv_nmos ad=0.2553p pd=2.17u as=0.1406p ps=1.12u w=0.74u l=0.13u
X685 r[5].t5 a_490_18984# VPWR.t116 VPWR.t17 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X686 a_490_17472# dr[7].t0 VPWR.t321 VPWR.t147 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X687 VGND.t417 VPWR.t496 VGND.t416 VGND.t415 sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
X688 VGND.t370 a_1066_5376# b[3].t2 VGND.t397 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X689 g[5].t0 a_490_11424# VGND.t356 VGND.t355 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X690 VGND.t127 VPWR.t478 VGND.t127 VGND.t126 sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
X691 VPWR.t415 a_490_13690# g[2].t4 VPWR.t52 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X692 b[3].t1 a_1066_5376# VGND.t396 VGND.t395 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X693 a_778_6888# db[1].t0 VGND.t314 VGND.t389 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X694 VGND.t394 a_1066_5376# b[3].t0 VGND.t393 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X695 VPWR.t151 VGND.t697 VPWR.t150 VPWR.t140 sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
X696 VPWR.t149 VGND.t698 VPWR.t149 VPWR.t147 sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
X697 VPWR.t148 VGND.t699 VPWR.t148 VPWR.t147 sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
X698 VGND.t310 a_778_6888# b[1].t1 VGND.t309 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X699 VPWR.t146 VGND.t700 VPWR.t146 VPWR.t106 sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
X700 r[4].t0 a_490_19738# VGND.t508 VGND.t241 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X701 VGND.t428 VPWR.t449 VGND.t428 VGND.t427 sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
X702 VGND.t114 a_490_22762# r[0].t0 VGND.t113 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X703 a_1066_21250# dr[2].t0 VPWR.t14 VPWR.t13 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X704 VGND.t221 a_1066_9912# g[7].t1 VGND.t220 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X705 a_1066_4618# db[4].t0 VGND.t462 VGND.t461 sg13_lv_nmos ad=0.2553p pd=2.17u as=0.1406p ps=1.12u w=0.74u l=0.13u
X706 VPWR.t145 VGND.t701 VPWR.t144 VPWR.t79 sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
X707 b[0].t4 a_490_7642# VPWR.t27 VPWR.t26 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X708 VPWR.t401 dg[7].t0 a_1066_9912# VPWR.t106 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X709 r[2].t5 a_1066_21250# VPWR.t99 VPWR.t13 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X710 VPWR.t143 VGND.t702 VPWR.t143 VPWR.t70 sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
X711 VGND.t219 a_1066_9912# g[7].t0 VGND.t218 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X712 VPWR.t423 a_490_2352# b[7].t4 VPWR.t91 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X713 g[7].t5 a_1066_9912# VPWR.t108 VPWR.t106 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X714 VPWR.t340 a_490_11424# g[5].t4 VPWR.t9 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X715 r[2].t4 a_1066_21250# VPWR.t98 VPWR.t13 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3864p ps=2.93u w=1.12u l=0.13u
X716 VPWR.t138 VGND.t703 VPWR.t138 VPWR.t106 sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
X717 a_490_18984# dr[5].t0 VGND.t151 VGND.t150 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X718 a_490_3864# db[5].t0 VGND.t244 VGND.t243 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X719 a_586_22008# dr[1].t0 VPWR.t412 VPWR.t13 sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
X720 VGND.t438 VPWR.t452 VGND.t438 VGND.t259 sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
X721 g[7].t4 a_1066_9912# VPWR.t107 VPWR.t106 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X722 VGND.t253 VPWR.t490 VGND.t253 VGND.t252 sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
X723 VGND.t269 VPWR.t484 VGND.t269 VGND.t268 sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
X724 VPWR.t141 VGND.t704 VPWR.t141 VPWR.t140 sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
X725 VPWR.t390 a_490_19738# r[4].t4 VPWR.t0 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X726 VGND.t442 VPWR.t453 VGND.t442 VGND.t441 sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
X727 a_1066_18226# dr[6].t0 VPWR.t130 VPWR.t17 sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
X728 VGND.t421 VPWR.t497 VGND.t420 VGND.t419 sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
X729 VGND.t491 a_586_22008# r[1].t0 VGND.t490 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X730 a_778_6888# db[1].t0 VPWR.t312 VPWR.t35 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X731 VGND.t308 a_778_6888# b[1].t0 VGND.t307 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X732 g[2].t0 a_490_13690# VGND.t561 VGND.t560 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1406p ps=1.12u w=0.74u l=0.13u
X733 a_490_22762# dr[0].t0 VPWR.t82 VPWR.t79 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X734 VPWR.t139 VGND.t705 VPWR.t138 VPWR.t106 sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
X735 a_1066_12936# dg[3].t0 VPWR.t370 VPWR.t180 sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
X736 VPWR.t137 VGND.t706 VPWR.t136 VPWR.t52 sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
X737 VPWR.t310 a_778_6888# b[1].t4 VPWR.t35 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X738 VPWR.t115 a_490_18984# r[5].t4 VPWR.t17 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X739 VPWR.t318 a_490_17472# r[7].t4 VPWR.t147 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X740 VGND.t144 VPWR.t482 VGND.t143 VGND.t142 sg13_lv_nmos ad=0.1428p pd=1.52u as=0 ps=0 w=0.42u l=1u
X741 VGND.t383 VPWR.t446 VGND.t383 VGND.t263 sg13_lv_nmos ad=79.8f pd=0.8u as=0 ps=0 w=0.42u l=1u
R0 VGND.n448 VGND.n364 11762.3
R1 VGND.n994 VGND.n993 11746.1
R2 VGND.n384 VGND.n319 11464.4
R3 VGND.n956 VGND.n955 11464.4
R4 VGND.n449 VGND.n448 10150
R5 VGND.n449 VGND.n310 10150
R6 VGND.n546 VGND.n310 10150
R7 VGND.n547 VGND.n546 10150
R8 VGND.n547 VGND.n210 10150
R9 VGND.n626 VGND.n210 10150
R10 VGND.n627 VGND.n626 10150
R11 VGND.n627 VGND.n112 10150
R12 VGND.n729 VGND.n112 10150
R13 VGND.n730 VGND.n729 10150
R14 VGND.n730 VGND.n24 10150
R15 VGND.n869 VGND.n24 10150
R16 VGND.n870 VGND.n869 10150
R17 VGND.n870 VGND.n17 10150
R18 VGND.n994 VGND.n17 10150
R19 VGND.n467 VGND.n319 9822.58
R20 VGND.n468 VGND.n467 9822.58
R21 VGND.n468 VGND.n263 9822.58
R22 VGND.n566 VGND.n263 9822.58
R23 VGND.n567 VGND.n566 9822.58
R24 VGND.n567 VGND.n163 9822.58
R25 VGND.n646 VGND.n163 9822.58
R26 VGND.n647 VGND.n646 9822.58
R27 VGND.n647 VGND.n75 9822.58
R28 VGND.n738 VGND.n75 9822.58
R29 VGND.n739 VGND.n738 9822.58
R30 VGND.n739 VGND.n22 9822.58
R31 VGND.n889 VGND.n22 9822.58
R32 VGND.n954 VGND.n889 9822.58
R33 VGND.n955 VGND.n954 9822.58
R34 VGND.n365 VGND.n319 958.561
R35 VGND.n467 VGND.n466 958.561
R36 VGND.n469 VGND.n468 958.561
R37 VGND.n311 VGND.n263 958.561
R38 VGND.n566 VGND.n565 958.561
R39 VGND.n568 VGND.n567 958.561
R40 VGND.n211 VGND.n163 958.561
R41 VGND.n646 VGND.n645 958.561
R42 VGND.n648 VGND.n647 958.561
R43 VGND.n113 VGND.n75 958.561
R44 VGND.n738 VGND.n737 958.561
R45 VGND.n740 VGND.n739 958.561
R46 VGND.n25 VGND.n22 958.561
R47 VGND.n889 VGND.n888 958.561
R48 VGND.n954 VGND.n953 958.561
R49 VGND.n955 VGND.n7 958.561
R50 VGND.n448 VGND.n447 941.418
R51 VGND.n450 VGND.n449 941.418
R52 VGND.n491 VGND.n310 941.418
R53 VGND.n546 VGND.n545 941.418
R54 VGND.n548 VGND.n547 941.418
R55 VGND.n578 VGND.n210 941.418
R56 VGND.n626 VGND.n625 941.418
R57 VGND.n628 VGND.n627 941.418
R58 VGND.n680 VGND.n112 941.418
R59 VGND.n729 VGND.n728 941.418
R60 VGND.n731 VGND.n730 941.418
R61 VGND.n763 VGND.n24 941.418
R62 VGND.n869 VGND.n868 941.418
R63 VGND.n871 VGND.n870 941.418
R64 VGND.n936 VGND.n17 941.418
R65 VGND.n995 VGND.n994 941.418
R66 VGND.n971 VGND.n970 725.962
R67 VGND.n993 VGND.n18 709.361
R68 VGND.n387 VGND.t128 423.017
R69 VGND.t518 VGND.n371 423.017
R70 VGND.n977 VGND.t425 423.017
R71 VGND.t177 VGND.n364 422.627
R72 VGND.n977 VGND.t427 408.238
R73 VGND.n387 VGND.t516 408.238
R74 VGND.t180 VGND.n371 408.238
R75 VGND.n970 VGND.t418 408.229
R76 VGND.t126 VGND.n384 407.849
R77 VGND.t423 VGND.n956 407.849
R78 VGND.t494 VGND.n455 407.144
R79 VGND.t2 VGND.n477 407.144
R80 VGND.t233 VGND.n522 407.144
R81 VGND.t324 VGND.n552 407.144
R82 VGND.t86 VGND.n232 407.144
R83 VGND.t560 VGND.n632 407.144
R84 VGND.t361 VGND.n670 407.144
R85 VGND.t68 VGND.n134 407.144
R86 VGND.t55 VGND.n46 407.144
R87 VGND.t456 VGND.n875 407.144
R88 VGND.t575 VGND.n940 407.144
R89 VGND.n971 VGND.t429 406.404
R90 VGND.t415 VGND.n18 406.404
R91 VGND.n457 VGND.t113 390
R92 VGND.n503 VGND.t12 390
R93 VGND.n534 VGND.t242 390
R94 VGND.n560 VGND.t35 390
R95 VGND.n614 VGND.t112 390
R96 VGND.n640 VGND.t342 390
R97 VGND.n696 VGND.t552 390
R98 VGND.n717 VGND.t227 390
R99 VGND.n857 VGND.t404 390
R100 VGND.n883 VGND.t99 390
R101 VGND.n948 VGND.t302 390
R102 VGND.t498 VGND.n454 381.43
R103 VGND.n501 VGND.t4 381.43
R104 VGND.n532 VGND.t238 381.43
R105 VGND.n458 VGND.t124 364.286
R106 VGND.t7 VGND.n475 364.286
R107 VGND.t239 VGND.n517 364.286
R108 VGND.n561 VGND.t30 364.286
R109 VGND.t107 VGND.n215 364.286
R110 VGND.n641 VGND.t337 364.286
R111 VGND.t547 VGND.n652 364.286
R112 VGND.t222 VGND.n117 364.286
R113 VGND.t402 VGND.n29 364.286
R114 VGND.n884 VGND.t97 364.286
R115 VGND.n949 VGND.t300 364.286
R116 VGND.t38 VGND.t311 360
R117 VGND.t317 VGND.t41 360
R118 VGND.t500 VGND.n453 355.714
R119 VGND.t9 VGND.n480 355.714
R120 VGND.t241 VGND.n525 355.714
R121 VGND.t332 VGND.n550 355.714
R122 VGND.t82 VGND.n234 355.714
R123 VGND.t569 VGND.n630 355.714
R124 VGND.t357 VGND.n672 355.714
R125 VGND.t64 VGND.n136 355.714
R126 VGND.n775 VGND.t319 355.714
R127 VGND.t36 VGND.n756 355.714
R128 VGND.t60 VGND.n48 355.714
R129 VGND.t448 VGND.n873 355.714
R130 VGND.t579 VGND.n938 355.714
R131 VGND.n459 VGND.t119 338.572
R132 VGND.n504 VGND.t5 338.572
R133 VGND.n535 VGND.t235 338.572
R134 VGND.n783 VGND.t47 338.572
R135 VGND.n385 VGND.t126 334.339
R136 VGND.t516 VGND.n374 334.339
R137 VGND.n403 VGND.t180 334.339
R138 VGND.n964 VGND.t423 334.337
R139 VGND.t427 VGND.n967 334.337
R140 VGND.t418 VGND.n969 334.337
R141 VGND.t502 VGND.n452 330
R142 VGND.n500 VGND.t11 330
R143 VGND.n531 VGND.t231 330
R144 VGND.t322 VGND.n549 330
R145 VGND.n242 VGND.t85 330
R146 VGND.t572 VGND.n629 330
R147 VGND.n681 VGND.t360 330
R148 VGND.n144 VGND.t67 330
R149 VGND.t307 VGND.n754 330
R150 VGND.n767 VGND.t40 330
R151 VGND.n56 VGND.t49 330
R152 VGND.t452 VGND.n872 330
R153 VGND.t583 VGND.n937 330
R154 VGND.t0 VGND.n483 320.613
R155 VGND.t121 VGND.n450 319.99
R156 VGND.n545 VGND.t236 319.99
R157 VGND.n969 VGND.t415 319.56
R158 VGND.t429 VGND.n967 319.56
R159 VGND.t425 VGND.n964 319.56
R160 VGND.t128 VGND.n385 319.558
R161 VGND.n374 VGND.t518 319.558
R162 VGND.n403 VGND.t177 319.558
R163 VGND.n460 VGND.t536 312.858
R164 VGND.t18 VGND.n471 312.858
R165 VGND.t150 VGND.n514 312.858
R166 VGND.n563 VGND.t287 312.858
R167 VGND.t588 VGND.n213 312.858
R168 VGND.n643 VGND.t460 312.858
R169 VGND.t506 VGND.n650 312.858
R170 VGND.t543 VGND.n115 312.858
R171 VGND.n788 VGND.t389 312.858
R172 VGND.t266 VGND.n748 312.858
R173 VGND.t369 VGND.n27 312.858
R174 VGND.n886 VGND.t464 312.858
R175 VGND.n951 VGND.t348 312.858
R176 VGND.t492 VGND.n451 304.286
R177 VGND.n771 VGND.t315 304.286
R178 VGND.n461 VGND.t539 287.144
R179 VGND.n505 VGND.t22 287.144
R180 VGND.n536 VGND.t154 287.144
R181 VGND.n564 VGND.t290 287.144
R182 VGND.n618 VGND.t591 287.144
R183 VGND.n644 VGND.t459 287.144
R184 VGND.n700 VGND.t505 287.144
R185 VGND.n721 VGND.t542 287.144
R186 VGND.t392 VGND.n743 287.144
R187 VGND.n787 VGND.t264 287.144
R188 VGND.n861 VGND.t367 287.144
R189 VGND.n887 VGND.t463 287.144
R190 VGND.n952 VGND.t346 287.144
R191 VGND.t25 VGND.t599 282.858
R192 VGND.t27 VGND.t596 282.858
R193 VGND.t32 VGND.t326 282.858
R194 VGND.t34 VGND.t331 282.858
R195 VGND.t23 VGND.t320 282.858
R196 VGND.t102 VGND.t208 282.858
R197 VGND.t209 VGND.t104 282.858
R198 VGND.t109 VGND.t74 282.858
R199 VGND.t80 VGND.t111 282.858
R200 VGND.t100 VGND.t84 282.858
R201 VGND.t345 VGND.t594 282.858
R202 VGND.t333 VGND.t595 282.858
R203 VGND.t339 VGND.t562 282.858
R204 VGND.t341 VGND.t567 282.858
R205 VGND.t343 VGND.t571 282.858
R206 VGND.t555 VGND.t352 282.858
R207 VGND.t353 VGND.t544 282.858
R208 VGND.t549 VGND.t363 282.858
R209 VGND.t355 VGND.t551 282.858
R210 VGND.t553 VGND.t359 282.858
R211 VGND.t230 VGND.t15 282.858
R212 VGND.t16 VGND.t218 282.858
R213 VGND.t224 VGND.t70 282.858
R214 VGND.t62 VGND.t226 282.858
R215 VGND.t228 VGND.t66 282.858
R216 VGND.t395 VGND.t465 282.858
R217 VGND.t467 VGND.t400 282.858
R218 VGND.t401 VGND.t58 282.858
R219 VGND.t61 VGND.t393 282.858
R220 VGND.t398 VGND.t51 282.858
R221 VGND.t89 VGND.t247 282.858
R222 VGND.t95 VGND.t243 282.858
R223 VGND.t96 VGND.t447 282.858
R224 VGND.t87 VGND.t450 282.858
R225 VGND.t93 VGND.t453 282.858
R226 VGND.t304 VGND.t205 282.858
R227 VGND.t296 VGND.t201 282.858
R228 VGND.t298 VGND.t578 282.858
R229 VGND.t303 VGND.t581 282.858
R230 VGND.t294 VGND.t584 282.858
R231 VGND.t152 VGND.n314 277.755
R232 VGND.n463 VGND.t556 277.132
R233 VGND.t20 VGND.n469 277.132
R234 VGND.n462 VGND.t537 261.43
R235 VGND.n559 VGND.t597 261.43
R236 VGND.t206 VGND.n219 261.43
R237 VGND.n639 VGND.t592 261.43
R238 VGND.t350 VGND.n656 261.43
R239 VGND.t13 VGND.n121 261.43
R240 VGND.t267 VGND.n746 261.43
R241 VGND.t468 VGND.n33 261.43
R242 VGND.n882 VGND.t245 261.43
R243 VGND.n947 VGND.t203 261.43
R244 VGND.t476 VGND.n438 252.065
R245 VGND.n415 VGND.t142 252.065
R246 VGND.t130 VGND.n595 252.065
R247 VGND.n572 VGND.t379 252.065
R248 VGND.t260 VGND.n735 252.065
R249 VGND.t256 VGND.n733 252.065
R250 VGND.t248 VGND.n1012 252.065
R251 VGND.n11 VGND.t283 252.065
R252 VGND.t195 VGND.n314 252.041
R253 VGND.n447 VGND.t377 251.417
R254 VGND.t185 VGND.n463 251.417
R255 VGND.t164 VGND.n491 251.417
R256 VGND.t485 VGND.n548 251.417
R257 VGND.t199 VGND.n578 251.417
R258 VGND.n625 VGND.t281 251.417
R259 VGND.t136 VGND.n628 251.417
R260 VGND.t254 VGND.n680 251.417
R261 VGND.n728 VGND.t520 251.417
R262 VGND.t166 VGND.n731 251.417
R263 VGND.n868 VGND.t173 251.417
R264 VGND.t405 VGND.n871 251.417
R265 VGND.t443 VGND.n936 251.417
R266 VGND.t419 VGND.n995 251.417
R267 VGND.n438 VGND.t145 243.494
R268 VGND.t375 VGND.n415 243.494
R269 VGND.n595 VGND.t382 243.494
R270 VGND.t197 VGND.n572 243.494
R271 VGND.n735 VGND.t259 243.494
R272 VGND.n733 VGND.t169 243.494
R273 VGND.n1012 VGND.t286 243.494
R274 VGND.t422 VGND.n11 243.494
R275 VGND.t162 VGND.n483 243.47
R276 VGND.t479 VGND.n365 242.846
R277 VGND.n466 VGND.t188 242.846
R278 VGND.t193 VGND.n311 242.846
R279 VGND.n565 VGND.t268 242.846
R280 VGND.t133 VGND.n568 242.846
R281 VGND.t434 VGND.n211 242.846
R282 VGND.n645 VGND.t278 242.846
R283 VGND.t472 VGND.n648 242.846
R284 VGND.t189 VGND.n113 242.846
R285 VGND.n737 VGND.t263 242.846
R286 VGND.t158 VGND.n25 242.846
R287 VGND.n888 VGND.t184 242.846
R288 VGND.n953 VGND.t149 242.846
R289 VGND.t251 VGND.n7 242.846
R290 VGND.n465 VGND.t530 221.417
R291 VGND.t527 VGND.n740 221.417
R292 VGND.t272 VGND.n763 221.417
R293 VGND.t530 VGND.n464 205.714
R294 VGND.n441 VGND.t479 200.613
R295 VGND.t145 VGND.n413 200.613
R296 VGND.n423 VGND.t375 200.613
R297 VGND.n494 VGND.t162 200.613
R298 VGND.n539 VGND.t193 200.613
R299 VGND.n598 VGND.t133 200.613
R300 VGND.t382 VGND.n570 200.613
R301 VGND.n581 VGND.t197 200.613
R302 VGND.t263 VGND.n736 200.613
R303 VGND.t259 VGND.n734 200.613
R304 VGND.t169 VGND.n732 200.613
R305 VGND.n796 VGND.t141 200.613
R306 VGND.n1015 VGND.t251 200.613
R307 VGND.t286 VGND.n9 200.613
R308 VGND.n998 VGND.t422 200.613
R309 VGND.t188 VGND.n465 199.989
R310 VGND.t330 VGND.t483 197.143
R311 VGND.t279 VGND.t78 197.143
R312 VGND.t566 VGND.t134 197.143
R313 VGND.t252 VGND.t366 197.143
R314 VGND.t523 VGND.t73 197.143
R315 VGND.t176 VGND.t57 197.143
R316 VGND.t445 VGND.t408 197.143
R317 VGND.t577 VGND.t441 197.143
R318 VGND.n423 VGND.t377 192.042
R319 VGND.t142 VGND.n413 192.042
R320 VGND.n441 VGND.t476 192.042
R321 VGND.n494 VGND.t164 192.042
R322 VGND.n539 VGND.t195 192.042
R323 VGND.n581 VGND.t199 192.042
R324 VGND.t379 VGND.n570 192.042
R325 VGND.n598 VGND.t130 192.042
R326 VGND.n732 VGND.t166 192.042
R327 VGND.n734 VGND.t256 192.042
R328 VGND.n736 VGND.t260 192.042
R329 VGND.n796 VGND.t138 192.042
R330 VGND.n998 VGND.t419 192.042
R331 VGND.t283 VGND.n9 192.042
R332 VGND.n1015 VGND.t248 192.042
R333 VGND.t483 VGND.n551 184.286
R334 VGND.n245 VGND.t279 184.286
R335 VGND.t134 VGND.n631 184.286
R336 VGND.n684 VGND.t252 184.286
R337 VGND.n147 VGND.t523 184.286
R338 VGND.n59 VGND.t176 184.286
R339 VGND.t408 VGND.n874 184.286
R340 VGND.t441 VGND.n939 184.286
R341 VGND.n464 VGND.t185 175.714
R342 VGND.n562 VGND.t270 175.714
R343 VGND.n615 VGND.t431 175.714
R344 VGND.n642 VGND.t275 175.714
R345 VGND.n697 VGND.t474 175.714
R346 VGND.n718 VGND.t191 175.714
R347 VGND.n858 VGND.t155 175.714
R348 VGND.n885 VGND.t181 175.714
R349 VGND.n950 VGND.t146 175.714
R350 VGND.t270 VGND.t28 162.857
R351 VGND.t431 VGND.t105 162.857
R352 VGND.t275 VGND.t335 162.857
R353 VGND.t474 VGND.t546 162.857
R354 VGND.t191 VGND.t220 162.857
R355 VGND.t155 VGND.t397 162.857
R356 VGND.t181 VGND.t91 162.857
R357 VGND.t146 VGND.t305 162.857
R358 VGND.t556 VGND.n462 150
R359 VGND.n505 VGND.t20 150
R360 VGND.n536 VGND.t152 150
R361 VGND.t288 VGND.n564 150
R362 VGND.t597 VGND.n558 150
R363 VGND.n618 VGND.t589 150
R364 VGND.n256 VGND.t206 150
R365 VGND.t457 VGND.n644 150
R366 VGND.t592 VGND.n638 150
R367 VGND.n700 VGND.t503 150
R368 VGND.n695 VGND.t350 150
R369 VGND.n721 VGND.t540 150
R370 VGND.n158 VGND.t13 150
R371 VGND.t390 VGND.n743 150
R372 VGND.n861 VGND.t371 150
R373 VGND.n70 VGND.t468 150
R374 VGND.t461 VGND.n887 150
R375 VGND.t245 VGND.n881 150
R376 VGND.t349 VGND.n952 150
R377 VGND.t203 VGND.n946 150
R378 VGND.t558 VGND.n461 124.287
R379 VGND.t22 VGND.n471 124.287
R380 VGND.t154 VGND.n514 124.287
R381 VGND.t290 VGND.n563 124.287
R382 VGND.t599 VGND.n557 124.287
R383 VGND.t591 VGND.n213 124.287
R384 VGND.t208 VGND.n221 124.287
R385 VGND.t459 VGND.n643 124.287
R386 VGND.t594 VGND.n637 124.287
R387 VGND.t505 VGND.n650 124.287
R388 VGND.t352 VGND.n659 124.287
R389 VGND.t542 VGND.n115 124.287
R390 VGND.t15 VGND.n123 124.287
R391 VGND.n788 VGND.t392 124.287
R392 VGND.t367 VGND.n27 124.287
R393 VGND.t465 VGND.n35 124.287
R394 VGND.t463 VGND.n886 124.287
R395 VGND.t247 VGND.n880 124.287
R396 VGND.t346 VGND.n951 124.287
R397 VGND.t205 VGND.n945 124.287
R398 VGND.n451 VGND.t121 107.144
R399 VGND.n500 VGND.t0 107.144
R400 VGND.n531 VGND.t236 107.144
R401 VGND.n554 VGND.t23 107.144
R402 VGND.n549 VGND.t328 107.144
R403 VGND.n254 VGND.t100 107.144
R404 VGND.n242 VGND.t76 107.144
R405 VGND.n634 VGND.t343 107.144
R406 VGND.n629 VGND.t564 107.144
R407 VGND.n693 VGND.t553 107.144
R408 VGND.n681 VGND.t364 107.144
R409 VGND.n156 VGND.t228 107.144
R410 VGND.n144 VGND.t71 107.144
R411 VGND.n767 VGND.t42 107.144
R412 VGND.n68 VGND.t398 107.144
R413 VGND.n56 VGND.t53 107.144
R414 VGND.n877 VGND.t93 107.144
R415 VGND.n872 VGND.t454 107.144
R416 VGND.n942 VGND.t294 107.144
R417 VGND.n937 VGND.t573 107.144
R418 VGND.t559 VGND.n460 98.5719
R419 VGND.n504 VGND.t18 98.5719
R420 VGND.n535 VGND.t150 98.5719
R421 VGND.t287 VGND.n562 98.5719
R422 VGND.t596 VGND.n556 98.5719
R423 VGND.n615 VGND.t588 98.5719
R424 VGND.n255 VGND.t209 98.5719
R425 VGND.t460 VGND.n642 98.5719
R426 VGND.t595 VGND.n636 98.5719
R427 VGND.n697 VGND.t506 98.5719
R428 VGND.n694 VGND.t353 98.5719
R429 VGND.n718 VGND.t543 98.5719
R430 VGND.n157 VGND.t16 98.5719
R431 VGND.t389 VGND.n746 98.5719
R432 VGND.t42 VGND.t272 98.5719
R433 VGND.n858 VGND.t369 98.5719
R434 VGND.n69 VGND.t467 98.5719
R435 VGND.t464 VGND.n885 98.5719
R436 VGND.t243 VGND.n879 98.5719
R437 VGND.t348 VGND.n950 98.5719
R438 VGND.t201 VGND.n944 98.5719
R439 VGND.t138 VGND.t390 85.7148
R440 VGND.n452 VGND.t115 81.4291
R441 VGND.t11 VGND.n480 81.4291
R442 VGND.t231 VGND.n525 81.4291
R443 VGND.n555 VGND.t34 81.4291
R444 VGND.n550 VGND.t322 81.4291
R445 VGND.t111 VGND.n225 81.4291
R446 VGND.t85 VGND.n234 81.4291
R447 VGND.n635 VGND.t341 81.4291
R448 VGND.n630 VGND.t572 81.4291
R449 VGND.t551 VGND.n663 81.4291
R450 VGND.t360 VGND.n672 81.4291
R451 VGND.t226 VGND.n127 81.4291
R452 VGND.t67 VGND.n136 81.4291
R453 VGND.t40 VGND.n756 81.4291
R454 VGND.t393 VGND.n39 81.4291
R455 VGND.t49 VGND.n48 81.4291
R456 VGND.n878 VGND.t87 81.4291
R457 VGND.n873 VGND.t452 81.4291
R458 VGND.n943 VGND.t303 81.4291
R459 VGND.n938 VGND.t583 81.4291
R460 VGND.t313 VGND.t267 77.1434
R461 VGND.t264 VGND.t318 77.1434
R462 VGND.t309 VGND.t266 77.1434
R463 VGND.t44 VGND.t307 77.1434
R464 VGND.t315 VGND.t46 77.1434
R465 VGND.t496 VGND.n459 72.8576
R466 VGND.t5 VGND.n475 72.8576
R467 VGND.t235 VGND.n517 72.8576
R468 VGND.t28 VGND.n561 72.8576
R469 VGND.t326 VGND.n555 72.8576
R470 VGND.t105 VGND.n215 72.8576
R471 VGND.t74 VGND.n225 72.8576
R472 VGND.t335 VGND.n641 72.8576
R473 VGND.t562 VGND.n635 72.8576
R474 VGND.t546 VGND.n652 72.8576
R475 VGND.t363 VGND.n663 72.8576
R476 VGND.t220 VGND.n117 72.8576
R477 VGND.t70 VGND.n127 72.8576
R478 VGND.n787 VGND.t313 72.8576
R479 VGND.t47 VGND.n750 72.8576
R480 VGND.t397 VGND.n29 72.8576
R481 VGND.t58 VGND.n39 72.8576
R482 VGND.t91 VGND.n884 72.8576
R483 VGND.t447 VGND.n878 72.8576
R484 VGND.t305 VGND.n949 72.8576
R485 VGND.t578 VGND.n943 72.8576
R486 VGND.t328 VGND.t485 68.5719
R487 VGND.t76 VGND.t281 68.5719
R488 VGND.t564 VGND.t136 68.5719
R489 VGND.t364 VGND.t254 68.5719
R490 VGND.t71 VGND.t520 68.5719
R491 VGND.t53 VGND.t173 68.5719
R492 VGND.t454 VGND.t405 68.5719
R493 VGND.t573 VGND.t443 68.5719
R494 VGND.n453 VGND.t125 55.7148
R495 VGND.n501 VGND.t9 55.7148
R496 VGND.n532 VGND.t241 55.7148
R497 VGND.n556 VGND.t32 55.7148
R498 VGND.n551 VGND.t332 55.7148
R499 VGND.n255 VGND.t109 55.7148
R500 VGND.n245 VGND.t82 55.7148
R501 VGND.n636 VGND.t339 55.7148
R502 VGND.n631 VGND.t569 55.7148
R503 VGND.n694 VGND.t549 55.7148
R504 VGND.n684 VGND.t357 55.7148
R505 VGND.n157 VGND.t224 55.7148
R506 VGND.n147 VGND.t64 55.7148
R507 VGND.t319 VGND.n752 55.7148
R508 VGND.n771 VGND.t36 55.7148
R509 VGND.n69 VGND.t401 55.7148
R510 VGND.n59 VGND.t60 55.7148
R511 VGND.n879 VGND.t96 55.7148
R512 VGND.n874 VGND.t448 55.7148
R513 VGND.n944 VGND.t298 55.7148
R514 VGND.n939 VGND.t579 55.7148
R515 VGND.t499 VGND.n458 47.1434
R516 VGND.n503 VGND.t7 47.1434
R517 VGND.n534 VGND.t239 47.1434
R518 VGND.t30 VGND.n560 47.1434
R519 VGND.t331 VGND.n554 47.1434
R520 VGND.n614 VGND.t107 47.1434
R521 VGND.n254 VGND.t80 47.1434
R522 VGND.t337 VGND.n640 47.1434
R523 VGND.t567 VGND.n634 47.1434
R524 VGND.n696 VGND.t547 47.1434
R525 VGND.n693 VGND.t355 47.1434
R526 VGND.n717 VGND.t222 47.1434
R527 VGND.n156 VGND.t62 47.1434
R528 VGND.t318 VGND.n748 47.1434
R529 VGND.n779 VGND.t38 47.1434
R530 VGND.n857 VGND.t402 47.1434
R531 VGND.n68 VGND.t61 47.1434
R532 VGND.t97 VGND.n883 47.1434
R533 VGND.t450 VGND.n877 47.1434
R534 VGND.t300 VGND.n948 47.1434
R535 VGND.t581 VGND.n942 47.1434
R536 VGND.t12 VGND.n502 37.1319
R537 VGND.t242 VGND.n533 37.1319
R538 VGND.t320 VGND.n553 37.1319
R539 VGND.t84 VGND.n253 37.1319
R540 VGND.t571 VGND.n633 37.1319
R541 VGND.t359 VGND.n692 37.1319
R542 VGND.t66 VGND.n155 37.1319
R543 VGND.t51 VGND.n67 37.1319
R544 VGND.t453 VGND.n876 37.1319
R545 VGND.t584 VGND.n941 37.1319
R546 VGND.t268 VGND.t288 34.2862
R547 VGND.t589 VGND.t434 34.2862
R548 VGND.t278 VGND.t457 34.2862
R549 VGND.t503 VGND.t472 34.2862
R550 VGND.t540 VGND.t189 34.2862
R551 VGND.t371 VGND.t158 34.2862
R552 VGND.t184 VGND.t461 34.2862
R553 VGND.t149 VGND.t349 34.2862
R554 VGND.n454 VGND.t123 30.0005
R555 VGND.t4 VGND.n477 30.0005
R556 VGND.t238 VGND.n522 30.0005
R557 VGND.n557 VGND.t27 30.0005
R558 VGND.n552 VGND.t330 30.0005
R559 VGND.t104 VGND.n221 30.0005
R560 VGND.t78 VGND.n232 30.0005
R561 VGND.n637 VGND.t333 30.0005
R562 VGND.n632 VGND.t566 30.0005
R563 VGND.t544 VGND.n659 30.0005
R564 VGND.t366 VGND.n670 30.0005
R565 VGND.t218 VGND.n123 30.0005
R566 VGND.t73 VGND.n134 30.0005
R567 VGND.n779 VGND.t317 30.0005
R568 VGND.t46 VGND.n754 30.0005
R569 VGND.t400 VGND.n35 30.0005
R570 VGND.t57 VGND.n46 30.0005
R571 VGND.n880 VGND.t95 30.0005
R572 VGND.n875 VGND.t445 30.0005
R573 VGND.n945 VGND.t296 30.0005
R574 VGND.n940 VGND.t577 30.0005
R575 VGND.t537 VGND.t558 25.7148
R576 VGND.t539 VGND.t559 25.7148
R577 VGND.t536 VGND.t496 25.7148
R578 VGND.t119 VGND.t499 25.7148
R579 VGND.t124 VGND.t490 25.7148
R580 VGND.t117 VGND.t498 25.7148
R581 VGND.t123 VGND.t500 25.7148
R582 VGND.t125 VGND.t502 25.7148
R583 VGND.t115 VGND.t492 25.7148
R584 VGND.t490 VGND.n457 21.4291
R585 VGND.t113 VGND.n456 21.4291
R586 VGND.t35 VGND.n559 21.4291
R587 VGND.t112 VGND.n219 21.4291
R588 VGND.t342 VGND.n639 21.4291
R589 VGND.t552 VGND.n656 21.4291
R590 VGND.t227 VGND.n121 21.4291
R591 VGND.t141 VGND.t527 21.4291
R592 VGND.n783 VGND.t309 21.4291
R593 VGND.t41 VGND.n752 21.4291
R594 VGND.t404 VGND.n33 21.4291
R595 VGND.t99 VGND.n882 21.4291
R596 VGND.t302 VGND.n947 21.4291
R597 VGND.n502 VGND.t2 19.9891
R598 VGND.n533 VGND.t233 19.9891
R599 VGND.n553 VGND.t324 19.9891
R600 VGND.n253 VGND.t86 19.9891
R601 VGND.n633 VGND.t560 19.9891
R602 VGND.n692 VGND.t361 19.9891
R603 VGND.n155 VGND.t68 19.9891
R604 VGND.n67 VGND.t55 19.9891
R605 VGND.n876 VGND.t456 19.9891
R606 VGND.n941 VGND.t575 19.9891
R607 VGND.n931 VGND.t347 17.2861
R608 VGND.n892 VGND.t306 17.2861
R609 VGND.n899 VGND.t202 17.2861
R610 VGND.n896 VGND.t204 17.2861
R611 VGND.n811 VGND.t462 17.2861
R612 VGND.n814 VGND.t92 17.2861
R613 VGND.n840 VGND.t244 17.2861
R614 VGND.n843 VGND.t246 17.2861
R615 VGND.n30 VGND.t370 17.2861
R616 VGND.n863 VGND.t368 17.2861
R617 VGND.n36 VGND.t466 17.2861
R618 VGND.n40 VGND.t59 17.2861
R619 VGND.n73 VGND.t391 17.2861
R620 VGND.n785 VGND.t265 17.2861
R621 VGND.n781 VGND.t48 17.2861
R622 VGND.n784 VGND.t314 17.2861
R623 VGND.n118 VGND.t221 17.2861
R624 VGND.n723 VGND.t541 17.2861
R625 VGND.n124 VGND.t14 17.2861
R626 VGND.n128 VGND.t17 17.2861
R627 VGND.n702 VGND.t504 17.2861
R628 VGND.n653 VGND.t507 17.2861
R629 VGND.n664 VGND.t354 17.2861
R630 VGND.n660 VGND.t351 17.2861
R631 VGND.n166 VGND.t336 17.2861
R632 VGND.n205 VGND.t458 17.2861
R633 VGND.n170 VGND.t593 17.2861
R634 VGND.n173 VGND.t563 17.2861
R635 VGND.n620 VGND.t590 17.2861
R636 VGND.n216 VGND.t106 17.2861
R637 VGND.n226 VGND.t75 17.2861
R638 VGND.n222 VGND.t207 17.2861
R639 VGND.n305 VGND.t289 17.2861
R640 VGND.n266 VGND.t29 17.2861
R641 VGND.n273 VGND.t327 17.2861
R642 VGND.n270 VGND.t598 17.2861
R643 VGND.n515 VGND.t586 17.2861
R644 VGND.n515 VGND.t153 17.2861
R645 VGND.n518 VGND.t512 17.2861
R646 VGND.n518 VGND.t151 17.2861
R647 VGND.n473 VGND.t21 17.2861
R648 VGND.n473 VGND.t292 17.2861
R649 VGND.n472 VGND.t19 17.2861
R650 VGND.n472 VGND.t6 17.2861
R651 VGND.n347 VGND.t538 17.2861
R652 VGND.n344 VGND.t120 17.2861
R653 VGND.n343 VGND.t497 17.2861
R654 VGND.n346 VGND.t557 17.2861
R655 VGND.n925 VGND.t301 17.2649
R656 VGND.n897 VGND.t297 17.2649
R657 VGND.n900 VGND.t299 17.2649
R658 VGND.n902 VGND.t582 17.2649
R659 VGND.n917 VGND.t576 17.2649
R660 VGND.n918 VGND.t580 17.2649
R661 VGND.n845 VGND.t98 17.2649
R662 VGND.n842 VGND.t90 17.2649
R663 VGND.n839 VGND.t88 17.2649
R664 VGND.n837 VGND.t451 17.2649
R665 VGND.n818 VGND.t446 17.2649
R666 VGND.n823 VGND.t449 17.2649
R667 VGND.n43 VGND.t52 17.2649
R668 VGND.n41 VGND.t394 17.2649
R669 VGND.n37 VGND.t396 17.2649
R670 VGND.n854 VGND.t403 17.2649
R671 VGND.n62 VGND.t56 17.2649
R672 VGND.n63 VGND.t50 17.2649
R673 VGND.n777 VGND.t39 17.2649
R674 VGND.n773 VGND.t45 17.2649
R675 VGND.n769 VGND.t37 17.2649
R676 VGND.n772 VGND.t308 17.2649
R677 VGND.n776 VGND.t312 17.2649
R678 VGND.n780 VGND.t310 17.2649
R679 VGND.n131 VGND.t63 17.2649
R680 VGND.n129 VGND.t225 17.2649
R681 VGND.n125 VGND.t219 17.2649
R682 VGND.n714 VGND.t223 17.2649
R683 VGND.n150 VGND.t69 17.2649
R684 VGND.n151 VGND.t65 17.2649
R685 VGND.n657 VGND.t548 17.2649
R686 VGND.n661 VGND.t545 17.2649
R687 VGND.n665 VGND.t550 17.2649
R688 VGND.n667 VGND.t356 17.2649
R689 VGND.n687 VGND.t362 17.2649
R690 VGND.n688 VGND.t358 17.2649
R691 VGND.n176 VGND.t568 17.2649
R692 VGND.n174 VGND.t340 17.2649
R693 VGND.n171 VGND.t334 17.2649
R694 VGND.n199 VGND.t338 17.2649
R695 VGND.n191 VGND.t561 17.2649
R696 VGND.n192 VGND.t570 17.2649
R697 VGND.n611 VGND.t108 17.2649
R698 VGND.n223 VGND.t103 17.2649
R699 VGND.n227 VGND.t110 17.2649
R700 VGND.n229 VGND.t81 17.2649
R701 VGND.n248 VGND.t79 17.2649
R702 VGND.n249 VGND.t83 17.2649
R703 VGND.n299 VGND.t31 17.2649
R704 VGND.n271 VGND.t26 17.2649
R705 VGND.n274 VGND.t33 17.2649
R706 VGND.n276 VGND.t321 17.2649
R707 VGND.n291 VGND.t325 17.2649
R708 VGND.n292 VGND.t323 17.2649
R709 VGND.n520 VGND.t509 17.2649
R710 VGND.n520 VGND.t240 17.2649
R711 VGND.n523 VGND.t511 17.2649
R712 VGND.n523 VGND.t234 17.2649
R713 VGND.n526 VGND.t508 17.2649
R714 VGND.n526 VGND.t232 17.2649
R715 VGND.n318 VGND.t214 17.2649
R716 VGND.n318 VGND.t8 17.2649
R717 VGND.n478 VGND.t211 17.2649
R718 VGND.n478 VGND.t3 17.2649
R719 VGND.n481 VGND.t215 17.2649
R720 VGND.n481 VGND.t10 17.2649
R721 VGND.n341 VGND.t114 17.2649
R722 VGND.n338 VGND.t118 17.2649
R723 VGND.n335 VGND.t116 17.2649
R724 VGND.n334 VGND.t501 17.2649
R725 VGND.n337 VGND.t495 17.2649
R726 VGND.n340 VGND.t491 17.2649
R727 VGND.n962 VGND.t424 17.2313
R728 VGND.t428 VGND.n972 17.2313
R729 VGND.n988 VGND.t416 17.2313
R730 VGND.n1017 VGND.t249 17.2313
R731 VGND.t412 VGND.n1017 17.2313
R732 VGND.n1007 VGND.t284 17.2313
R733 VGND.n1007 VGND.t409 17.2313
R734 VGND.n1000 VGND.t420 17.2313
R735 VGND.t487 VGND.n1000 17.2313
R736 VGND.t147 VGND.n932 17.2313
R737 VGND.t442 VGND.n919 17.2313
R738 VGND.n812 VGND.t182 17.2313
R739 VGND.t406 VGND.n831 17.2313
R740 VGND.t156 VGND.n864 17.2313
R741 VGND.t174 VGND.n64 17.2313
R742 VGND.t139 VGND.n742 17.2313
R743 VGND.n108 VGND.t261 17.2313
R744 VGND.t383 VGND.n108 17.2313
R745 VGND.n100 VGND.t257 17.2313
R746 VGND.t438 VGND.n100 17.2313
R747 VGND.n92 VGND.t372 17.2313
R748 VGND.t167 VGND.n92 17.2313
R749 VGND.t190 VGND.n724 17.2313
R750 VGND.t521 VGND.n152 17.2313
R751 VGND.t473 VGND.n703 17.2313
R752 VGND.t253 VGND.n689 17.2313
R753 VGND.t276 VGND.n206 17.2313
R754 VGND.t135 VGND.n193 17.2313
R755 VGND.t432 VGND.n621 17.2313
R756 VGND.t280 VGND.n250 17.2313
R757 VGND.n600 VGND.t170 17.2313
R758 VGND.t131 VGND.n600 17.2313
R759 VGND.n590 VGND.t469 17.2313
R760 VGND.n590 VGND.t380 17.2313
R761 VGND.n583 VGND.t524 17.2313
R762 VGND.t198 VGND.n583 17.2313
R763 VGND.t269 VGND.n306 17.2313
R764 VGND.t484 VGND.n293 17.2313
R765 VGND.n541 VGND.t194 17.2313
R766 VGND.t386 VGND.n541 17.2313
R767 VGND.n497 VGND.t435 17.2313
R768 VGND.t163 VGND.n497 17.2313
R769 VGND.t186 VGND.n321 17.2313
R770 VGND.n443 VGND.t533 17.2313
R771 VGND.t477 VGND.n443 17.2313
R772 VGND.n433 VGND.t143 17.2313
R773 VGND.t159 VGND.n433 17.2313
R774 VGND.n425 VGND.t480 17.2313
R775 VGND.t376 VGND.n425 17.2313
R776 VGND.n399 VGND.t178 17.2313
R777 VGND.n391 VGND.t517 17.2313
R778 VGND.t127 VGND.n369 17.2313
R779 VGND.n799 VGND.t528 17.2284
R780 VGND.n764 VGND.t273 17.2284
R781 VGND.n358 VGND.t531 17.2284
R782 VGND.n800 VGND.n799 17.008
R783 VGND.n993 VGND.n992 17.001
R784 VGND.t424 VGND.n961 17.0005
R785 VGND.n1018 VGND.t249 17.0005
R786 VGND.n1018 VGND.t412 17.0005
R787 VGND.n5 VGND.t250 17.0005
R788 VGND.n3 VGND.t413 17.0005
R789 VGND.t284 VGND.n6 17.0005
R790 VGND.t409 VGND.n6 17.0005
R791 VGND.n1004 VGND.t285 17.0005
R792 VGND.n1003 VGND.t410 17.0005
R793 VGND.n1001 VGND.t420 17.0005
R794 VGND.n1001 VGND.t487 17.0005
R795 VGND.n14 VGND.t421 17.0005
R796 VGND.n13 VGND.t488 17.0005
R797 VGND.n933 VGND.t147 17.0005
R798 VGND.n924 VGND.t148 17.0005
R799 VGND.n920 VGND.t442 17.0005
R800 VGND.n909 VGND.t444 17.0005
R801 VGND.n806 VGND.t182 17.0005
R802 VGND.n848 VGND.t183 17.0005
R803 VGND.n832 VGND.t406 17.0005
R804 VGND.n824 VGND.t407 17.0005
R805 VGND.n865 VGND.t156 17.0005
R806 VGND.n853 VGND.t157 17.0005
R807 VGND.n65 VGND.t174 17.0005
R808 VGND.n52 VGND.t175 17.0005
R809 VGND.n797 VGND.t139 17.0005
R810 VGND.n793 VGND.t529 17.0005
R811 VGND.n802 VGND.t140 17.0005
R812 VGND.n759 VGND.t274 17.0005
R813 VGND.n109 VGND.t261 17.0005
R814 VGND.n109 VGND.t383 17.0005
R815 VGND.n79 VGND.t262 17.0005
R816 VGND.n78 VGND.t385 17.0005
R817 VGND.n101 VGND.t257 17.0005
R818 VGND.n101 VGND.t438 17.0005
R819 VGND.n96 VGND.t258 17.0005
R820 VGND.n95 VGND.t440 17.0005
R821 VGND.n93 VGND.t372 17.0005
R822 VGND.n93 VGND.t167 17.0005
R823 VGND.n86 VGND.t373 17.0005
R824 VGND.n85 VGND.t168 17.0005
R825 VGND.n725 VGND.t190 17.0005
R826 VGND.n713 VGND.t192 17.0005
R827 VGND.n153 VGND.t521 17.0005
R828 VGND.n140 VGND.t522 17.0005
R829 VGND.n704 VGND.t473 17.0005
R830 VGND.n708 VGND.t475 17.0005
R831 VGND.n690 VGND.t253 17.0005
R832 VGND.n676 VGND.t255 17.0005
R833 VGND.n207 VGND.t276 17.0005
R834 VGND.n198 VGND.t277 17.0005
R835 VGND.n194 VGND.t135 17.0005
R836 VGND.n183 VGND.t137 17.0005
R837 VGND.n622 VGND.t432 17.0005
R838 VGND.n610 VGND.t433 17.0005
R839 VGND.n251 VGND.t280 17.0005
R840 VGND.n238 VGND.t282 17.0005
R841 VGND.n601 VGND.t170 17.0005
R842 VGND.n601 VGND.t131 17.0005
R843 VGND.n261 VGND.t172 17.0005
R844 VGND.n259 VGND.t132 17.0005
R845 VGND.t469 VGND.n262 17.0005
R846 VGND.t380 VGND.n262 17.0005
R847 VGND.n587 VGND.t471 17.0005
R848 VGND.n586 VGND.t381 17.0005
R849 VGND.n584 VGND.t524 17.0005
R850 VGND.n584 VGND.t198 17.0005
R851 VGND.n575 VGND.t525 17.0005
R852 VGND.n574 VGND.t200 17.0005
R853 VGND.n307 VGND.t269 17.0005
R854 VGND.n298 VGND.t271 17.0005
R855 VGND.n294 VGND.t484 17.0005
R856 VGND.n283 VGND.t486 17.0005
R857 VGND.n542 VGND.t194 17.0005
R858 VGND.n542 VGND.t386 17.0005
R859 VGND.n511 VGND.t196 17.0005
R860 VGND.n315 VGND.t387 17.0005
R861 VGND.n498 VGND.t435 17.0005
R862 VGND.n498 VGND.t163 17.0005
R863 VGND.n488 VGND.t437 17.0005
R864 VGND.n487 VGND.t165 17.0005
R865 VGND.n361 VGND.t186 17.0005
R866 VGND.n349 VGND.t187 17.0005
R867 VGND.n354 VGND.t532 17.0005
R868 VGND.n444 VGND.t533 17.0005
R869 VGND.n444 VGND.t477 17.0005
R870 VGND.n409 VGND.t535 17.0005
R871 VGND.n368 VGND.t478 17.0005
R872 VGND.n434 VGND.t143 17.0005
R873 VGND.n434 VGND.t159 17.0005
R874 VGND.n429 VGND.t144 17.0005
R875 VGND.n428 VGND.t161 17.0005
R876 VGND.n426 VGND.t480 17.0005
R877 VGND.n426 VGND.t376 17.0005
R878 VGND.n418 VGND.t481 17.0005
R879 VGND.n417 VGND.t378 17.0005
R880 VGND.n382 VGND.t127 17.0005
R881 VGND.n400 VGND.t179 17.0005
R882 VGND.t178 VGND.n398 17.0005
R883 VGND.n393 VGND.t519 17.0005
R884 VGND.t517 VGND.n390 17.0005
R885 VGND.n406 VGND.t129 17.0005
R886 VGND.n404 VGND.n383 17.0005
R887 VGND.n404 VGND.n380 17.0005
R888 VGND.n404 VGND.n377 17.0005
R889 VGND.n404 VGND.n386 17.0005
R890 VGND.n404 VGND.n396 17.0005
R891 VGND.n404 VGND.n373 17.0005
R892 VGND.n446 VGND.n422 17.0005
R893 VGND.n446 VGND.n416 17.0005
R894 VGND.n446 VGND.n427 17.0005
R895 VGND.n446 VGND.n414 17.0005
R896 VGND.n446 VGND.n437 17.0005
R897 VGND.n446 VGND.n412 17.0005
R898 VGND.n446 VGND.n440 17.0005
R899 VGND.n446 VGND.n366 17.0005
R900 VGND.n446 VGND.n445 17.0005
R901 VGND.n363 VGND.n330 17.0005
R902 VGND.n363 VGND.n329 17.0005
R903 VGND.n363 VGND.n333 17.0005
R904 VGND.n451 VGND.n363 17.0005
R905 VGND.n363 VGND.n328 17.0005
R906 VGND.n452 VGND.n363 17.0005
R907 VGND.n363 VGND.n336 17.0005
R908 VGND.n453 VGND.n363 17.0005
R909 VGND.n363 VGND.n327 17.0005
R910 VGND.n454 VGND.n363 17.0005
R911 VGND.n363 VGND.n339 17.0005
R912 VGND.n455 VGND.n363 17.0005
R913 VGND.n363 VGND.n326 17.0005
R914 VGND.n456 VGND.n363 17.0005
R915 VGND.n363 VGND.n342 17.0005
R916 VGND.n457 VGND.n363 17.0005
R917 VGND.n363 VGND.n325 17.0005
R918 VGND.n458 VGND.n363 17.0005
R919 VGND.n363 VGND.n345 17.0005
R920 VGND.n459 VGND.n363 17.0005
R921 VGND.n363 VGND.n324 17.0005
R922 VGND.n460 VGND.n363 17.0005
R923 VGND.n363 VGND.n348 17.0005
R924 VGND.n461 VGND.n363 17.0005
R925 VGND.n363 VGND.n323 17.0005
R926 VGND.n462 VGND.n363 17.0005
R927 VGND.n363 VGND.n352 17.0005
R928 VGND.n363 VGND.n322 17.0005
R929 VGND.n363 VGND.n356 17.0005
R930 VGND.n464 VGND.n363 17.0005
R931 VGND.n363 VGND.n321 17.0005
R932 VGND.n363 VGND.n359 17.0005
R933 VGND.n363 VGND.n320 17.0005
R934 VGND.n363 VGND.n362 17.0005
R935 VGND.n506 VGND.n493 17.0005
R936 VGND.n506 VGND.n486 17.0005
R937 VGND.n506 VGND.n499 17.0005
R938 VGND.n506 VGND.n485 17.0005
R939 VGND.n506 VGND.n500 17.0005
R940 VGND.n506 VGND.n480 17.0005
R941 VGND.n506 VGND.n501 17.0005
R942 VGND.n506 VGND.n477 17.0005
R943 VGND.n507 VGND.n506 17.0005
R944 VGND.n506 VGND.n503 17.0005
R945 VGND.n506 VGND.n317 17.0005
R946 VGND.n506 VGND.n475 17.0005
R947 VGND.n506 VGND.n504 17.0005
R948 VGND.n506 VGND.n471 17.0005
R949 VGND.n506 VGND.n505 17.0005
R950 VGND.n544 VGND.n530 17.0005
R951 VGND.n544 VGND.n529 17.0005
R952 VGND.n544 VGND.n531 17.0005
R953 VGND.n544 VGND.n525 17.0005
R954 VGND.n544 VGND.n532 17.0005
R955 VGND.n544 VGND.n522 17.0005
R956 VGND.n544 VGND.n534 17.0005
R957 VGND.n544 VGND.n517 17.0005
R958 VGND.n544 VGND.n535 17.0005
R959 VGND.n544 VGND.n514 17.0005
R960 VGND.n544 VGND.n536 17.0005
R961 VGND.n544 VGND.n538 17.0005
R962 VGND.n544 VGND.n312 17.0005
R963 VGND.n544 VGND.n543 17.0005
R964 VGND.n309 VGND.n286 17.0005
R965 VGND.n309 VGND.n282 17.0005
R966 VGND.n549 VGND.n309 17.0005
R967 VGND.n550 VGND.n309 17.0005
R968 VGND.n309 VGND.n288 17.0005
R969 VGND.n551 VGND.n309 17.0005
R970 VGND.n309 VGND.n279 17.0005
R971 VGND.n552 VGND.n309 17.0005
R972 VGND.n309 VGND.n295 17.0005
R973 VGND.n309 VGND.n278 17.0005
R974 VGND.n554 VGND.n309 17.0005
R975 VGND.n555 VGND.n309 17.0005
R976 VGND.n556 VGND.n309 17.0005
R977 VGND.n557 VGND.n309 17.0005
R978 VGND.n558 VGND.n309 17.0005
R979 VGND.n559 VGND.n309 17.0005
R980 VGND.n309 VGND.n301 17.0005
R981 VGND.n560 VGND.n309 17.0005
R982 VGND.n309 VGND.n268 17.0005
R983 VGND.n561 VGND.n309 17.0005
R984 VGND.n562 VGND.n309 17.0005
R985 VGND.n563 VGND.n309 17.0005
R986 VGND.n309 VGND.n303 17.0005
R987 VGND.n564 VGND.n309 17.0005
R988 VGND.n309 VGND.n264 17.0005
R989 VGND.n309 VGND.n308 17.0005
R990 VGND.n603 VGND.n580 17.0005
R991 VGND.n603 VGND.n573 17.0005
R992 VGND.n603 VGND.n585 17.0005
R993 VGND.n603 VGND.n571 17.0005
R994 VGND.n603 VGND.n594 17.0005
R995 VGND.n604 VGND.n603 17.0005
R996 VGND.n603 VGND.n597 17.0005
R997 VGND.n603 VGND.n569 17.0005
R998 VGND.n603 VGND.n602 17.0005
R999 VGND.n624 VGND.n241 17.0005
R1000 VGND.n624 VGND.n237 17.0005
R1001 VGND.n624 VGND.n242 17.0005
R1002 VGND.n624 VGND.n234 17.0005
R1003 VGND.n624 VGND.n244 17.0005
R1004 VGND.n624 VGND.n245 17.0005
R1005 VGND.n624 VGND.n233 17.0005
R1006 VGND.n624 VGND.n232 17.0005
R1007 VGND.n624 VGND.n252 17.0005
R1008 VGND.n624 VGND.n231 17.0005
R1009 VGND.n624 VGND.n254 17.0005
R1010 VGND.n624 VGND.n225 17.0005
R1011 VGND.n624 VGND.n255 17.0005
R1012 VGND.n624 VGND.n221 17.0005
R1013 VGND.n624 VGND.n256 17.0005
R1014 VGND.n624 VGND.n219 17.0005
R1015 VGND.n624 VGND.n613 17.0005
R1016 VGND.n624 VGND.n614 17.0005
R1017 VGND.n624 VGND.n218 17.0005
R1018 VGND.n624 VGND.n215 17.0005
R1019 VGND.n624 VGND.n615 17.0005
R1020 VGND.n624 VGND.n213 17.0005
R1021 VGND.n624 VGND.n617 17.0005
R1022 VGND.n624 VGND.n618 17.0005
R1023 VGND.n624 VGND.n212 17.0005
R1024 VGND.n624 VGND.n623 17.0005
R1025 VGND.n209 VGND.n186 17.0005
R1026 VGND.n209 VGND.n182 17.0005
R1027 VGND.n629 VGND.n209 17.0005
R1028 VGND.n630 VGND.n209 17.0005
R1029 VGND.n209 VGND.n188 17.0005
R1030 VGND.n631 VGND.n209 17.0005
R1031 VGND.n209 VGND.n179 17.0005
R1032 VGND.n632 VGND.n209 17.0005
R1033 VGND.n209 VGND.n195 17.0005
R1034 VGND.n209 VGND.n178 17.0005
R1035 VGND.n634 VGND.n209 17.0005
R1036 VGND.n635 VGND.n209 17.0005
R1037 VGND.n636 VGND.n209 17.0005
R1038 VGND.n637 VGND.n209 17.0005
R1039 VGND.n638 VGND.n209 17.0005
R1040 VGND.n639 VGND.n209 17.0005
R1041 VGND.n209 VGND.n201 17.0005
R1042 VGND.n640 VGND.n209 17.0005
R1043 VGND.n209 VGND.n168 17.0005
R1044 VGND.n641 VGND.n209 17.0005
R1045 VGND.n642 VGND.n209 17.0005
R1046 VGND.n643 VGND.n209 17.0005
R1047 VGND.n209 VGND.n203 17.0005
R1048 VGND.n644 VGND.n209 17.0005
R1049 VGND.n209 VGND.n164 17.0005
R1050 VGND.n209 VGND.n208 17.0005
R1051 VGND.n706 VGND.n679 17.0005
R1052 VGND.n706 VGND.n675 17.0005
R1053 VGND.n706 VGND.n681 17.0005
R1054 VGND.n706 VGND.n672 17.0005
R1055 VGND.n706 VGND.n683 17.0005
R1056 VGND.n706 VGND.n684 17.0005
R1057 VGND.n706 VGND.n671 17.0005
R1058 VGND.n706 VGND.n670 17.0005
R1059 VGND.n706 VGND.n691 17.0005
R1060 VGND.n706 VGND.n669 17.0005
R1061 VGND.n706 VGND.n693 17.0005
R1062 VGND.n706 VGND.n663 17.0005
R1063 VGND.n706 VGND.n694 17.0005
R1064 VGND.n706 VGND.n659 17.0005
R1065 VGND.n706 VGND.n695 17.0005
R1066 VGND.n706 VGND.n656 17.0005
R1067 VGND.n707 VGND.n706 17.0005
R1068 VGND.n706 VGND.n696 17.0005
R1069 VGND.n706 VGND.n655 17.0005
R1070 VGND.n706 VGND.n652 17.0005
R1071 VGND.n706 VGND.n697 17.0005
R1072 VGND.n706 VGND.n650 17.0005
R1073 VGND.n706 VGND.n699 17.0005
R1074 VGND.n706 VGND.n700 17.0005
R1075 VGND.n706 VGND.n649 17.0005
R1076 VGND.n706 VGND.n705 17.0005
R1077 VGND.n727 VGND.n143 17.0005
R1078 VGND.n727 VGND.n139 17.0005
R1079 VGND.n727 VGND.n144 17.0005
R1080 VGND.n727 VGND.n136 17.0005
R1081 VGND.n727 VGND.n146 17.0005
R1082 VGND.n727 VGND.n147 17.0005
R1083 VGND.n727 VGND.n135 17.0005
R1084 VGND.n727 VGND.n134 17.0005
R1085 VGND.n727 VGND.n154 17.0005
R1086 VGND.n727 VGND.n133 17.0005
R1087 VGND.n727 VGND.n156 17.0005
R1088 VGND.n727 VGND.n127 17.0005
R1089 VGND.n727 VGND.n157 17.0005
R1090 VGND.n727 VGND.n123 17.0005
R1091 VGND.n727 VGND.n158 17.0005
R1092 VGND.n727 VGND.n121 17.0005
R1093 VGND.n727 VGND.n716 17.0005
R1094 VGND.n727 VGND.n717 17.0005
R1095 VGND.n727 VGND.n120 17.0005
R1096 VGND.n727 VGND.n117 17.0005
R1097 VGND.n727 VGND.n718 17.0005
R1098 VGND.n727 VGND.n115 17.0005
R1099 VGND.n727 VGND.n720 17.0005
R1100 VGND.n727 VGND.n721 17.0005
R1101 VGND.n727 VGND.n114 17.0005
R1102 VGND.n727 VGND.n726 17.0005
R1103 VGND.n111 VGND.n90 17.0005
R1104 VGND.n111 VGND.n84 17.0005
R1105 VGND.n111 VGND.n94 17.0005
R1106 VGND.n111 VGND.n83 17.0005
R1107 VGND.n111 VGND.n104 17.0005
R1108 VGND.n111 VGND.n82 17.0005
R1109 VGND.n111 VGND.n106 17.0005
R1110 VGND.n111 VGND.n76 17.0005
R1111 VGND.n111 VGND.n110 17.0005
R1112 VGND.n800 VGND.n762 17.0005
R1113 VGND.n800 VGND.n758 17.0005
R1114 VGND.n800 VGND.n766 17.0005
R1115 VGND.n800 VGND.n767 17.0005
R1116 VGND.n800 VGND.n757 17.0005
R1117 VGND.n800 VGND.n756 17.0005
R1118 VGND.n800 VGND.n770 17.0005
R1119 VGND.n800 VGND.n771 17.0005
R1120 VGND.n800 VGND.n755 17.0005
R1121 VGND.n800 VGND.n754 17.0005
R1122 VGND.n800 VGND.n774 17.0005
R1123 VGND.n800 VGND.n775 17.0005
R1124 VGND.n800 VGND.n753 17.0005
R1125 VGND.n800 VGND.n752 17.0005
R1126 VGND.n800 VGND.n778 17.0005
R1127 VGND.n800 VGND.n779 17.0005
R1128 VGND.n800 VGND.n751 17.0005
R1129 VGND.n800 VGND.n750 17.0005
R1130 VGND.n800 VGND.n782 17.0005
R1131 VGND.n800 VGND.n783 17.0005
R1132 VGND.n800 VGND.n749 17.0005
R1133 VGND.n800 VGND.n748 17.0005
R1134 VGND.n800 VGND.n786 17.0005
R1135 VGND.n800 VGND.n787 17.0005
R1136 VGND.n800 VGND.n747 17.0005
R1137 VGND.n800 VGND.n746 17.0005
R1138 VGND.n801 VGND.n800 17.0005
R1139 VGND.n800 VGND.n788 17.0005
R1140 VGND.n800 VGND.n745 17.0005
R1141 VGND.n800 VGND.n743 17.0005
R1142 VGND.n800 VGND.n790 17.0005
R1143 VGND.n800 VGND.n742 17.0005
R1144 VGND.n800 VGND.n795 17.0005
R1145 VGND.n800 VGND.n741 17.0005
R1146 VGND.n867 VGND.n55 17.0005
R1147 VGND.n867 VGND.n51 17.0005
R1148 VGND.n867 VGND.n56 17.0005
R1149 VGND.n867 VGND.n48 17.0005
R1150 VGND.n867 VGND.n58 17.0005
R1151 VGND.n867 VGND.n59 17.0005
R1152 VGND.n867 VGND.n47 17.0005
R1153 VGND.n867 VGND.n46 17.0005
R1154 VGND.n867 VGND.n66 17.0005
R1155 VGND.n867 VGND.n45 17.0005
R1156 VGND.n867 VGND.n68 17.0005
R1157 VGND.n867 VGND.n39 17.0005
R1158 VGND.n867 VGND.n69 17.0005
R1159 VGND.n867 VGND.n35 17.0005
R1160 VGND.n867 VGND.n70 17.0005
R1161 VGND.n867 VGND.n33 17.0005
R1162 VGND.n867 VGND.n856 17.0005
R1163 VGND.n867 VGND.n857 17.0005
R1164 VGND.n867 VGND.n32 17.0005
R1165 VGND.n867 VGND.n29 17.0005
R1166 VGND.n867 VGND.n858 17.0005
R1167 VGND.n867 VGND.n27 17.0005
R1168 VGND.n867 VGND.n860 17.0005
R1169 VGND.n867 VGND.n861 17.0005
R1170 VGND.n867 VGND.n26 17.0005
R1171 VGND.n867 VGND.n866 17.0005
R1172 VGND.n826 VGND.n23 17.0005
R1173 VGND.n828 VGND.n23 17.0005
R1174 VGND.n872 VGND.n23 17.0005
R1175 VGND.n873 VGND.n23 17.0005
R1176 VGND.n822 VGND.n23 17.0005
R1177 VGND.n874 VGND.n23 17.0005
R1178 VGND.n820 VGND.n23 17.0005
R1179 VGND.n875 VGND.n23 17.0005
R1180 VGND.n833 VGND.n23 17.0005
R1181 VGND.n835 VGND.n23 17.0005
R1182 VGND.n877 VGND.n23 17.0005
R1183 VGND.n878 VGND.n23 17.0005
R1184 VGND.n879 VGND.n23 17.0005
R1185 VGND.n880 VGND.n23 17.0005
R1186 VGND.n881 VGND.n23 17.0005
R1187 VGND.n882 VGND.n23 17.0005
R1188 VGND.n847 VGND.n23 17.0005
R1189 VGND.n883 VGND.n23 17.0005
R1190 VGND.n816 VGND.n23 17.0005
R1191 VGND.n884 VGND.n23 17.0005
R1192 VGND.n885 VGND.n23 17.0005
R1193 VGND.n886 VGND.n23 17.0005
R1194 VGND.n810 VGND.n23 17.0005
R1195 VGND.n887 VGND.n23 17.0005
R1196 VGND.n808 VGND.n23 17.0005
R1197 VGND.n805 VGND.n23 17.0005
R1198 VGND.n935 VGND.n912 17.0005
R1199 VGND.n935 VGND.n908 17.0005
R1200 VGND.n937 VGND.n935 17.0005
R1201 VGND.n938 VGND.n935 17.0005
R1202 VGND.n935 VGND.n914 17.0005
R1203 VGND.n939 VGND.n935 17.0005
R1204 VGND.n935 VGND.n905 17.0005
R1205 VGND.n940 VGND.n935 17.0005
R1206 VGND.n935 VGND.n921 17.0005
R1207 VGND.n935 VGND.n904 17.0005
R1208 VGND.n942 VGND.n935 17.0005
R1209 VGND.n943 VGND.n935 17.0005
R1210 VGND.n944 VGND.n935 17.0005
R1211 VGND.n945 VGND.n935 17.0005
R1212 VGND.n946 VGND.n935 17.0005
R1213 VGND.n947 VGND.n935 17.0005
R1214 VGND.n935 VGND.n927 17.0005
R1215 VGND.n948 VGND.n935 17.0005
R1216 VGND.n935 VGND.n894 17.0005
R1217 VGND.n949 VGND.n935 17.0005
R1218 VGND.n950 VGND.n935 17.0005
R1219 VGND.n951 VGND.n935 17.0005
R1220 VGND.n935 VGND.n929 17.0005
R1221 VGND.n952 VGND.n935 17.0005
R1222 VGND.n935 VGND.n890 17.0005
R1223 VGND.n935 VGND.n934 17.0005
R1224 VGND.n1020 VGND.n997 17.0005
R1225 VGND.n1020 VGND.n12 17.0005
R1226 VGND.n1020 VGND.n1002 17.0005
R1227 VGND.n1020 VGND.n10 17.0005
R1228 VGND.n1020 VGND.n1011 17.0005
R1229 VGND.n1021 VGND.n1020 17.0005
R1230 VGND.n1020 VGND.n1014 17.0005
R1231 VGND.n1020 VGND.n8 17.0005
R1232 VGND.n1020 VGND.n1019 17.0005
R1233 VGND.n973 VGND.t428 17.0005
R1234 VGND.n21 VGND.t430 17.0005
R1235 VGND.n983 VGND.t416 17.0005
R1236 VGND.n990 VGND.t417 17.0005
R1237 VGND.n19 VGND.n18 17.0005
R1238 VGND.n987 VGND.n19 17.0005
R1239 VGND.n985 VGND.n19 17.0005
R1240 VGND.n982 VGND.n19 17.0005
R1241 VGND.n978 VGND.n971 17.0005
R1242 VGND.n978 VGND.n968 17.0005
R1243 VGND.n978 VGND.n976 17.0005
R1244 VGND.n978 VGND.n966 17.0005
R1245 VGND.n978 VGND.n963 17.0005
R1246 VGND.n978 VGND.n958 17.0005
R1247 VGND.n978 VGND.n957 17.0005
R1248 VGND.n0 VGND.t426 17.0005
R1249 VGND.n797 VGND.t640 15.3099
R1250 VGND.n960 VGND.t657 15.2865
R1251 VGND.n1016 VGND.t686 15.2865
R1252 VGND.n1016 VGND.t647 15.2865
R1253 VGND.n1009 VGND.t680 15.2865
R1254 VGND.n1009 VGND.t665 15.2865
R1255 VGND.n999 VGND.t611 15.2865
R1256 VGND.n999 VGND.t655 15.2865
R1257 VGND.n930 VGND.t672 15.2865
R1258 VGND.n916 VGND.t624 15.2865
R1259 VGND.n807 VGND.t650 15.2865
R1260 VGND.n819 VGND.t605 15.2865
R1261 VGND.n862 VGND.t658 15.2865
R1262 VGND.n61 VGND.t674 15.2865
R1263 VGND.n107 VGND.t703 15.2865
R1264 VGND.n107 VGND.t604 15.2865
R1265 VGND.n102 VGND.t700 15.2865
R1266 VGND.n102 VGND.t601 15.2865
R1267 VGND.n91 VGND.t629 15.2865
R1268 VGND.n91 VGND.t638 15.2865
R1269 VGND.n722 VGND.t606 15.2865
R1270 VGND.n149 VGND.t614 15.2865
R1271 VGND.n701 VGND.t662 15.2865
R1272 VGND.n686 VGND.t616 15.2865
R1273 VGND.n204 VGND.t671 15.2865
R1274 VGND.n190 VGND.t602 15.2865
R1275 VGND.n619 VGND.t656 15.2865
R1276 VGND.n247 VGND.t688 15.2865
R1277 VGND.n599 VGND.t635 15.2865
R1278 VGND.n599 VGND.t636 15.2865
R1279 VGND.n592 VGND.t699 15.2865
R1280 VGND.n592 VGND.t702 15.2865
R1281 VGND.n582 VGND.t664 15.2865
R1282 VGND.n582 VGND.t667 15.2865
R1283 VGND.n304 VGND.t698 15.2865
R1284 VGND.n290 VGND.t677 15.2865
R1285 VGND.n540 VGND.t687 15.2865
R1286 VGND.n540 VGND.t684 15.2865
R1287 VGND.n496 VGND.t668 15.2865
R1288 VGND.n496 VGND.t675 15.2865
R1289 VGND.n360 VGND.t617 15.2865
R1290 VGND.n442 VGND.t704 15.2865
R1291 VGND.n442 VGND.t607 15.2865
R1292 VGND.n435 VGND.t660 15.2865
R1293 VGND.n435 VGND.t670 15.2865
R1294 VGND.n424 VGND.t631 15.2865
R1295 VGND.n424 VGND.t641 15.2865
R1296 VGND.n381 VGND.t696 15.2865
R1297 VGND.n397 VGND.t618 15.2865
R1298 VGND.n389 VGND.t653 15.2865
R1299 VGND.n974 VGND.t683 15.2865
R1300 VGND.n984 VGND.t669 15.2865
R1301 VGND.n3 VGND.t690 15.2696
R1302 VGND.n5 VGND.t678 15.2696
R1303 VGND.n1003 VGND.t612 15.2696
R1304 VGND.n1004 VGND.t673 15.2696
R1305 VGND.n13 VGND.t619 15.2696
R1306 VGND.n14 VGND.t663 15.2696
R1307 VGND.n909 VGND.t639 15.2696
R1308 VGND.n824 VGND.t615 15.2696
R1309 VGND.n52 VGND.t691 15.2696
R1310 VGND.n78 VGND.t705 15.2696
R1311 VGND.n79 VGND.t608 15.2696
R1312 VGND.n95 VGND.t632 15.2696
R1313 VGND.n96 VGND.t642 15.2696
R1314 VGND.n85 VGND.t645 15.2696
R1315 VGND.n86 VGND.t649 15.2696
R1316 VGND.n140 VGND.t626 15.2696
R1317 VGND.n676 VGND.t679 15.2696
R1318 VGND.n183 VGND.t661 15.2696
R1319 VGND.n238 VGND.t643 15.2696
R1320 VGND.n259 VGND.t682 15.2696
R1321 VGND.n261 VGND.t685 15.2696
R1322 VGND.n586 VGND.t628 15.2696
R1323 VGND.n587 VGND.t630 15.2696
R1324 VGND.n574 VGND.t620 15.2696
R1325 VGND.n575 VGND.t622 15.2696
R1326 VGND.n283 VGND.t634 15.2696
R1327 VGND.n315 VGND.t623 15.2696
R1328 VGND.n511 VGND.t621 15.2696
R1329 VGND.n487 VGND.t625 15.2696
R1330 VGND.n488 VGND.t633 15.2696
R1331 VGND.n349 VGND.t666 15.2696
R1332 VGND.n368 VGND.t648 15.2696
R1333 VGND.n409 VGND.t652 15.2696
R1334 VGND.n428 VGND.t697 15.2696
R1335 VGND.n429 VGND.t600 15.2696
R1336 VGND.n417 VGND.t695 15.2696
R1337 VGND.n418 VGND.t701 15.2696
R1338 VGND.n400 VGND.t689 15.2696
R1339 VGND.n393 VGND.t693 15.2696
R1340 VGND.n406 VGND.t637 15.2696
R1341 VGND.n21 VGND.t692 15.2696
R1342 VGND.n990 VGND.t681 15.2696
R1343 VGND.n0 VGND.t694 15.2696
R1344 VGND.n793 VGND.t603 15.2596
R1345 VGND.n759 VGND.t627 15.2596
R1346 VGND.n354 VGND.t610 15.2596
R1347 VGND.n922 VGND.t676 15.2471
R1348 VGND.n817 VGND.t654 15.2471
R1349 VGND.n71 VGND.t659 15.2471
R1350 VGND.n744 VGND.t644 15.2471
R1351 VGND.n159 VGND.t651 15.2471
R1352 VGND.n161 VGND.t609 15.2471
R1353 VGND.n196 VGND.t613 15.2471
R1354 VGND.n257 VGND.t706 15.2471
R1355 VGND.n296 VGND.t646 15.2471
R1356 VGND.n903 VGND.t295 8.76785
R1357 VGND.n907 VGND.t574 8.76785
R1358 VGND.n836 VGND.t94 8.76785
R1359 VGND.n829 VGND.t455 8.76785
R1360 VGND.n44 VGND.t399 8.76785
R1361 VGND.n50 VGND.t54 8.76785
R1362 VGND.n765 VGND.t43 8.76785
R1363 VGND.n768 VGND.t316 8.76785
R1364 VGND.n132 VGND.t229 8.76785
R1365 VGND.n138 VGND.t72 8.76785
R1366 VGND.n668 VGND.t554 8.76785
R1367 VGND.n674 VGND.t365 8.76785
R1368 VGND.n177 VGND.t344 8.76785
R1369 VGND.n181 VGND.t565 8.76785
R1370 VGND.n230 VGND.t101 8.76785
R1371 VGND.n236 VGND.t77 8.76785
R1372 VGND.n277 VGND.t24 8.76785
R1373 VGND.n281 VGND.t329 8.76785
R1374 VGND.n528 VGND.t513 8.76785
R1375 VGND.n528 VGND.t237 8.76785
R1376 VGND.n484 VGND.t210 8.76785
R1377 VGND.n484 VGND.t1 8.76785
R1378 VGND.n332 VGND.t122 8.76785
R1379 VGND.n331 VGND.t493 8.76785
R1380 VGND.n992 VGND.n991 8.501
R1381 VGND.n980 VGND.n979 8.501
R1382 VGND.n404 VGND.n378 8.47111
R1383 VGND.n404 VGND.n392 8.47111
R1384 VGND.n404 VGND.n370 8.47111
R1385 VGND.n506 VGND.n482 8.47111
R1386 VGND.n506 VGND.n479 8.47111
R1387 VGND.n506 VGND.n476 8.47111
R1388 VGND.n506 VGND.n474 8.47111
R1389 VGND.n544 VGND.n527 8.47111
R1390 VGND.n544 VGND.n524 8.47111
R1391 VGND.n544 VGND.n521 8.47111
R1392 VGND.n544 VGND.n519 8.47111
R1393 VGND.n544 VGND.n516 8.47111
R1394 VGND.n544 VGND.n513 8.47111
R1395 VGND.n309 VGND.n280 8.47111
R1396 VGND.n309 VGND.n275 8.47111
R1397 VGND.n309 VGND.n272 8.47111
R1398 VGND.n309 VGND.n269 8.47111
R1399 VGND.n309 VGND.n265 8.47111
R1400 VGND.n624 VGND.n235 8.47111
R1401 VGND.n624 VGND.n228 8.47111
R1402 VGND.n624 VGND.n224 8.47111
R1403 VGND.n624 VGND.n220 8.47111
R1404 VGND.n624 VGND.n214 8.47111
R1405 VGND.n209 VGND.n180 8.47111
R1406 VGND.n209 VGND.n175 8.47111
R1407 VGND.n209 VGND.n172 8.47111
R1408 VGND.n209 VGND.n169 8.47111
R1409 VGND.n209 VGND.n165 8.47111
R1410 VGND.n706 VGND.n673 8.47111
R1411 VGND.n706 VGND.n666 8.47111
R1412 VGND.n706 VGND.n662 8.47111
R1413 VGND.n706 VGND.n658 8.47111
R1414 VGND.n706 VGND.n651 8.47111
R1415 VGND.n727 VGND.n137 8.47111
R1416 VGND.n727 VGND.n130 8.47111
R1417 VGND.n727 VGND.n126 8.47111
R1418 VGND.n727 VGND.n122 8.47111
R1419 VGND.n727 VGND.n116 8.47111
R1420 VGND.n867 VGND.n49 8.47111
R1421 VGND.n867 VGND.n42 8.47111
R1422 VGND.n867 VGND.n38 8.47111
R1423 VGND.n867 VGND.n34 8.47111
R1424 VGND.n867 VGND.n28 8.47111
R1425 VGND.n830 VGND.n23 8.47111
R1426 VGND.n838 VGND.n23 8.47111
R1427 VGND.n841 VGND.n23 8.47111
R1428 VGND.n844 VGND.n23 8.47111
R1429 VGND.n813 VGND.n23 8.47111
R1430 VGND.n935 VGND.n906 8.47111
R1431 VGND.n935 VGND.n901 8.47111
R1432 VGND.n935 VGND.n898 8.47111
R1433 VGND.n935 VGND.n895 8.47111
R1434 VGND.n935 VGND.n891 8.47111
R1435 VGND.n989 VGND.n19 8.47111
R1436 VGND.n978 VGND.n20 8.47111
R1437 VGND.n408 VGND.n407 7.5029
R1438 VGND.n1026 VGND.n1025 7.2005
R1439 VGND.n1024 VGND.n1023 7.2005
R1440 VGND.n923 VGND.n2 7.2005
R1441 VGND.n850 VGND.n849 7.2005
R1442 VGND.n852 VGND.n851 7.2005
R1443 VGND.n804 VGND.n803 7.2005
R1444 VGND.n80 VGND.n72 7.2005
R1445 VGND.n712 VGND.n711 7.2005
R1446 VGND.n710 VGND.n709 7.2005
R1447 VGND.n197 VGND.n160 7.2005
R1448 VGND.n609 VGND.n608 7.2005
R1449 VGND.n607 VGND.n606 7.2005
R1450 VGND.n297 VGND.n258 7.2005
R1451 VGND.n512 VGND.n510 7.2005
R1452 VGND.n509 VGND.n508 7.2005
R1453 VGND VGND.n316 7.2005
R1454 VGND.n410 VGND.n408 7.2005
R1455 VGND.n405 VGND.n404 5.64608
R1456 VGND.n404 VGND.n375 5.64608
R1457 VGND.n404 VGND.n402 5.64608
R1458 VGND.n506 VGND.n470 5.63466
R1459 VGND.n456 VGND.t494 4.28621
R1460 VGND.n455 VGND.t117 4.28621
R1461 VGND.n558 VGND.t25 4.28621
R1462 VGND.n256 VGND.t102 4.28621
R1463 VGND.n638 VGND.t345 4.28621
R1464 VGND.n695 VGND.t555 4.28621
R1465 VGND.n158 VGND.t230 4.28621
R1466 VGND.t311 VGND.n750 4.28621
R1467 VGND.n775 VGND.t44 4.28621
R1468 VGND.n70 VGND.t395 4.28621
R1469 VGND.n881 VGND.t89 4.28621
R1470 VGND.n946 VGND.t304 4.28621
R1471 VGND.n446 VGND.n420 4.20468
R1472 VGND.n446 VGND.n432 4.20468
R1473 VGND.n446 VGND.n367 4.20468
R1474 VGND.n506 VGND.n490 4.20468
R1475 VGND.n544 VGND.n313 4.20468
R1476 VGND.n603 VGND.n577 4.20468
R1477 VGND.n603 VGND.n591 4.20468
R1478 VGND.n603 VGND.n260 4.20468
R1479 VGND.n111 VGND.n88 4.20468
R1480 VGND.n111 VGND.n99 4.20468
R1481 VGND.n111 VGND.n77 4.20468
R1482 VGND.n1020 VGND.n16 4.20468
R1483 VGND.n1020 VGND.n1008 4.20468
R1484 VGND.n1020 VGND.n4 4.20468
R1485 VGND.n978 VGND.n1 4.20455
R1486 VGND.n957 VGND 0.806068
R1487 VGND.n383 VGND 0.806068
R1488 VGND.n1019 VGND 0.803417
R1489 VGND.n110 VGND 0.803417
R1490 VGND.n602 VGND 0.803417
R1491 VGND.n543 VGND 0.803417
R1492 VGND.n445 VGND 0.803417
R1493 VGND.n1022 VGND 0.79925
R1494 VGND.n1005 VGND 0.79925
R1495 VGND.n81 VGND 0.79925
R1496 VGND.n97 VGND 0.79925
R1497 VGND.n605 VGND 0.79925
R1498 VGND.n588 VGND 0.79925
R1499 VGND.n495 VGND 0.79925
R1500 VGND.n411 VGND 0.79925
R1501 VGND.n430 VGND 0.79925
R1502 VGND.n395 VGND 0.79925
R1503 VGND.n376 VGND 0.79925
R1504 VGND.n965 VGND 0.79925
R1505 VGND.n981 VGND 0.79925
R1506 VGND.n915 VGND 0.67925
R1507 VGND.n834 VGND 0.67925
R1508 VGND.n60 VGND 0.67925
R1509 VGND.n148 VGND 0.67925
R1510 VGND.n685 VGND 0.67925
R1511 VGND.n189 VGND 0.67925
R1512 VGND.n246 VGND 0.67925
R1513 VGND.n289 VGND 0.67925
R1514 VGND.n447 VGND.n446 0.649813
R1515 VGND.n446 VGND.n365 0.649813
R1516 VGND.n450 VGND.n363 0.649813
R1517 VGND.n463 VGND.n363 0.649813
R1518 VGND.n465 VGND.n363 0.649813
R1519 VGND.n466 VGND.n363 0.649813
R1520 VGND.n506 VGND.n491 0.649813
R1521 VGND.n506 VGND.n502 0.649813
R1522 VGND.n506 VGND.n469 0.649813
R1523 VGND.n545 VGND.n544 0.649813
R1524 VGND.n544 VGND.n533 0.649813
R1525 VGND.n544 VGND.n311 0.649813
R1526 VGND.n548 VGND.n309 0.649813
R1527 VGND.n553 VGND.n309 0.649813
R1528 VGND.n565 VGND.n309 0.649813
R1529 VGND.n603 VGND.n578 0.649813
R1530 VGND.n603 VGND.n568 0.649813
R1531 VGND.n625 VGND.n624 0.649813
R1532 VGND.n624 VGND.n253 0.649813
R1533 VGND.n624 VGND.n211 0.649813
R1534 VGND.n628 VGND.n209 0.649813
R1535 VGND.n633 VGND.n209 0.649813
R1536 VGND.n645 VGND.n209 0.649813
R1537 VGND.n706 VGND.n680 0.649813
R1538 VGND.n706 VGND.n692 0.649813
R1539 VGND.n706 VGND.n648 0.649813
R1540 VGND.n728 VGND.n727 0.649813
R1541 VGND.n727 VGND.n155 0.649813
R1542 VGND.n727 VGND.n113 0.649813
R1543 VGND.n731 VGND.n111 0.649813
R1544 VGND.n737 VGND.n111 0.649813
R1545 VGND.n800 VGND.n763 0.649813
R1546 VGND.n800 VGND.n740 0.649813
R1547 VGND.n868 VGND.n867 0.649813
R1548 VGND.n867 VGND.n67 0.649813
R1549 VGND.n867 VGND.n25 0.649813
R1550 VGND.n871 VGND.n23 0.649813
R1551 VGND.n876 VGND.n23 0.649813
R1552 VGND.n888 VGND.n23 0.649813
R1553 VGND.n936 VGND.n935 0.649813
R1554 VGND.n941 VGND.n935 0.649813
R1555 VGND.n953 VGND.n935 0.649813
R1556 VGND.n1020 VGND.n995 0.649813
R1557 VGND.n1020 VGND.n7 0.649813
R1558 VGND.n404 VGND.n384 0.389775
R1559 VGND.n404 VGND.n364 0.389775
R1560 VGND.n978 VGND.n956 0.389775
R1561 VGND.n408 VGND.n316 0.3029
R1562 VGND.n509 VGND.n316 0.3029
R1563 VGND.n510 VGND.n509 0.3029
R1564 VGND.n510 VGND.n258 0.3029
R1565 VGND.n607 VGND.n258 0.3029
R1566 VGND.n608 VGND.n607 0.3029
R1567 VGND.n608 VGND.n160 0.3029
R1568 VGND.n710 VGND.n160 0.3029
R1569 VGND.n711 VGND.n710 0.3029
R1570 VGND.n711 VGND.n72 0.3029
R1571 VGND.n804 VGND.n72 0.3029
R1572 VGND.n851 VGND.n804 0.3029
R1573 VGND.n851 VGND.n850 0.3029
R1574 VGND.n850 VGND.n2 0.3029
R1575 VGND.n1024 VGND.n2 0.3029
R1576 VGND.n1025 VGND.n1024 0.3029
R1577 VGND.n791 VGND 0.28675
R1578 VGND.n959 VGND 0.2355
R1579 VGND.n928 VGND 0.2355
R1580 VGND.n809 VGND 0.2355
R1581 VGND.n859 VGND 0.2355
R1582 VGND.n719 VGND 0.2355
R1583 VGND.n698 VGND 0.2355
R1584 VGND.n202 VGND 0.2355
R1585 VGND.n616 VGND 0.2355
R1586 VGND.n302 VGND 0.2355
R1587 VGND.n379 VGND 0.2355
R1588 VGND.n372 VGND 0.2355
R1589 VGND.n388 VGND 0.2355
R1590 VGND.n975 VGND 0.2355
R1591 VGND.n986 VGND 0.2355
R1592 VGND.n792 VGND 0.21425
R1593 VGND.n353 VGND 0.21425
R1594 VGND.n362 VGND 0.206068
R1595 VGND.n1026 VGND 0.203
R1596 VGND.n1023 VGND 0.203
R1597 VGND.n1006 VGND 0.203
R1598 VGND.n15 VGND 0.203
R1599 VGND.n893 VGND 0.203
R1600 VGND.n815 VGND 0.203
R1601 VGND.n31 VGND 0.203
R1602 VGND.n789 VGND 0.203
R1603 VGND.n80 VGND 0.203
R1604 VGND.n98 VGND 0.203
R1605 VGND.n87 VGND 0.203
R1606 VGND.n119 VGND 0.203
R1607 VGND.n654 VGND 0.203
R1608 VGND.n167 VGND 0.203
R1609 VGND.n217 VGND 0.203
R1610 VGND.n606 VGND 0.203
R1611 VGND.n589 VGND 0.203
R1612 VGND.n576 VGND 0.203
R1613 VGND.n267 VGND 0.203
R1614 VGND.n512 VGND 0.203
R1615 VGND.n489 VGND 0.203
R1616 VGND.n410 VGND 0.203
R1617 VGND.n431 VGND 0.203
R1618 VGND.n419 VGND 0.203
R1619 VGND.n401 VGND 0.203
R1620 VGND.n394 VGND 0.203
R1621 VGND.n407 VGND 0.203
R1622 VGND.n980 VGND 0.203
R1623 VGND.n991 VGND 0.203
R1624 VGND.n913 VGND 0.191864
R1625 VGND.n821 VGND 0.191864
R1626 VGND.n57 VGND 0.191864
R1627 VGND.n145 VGND 0.191864
R1628 VGND.n682 VGND 0.191864
R1629 VGND.n187 VGND 0.191864
R1630 VGND.n243 VGND 0.191864
R1631 VGND.n287 VGND 0.191864
R1632 VGND.n761 VGND 0.186654
R1633 VGND.n402 VGND.n399 0.185752
R1634 VGND.n391 VGND.n375 0.185752
R1635 VGND.n405 VGND.n369 0.185752
R1636 VGND.n372 VGND.n370 0.167039
R1637 VGND.n392 VGND.n388 0.167039
R1638 VGND.n379 VGND.n378 0.167039
R1639 VGND.n516 VGND.n515 0.160789
R1640 VGND.n474 VGND.n473 0.160789
R1641 VGND.n980 VGND.n20 0.158289
R1642 VGND.n991 VGND.n989 0.158289
R1643 VGND.n907 VGND.n906 0.155789
R1644 VGND.n830 VGND.n829 0.155789
R1645 VGND.n50 VGND.n49 0.155789
R1646 VGND.n138 VGND.n137 0.155789
R1647 VGND.n674 VGND.n673 0.155789
R1648 VGND.n181 VGND.n180 0.155789
R1649 VGND.n236 VGND.n235 0.155789
R1650 VGND.n281 VGND.n280 0.155789
R1651 VGND.n528 VGND.n527 0.155789
R1652 VGND.n484 VGND.n482 0.155789
R1653 VGND.n1023 VGND.n3 0.149476
R1654 VGND.n1006 VGND.n1003 0.149476
R1655 VGND.n15 VGND.n13 0.149476
R1656 VGND.n80 VGND.n78 0.149476
R1657 VGND.n98 VGND.n95 0.149476
R1658 VGND.n87 VGND.n85 0.149476
R1659 VGND.n606 VGND.n259 0.149476
R1660 VGND.n589 VGND.n586 0.149476
R1661 VGND.n576 VGND.n574 0.149476
R1662 VGND.n512 VGND.n315 0.149476
R1663 VGND.n489 VGND.n487 0.149476
R1664 VGND.n410 VGND.n368 0.149476
R1665 VGND.n431 VGND.n428 0.149476
R1666 VGND.n419 VGND.n417 0.149476
R1667 VGND.n980 VGND.n21 0.149476
R1668 VGND.n991 VGND.n990 0.149476
R1669 VGND.n1026 VGND.n0 0.149476
R1670 VGND.n519 VGND.n518 0.145789
R1671 VGND.n1013 VGND 0.144111
R1672 VGND.n1010 VGND 0.144111
R1673 VGND.n996 VGND 0.144111
R1674 VGND.n105 VGND 0.144111
R1675 VGND.n103 VGND 0.144111
R1676 VGND.n89 VGND 0.144111
R1677 VGND.n596 VGND 0.144111
R1678 VGND.n593 VGND 0.144111
R1679 VGND.n579 VGND 0.144111
R1680 VGND.n537 VGND 0.144111
R1681 VGND.n492 VGND 0.144111
R1682 VGND.n439 VGND 0.144111
R1683 VGND.n436 VGND 0.144111
R1684 VGND.n421 VGND 0.144111
R1685 VGND.n526 VGND.n524 0.140789
R1686 VGND.n481 VGND.n479 0.140789
R1687 VGND.n425 VGND.n420 0.139432
R1688 VGND.n433 VGND.n432 0.139432
R1689 VGND.n443 VGND.n367 0.139432
R1690 VGND.n497 VGND.n490 0.139432
R1691 VGND.n541 VGND.n313 0.139432
R1692 VGND.n583 VGND.n577 0.139432
R1693 VGND.n591 VGND.n590 0.139432
R1694 VGND.n600 VGND.n260 0.139432
R1695 VGND.n92 VGND.n88 0.139432
R1696 VGND.n100 VGND.n99 0.139432
R1697 VGND.n108 VGND.n77 0.139432
R1698 VGND.n1000 VGND.n16 0.139432
R1699 VGND.n1008 VGND.n1007 0.139432
R1700 VGND.n1017 VGND.n4 0.139432
R1701 VGND.n962 VGND.n1 0.139321
R1702 VGND.n15 VGND 0.138786
R1703 VGND.n911 VGND 0.138786
R1704 VGND.n825 VGND 0.138786
R1705 VGND.n54 VGND 0.138786
R1706 VGND.n87 VGND 0.138786
R1707 VGND.n142 VGND 0.138786
R1708 VGND.n678 VGND 0.138786
R1709 VGND.n185 VGND 0.138786
R1710 VGND.n240 VGND 0.138786
R1711 VGND.n576 VGND 0.138786
R1712 VGND.n285 VGND 0.138786
R1713 VGND.n489 VGND 0.138786
R1714 VGND.n419 VGND 0.138786
R1715 VGND.n401 VGND 0.138786
R1716 VGND.n991 VGND 0.138786
R1717 VGND.n521 VGND.n520 0.130789
R1718 VGND.n476 VGND.n318 0.130789
R1719 VGND.n523 VGND.n521 0.125789
R1720 VGND.n478 VGND.n476 0.125789
R1721 VGND.n473 VGND.n470 0.121012
R1722 VGND VGND.n895 0.120789
R1723 VGND VGND.n844 0.120789
R1724 VGND VGND.n34 0.120789
R1725 VGND VGND.n122 0.120789
R1726 VGND.n658 VGND 0.120789
R1727 VGND VGND.n169 0.120789
R1728 VGND VGND.n220 0.120789
R1729 VGND VGND.n269 0.120789
R1730 VGND.n513 VGND 0.120789
R1731 VGND.n963 VGND.n962 0.1205
R1732 VGND.n1017 VGND.n1014 0.1205
R1733 VGND.n1007 VGND.n10 0.1205
R1734 VGND.n1000 VGND.n997 0.1205
R1735 VGND.n108 VGND.n106 0.1205
R1736 VGND.n100 VGND.n83 0.1205
R1737 VGND.n92 VGND.n90 0.1205
R1738 VGND.n600 VGND.n597 0.1205
R1739 VGND.n590 VGND.n571 0.1205
R1740 VGND.n583 VGND.n580 0.1205
R1741 VGND.n541 VGND.n538 0.1205
R1742 VGND.n497 VGND.n493 0.1205
R1743 VGND.n443 VGND.n440 0.1205
R1744 VGND.n433 VGND.n414 0.1205
R1745 VGND.n425 VGND.n422 0.1205
R1746 VGND.n972 VGND.n968 0.1205
R1747 VGND.n988 VGND.n987 0.1205
R1748 VGND.n798 VGND.n797 0.11591
R1749 VGND.n898 VGND.n897 0.115789
R1750 VGND.n842 VGND.n841 0.115789
R1751 VGND.n38 VGND.n37 0.115789
R1752 VGND.n126 VGND.n125 0.115789
R1753 VGND.n662 VGND.n661 0.115789
R1754 VGND.n172 VGND.n171 0.115789
R1755 VGND.n224 VGND.n223 0.115789
R1756 VGND.n272 VGND.n271 0.115789
R1757 VGND.n524 VGND.n523 0.115789
R1758 VGND.n479 VGND.n478 0.115789
R1759 VGND.n766 VGND.n764 0.113
R1760 VGND.n358 VGND.n321 0.113
R1761 VGND VGND.n5 0.111366
R1762 VGND VGND.n1004 0.111366
R1763 VGND VGND.n14 0.111366
R1764 VGND.n910 VGND.n909 0.111366
R1765 VGND.n827 VGND.n824 0.111366
R1766 VGND.n53 VGND.n52 0.111366
R1767 VGND VGND.n79 0.111366
R1768 VGND VGND.n96 0.111366
R1769 VGND VGND.n86 0.111366
R1770 VGND.n141 VGND.n140 0.111366
R1771 VGND.n677 VGND.n676 0.111366
R1772 VGND.n184 VGND.n183 0.111366
R1773 VGND.n239 VGND.n238 0.111366
R1774 VGND VGND.n261 0.111366
R1775 VGND VGND.n587 0.111366
R1776 VGND VGND.n575 0.111366
R1777 VGND.n284 VGND.n283 0.111366
R1778 VGND VGND.n511 0.111366
R1779 VGND VGND.n488 0.111366
R1780 VGND.n350 VGND.n349 0.111366
R1781 VGND VGND.n409 0.111366
R1782 VGND VGND.n429 0.111366
R1783 VGND VGND.n418 0.111366
R1784 VGND VGND.n400 0.111366
R1785 VGND VGND.n393 0.111366
R1786 VGND VGND.n406 0.111366
R1787 VGND.n902 VGND.n901 0.110789
R1788 VGND.n838 VGND.n837 0.110789
R1789 VGND.n43 VGND.n42 0.110789
R1790 VGND.n131 VGND.n130 0.110789
R1791 VGND.n667 VGND.n666 0.110789
R1792 VGND.n176 VGND.n175 0.110789
R1793 VGND.n229 VGND.n228 0.110789
R1794 VGND.n276 VGND.n275 0.110789
R1795 VGND.n520 VGND.n519 0.110789
R1796 VGND.n963 VGND.n959 0.10675
R1797 VGND.n1014 VGND.n1013 0.10675
R1798 VGND.n1010 VGND.n10 0.10675
R1799 VGND.n997 VGND.n996 0.10675
R1800 VGND.n929 VGND.n928 0.10675
R1801 VGND.n914 VGND.n913 0.10675
R1802 VGND.n810 VGND.n809 0.10675
R1803 VGND.n822 VGND.n821 0.10675
R1804 VGND.n860 VGND.n859 0.10675
R1805 VGND.n58 VGND.n57 0.10675
R1806 VGND.n106 VGND.n105 0.10675
R1807 VGND.n103 VGND.n83 0.10675
R1808 VGND.n90 VGND.n89 0.10675
R1809 VGND.n720 VGND.n719 0.10675
R1810 VGND.n146 VGND.n145 0.10675
R1811 VGND.n699 VGND.n698 0.10675
R1812 VGND.n683 VGND.n682 0.10675
R1813 VGND.n203 VGND.n202 0.10675
R1814 VGND.n188 VGND.n187 0.10675
R1815 VGND.n617 VGND.n616 0.10675
R1816 VGND.n244 VGND.n243 0.10675
R1817 VGND.n597 VGND.n596 0.10675
R1818 VGND.n593 VGND.n571 0.10675
R1819 VGND.n580 VGND.n579 0.10675
R1820 VGND.n303 VGND.n302 0.10675
R1821 VGND.n288 VGND.n287 0.10675
R1822 VGND.n538 VGND.n537 0.10675
R1823 VGND.n493 VGND.n492 0.10675
R1824 VGND.n440 VGND.n439 0.10675
R1825 VGND.n436 VGND.n414 0.10675
R1826 VGND.n422 VGND.n421 0.10675
R1827 VGND.n975 VGND.n968 0.10675
R1828 VGND.n987 VGND.n986 0.10675
R1829 VGND.n901 VGND.n900 0.100789
R1830 VGND.n839 VGND.n838 0.100789
R1831 VGND.n42 VGND.n41 0.100789
R1832 VGND.n130 VGND.n129 0.100789
R1833 VGND.n666 VGND.n665 0.100789
R1834 VGND.n175 VGND.n174 0.100789
R1835 VGND.n228 VGND.n227 0.100789
R1836 VGND.n275 VGND.n274 0.100789
R1837 VGND.n527 VGND.n526 0.100789
R1838 VGND.n482 VGND.n481 0.100789
R1839 VGND.n932 VGND.n931 0.1005
R1840 VGND.n812 VGND.n811 0.1005
R1841 VGND.n864 VGND.n863 0.1005
R1842 VGND.n785 VGND.n749 0.1005
R1843 VGND.n724 VGND.n723 0.1005
R1844 VGND.n703 VGND.n702 0.1005
R1845 VGND.n206 VGND.n205 0.1005
R1846 VGND.n621 VGND.n620 0.1005
R1847 VGND.n306 VGND.n305 0.1005
R1848 VGND.n348 VGND.n346 0.1005
R1849 VGND.n347 VGND.n324 0.1005
R1850 VGND.n790 VGND.n789 0.098
R1851 VGND.n892 VGND.n891 0.095789
R1852 VGND.n899 VGND.n898 0.095789
R1853 VGND.n814 VGND.n813 0.095789
R1854 VGND.n841 VGND.n840 0.095789
R1855 VGND.n30 VGND.n28 0.095789
R1856 VGND.n40 VGND.n38 0.095789
R1857 VGND.n118 VGND.n116 0.095789
R1858 VGND.n128 VGND.n126 0.095789
R1859 VGND.n653 VGND.n651 0.095789
R1860 VGND.n664 VGND.n662 0.095789
R1861 VGND.n166 VGND.n165 0.095789
R1862 VGND.n173 VGND.n172 0.095789
R1863 VGND.n216 VGND.n214 0.095789
R1864 VGND.n226 VGND.n224 0.095789
R1865 VGND.n266 VGND.n265 0.095789
R1866 VGND.n273 VGND.n272 0.095789
R1867 VGND.n518 VGND.n516 0.095789
R1868 VGND.n474 VGND.n472 0.095789
R1869 VGND.n768 VGND.n755 0.0955
R1870 VGND.n766 VGND.n765 0.0955
R1871 VGND.n331 VGND.n328 0.0955
R1872 VGND.n794 VGND.n793 0.0885
R1873 VGND.n760 VGND.n759 0.0885
R1874 VGND.n355 VGND.n354 0.0885
R1875 VGND.n353 VGND.n321 0.08675
R1876 VGND.n934 VGND 0.0860682
R1877 VGND.n805 VGND 0.0860682
R1878 VGND.n866 VGND 0.0860682
R1879 VGND.n726 VGND 0.0860682
R1880 VGND.n705 VGND 0.0860682
R1881 VGND.n208 VGND 0.0860682
R1882 VGND.n623 VGND 0.0860682
R1883 VGND.n308 VGND 0.0860682
R1884 VGND.n786 VGND.n784 0.0855
R1885 VGND.n781 VGND.n751 0.0855
R1886 VGND.n472 VGND.n317 0.0855
R1887 VGND.n345 VGND.n343 0.0855
R1888 VGND.n344 VGND.n325 0.0855
R1889 VGND.n470 VGND 0.0810023
R1890 VGND.n896 VGND.n895 0.080789
R1891 VGND.n844 VGND.n843 0.080789
R1892 VGND.n36 VGND.n34 0.080789
R1893 VGND.n124 VGND.n122 0.080789
R1894 VGND.n660 VGND.n658 0.080789
R1895 VGND.n170 VGND.n169 0.080789
R1896 VGND.n222 VGND.n220 0.080789
R1897 VGND.n270 VGND.n269 0.080789
R1898 VGND.n515 VGND.n513 0.080789
R1899 VGND.n918 VGND.n914 0.0805
R1900 VGND.n823 VGND.n822 0.0805
R1901 VGND.n63 VGND.n58 0.0805
R1902 VGND.n772 VGND.n753 0.0805
R1903 VGND.n151 VGND.n146 0.0805
R1904 VGND.n688 VGND.n683 0.0805
R1905 VGND.n192 VGND.n188 0.0805
R1906 VGND.n249 VGND.n244 0.0805
R1907 VGND.n292 VGND.n288 0.0805
R1908 VGND.n334 VGND.n327 0.0805
R1909 VGND.n336 VGND.n335 0.0805
R1910 VGND.n420 VGND.n419 0.0801811
R1911 VGND.n432 VGND.n431 0.0801811
R1912 VGND.n410 VGND.n367 0.0801811
R1913 VGND.n490 VGND.n489 0.0801811
R1914 VGND.n512 VGND.n313 0.0801811
R1915 VGND.n577 VGND.n576 0.0801811
R1916 VGND.n591 VGND.n589 0.0801811
R1917 VGND.n606 VGND.n260 0.0801811
R1918 VGND.n88 VGND.n87 0.0801811
R1919 VGND.n99 VGND.n98 0.0801811
R1920 VGND.n80 VGND.n77 0.0801811
R1921 VGND.n16 VGND.n15 0.0801811
R1922 VGND.n1008 VGND.n1006 0.0801811
R1923 VGND.n1023 VGND.n4 0.0801811
R1924 VGND.n1026 VGND.n1 0.0793031
R1925 VGND.n792 VGND.n791 0.073
R1926 VGND.n782 VGND.n780 0.0705
R1927 VGND.n777 VGND.n753 0.0705
R1928 VGND.n342 VGND.n340 0.0705
R1929 VGND.n341 VGND.n326 0.0705
R1930 VGND.n776 VGND.n751 0.0655
R1931 VGND.n774 VGND.n773 0.0655
R1932 VGND.n337 VGND.n326 0.0655
R1933 VGND.n339 VGND.n338 0.0655
R1934 VGND.n893 VGND.n892 0.063
R1935 VGND.n815 VGND.n814 0.063
R1936 VGND.n31 VGND.n30 0.063
R1937 VGND.n798 VGND.n741 0.063
R1938 VGND.n794 VGND.n742 0.063
R1939 VGND.n119 VGND.n118 0.063
R1940 VGND.n654 VGND.n653 0.063
R1941 VGND.n167 VGND.n166 0.063
R1942 VGND.n217 VGND.n216 0.063
R1943 VGND.n267 VGND.n266 0.063
R1944 VGND.n355 VGND.n322 0.063
R1945 VGND.n932 VGND.n891 0.060789
R1946 VGND.n919 VGND.n906 0.060789
R1947 VGND.n813 VGND.n812 0.060789
R1948 VGND.n831 VGND.n830 0.060789
R1949 VGND.n864 VGND.n28 0.060789
R1950 VGND.n64 VGND.n49 0.060789
R1951 VGND.n724 VGND.n116 0.060789
R1952 VGND.n152 VGND.n137 0.060789
R1953 VGND.n703 VGND.n651 0.060789
R1954 VGND.n689 VGND.n673 0.060789
R1955 VGND.n206 VGND.n165 0.060789
R1956 VGND.n193 VGND.n180 0.060789
R1957 VGND.n621 VGND.n214 0.060789
R1958 VGND.n250 VGND.n235 0.060789
R1959 VGND.n306 VGND.n265 0.060789
R1960 VGND.n293 VGND.n280 0.060789
R1961 VGND.n399 VGND.n370 0.060789
R1962 VGND.n392 VGND.n391 0.060789
R1963 VGND.n378 VGND.n369 0.060789
R1964 VGND.n972 VGND.n20 0.060789
R1965 VGND.n989 VGND.n988 0.060789
R1966 VGND VGND.n904 0.0605
R1967 VGND.n912 VGND 0.0605
R1968 VGND.n835 VGND 0.0605
R1969 VGND VGND.n826 0.0605
R1970 VGND VGND.n45 0.0605
R1971 VGND.n55 VGND 0.0605
R1972 VGND VGND.n742 0.0605
R1973 VGND.n790 VGND 0.0605
R1974 VGND.n747 VGND 0.0605
R1975 VGND.n770 VGND 0.0605
R1976 VGND.n762 VGND 0.0605
R1977 VGND VGND.n133 0.0605
R1978 VGND.n143 VGND 0.0605
R1979 VGND VGND.n669 0.0605
R1980 VGND.n679 VGND 0.0605
R1981 VGND VGND.n178 0.0605
R1982 VGND.n186 VGND 0.0605
R1983 VGND VGND.n231 0.0605
R1984 VGND.n241 VGND 0.0605
R1985 VGND VGND.n278 0.0605
R1986 VGND.n286 VGND 0.0605
R1987 VGND VGND.n529 0.0605
R1988 VGND.n530 VGND 0.0605
R1989 VGND.n530 VGND 0.0605
R1990 VGND.n508 VGND.n317 0.0605
R1991 VGND.n508 VGND.n507 0.0605
R1992 VGND VGND.n485 0.0605
R1993 VGND.n359 VGND 0.0605
R1994 VGND.n352 VGND 0.0605
R1995 VGND VGND.n323 0.0605
R1996 VGND.n333 VGND 0.0605
R1997 VGND VGND.n329 0.0605
R1998 VGND.n330 VGND 0.0605
R1999 VGND.n330 VGND 0.0605
R2000 VGND.n910 VGND.n908 0.058
R2001 VGND.n828 VGND.n827 0.058
R2002 VGND.n53 VGND.n51 0.058
R2003 VGND.n795 VGND.n794 0.058
R2004 VGND.n760 VGND.n758 0.058
R2005 VGND.n141 VGND.n139 0.058
R2006 VGND.n677 VGND.n675 0.058
R2007 VGND.n184 VGND.n182 0.058
R2008 VGND.n239 VGND.n237 0.058
R2009 VGND.n284 VGND.n282 0.058
R2010 VGND.n356 VGND.n355 0.058
R2011 VGND.n350 VGND.n322 0.058
R2012 VGND.n778 VGND.n776 0.0555
R2013 VGND.n773 VGND.n755 0.0555
R2014 VGND.n339 VGND.n337 0.0555
R2015 VGND.n338 VGND.n327 0.0555
R2016 VGND.n799 VGND.n798 0.0505
R2017 VGND.n780 VGND.n749 0.0505
R2018 VGND.n778 VGND.n777 0.0505
R2019 VGND.n507 VGND.n318 0.0505
R2020 VGND.n340 VGND.n325 0.0505
R2021 VGND.n342 VGND.n341 0.0505
R2022 VGND VGND.n357 0.04675
R2023 VGND.n897 VGND.n896 0.0455
R2024 VGND.n900 VGND.n899 0.0455
R2025 VGND.n903 VGND.n902 0.0455
R2026 VGND.n843 VGND.n842 0.0455
R2027 VGND.n840 VGND.n839 0.0455
R2028 VGND.n837 VGND.n836 0.0455
R2029 VGND.n37 VGND.n36 0.0455
R2030 VGND.n41 VGND.n40 0.0455
R2031 VGND.n44 VGND.n43 0.0455
R2032 VGND.n125 VGND.n124 0.0455
R2033 VGND.n129 VGND.n128 0.0455
R2034 VGND.n132 VGND.n131 0.0455
R2035 VGND.n661 VGND.n660 0.0455
R2036 VGND.n665 VGND.n664 0.0455
R2037 VGND.n668 VGND.n667 0.0455
R2038 VGND.n171 VGND.n170 0.0455
R2039 VGND.n174 VGND.n173 0.0455
R2040 VGND.n177 VGND.n176 0.0455
R2041 VGND.n223 VGND.n222 0.0455
R2042 VGND.n227 VGND.n226 0.0455
R2043 VGND.n230 VGND.n229 0.0455
R2044 VGND.n271 VGND.n270 0.0455
R2045 VGND.n274 VGND.n273 0.0455
R2046 VGND.n277 VGND.n276 0.0455
R2047 VGND.n1023 VGND 0.04425
R2048 VGND.n1006 VGND 0.04425
R2049 VGND.n911 VGND 0.04425
R2050 VGND.n825 VGND 0.04425
R2051 VGND.n54 VGND 0.04425
R2052 VGND VGND.n74 0.04425
R2053 VGND VGND.n80 0.04425
R2054 VGND.n98 VGND 0.04425
R2055 VGND.n142 VGND 0.04425
R2056 VGND.n678 VGND 0.04425
R2057 VGND.n185 VGND 0.04425
R2058 VGND.n240 VGND 0.04425
R2059 VGND.n606 VGND 0.04425
R2060 VGND.n589 VGND 0.04425
R2061 VGND.n285 VGND 0.04425
R2062 VGND VGND.n512 0.04425
R2063 VGND.n351 VGND 0.04425
R2064 VGND.n351 VGND 0.04425
R2065 VGND VGND.n410 0.04425
R2066 VGND.n431 VGND 0.04425
R2067 VGND VGND.n394 0.04425
R2068 VGND.n407 VGND 0.04425
R2069 VGND.n1026 VGND 0.04425
R2070 VGND VGND.n980 0.04425
R2071 VGND VGND.n1022 0.04175
R2072 VGND VGND.n1005 0.04175
R2073 VGND.n915 VGND 0.04175
R2074 VGND VGND.n834 0.04175
R2075 VGND.n60 VGND 0.04175
R2076 VGND.n81 VGND 0.04175
R2077 VGND VGND.n97 0.04175
R2078 VGND.n148 VGND 0.04175
R2079 VGND.n685 VGND 0.04175
R2080 VGND.n189 VGND 0.04175
R2081 VGND.n246 VGND 0.04175
R2082 VGND VGND.n605 0.04175
R2083 VGND VGND.n588 0.04175
R2084 VGND.n289 VGND 0.04175
R2085 VGND.n495 VGND 0.04175
R2086 VGND.n411 VGND 0.04175
R2087 VGND VGND.n430 0.04175
R2088 VGND.n395 VGND 0.04175
R2089 VGND.n376 VGND 0.04175
R2090 VGND.n965 VGND 0.04175
R2091 VGND.n981 VGND 0.04175
R2092 VGND.n919 VGND.n918 0.0405
R2093 VGND.n831 VGND.n823 0.0405
R2094 VGND.n64 VGND.n63 0.0405
R2095 VGND.n774 VGND.n772 0.0405
R2096 VGND.n769 VGND.n757 0.0405
R2097 VGND.n152 VGND.n151 0.0405
R2098 VGND.n689 VGND.n688 0.0405
R2099 VGND.n193 VGND.n192 0.0405
R2100 VGND.n250 VGND.n249 0.0405
R2101 VGND.n293 VGND.n292 0.0405
R2102 VGND.n336 VGND.n334 0.0405
R2103 VGND.n335 VGND.n328 0.0405
R2104 VGND.n1023 VGND 0.0386102
R2105 VGND.n1006 VGND 0.0386102
R2106 VGND.n15 VGND 0.0386102
R2107 VGND.n80 VGND 0.0386102
R2108 VGND.n98 VGND 0.0386102
R2109 VGND.n87 VGND 0.0386102
R2110 VGND.n606 VGND 0.0386102
R2111 VGND.n589 VGND 0.0386102
R2112 VGND.n576 VGND 0.0386102
R2113 VGND.n512 VGND 0.0386102
R2114 VGND.n489 VGND 0.0386102
R2115 VGND.n410 VGND 0.0386102
R2116 VGND.n431 VGND 0.0386102
R2117 VGND.n419 VGND 0.0386102
R2118 VGND.n401 VGND 0.0386102
R2119 VGND.n394 VGND 0.0386102
R2120 VGND.n407 VGND 0.0386102
R2121 VGND.n980 VGND 0.0386102
R2122 VGND.n991 VGND 0.0386102
R2123 VGND VGND.n1026 0.0386102
R2124 VGND.n784 VGND.n747 0.0355
R2125 VGND.n782 VGND.n781 0.0355
R2126 VGND.n343 VGND.n324 0.0355
R2127 VGND.n345 VGND.n344 0.0355
R2128 VGND VGND.n332 0.0355
R2129 VGND.n926 VGND.n925 0.03425
R2130 VGND.n846 VGND.n845 0.03425
R2131 VGND.n855 VGND.n854 0.03425
R2132 VGND.n795 VGND.n792 0.03425
R2133 VGND.n715 VGND.n714 0.03425
R2134 VGND.n657 VGND.n162 0.03425
R2135 VGND.n200 VGND.n199 0.03425
R2136 VGND.n612 VGND.n611 0.03425
R2137 VGND.n300 VGND.n299 0.03425
R2138 VGND.n356 VGND.n353 0.03425
R2139 VGND.n407 VGND.n405 0.0333762
R2140 VGND.n394 VGND.n375 0.0333762
R2141 VGND.n402 VGND.n401 0.0333762
R2142 VGND.n761 VGND 0.033
R2143 VGND.n961 VGND.n960 0.0327727
R2144 VGND.n361 VGND.n360 0.0327727
R2145 VGND.n382 VGND.n381 0.0327727
R2146 VGND.n398 VGND.n397 0.0327727
R2147 VGND.n390 VGND.n389 0.0327727
R2148 VGND.n974 VGND.n973 0.0327727
R2149 VGND.n984 VGND.n983 0.0327727
R2150 VGND.n762 VGND.n761 0.028
R2151 VGND.n446 VGND.n423 0.0258175
R2152 VGND.n446 VGND.n413 0.0258175
R2153 VGND.n446 VGND.n441 0.0258175
R2154 VGND.n506 VGND.n494 0.0258175
R2155 VGND.n506 VGND.n483 0.0258175
R2156 VGND.n544 VGND.n314 0.0258175
R2157 VGND.n544 VGND.n539 0.0258175
R2158 VGND.n603 VGND.n581 0.0258175
R2159 VGND.n603 VGND.n570 0.0258175
R2160 VGND.n603 VGND.n598 0.0258175
R2161 VGND.n732 VGND.n111 0.0258175
R2162 VGND.n734 VGND.n111 0.0258175
R2163 VGND.n736 VGND.n111 0.0258175
R2164 VGND.n800 VGND.n796 0.0258175
R2165 VGND.n1020 VGND.n998 0.0258175
R2166 VGND.n1020 VGND.n9 0.0258175
R2167 VGND.n1020 VGND.n1015 0.0258175
R2168 VGND.n904 VGND.n903 0.0255
R2169 VGND.n908 VGND.n907 0.0255
R2170 VGND.n836 VGND.n835 0.0255
R2171 VGND.n829 VGND.n828 0.0255
R2172 VGND.n45 VGND.n44 0.0255
R2173 VGND.n51 VGND.n50 0.0255
R2174 VGND.n770 VGND.n768 0.0255
R2175 VGND.n765 VGND.n758 0.0255
R2176 VGND.n133 VGND.n132 0.0255
R2177 VGND.n139 VGND.n138 0.0255
R2178 VGND.n669 VGND.n668 0.0255
R2179 VGND.n675 VGND.n674 0.0255
R2180 VGND.n178 VGND.n177 0.0255
R2181 VGND.n182 VGND.n181 0.0255
R2182 VGND.n231 VGND.n230 0.0255
R2183 VGND.n237 VGND.n236 0.0255
R2184 VGND.n278 VGND.n277 0.0255
R2185 VGND.n282 VGND.n281 0.0255
R2186 VGND.n529 VGND.n528 0.0255
R2187 VGND.n485 VGND.n484 0.0255
R2188 VGND.n333 VGND.n331 0.0255
R2189 VGND.n332 VGND.n329 0.0255
R2190 VGND.n931 VGND.n929 0.0205
R2191 VGND.n811 VGND.n810 0.0205
R2192 VGND.n863 VGND.n860 0.0205
R2193 VGND.n786 VGND.n785 0.0205
R2194 VGND VGND.n769 0.0205
R2195 VGND.n723 VGND.n720 0.0205
R2196 VGND.n702 VGND.n699 0.0205
R2197 VGND.n205 VGND.n203 0.0205
R2198 VGND.n620 VGND.n617 0.0205
R2199 VGND.n305 VGND.n303 0.0205
R2200 VGND.n346 VGND.n323 0.0205
R2201 VGND.n348 VGND.n347 0.0205
R2202 VGND.n1018 VGND.n1016 0.0202222
R2203 VGND.n1009 VGND.n6 0.0202222
R2204 VGND.n1001 VGND.n999 0.0202222
R2205 VGND.n109 VGND.n107 0.0202222
R2206 VGND.n102 VGND.n101 0.0202222
R2207 VGND.n93 VGND.n91 0.0202222
R2208 VGND.n601 VGND.n599 0.0202222
R2209 VGND.n592 VGND.n262 0.0202222
R2210 VGND.n584 VGND.n582 0.0202222
R2211 VGND.n542 VGND.n540 0.0202222
R2212 VGND.n498 VGND.n496 0.0202222
R2213 VGND.n444 VGND.n442 0.0202222
R2214 VGND.n435 VGND.n434 0.0202222
R2215 VGND.n426 VGND.n424 0.0202222
R2216 VGND.n920 VGND.n917 0.0191364
R2217 VGND.n832 VGND.n818 0.0191364
R2218 VGND.n65 VGND.n62 0.0191364
R2219 VGND.n153 VGND.n150 0.0191364
R2220 VGND.n690 VGND.n687 0.0191364
R2221 VGND.n194 VGND.n191 0.0191364
R2222 VGND.n251 VGND.n248 0.0191364
R2223 VGND.n294 VGND.n291 0.0191364
R2224 VGND.n933 VGND 0.0173182
R2225 VGND.n923 VGND.n922 0.0173182
R2226 VGND VGND.n806 0.0173182
R2227 VGND.n849 VGND.n817 0.0173182
R2228 VGND.n865 VGND 0.0173182
R2229 VGND.n852 VGND.n71 0.0173182
R2230 VGND.n725 VGND 0.0173182
R2231 VGND.n712 VGND.n159 0.0173182
R2232 VGND.n704 VGND 0.0173182
R2233 VGND.n709 VGND.n161 0.0173182
R2234 VGND.n207 VGND 0.0173182
R2235 VGND.n197 VGND.n196 0.0173182
R2236 VGND.n622 VGND 0.0173182
R2237 VGND.n609 VGND.n257 0.0173182
R2238 VGND.n307 VGND 0.0173182
R2239 VGND.n297 VGND.n296 0.0173182
R2240 VGND.n357 VGND 0.0173182
R2241 VGND.n912 VGND.n911 0.01675
R2242 VGND.n826 VGND.n825 0.01675
R2243 VGND.n55 VGND.n54 0.01675
R2244 VGND.n143 VGND.n142 0.01675
R2245 VGND.n679 VGND.n678 0.01675
R2246 VGND.n186 VGND.n185 0.01675
R2247 VGND.n241 VGND.n240 0.01675
R2248 VGND.n286 VGND.n285 0.01675
R2249 VGND.n352 VGND.n351 0.01675
R2250 VGND.n924 VGND.n923 0.0164091
R2251 VGND.n926 VGND 0.0164091
R2252 VGND.n849 VGND.n848 0.0164091
R2253 VGND.n846 VGND 0.0164091
R2254 VGND.n853 VGND.n852 0.0164091
R2255 VGND.n855 VGND 0.0164091
R2256 VGND.n803 VGND.n802 0.0164091
R2257 VGND.n74 VGND 0.0164091
R2258 VGND.n713 VGND.n712 0.0164091
R2259 VGND.n715 VGND 0.0164091
R2260 VGND.n709 VGND.n708 0.0164091
R2261 VGND.n162 VGND 0.0164091
R2262 VGND.n198 VGND.n197 0.0164091
R2263 VGND.n200 VGND 0.0164091
R2264 VGND.n610 VGND.n609 0.0164091
R2265 VGND.n612 VGND 0.0164091
R2266 VGND.n298 VGND.n297 0.0164091
R2267 VGND.n300 VGND 0.0164091
R2268 VGND VGND.n930 0.0159545
R2269 VGND.n807 VGND 0.0159545
R2270 VGND VGND.n862 0.0159545
R2271 VGND VGND.n722 0.0159545
R2272 VGND VGND.n701 0.0159545
R2273 VGND VGND.n204 0.0159545
R2274 VGND VGND.n619 0.0159545
R2275 VGND VGND.n304 0.0159545
R2276 VGND.n803 VGND.n73 0.0150455
R2277 VGND.n791 VGND.n741 0.01425
R2278 VGND.n917 VGND.n916 0.0141364
R2279 VGND.n819 VGND.n818 0.0141364
R2280 VGND.n62 VGND.n61 0.0141364
R2281 VGND.n150 VGND.n149 0.0141364
R2282 VGND.n687 VGND.n686 0.0141364
R2283 VGND.n191 VGND.n190 0.0141364
R2284 VGND.n248 VGND.n247 0.0141364
R2285 VGND.n291 VGND.n290 0.0141364
R2286 VGND.n925 VGND 0.0105
R2287 VGND.n845 VGND 0.0105
R2288 VGND.n854 VGND 0.0105
R2289 VGND.n714 VGND 0.0105
R2290 VGND VGND.n657 0.0105
R2291 VGND.n199 VGND 0.0105
R2292 VGND.n611 VGND 0.0105
R2293 VGND.n299 VGND 0.0105
R2294 VGND.n404 VGND.n385 0.00990704
R2295 VGND.n404 VGND.n374 0.00990704
R2296 VGND.n404 VGND.n403 0.00990704
R2297 VGND.n969 VGND.n19 0.00990704
R2298 VGND.n970 VGND.n19 0.00990704
R2299 VGND.n978 VGND.n967 0.00990704
R2300 VGND.n978 VGND.n964 0.00990704
R2301 VGND.n1025 VGND 0.0093
R2302 VGND.n894 VGND.n893 0.00868182
R2303 VGND.n816 VGND.n815 0.00868182
R2304 VGND.n32 VGND.n31 0.00868182
R2305 VGND.n789 VGND.n745 0.00868182
R2306 VGND.n120 VGND.n119 0.00868182
R2307 VGND.n655 VGND.n654 0.00868182
R2308 VGND.n168 VGND.n167 0.00868182
R2309 VGND.n218 VGND.n217 0.00868182
R2310 VGND.n268 VGND.n267 0.00868182
R2311 VGND.n764 VGND.n757 0.008
R2312 VGND.n359 VGND.n358 0.008
R2313 VGND.n921 VGND.n915 0.00731818
R2314 VGND.n834 VGND.n833 0.00731818
R2315 VGND.n66 VGND.n60 0.00731818
R2316 VGND.n154 VGND.n148 0.00731818
R2317 VGND.n691 VGND.n685 0.00731818
R2318 VGND.n195 VGND.n189 0.00731818
R2319 VGND.n252 VGND.n246 0.00731818
R2320 VGND.n295 VGND.n289 0.00731818
R2321 VGND.n396 VGND.n395 0.00731818
R2322 VGND.n377 VGND.n376 0.00731818
R2323 VGND.n966 VGND.n965 0.00731818
R2324 VGND.n982 VGND.n981 0.00731818
R2325 VGND.n960 VGND.n958 0.00686364
R2326 VGND.n930 VGND.n890 0.00686364
R2327 VGND.n916 VGND.n905 0.00686364
R2328 VGND.n808 VGND.n807 0.00686364
R2329 VGND.n820 VGND.n819 0.00686364
R2330 VGND.n862 VGND.n26 0.00686364
R2331 VGND.n61 VGND.n47 0.00686364
R2332 VGND.n722 VGND.n114 0.00686364
R2333 VGND.n149 VGND.n135 0.00686364
R2334 VGND.n701 VGND.n649 0.00686364
R2335 VGND.n686 VGND.n671 0.00686364
R2336 VGND.n204 VGND.n164 0.00686364
R2337 VGND.n190 VGND.n179 0.00686364
R2338 VGND.n619 VGND.n212 0.00686364
R2339 VGND.n247 VGND.n233 0.00686364
R2340 VGND.n304 VGND.n264 0.00686364
R2341 VGND.n290 VGND.n279 0.00686364
R2342 VGND.n360 VGND.n320 0.00686364
R2343 VGND.n381 VGND.n380 0.00686364
R2344 VGND.n397 VGND.n373 0.00686364
R2345 VGND.n389 VGND.n386 0.00686364
R2346 VGND.n976 VGND.n974 0.00686364
R2347 VGND.n985 VGND.n984 0.00686364
R2348 VGND.n927 VGND.n924 0.00640909
R2349 VGND.n927 VGND.n926 0.00640909
R2350 VGND.n848 VGND.n847 0.00640909
R2351 VGND.n847 VGND.n846 0.00640909
R2352 VGND.n856 VGND.n853 0.00640909
R2353 VGND.n856 VGND.n855 0.00640909
R2354 VGND.n802 VGND.n801 0.00640909
R2355 VGND.n801 VGND.n74 0.00640909
R2356 VGND.n716 VGND.n713 0.00640909
R2357 VGND.n716 VGND.n715 0.00640909
R2358 VGND.n708 VGND.n707 0.00640909
R2359 VGND.n707 VGND.n162 0.00640909
R2360 VGND.n201 VGND.n198 0.00640909
R2361 VGND.n201 VGND.n200 0.00640909
R2362 VGND.n613 VGND.n610 0.00640909
R2363 VGND.n613 VGND.n612 0.00640909
R2364 VGND.n301 VGND.n298 0.00640909
R2365 VGND.n301 VGND.n300 0.00640909
R2366 VGND.n961 VGND.n957 0.0055
R2367 VGND.n959 VGND.n958 0.0055
R2368 VGND.n934 VGND.n933 0.0055
R2369 VGND.n928 VGND.n890 0.0055
R2370 VGND.n922 VGND.n894 0.0055
R2371 VGND.n921 VGND.n920 0.0055
R2372 VGND.n913 VGND.n905 0.0055
R2373 VGND.n806 VGND.n805 0.0055
R2374 VGND.n809 VGND.n808 0.0055
R2375 VGND.n817 VGND.n816 0.0055
R2376 VGND.n833 VGND.n832 0.0055
R2377 VGND.n821 VGND.n820 0.0055
R2378 VGND.n866 VGND.n865 0.0055
R2379 VGND.n859 VGND.n26 0.0055
R2380 VGND.n71 VGND.n32 0.0055
R2381 VGND.n66 VGND.n65 0.0055
R2382 VGND.n57 VGND.n47 0.0055
R2383 VGND.n745 VGND.n744 0.0055
R2384 VGND.n726 VGND.n725 0.0055
R2385 VGND.n719 VGND.n114 0.0055
R2386 VGND.n159 VGND.n120 0.0055
R2387 VGND.n154 VGND.n153 0.0055
R2388 VGND.n145 VGND.n135 0.0055
R2389 VGND.n705 VGND.n704 0.0055
R2390 VGND.n698 VGND.n649 0.0055
R2391 VGND.n655 VGND.n161 0.0055
R2392 VGND.n691 VGND.n690 0.0055
R2393 VGND.n682 VGND.n671 0.0055
R2394 VGND.n208 VGND.n207 0.0055
R2395 VGND.n202 VGND.n164 0.0055
R2396 VGND.n196 VGND.n168 0.0055
R2397 VGND.n195 VGND.n194 0.0055
R2398 VGND.n187 VGND.n179 0.0055
R2399 VGND.n623 VGND.n622 0.0055
R2400 VGND.n616 VGND.n212 0.0055
R2401 VGND.n257 VGND.n218 0.0055
R2402 VGND.n252 VGND.n251 0.0055
R2403 VGND.n243 VGND.n233 0.0055
R2404 VGND.n308 VGND.n307 0.0055
R2405 VGND.n302 VGND.n264 0.0055
R2406 VGND.n296 VGND.n268 0.0055
R2407 VGND.n295 VGND.n294 0.0055
R2408 VGND.n287 VGND.n279 0.0055
R2409 VGND.n362 VGND.n361 0.0055
R2410 VGND.n357 VGND.n320 0.0055
R2411 VGND.n383 VGND.n382 0.0055
R2412 VGND.n380 VGND.n379 0.0055
R2413 VGND.n398 VGND.n396 0.0055
R2414 VGND.n373 VGND.n372 0.0055
R2415 VGND.n390 VGND.n377 0.0055
R2416 VGND.n388 VGND.n386 0.0055
R2417 VGND.n973 VGND.n966 0.0055
R2418 VGND.n976 VGND.n975 0.0055
R2419 VGND.n983 VGND.n982 0.0055
R2420 VGND.n986 VGND.n985 0.0055
R2421 VGND.n1022 VGND.n1021 0.00466667
R2422 VGND.n1005 VGND.n1002 0.00466667
R2423 VGND.n82 VGND.n81 0.00466667
R2424 VGND.n97 VGND.n94 0.00466667
R2425 VGND.n605 VGND.n604 0.00466667
R2426 VGND.n588 VGND.n585 0.00466667
R2427 VGND.n499 VGND.n495 0.00466667
R2428 VGND.n412 VGND.n411 0.00466667
R2429 VGND.n430 VGND.n427 0.00466667
R2430 VGND.n1016 VGND.n8 0.00438889
R2431 VGND.n1011 VGND.n1009 0.00438889
R2432 VGND.n999 VGND.n12 0.00438889
R2433 VGND.n107 VGND.n76 0.00438889
R2434 VGND.n104 VGND.n102 0.00438889
R2435 VGND.n91 VGND.n84 0.00438889
R2436 VGND.n599 VGND.n569 0.00438889
R2437 VGND.n594 VGND.n592 0.00438889
R2438 VGND.n582 VGND.n573 0.00438889
R2439 VGND.n540 VGND.n312 0.00438889
R2440 VGND.n496 VGND.n486 0.00438889
R2441 VGND.n442 VGND.n366 0.00438889
R2442 VGND.n437 VGND.n435 0.00438889
R2443 VGND.n424 VGND.n416 0.00438889
R2444 VGND.n1019 VGND.n1018 0.00355556
R2445 VGND.n1013 VGND.n8 0.00355556
R2446 VGND.n1021 VGND.n6 0.00355556
R2447 VGND.n1011 VGND.n1010 0.00355556
R2448 VGND.n1002 VGND.n1001 0.00355556
R2449 VGND.n996 VGND.n12 0.00355556
R2450 VGND.n110 VGND.n109 0.00355556
R2451 VGND.n105 VGND.n76 0.00355556
R2452 VGND.n101 VGND.n82 0.00355556
R2453 VGND.n104 VGND.n103 0.00355556
R2454 VGND.n94 VGND.n93 0.00355556
R2455 VGND.n89 VGND.n84 0.00355556
R2456 VGND.n602 VGND.n601 0.00355556
R2457 VGND.n596 VGND.n569 0.00355556
R2458 VGND.n604 VGND.n262 0.00355556
R2459 VGND.n594 VGND.n593 0.00355556
R2460 VGND.n585 VGND.n584 0.00355556
R2461 VGND.n579 VGND.n573 0.00355556
R2462 VGND.n543 VGND.n542 0.00355556
R2463 VGND.n537 VGND.n312 0.00355556
R2464 VGND.n499 VGND.n498 0.00355556
R2465 VGND.n492 VGND.n486 0.00355556
R2466 VGND.n445 VGND.n444 0.00355556
R2467 VGND.n439 VGND.n366 0.00355556
R2468 VGND.n434 VGND.n412 0.00355556
R2469 VGND.n437 VGND.n436 0.00355556
R2470 VGND.n427 VGND.n426 0.00355556
R2471 VGND.n421 VGND.n416 0.00355556
R2472 VGND VGND.n910 0.003
R2473 VGND.n827 VGND 0.003
R2474 VGND VGND.n53 0.003
R2475 VGND VGND.n760 0.003
R2476 VGND VGND.n141 0.003
R2477 VGND VGND.n677 0.003
R2478 VGND VGND.n184 0.003
R2479 VGND VGND.n239 0.003
R2480 VGND VGND.n284 0.003
R2481 VGND VGND.n350 0.003
R2482 VGND.n744 VGND.n73 0.00277273
R2483 VGND.n446 VGND.n415 0.00194928
R2484 VGND.n446 VGND.n438 0.00194928
R2485 VGND.n603 VGND.n572 0.00194928
R2486 VGND.n603 VGND.n595 0.00194928
R2487 VGND.n733 VGND.n111 0.00194928
R2488 VGND.n735 VGND.n111 0.00194928
R2489 VGND.n1020 VGND.n11 0.00194928
R2490 VGND.n1020 VGND.n1012 0.00194928
R2491 VGND.n404 VGND.n387 0.00121524
R2492 VGND.n404 VGND.n371 0.00121524
R2493 VGND.n978 VGND.n977 0.00120406
R2494 VGND.n979 VGND.n978 0.001
R2495 VGND.n992 VGND.n19 0.001
R2496 VGND.n979 VGND.n19 0.001
R2497 b[5].n9 b[5] 10.8542
R2498 b[5].n7 b[5].t3 8.56366
R2499 b[5].n0 b[5].t2 8.52233
R2500 b[5].n2 b[5].t4 8.5005
R2501 b[5].n5 b[5].t1 8.5005
R2502 b[5].n8 b[5].t0 6.31291
R2503 b[5].n8 b[5].t6 5.79041
R2504 b[5].n11 b[5].t7 5.79041
R2505 b[5].n9 b[5].t5 5.60428
R2506 b[5].n1 b[5] 1.48874
R2507 b[5].n4 b[5] 0.828735
R2508 b[5].n11 b[5].n10 0.523
R2509 b[5].n10 b[5].n8 0.523
R2510 b[5].n0 b[5] 0.514393
R2511 b[5].n1 b[5].n0 0.492265
R2512 b[5].n4 b[5].n3 0.492265
R2513 b[5].n7 b[5].n6 0.492265
R2514 b[5] b[5].n11 0.360115
R2515 b[5].n3 b[5] 0.3405
R2516 b[5].n10 b[5].n9 0.186974
R2517 b[5].n6 b[5] 0.171798
R2518 b[5].n7 b[5] 0.168735
R2519 b[5] b[5].n7 0.0364615
R2520 b[5].n5 b[5].n4 0.0223321
R2521 b[5].n6 b[5].n5 0.0223321
R2522 b[5].n2 b[5].n1 0.0221667
R2523 b[5].n3 b[5].n2 0.0221667
R2524 VPWR.n169 VPWR.n140 17.0117
R2525 VPWR.n206 VPWR.n177 17.0117
R2526 VPWR.n282 VPWR.n252 17.0117
R2527 VPWR.n395 VPWR.n365 17.0117
R2528 VPWR.n545 VPWR.n516 17.0117
R2529 VPWR.n51 VPWR.n45 17.0005
R2530 VPWR.n51 VPWR.n44 17.0005
R2531 VPWR.n51 VPWR.n36 17.0005
R2532 VPWR.n51 VPWR.n35 17.0005
R2533 VPWR.n51 VPWR.n27 17.0005
R2534 VPWR.n52 VPWR.n51 17.0005
R2535 VPWR.n51 VPWR.n25 17.0005
R2536 VPWR.n87 VPWR.n81 17.0005
R2537 VPWR.n87 VPWR.n80 17.0005
R2538 VPWR.n87 VPWR.n69 17.0005
R2539 VPWR.n87 VPWR.n68 17.0005
R2540 VPWR.n87 VPWR.n66 17.0005
R2541 VPWR.n87 VPWR.n65 17.0005
R2542 VPWR.n87 VPWR.n64 17.0005
R2543 VPWR.n87 VPWR.n56 17.0005
R2544 VPWR.n88 VPWR.n87 17.0005
R2545 VPWR.n87 VPWR.n54 17.0005
R2546 VPWR.n133 VPWR.n97 17.0005
R2547 VPWR.n133 VPWR.n103 17.0005
R2548 VPWR.n133 VPWR.n126 17.0005
R2549 VPWR.n133 VPWR.n124 17.0005
R2550 VPWR.n133 VPWR.n123 17.0005
R2551 VPWR.n133 VPWR.n121 17.0005
R2552 VPWR.n133 VPWR.n119 17.0005
R2553 VPWR.n133 VPWR.n117 17.0005
R2554 VPWR.n133 VPWR.n115 17.0005
R2555 VPWR.n133 VPWR.n113 17.0005
R2556 VPWR.n133 VPWR.n111 17.0005
R2557 VPWR.n133 VPWR.n109 17.0005
R2558 VPWR.n133 VPWR.n107 17.0005
R2559 VPWR.n133 VPWR.n106 17.0005
R2560 VPWR.n133 VPWR.n95 17.0005
R2561 VPWR.n133 VPWR.n94 17.0005
R2562 VPWR.n134 VPWR.n133 17.0005
R2563 VPWR.n133 VPWR.n92 17.0005
R2564 VPWR.n133 VPWR.n132 17.0005
R2565 VPWR.n169 VPWR.n163 17.0005
R2566 VPWR.n169 VPWR.n162 17.0005
R2567 VPWR.n169 VPWR.n151 17.0005
R2568 VPWR.n169 VPWR.n149 17.0005
R2569 VPWR.n169 VPWR.n147 17.0005
R2570 VPWR.n169 VPWR.n145 17.0005
R2571 VPWR.n169 VPWR.n139 17.0005
R2572 VPWR.n170 VPWR.n169 17.0005
R2573 VPWR.n169 VPWR.n137 17.0005
R2574 VPWR.n206 VPWR.n200 17.0005
R2575 VPWR.n206 VPWR.n199 17.0005
R2576 VPWR.n206 VPWR.n188 17.0005
R2577 VPWR.n206 VPWR.n186 17.0005
R2578 VPWR.n206 VPWR.n184 17.0005
R2579 VPWR.n206 VPWR.n182 17.0005
R2580 VPWR.n206 VPWR.n176 17.0005
R2581 VPWR.n207 VPWR.n206 17.0005
R2582 VPWR.n206 VPWR.n174 17.0005
R2583 VPWR.n244 VPWR.n238 17.0005
R2584 VPWR.n244 VPWR.n237 17.0005
R2585 VPWR.n244 VPWR.n226 17.0005
R2586 VPWR.n244 VPWR.n225 17.0005
R2587 VPWR.n244 VPWR.n223 17.0005
R2588 VPWR.n244 VPWR.n222 17.0005
R2589 VPWR.n244 VPWR.n221 17.0005
R2590 VPWR.n244 VPWR.n213 17.0005
R2591 VPWR.n245 VPWR.n244 17.0005
R2592 VPWR.n244 VPWR.n211 17.0005
R2593 VPWR.n282 VPWR.n276 17.0005
R2594 VPWR.n282 VPWR.n275 17.0005
R2595 VPWR.n282 VPWR.n266 17.0005
R2596 VPWR.n282 VPWR.n265 17.0005
R2597 VPWR.n282 VPWR.n263 17.0005
R2598 VPWR.n282 VPWR.n261 17.0005
R2599 VPWR.n282 VPWR.n259 17.0005
R2600 VPWR.n282 VPWR.n257 17.0005
R2601 VPWR.n282 VPWR.n251 17.0005
R2602 VPWR.n283 VPWR.n282 17.0005
R2603 VPWR.n282 VPWR.n249 17.0005
R2604 VPWR.n306 VPWR.n297 17.0005
R2605 VPWR.n307 VPWR.n306 17.0005
R2606 VPWR.n306 VPWR.n298 17.0005
R2607 VPWR.n333 VPWR.n327 17.0005
R2608 VPWR.n333 VPWR.n326 17.0005
R2609 VPWR.n333 VPWR.n313 17.0005
R2610 VPWR.n334 VPWR.n333 17.0005
R2611 VPWR.n333 VPWR.n311 17.0005
R2612 VPWR.n357 VPWR.n348 17.0005
R2613 VPWR.n358 VPWR.n357 17.0005
R2614 VPWR.n357 VPWR.n349 17.0005
R2615 VPWR.n395 VPWR.n389 17.0005
R2616 VPWR.n395 VPWR.n388 17.0005
R2617 VPWR.n395 VPWR.n379 17.0005
R2618 VPWR.n395 VPWR.n378 17.0005
R2619 VPWR.n395 VPWR.n376 17.0005
R2620 VPWR.n395 VPWR.n374 17.0005
R2621 VPWR.n395 VPWR.n372 17.0005
R2622 VPWR.n395 VPWR.n370 17.0005
R2623 VPWR.n395 VPWR.n364 17.0005
R2624 VPWR.n396 VPWR.n395 17.0005
R2625 VPWR.n395 VPWR.n362 17.0005
R2626 VPWR.n432 VPWR.n426 17.0005
R2627 VPWR.n432 VPWR.n425 17.0005
R2628 VPWR.n432 VPWR.n414 17.0005
R2629 VPWR.n432 VPWR.n413 17.0005
R2630 VPWR.n432 VPWR.n411 17.0005
R2631 VPWR.n432 VPWR.n410 17.0005
R2632 VPWR.n432 VPWR.n409 17.0005
R2633 VPWR.n432 VPWR.n401 17.0005
R2634 VPWR.n433 VPWR.n432 17.0005
R2635 VPWR.n432 VPWR.n399 17.0005
R2636 VPWR.n482 VPWR.n443 17.0005
R2637 VPWR.n482 VPWR.n444 17.0005
R2638 VPWR.n482 VPWR.n441 17.0005
R2639 VPWR.n482 VPWR.n454 17.0005
R2640 VPWR.n482 VPWR.n481 17.0005
R2641 VPWR.n482 VPWR.n478 17.0005
R2642 VPWR.n482 VPWR.n476 17.0005
R2643 VPWR.n482 VPWR.n474 17.0005
R2644 VPWR.n482 VPWR.n472 17.0005
R2645 VPWR.n482 VPWR.n470 17.0005
R2646 VPWR.n482 VPWR.n468 17.0005
R2647 VPWR.n482 VPWR.n466 17.0005
R2648 VPWR.n482 VPWR.n464 17.0005
R2649 VPWR.n482 VPWR.n462 17.0005
R2650 VPWR.n482 VPWR.n460 17.0005
R2651 VPWR.n482 VPWR.n458 17.0005
R2652 VPWR.n482 VPWR.n457 17.0005
R2653 VPWR.n482 VPWR.n439 17.0005
R2654 VPWR.n483 VPWR.n482 17.0005
R2655 VPWR.n509 VPWR.n503 17.0005
R2656 VPWR.n509 VPWR.n502 17.0005
R2657 VPWR.n509 VPWR.n489 17.0005
R2658 VPWR.n510 VPWR.n509 17.0005
R2659 VPWR.n509 VPWR.n487 17.0005
R2660 VPWR.n545 VPWR.n539 17.0005
R2661 VPWR.n545 VPWR.n538 17.0005
R2662 VPWR.n545 VPWR.n527 17.0005
R2663 VPWR.n545 VPWR.n525 17.0005
R2664 VPWR.n545 VPWR.n523 17.0005
R2665 VPWR.n545 VPWR.n521 17.0005
R2666 VPWR.n545 VPWR.n515 17.0005
R2667 VPWR.n546 VPWR.n545 17.0005
R2668 VPWR.n545 VPWR.n513 17.0005
R2669 VPWR.n583 VPWR.n577 17.0005
R2670 VPWR.n583 VPWR.n576 17.0005
R2671 VPWR.n583 VPWR.n565 17.0005
R2672 VPWR.n583 VPWR.n564 17.0005
R2673 VPWR.n583 VPWR.n562 17.0005
R2674 VPWR.n583 VPWR.n561 17.0005
R2675 VPWR.n583 VPWR.n560 17.0005
R2676 VPWR.n583 VPWR.n552 17.0005
R2677 VPWR.n584 VPWR.n583 17.0005
R2678 VPWR.n583 VPWR.n550 17.0005
R2679 VPWR.n591 VPWR.n19 17.0005
R2680 VPWR.n591 VPWR.n18 17.0005
R2681 VPWR.n591 VPWR.n10 17.0005
R2682 VPWR.n591 VPWR.n9 17.0005
R2683 VPWR.n592 VPWR.n591 17.0005
R2684 VPWR.n591 VPWR.n1 17.0005
R2685 VPWR.n591 VPWR.n590 17.0005
R2686 VPWR.n479 VPWR.t485 15.3408
R2687 VPWR.n100 VPWR.t464 15.2933
R2688 VPWR.n446 VPWR.t463 15.2933
R2689 VPWR.n75 VPWR.t482 15.0005
R2690 VPWR.t482 VPWR.n74 15.0005
R2691 VPWR.n232 VPWR.t445 15.0005
R2692 VPWR.t445 VPWR.n231 15.0005
R2693 VPWR.n420 VPWR.t491 15.0005
R2694 VPWR.t491 VPWR.n419 15.0005
R2695 VPWR.n453 VPWR.t472 15.0005
R2696 VPWR.t472 VPWR.n452 15.0005
R2697 VPWR.n571 VPWR.t494 15.0005
R2698 VPWR.t494 VPWR.n570 15.0005
R2699 VPWR.n204 VPWR.t115 8.80529
R2700 VPWR.n242 VPWR.t319 8.80529
R2701 VPWR.n384 VPWR.t107 8.80529
R2702 VPWR.n543 VPWR.t364 8.80529
R2703 VPWR.n581 VPWR.t425 8.80529
R2704 VPWR.n82 VPWR.t81 8.7794
R2705 VPWR.n78 VPWR.t85 8.7794
R2706 VPWR VPWR.t80 8.7794
R2707 VPWR.n118 VPWR.t380 8.7794
R2708 VPWR.n122 VPWR.t379 8.7794
R2709 VPWR.n125 VPWR.t381 8.7794
R2710 VPWR.n116 VPWR.t103 8.7794
R2711 VPWR.n112 VPWR.t99 8.7794
R2712 VPWR.n108 VPWR.t102 8.7794
R2713 VPWR.n152 VPWR.t3 8.7794
R2714 VPWR.n155 VPWR.t1 8.7794
R2715 VPWR.n158 VPWR.t4 8.7794
R2716 VPWR.n164 VPWR.t391 8.7794
R2717 VPWR.n160 VPWR.t395 8.7794
R2718 VPWR VPWR.t390 8.7794
R2719 VPWR.n197 VPWR.t120 8.7794
R2720 VPWR.n201 VPWR.t116 8.7794
R2721 VPWR.n195 VPWR.t18 8.7794
R2722 VPWR.n192 VPWR.t22 8.7794
R2723 VPWR.n189 VPWR.t20 8.7794
R2724 VPWR.n235 VPWR.t318 8.7794
R2725 VPWR.n239 VPWR.t320 8.7794
R2726 VPWR.n267 VPWR.t72 8.7794
R2727 VPWR.n264 VPWR.t75 8.7794
R2728 VPWR VPWR.t76 8.7794
R2729 VPWR.n292 VPWR.t53 8.7794
R2730 VPWR.n292 VPWR.t418 8.7794
R2731 VPWR.n295 VPWR.t57 8.7794
R2732 VPWR.n295 VPWR.t417 8.7794
R2733 VPWR.n294 VPWR.t54 8.7794
R2734 VPWR.n294 VPWR.t419 8.7794
R2735 VPWR.n319 VPWR.t328 8.7794
R2736 VPWR.n319 VPWR.t408 8.7794
R2737 VPWR.n321 VPWR.t330 8.7794
R2738 VPWR.n321 VPWR.t405 8.7794
R2739 VPWR.n323 VPWR.t326 8.7794
R2740 VPWR.n323 VPWR.t409 8.7794
R2741 VPWR.n343 VPWR.t340 8.7794
R2742 VPWR.n343 VPWR.t44 8.7794
R2743 VPWR.n346 VPWR.t342 8.7794
R2744 VPWR.n346 VPWR.t48 8.7794
R2745 VPWR.n345 VPWR.t341 8.7794
R2746 VPWR.n345 VPWR.t45 8.7794
R2747 VPWR.n377 VPWR.t108 8.7794
R2748 VPWR.n380 VPWR.t111 8.7794
R2749 VPWR.n427 VPWR.t32 8.7794
R2750 VPWR.n423 VPWR.t28 8.7794
R2751 VPWR VPWR.t27 8.7794
R2752 VPWR.n463 VPWR.t310 8.7794
R2753 VPWR.n467 VPWR.t311 8.7794
R2754 VPWR.n471 VPWR.t316 8.7794
R2755 VPWR.n477 VPWR.t36 8.7794
R2756 VPWR.n473 VPWR.t39 8.7794
R2757 VPWR.n469 VPWR.t37 8.7794
R2758 VPWR.n495 VPWR.t357 8.7794
R2759 VPWR.n495 VPWR.t62 8.7794
R2760 VPWR.n497 VPWR.t355 8.7794
R2761 VPWR.n497 VPWR.t64 8.7794
R2762 VPWR.n499 VPWR.t356 8.7794
R2763 VPWR.n499 VPWR.t63 8.7794
R2764 VPWR.n536 VPWR.t365 8.7794
R2765 VPWR.n540 VPWR.t362 8.7794
R2766 VPWR.n534 VPWR.t302 8.7794
R2767 VPWR.n531 VPWR.t303 8.7794
R2768 VPWR.n528 VPWR.t308 8.7794
R2769 VPWR.n574 VPWR.t426 8.7794
R2770 VPWR.n578 VPWR.t423 8.7794
R2771 VPWR.n70 VPWR.t82 8.76423
R2772 VPWR.n114 VPWR.t386 8.76423
R2773 VPWR.n104 VPWR.t14 8.76423
R2774 VPWR.n148 VPWR.t2 8.76423
R2775 VPWR.n157 VPWR.t392 8.76423
R2776 VPWR.n194 VPWR.t90 8.76423
R2777 VPWR.n185 VPWR.t24 8.76423
R2778 VPWR.n227 VPWR.t321 8.76423
R2779 VPWR.n260 VPWR.t74 8.76423
R2780 VPWR.n290 VPWR.t58 8.76423
R2781 VPWR.n290 VPWR.t415 8.76423
R2782 VPWR.n317 VPWR.t332 8.76423
R2783 VPWR.n317 VPWR.t387 8.76423
R2784 VPWR.n341 VPWR.t337 8.76423
R2785 VPWR.n341 VPWR.t12 8.76423
R2786 VPWR.n373 VPWR.t112 8.76423
R2787 VPWR.n415 VPWR.t34 8.76423
R2788 VPWR.n459 VPWR.t312 8.76423
R2789 VPWR.n465 VPWR.t41 8.76423
R2790 VPWR.n493 VPWR.t349 8.76423
R2791 VPWR.n493 VPWR.t65 8.76423
R2792 VPWR.n533 VPWR.t126 8.76423
R2793 VPWR.n524 VPWR.t304 8.76423
R2794 VPWR.n566 VPWR.t94 8.76423
R2795 VPWR.n67 VPWR.t399 8.7637
R2796 VPWR.n101 VPWR.t15 8.7637
R2797 VPWR.n110 VPWR.t412 8.7637
R2798 VPWR.n143 VPWR.t133 8.7637
R2799 VPWR.n154 VPWR.t431 8.7637
R2800 VPWR.n180 VPWR.t130 8.7637
R2801 VPWR.n191 VPWR.t88 8.7637
R2802 VPWR.n224 VPWR.t441 8.7637
R2803 VPWR.n255 VPWR.t435 8.7637
R2804 VPWR.n288 VPWR.t95 8.7637
R2805 VPWR.n288 VPWR.t437 8.7637
R2806 VPWR.n315 VPWR.t370 8.7637
R2807 VPWR.n315 VPWR.t388 8.7637
R2808 VPWR.n339 VPWR.t338 8.7637
R2809 VPWR.n339 VPWR.t10 8.7637
R2810 VPWR.n368 VPWR.t401 8.7637
R2811 VPWR.n412 VPWR.t127 8.7637
R2812 VPWR.n455 VPWR.t352 8.7637
R2813 VPWR.n461 VPWR.t376 8.7637
R2814 VPWR.n491 VPWR.t348 8.7637
R2815 VPWR.n491 VPWR.t374 8.7637
R2816 VPWR.n519 VPWR.t334 8.7637
R2817 VPWR.n530 VPWR.t124 8.7637
R2818 VPWR.n563 VPWR.t92 8.7637
R2819 VPWR.n105 VPWR.t287 8.75396
R2820 VPWR.n451 VPWR.t297 8.75396
R2821 VPWR.n438 VPWR.t259 8.75396
R2822 VPWR.n133 VPWR.n98 8.501
R2823 VPWR.n282 VPWR.n268 8.50069
R2824 VPWR.n395 VPWR.n381 8.50069
R2825 VPWR.n102 VPWR.t286 8.5005
R2826 VPWR.n445 VPWR.t296 8.5005
R2827 VPWR.n479 VPWR.t258 8.48775
R2828 VPWR.n51 VPWR.n37 8.47111
R2829 VPWR.n51 VPWR.n33 8.47111
R2830 VPWR.n87 VPWR.n77 8.47111
R2831 VPWR.n87 VPWR.n62 8.47111
R2832 VPWR.n169 VPWR.n159 8.47111
R2833 VPWR.n169 VPWR.n156 8.47111
R2834 VPWR.n169 VPWR.n153 8.47111
R2835 VPWR.n169 VPWR.n141 8.47111
R2836 VPWR.n206 VPWR.n196 8.47111
R2837 VPWR.n206 VPWR.n193 8.47111
R2838 VPWR.n206 VPWR.n190 8.47111
R2839 VPWR.n206 VPWR.n178 8.47111
R2840 VPWR.n244 VPWR.n234 8.47111
R2841 VPWR.n244 VPWR.n219 8.47111
R2842 VPWR.n282 VPWR.n272 8.47111
R2843 VPWR.n282 VPWR.n253 8.47111
R2844 VPWR.n306 VPWR.n286 8.47111
R2845 VPWR.n306 VPWR.n296 8.47111
R2846 VPWR.n306 VPWR.n293 8.47111
R2847 VPWR.n306 VPWR.n291 8.47111
R2848 VPWR.n306 VPWR.n289 8.47111
R2849 VPWR.n306 VPWR.n287 8.47111
R2850 VPWR.n306 VPWR.n305 8.47111
R2851 VPWR.n333 VPWR.n324 8.47111
R2852 VPWR.n333 VPWR.n322 8.47111
R2853 VPWR.n333 VPWR.n320 8.47111
R2854 VPWR.n333 VPWR.n318 8.47111
R2855 VPWR.n333 VPWR.n316 8.47111
R2856 VPWR.n357 VPWR.n337 8.47111
R2857 VPWR.n357 VPWR.n347 8.47111
R2858 VPWR.n357 VPWR.n344 8.47111
R2859 VPWR.n357 VPWR.n342 8.47111
R2860 VPWR.n357 VPWR.n340 8.47111
R2861 VPWR.n357 VPWR.n338 8.47111
R2862 VPWR.n357 VPWR.n356 8.47111
R2863 VPWR.n395 VPWR.n385 8.47111
R2864 VPWR.n395 VPWR.n366 8.47111
R2865 VPWR.n432 VPWR.n422 8.47111
R2866 VPWR.n432 VPWR.n407 8.47111
R2867 VPWR.n482 VPWR.n440 8.47111
R2868 VPWR.n509 VPWR.n500 8.47111
R2869 VPWR.n509 VPWR.n498 8.47111
R2870 VPWR.n509 VPWR.n496 8.47111
R2871 VPWR.n509 VPWR.n494 8.47111
R2872 VPWR.n509 VPWR.n492 8.47111
R2873 VPWR.n545 VPWR.n535 8.47111
R2874 VPWR.n545 VPWR.n532 8.47111
R2875 VPWR.n545 VPWR.n529 8.47111
R2876 VPWR.n545 VPWR.n517 8.47111
R2877 VPWR.n583 VPWR.n573 8.47111
R2878 VPWR.n583 VPWR.n558 8.47111
R2879 VPWR.n591 VPWR.n11 8.47111
R2880 VPWR.n591 VPWR.n7 8.47111
R2881 VPWR.n142 VPWR.t447 7.62628
R2882 VPWR.n367 VPWR.t446 7.62628
R2883 VPWR.n47 VPWR.t466 7.62628
R2884 VPWR.n84 VPWR.t457 7.62628
R2885 VPWR.n166 VPWR.t451 7.62628
R2886 VPWR.n278 VPWR.t462 7.62628
R2887 VPWR.n301 VPWR.t450 7.62628
R2888 VPWR.n329 VPWR.t480 7.62628
R2889 VPWR.n352 VPWR.t455 7.62628
R2890 VPWR.n391 VPWR.t461 7.62628
R2891 VPWR.n429 VPWR.t443 7.62628
R2892 VPWR.n505 VPWR.t477 7.62628
R2893 VPWR.n21 VPWR.t497 7.62628
R2894 VPWR.n31 VPWR.t456 7.62594
R2895 VPWR.n40 VPWR.t473 7.62594
R2896 VPWR.n48 VPWR.t444 7.62594
R2897 VPWR.n60 VPWR.t468 7.62594
R2898 VPWR.n128 VPWR.t474 7.62594
R2899 VPWR.n203 VPWR.t458 7.62594
R2900 VPWR.n217 VPWR.t479 7.62594
R2901 VPWR.n241 VPWR.t471 7.62594
R2902 VPWR.n279 VPWR.t487 7.62594
R2903 VPWR.n303 VPWR.t486 7.62594
R2904 VPWR.n330 VPWR.t490 7.62594
R2905 VPWR.n354 VPWR.t469 7.62594
R2906 VPWR.n383 VPWR.t452 7.62594
R2907 VPWR.n392 VPWR.t475 7.62594
R2908 VPWR.n405 VPWR.t481 7.62594
R2909 VPWR.n506 VPWR.t493 7.62594
R2910 VPWR.n542 VPWR.t453 7.62594
R2911 VPWR.n556 VPWR.t495 7.62594
R2912 VPWR.n580 VPWR.t459 7.62594
R2913 VPWR.n5 VPWR.t448 7.62594
R2914 VPWR.n14 VPWR.t449 7.62594
R2915 VPWR.n23 VPWR.t496 7.62594
R2916 VPWR.n29 VPWR.t478 7.62594
R2917 VPWR.n38 VPWR.t460 7.62594
R2918 VPWR.n58 VPWR.t465 7.62594
R2919 VPWR.n179 VPWR.t470 7.62594
R2920 VPWR.n215 VPWR.t484 7.62594
R2921 VPWR.n254 VPWR.t476 7.62594
R2922 VPWR.n270 VPWR.t454 7.62594
R2923 VPWR.n403 VPWR.t492 7.62594
R2924 VPWR.n518 VPWR.t467 7.62594
R2925 VPWR.n554 VPWR.t483 7.62594
R2926 VPWR.n3 VPWR.t489 7.62594
R2927 VPWR.n12 VPWR.t488 7.62594
R2928 VPWR.n91 VPWR.n53 7.5029
R2929 VPWR.n91 VPWR.n90 7.2005
R2930 VPWR.n136 VPWR.n135 7.2005
R2931 VPWR.n173 VPWR.n172 7.2005
R2932 VPWR.n210 VPWR.n209 7.2005
R2933 VPWR.n248 VPWR.n247 7.2005
R2934 VPWR.n285 VPWR.n284 7.2005
R2935 VPWR.n310 VPWR.n309 7.2005
R2936 VPWR.n336 VPWR.n335 7.2005
R2937 VPWR.n361 VPWR.n360 7.2005
R2938 VPWR.n398 VPWR.n397 7.2005
R2939 VPWR.n436 VPWR.n435 7.2005
R2940 VPWR.n486 VPWR.n485 7.2005
R2941 VPWR.n512 VPWR.n511 7.2005
R2942 VPWR.n549 VPWR.n548 7.2005
R2943 VPWR.n587 VPWR.n586 7.2005
R2944 VPWR.n589 VPWR.n588 7.2005
R2945 VPWR.n131 VPWR.t384 5.98882
R2946 VPWR.n161 VPWR.t7 5.98882
R2947 VPWR.n208 VPWR.t118 5.98882
R2948 VPWR.n246 VPWR.t322 5.98882
R2949 VPWR.n308 VPWR.t59 5.98882
R2950 VPWR.n325 VPWR.t329 5.98882
R2951 VPWR.n359 VPWR.t344 5.98882
R2952 VPWR.n386 VPWR.t113 5.98882
R2953 VPWR.n475 VPWR.t313 5.98882
R2954 VPWR.n501 VPWR.t354 5.98882
R2955 VPWR.n547 VPWR.t368 5.98882
R2956 VPWR.n585 VPWR.t429 5.98882
R2957 VPWR.n89 VPWR.t83 5.9886
R2958 VPWR.n120 VPWR.t98 5.9886
R2959 VPWR.n171 VPWR.t393 5.9886
R2960 VPWR.n198 VPWR.t21 5.9886
R2961 VPWR.n273 VPWR.t71 5.9886
R2962 VPWR.n308 VPWR.t416 5.9886
R2963 VPWR.n325 VPWR.t404 5.9886
R2964 VPWR.n359 VPWR.t50 5.9886
R2965 VPWR.n434 VPWR.t31 5.9886
R2966 VPWR.n484 VPWR.t38 5.9886
R2967 VPWR.n501 VPWR.t66 5.9886
R2968 VPWR.n537 VPWR.t305 5.9886
R2969 VPWR.n34 VPWR.t243 5.97235
R2970 VPWR.n43 VPWR.t159 5.97235
R2971 VPWR.t166 VPWR.n46 5.97235
R2972 VPWR.n26 VPWR.t167 5.97235
R2973 VPWR.n63 VPWR.t218 5.97235
R2974 VPWR.t194 VPWR.n72 5.97235
R2975 VPWR.n79 VPWR.t301 5.97235
R2976 VPWR.t144 VPWR.n83 5.97235
R2977 VPWR.n55 VPWR.t145 5.97235
R2978 VPWR.t188 VPWR.n165 5.97235
R2979 VPWR.n138 VPWR.t249 5.97235
R2980 VPWR.n187 VPWR.t270 5.97235
R2981 VPWR.n220 VPWR.t228 5.97235
R2982 VPWR.n262 VPWR.t172 5.97235
R2983 VPWR.n274 VPWR.t254 5.97235
R2984 VPWR.t197 VPWR.n277 5.97235
R2985 VPWR.n250 VPWR.t268 5.97235
R2986 VPWR.n302 VPWR.t136 5.97235
R2987 VPWR.n300 VPWR.t137 5.97235
R2988 VPWR.t205 VPWR.n328 5.97235
R2989 VPWR.n312 VPWR.t206 5.97235
R2990 VPWR.n353 VPWR.t204 5.97235
R2991 VPWR.n351 VPWR.t289 5.97235
R2992 VPWR.t260 VPWR.n390 5.97235
R2993 VPWR.n363 VPWR.t261 5.97235
R2994 VPWR.n408 VPWR.t291 5.97235
R2995 VPWR.t235 VPWR.n417 5.97235
R2996 VPWR.n424 VPWR.t236 5.97235
R2997 VPWR.t222 VPWR.n428 5.97235
R2998 VPWR.n400 VPWR.t223 5.97235
R2999 VPWR.t162 VPWR.n504 5.97235
R3000 VPWR.n488 VPWR.t163 5.97235
R3001 VPWR.n526 VPWR.t215 5.97235
R3002 VPWR.n559 VPWR.t187 5.97235
R3003 VPWR.n8 VPWR.t184 5.97235
R3004 VPWR.n17 VPWR.t191 5.97235
R3005 VPWR.n22 VPWR.t202 5.97235
R3006 VPWR.n0 VPWR.t203 5.97235
R3007 VPWR.n34 VPWR.t225 5.97213
R3008 VPWR.n43 VPWR.t151 5.97213
R3009 VPWR.n26 VPWR.t154 5.97213
R3010 VPWR.n63 VPWR.t199 5.97213
R3011 VPWR.n93 VPWR.t263 5.97213
R3012 VPWR.t169 VPWR.n140 5.97213
R3013 VPWR.n150 VPWR.t266 5.97213
R3014 VPWR.n175 VPWR.t247 5.97213
R3015 VPWR.n220 VPWR.t176 5.97213
R3016 VPWR.t148 VPWR.n229 5.97213
R3017 VPWR.n236 VPWR.t257 5.97213
R3018 VPWR.n212 VPWR.t272 5.97213
R3019 VPWR.n250 VPWR.t234 5.97213
R3020 VPWR.n300 VPWR.t282 5.97213
R3021 VPWR.n312 VPWR.t182 5.97213
R3022 VPWR.n351 VPWR.t220 5.97213
R3023 VPWR.t138 VPWR.n365 5.97213
R3024 VPWR.n375 VPWR.t139 5.97213
R3025 VPWR.n387 VPWR.t251 5.97213
R3026 VPWR.n363 VPWR.t230 5.97213
R3027 VPWR.n408 VPWR.t232 5.97213
R3028 VPWR.t208 VPWR.n447 5.97213
R3029 VPWR.n456 VPWR.t209 5.97213
R3030 VPWR.n488 VPWR.t279 5.97213
R3031 VPWR.n514 VPWR.t240 5.97213
R3032 VPWR.n559 VPWR.t165 5.97213
R3033 VPWR.t179 VPWR.n568 5.97213
R3034 VPWR.n575 VPWR.t284 5.97213
R3035 VPWR.n551 VPWR.t274 5.97213
R3036 VPWR.n8 VPWR.t157 5.97213
R3037 VPWR.n17 VPWR.t161 5.97213
R3038 VPWR.n0 VPWR.t178 5.97213
R3039 VPWR.n30 VPWR.t152 5.97135
R3040 VPWR.t141 VPWR.n30 5.97135
R3041 VPWR.n39 VPWR.t158 5.97135
R3042 VPWR.t150 VPWR.n39 5.97135
R3043 VPWR.t153 VPWR.n46 5.97135
R3044 VPWR.n59 VPWR.t217 5.97135
R3045 VPWR.t198 VPWR.n59 5.97135
R3046 VPWR.t196 VPWR.n127 5.97135
R3047 VPWR.t173 VPWR.n177 5.97135
R3048 VPWR.t185 VPWR.n202 5.97135
R3049 VPWR.n216 VPWR.t149 5.97135
R3050 VPWR.t175 VPWR.n216 5.97135
R3051 VPWR.t201 VPWR.n240 5.97135
R3052 VPWR.t171 VPWR.n252 5.97135
R3053 VPWR.t143 VPWR.n269 5.97135
R3054 VPWR.t168 VPWR.n277 5.97135
R3055 VPWR.t193 VPWR.n302 5.97135
R3056 VPWR.t181 VPWR.n328 5.97135
R3057 VPWR.t219 VPWR.n353 5.97135
R3058 VPWR.t146 VPWR.n382 5.97135
R3059 VPWR.t229 VPWR.n390 5.97135
R3060 VPWR.n404 VPWR.t290 5.97135
R3061 VPWR.t231 VPWR.n404 5.97135
R3062 VPWR.t278 VPWR.n504 5.97135
R3063 VPWR.t214 VPWR.n516 5.97135
R3064 VPWR.t239 VPWR.n541 5.97135
R3065 VPWR.n555 VPWR.t186 5.97135
R3066 VPWR.t164 VPWR.n555 5.97135
R3067 VPWR.t273 VPWR.n579 5.97135
R3068 VPWR.n4 VPWR.t183 5.97135
R3069 VPWR.t156 VPWR.n4 5.97135
R3070 VPWR.n13 VPWR.t190 5.97135
R3071 VPWR.t160 VPWR.n13 5.97135
R3072 VPWR.t177 VPWR.n22 5.97135
R3073 VPWR.n73 VPWR.t194 5.66717
R3074 VPWR.n230 VPWR.t148 5.66717
R3075 VPWR.n418 VPWR.t235 5.66717
R3076 VPWR.n448 VPWR.t208 5.66717
R3077 VPWR.n569 VPWR.t179 5.66717
R3078 VPWR.n31 VPWR.t141 5.65005
R3079 VPWR.t152 VPWR.n29 5.65005
R3080 VPWR.n40 VPWR.t150 5.65005
R3081 VPWR.t158 VPWR.n38 5.65005
R3082 VPWR.n48 VPWR.t153 5.65005
R3083 VPWR.n47 VPWR.t166 5.65005
R3084 VPWR.n60 VPWR.t198 5.65005
R3085 VPWR.t217 VPWR.n58 5.65005
R3086 VPWR.n84 VPWR.t144 5.65005
R3087 VPWR.n128 VPWR.t196 5.65005
R3088 VPWR.n142 VPWR.t169 5.65005
R3089 VPWR.n166 VPWR.t188 5.65005
R3090 VPWR.n179 VPWR.t173 5.65005
R3091 VPWR.n203 VPWR.t185 5.65005
R3092 VPWR.n217 VPWR.t175 5.65005
R3093 VPWR.t149 VPWR.n215 5.65005
R3094 VPWR.n241 VPWR.t201 5.65005
R3095 VPWR.n254 VPWR.t171 5.65005
R3096 VPWR.n270 VPWR.t143 5.65005
R3097 VPWR.n279 VPWR.t168 5.65005
R3098 VPWR.n278 VPWR.t197 5.65005
R3099 VPWR.n303 VPWR.t193 5.65005
R3100 VPWR.t136 VPWR.n301 5.65005
R3101 VPWR.n330 VPWR.t181 5.65005
R3102 VPWR.n329 VPWR.t205 5.65005
R3103 VPWR.n354 VPWR.t219 5.65005
R3104 VPWR.t204 VPWR.n352 5.65005
R3105 VPWR.n367 VPWR.t138 5.65005
R3106 VPWR.n383 VPWR.t146 5.65005
R3107 VPWR.n392 VPWR.t229 5.65005
R3108 VPWR.n391 VPWR.t260 5.65005
R3109 VPWR.n405 VPWR.t231 5.65005
R3110 VPWR.t290 VPWR.n403 5.65005
R3111 VPWR.n429 VPWR.t222 5.65005
R3112 VPWR.n506 VPWR.t278 5.65005
R3113 VPWR.n505 VPWR.t162 5.65005
R3114 VPWR.n518 VPWR.t214 5.65005
R3115 VPWR.n542 VPWR.t239 5.65005
R3116 VPWR.n556 VPWR.t164 5.65005
R3117 VPWR.t186 VPWR.n554 5.65005
R3118 VPWR.n580 VPWR.t273 5.65005
R3119 VPWR.n5 VPWR.t156 5.65005
R3120 VPWR.t183 VPWR.n3 5.65005
R3121 VPWR.n14 VPWR.t160 5.65005
R3122 VPWR.t190 VPWR.n12 5.65005
R3123 VPWR.n23 VPWR.t177 5.65005
R3124 VPWR.t202 VPWR.n21 5.65005
R3125 VPWR.n51 VPWR.n50 5.64096
R3126 VPWR.n87 VPWR.n86 5.64096
R3127 VPWR.n169 VPWR.n168 5.64096
R3128 VPWR.n206 VPWR.n205 5.64096
R3129 VPWR.n244 VPWR.n243 5.64096
R3130 VPWR.n282 VPWR.n281 5.64096
R3131 VPWR.n333 VPWR.n332 5.64096
R3132 VPWR.n395 VPWR.n394 5.64096
R3133 VPWR.n432 VPWR.n431 5.64096
R3134 VPWR.n509 VPWR.n508 5.64096
R3135 VPWR.n545 VPWR.n544 5.64096
R3136 VPWR.n583 VPWR.n582 5.64096
R3137 VPWR.n591 VPWR.n20 5.64096
R3138 VPWR.n51 VPWR.n42 5.64013
R3139 VPWR.n591 VPWR.n16 5.64013
R3140 VPWR.n333 VPWR.n314 5.63466
R3141 VPWR.n509 VPWR.n490 5.63466
R3142 VPWR.n51 VPWR.n28 4.20159
R3143 VPWR.n87 VPWR.n57 4.20159
R3144 VPWR.n244 VPWR.n214 4.20159
R3145 VPWR.n306 VPWR.n299 4.20159
R3146 VPWR.n357 VPWR.n350 4.20159
R3147 VPWR.n432 VPWR.n402 4.20159
R3148 VPWR.n583 VPWR.n553 4.20159
R3149 VPWR.n591 VPWR.n2 4.20159
R3150 VPWR.n51 VPWR.t140 0.810024
R3151 VPWR.n87 VPWR.t79 0.810024
R3152 VPWR.n133 VPWR.t13 0.810024
R3153 VPWR.n169 VPWR.t0 0.810024
R3154 VPWR.n206 VPWR.t17 0.810024
R3155 VPWR.n244 VPWR.t147 0.810024
R3156 VPWR.n282 VPWR.t70 0.810024
R3157 VPWR.n306 VPWR.t52 0.810024
R3158 VPWR.n333 VPWR.t180 0.810024
R3159 VPWR.n357 VPWR.t9 0.810024
R3160 VPWR.n395 VPWR.t106 0.810024
R3161 VPWR.n432 VPWR.t26 0.810024
R3162 VPWR.n482 VPWR.t35 0.810024
R3163 VPWR.n509 VPWR.t61 0.810024
R3164 VPWR.n545 VPWR.t123 0.810024
R3165 VPWR.n583 VPWR.t91 0.810024
R3166 VPWR.n591 VPWR.t155 0.810024
R3167 VPWR.n32 VPWR 0.53925
R3168 VPWR.n41 VPWR 0.53925
R3169 VPWR.n49 VPWR 0.53925
R3170 VPWR.n61 VPWR 0.53925
R3171 VPWR.n71 VPWR 0.53925
R3172 VPWR.n218 VPWR 0.53925
R3173 VPWR.n228 VPWR 0.53925
R3174 VPWR.n271 VPWR 0.53925
R3175 VPWR.n280 VPWR 0.53925
R3176 VPWR.n304 VPWR 0.53925
R3177 VPWR.n331 VPWR 0.53925
R3178 VPWR.n355 VPWR 0.53925
R3179 VPWR.n384 VPWR 0.53925
R3180 VPWR.n393 VPWR 0.53925
R3181 VPWR.n406 VPWR 0.53925
R3182 VPWR.n416 VPWR 0.53925
R3183 VPWR.n507 VPWR 0.53925
R3184 VPWR.n557 VPWR 0.53925
R3185 VPWR.n567 VPWR 0.53925
R3186 VPWR.n6 VPWR 0.53925
R3187 VPWR.n15 VPWR 0.53925
R3188 VPWR.n24 VPWR 0.53925
R3189 VPWR.n444 VPWR 0.456288
R3190 VPWR.n99 VPWR 0.448
R3191 VPWR.n85 VPWR 0.41925
R3192 VPWR.n167 VPWR 0.41925
R3193 VPWR.n204 VPWR 0.41925
R3194 VPWR.n242 VPWR 0.41925
R3195 VPWR.n430 VPWR 0.41925
R3196 VPWR.n543 VPWR 0.41925
R3197 VPWR.n581 VPWR 0.41925
R3198 VPWR.n146 VPWR 0.3055
R3199 VPWR.n183 VPWR 0.3055
R3200 VPWR.n258 VPWR 0.3055
R3201 VPWR.n371 VPWR 0.3055
R3202 VPWR.n522 VPWR 0.3055
R3203 VPWR.n136 VPWR.n91 0.3029
R3204 VPWR.n173 VPWR.n136 0.3029
R3205 VPWR.n210 VPWR.n173 0.3029
R3206 VPWR.n248 VPWR.n210 0.3029
R3207 VPWR.n285 VPWR.n248 0.3029
R3208 VPWR.n310 VPWR.n285 0.3029
R3209 VPWR.n336 VPWR.n310 0.3029
R3210 VPWR.n361 VPWR.n336 0.3029
R3211 VPWR.n398 VPWR.n361 0.3029
R3212 VPWR.n436 VPWR.n398 0.3029
R3213 VPWR.n486 VPWR.n436 0.3029
R3214 VPWR.n512 VPWR.n486 0.3029
R3215 VPWR.n549 VPWR.n512 0.3029
R3216 VPWR.n587 VPWR.n549 0.3029
R3217 VPWR.n588 VPWR.n587 0.3029
R3218 VPWR.n129 VPWR 0.29925
R3219 VPWR.n50 VPWR.n46 0.190118
R3220 VPWR.n281 VPWR.n277 0.190118
R3221 VPWR.n332 VPWR.n328 0.190118
R3222 VPWR.n394 VPWR.n390 0.190118
R3223 VPWR.n508 VPWR.n504 0.190118
R3224 VPWR.n22 VPWR.n20 0.190118
R3225 VPWR.n43 VPWR.n42 0.183859
R3226 VPWR.n17 VPWR.n16 0.183859
R3227 VPWR.n450 VPWR 0.17925
R3228 VPWR.n39 VPWR.n37 0.169539
R3229 VPWR.n13 VPWR.n11 0.169539
R3230 VPWR.n34 VPWR.n33 0.162039
R3231 VPWR.n63 VPWR.n62 0.162039
R3232 VPWR.n220 VPWR.n219 0.162039
R3233 VPWR.n305 VPWR.n300 0.162039
R3234 VPWR.n356 VPWR.n351 0.162039
R3235 VPWR.n408 VPWR.n407 0.162039
R3236 VPWR.n559 VPWR.n558 0.162039
R3237 VPWR.n8 VPWR.n7 0.162039
R3238 VPWR.n289 VPWR.n288 0.160789
R3239 VPWR.n316 VPWR.n315 0.160789
R3240 VPWR.n340 VPWR.n339 0.160789
R3241 VPWR.n492 VPWR.n491 0.160789
R3242 VPWR.n588 VPWR 0.1605
R3243 VPWR.n273 VPWR.n272 0.155789
R3244 VPWR.n325 VPWR.n324 0.155789
R3245 VPWR.n386 VPWR.n385 0.155789
R3246 VPWR.n501 VPWR.n500 0.155789
R3247 VPWR.n437 VPWR 0.14675
R3248 VPWR.n291 VPWR.n290 0.145789
R3249 VPWR.n318 VPWR.n317 0.145789
R3250 VPWR.n342 VPWR.n341 0.145789
R3251 VPWR.n494 VPWR.n493 0.145789
R3252 VPWR.n30 VPWR.n28 0.1426
R3253 VPWR.n59 VPWR.n57 0.1426
R3254 VPWR.n216 VPWR.n214 0.1426
R3255 VPWR.n302 VPWR.n299 0.1426
R3256 VPWR.n353 VPWR.n350 0.1426
R3257 VPWR.n404 VPWR.n402 0.1426
R3258 VPWR.n555 VPWR.n553 0.1426
R3259 VPWR.n4 VPWR.n2 0.1426
R3260 VPWR.n296 VPWR.n294 0.140789
R3261 VPWR.n323 VPWR.n322 0.140789
R3262 VPWR.n347 VPWR.n345 0.140789
R3263 VPWR.n499 VPWR.n498 0.140789
R3264 VPWR.n86 VPWR.n82 0.136368
R3265 VPWR.n168 VPWR.n164 0.136368
R3266 VPWR.n205 VPWR.n201 0.136368
R3267 VPWR.n243 VPWR.n239 0.136368
R3268 VPWR.n431 VPWR.n427 0.136368
R3269 VPWR.n544 VPWR.n540 0.136368
R3270 VPWR.n582 VPWR.n578 0.136368
R3271 VPWR.n293 VPWR.n292 0.130789
R3272 VPWR.n320 VPWR.n319 0.130789
R3273 VPWR.n344 VPWR.n343 0.130789
R3274 VPWR.n496 VPWR.n495 0.130789
R3275 VPWR.n32 VPWR.n29 0.12922
R3276 VPWR.n41 VPWR.n38 0.12922
R3277 VPWR.n61 VPWR.n58 0.12922
R3278 VPWR.n218 VPWR.n215 0.12922
R3279 VPWR.n271 VPWR.n270 0.12922
R3280 VPWR.n406 VPWR.n403 0.12922
R3281 VPWR.n557 VPWR.n554 0.12922
R3282 VPWR.n6 VPWR.n3 0.12922
R3283 VPWR.n15 VPWR.n12 0.12922
R3284 VPWR.n49 VPWR.n47 0.128884
R3285 VPWR.n85 VPWR.n84 0.128884
R3286 VPWR.n167 VPWR.n166 0.128884
R3287 VPWR.n280 VPWR.n278 0.128884
R3288 VPWR.n304 VPWR.n301 0.128884
R3289 VPWR.n331 VPWR.n329 0.128884
R3290 VPWR.n355 VPWR.n352 0.128884
R3291 VPWR.n393 VPWR.n391 0.128884
R3292 VPWR.n430 VPWR.n429 0.128884
R3293 VPWR.n507 VPWR.n505 0.128884
R3294 VPWR.n24 VPWR.n21 0.128884
R3295 VPWR.n295 VPWR.n293 0.125789
R3296 VPWR.n321 VPWR.n320 0.125789
R3297 VPWR.n346 VPWR.n344 0.125789
R3298 VPWR.n497 VPWR.n496 0.125789
R3299 VPWR.n141 VPWR 0.120789
R3300 VPWR.n153 VPWR 0.120789
R3301 VPWR.n178 VPWR 0.120789
R3302 VPWR.n190 VPWR 0.120789
R3303 VPWR.n253 VPWR 0.120789
R3304 VPWR VPWR.n287 0.120789
R3305 VPWR VPWR.n338 0.120789
R3306 VPWR.n366 VPWR 0.120789
R3307 VPWR.n517 VPWR 0.120789
R3308 VPWR.n529 VPWR 0.120789
R3309 VPWR.n315 VPWR.n314 0.120673
R3310 VPWR.n491 VPWR.n490 0.120673
R3311 VPWR.n130 VPWR.n129 0.118
R3312 VPWR.n156 VPWR.n155 0.115789
R3313 VPWR.n193 VPWR.n192 0.115789
R3314 VPWR.n296 VPWR.n295 0.115789
R3315 VPWR.n322 VPWR.n321 0.115789
R3316 VPWR.n347 VPWR.n346 0.115789
R3317 VPWR.n498 VPWR.n497 0.115789
R3318 VPWR.n532 VPWR.n531 0.115789
R3319 VPWR.n146 VPWR.n145 0.1155
R3320 VPWR.n183 VPWR.n182 0.1155
R3321 VPWR.n258 VPWR.n257 0.1155
R3322 VPWR.n371 VPWR.n370 0.1155
R3323 VPWR.n522 VPWR.n521 0.1155
R3324 VPWR.n78 VPWR.n77 0.110789
R3325 VPWR.n160 VPWR.n159 0.110789
R3326 VPWR.n197 VPWR.n196 0.110789
R3327 VPWR.n235 VPWR.n234 0.110789
R3328 VPWR.n292 VPWR.n291 0.110789
R3329 VPWR.n309 VPWR.n286 0.110789
R3330 VPWR.n319 VPWR.n318 0.110789
R3331 VPWR.n343 VPWR.n342 0.110789
R3332 VPWR.n360 VPWR.n337 0.110789
R3333 VPWR.n423 VPWR.n422 0.110789
R3334 VPWR.n495 VPWR.n494 0.110789
R3335 VPWR.n536 VPWR.n535 0.110789
R3336 VPWR.n574 VPWR.n573 0.110789
R3337 VPWR.n72 VPWR.n66 0.10925
R3338 VPWR.n127 VPWR.n124 0.10925
R3339 VPWR.n229 VPWR.n223 0.10925
R3340 VPWR.n269 VPWR.n266 0.10925
R3341 VPWR.n382 VPWR.n379 0.10925
R3342 VPWR.n417 VPWR.n411 0.10925
R3343 VPWR.n568 VPWR.n562 0.10925
R3344 VPWR.n480 VPWR.n479 0.108683
R3345 VPWR VPWR.n31 0.103337
R3346 VPWR VPWR.n40 0.103337
R3347 VPWR VPWR.n48 0.103337
R3348 VPWR VPWR.n60 0.103337
R3349 VPWR.n130 VPWR.n128 0.103337
R3350 VPWR.n181 VPWR.n179 0.103337
R3351 VPWR VPWR.n203 0.103337
R3352 VPWR VPWR.n217 0.103337
R3353 VPWR VPWR.n241 0.103337
R3354 VPWR.n256 VPWR.n254 0.103337
R3355 VPWR VPWR.n279 0.103337
R3356 VPWR VPWR.n303 0.103337
R3357 VPWR VPWR.n330 0.103337
R3358 VPWR VPWR.n354 0.103337
R3359 VPWR VPWR.n383 0.103337
R3360 VPWR VPWR.n392 0.103337
R3361 VPWR VPWR.n405 0.103337
R3362 VPWR VPWR.n506 0.103337
R3363 VPWR.n520 VPWR.n518 0.103337
R3364 VPWR VPWR.n542 0.103337
R3365 VPWR VPWR.n556 0.103337
R3366 VPWR VPWR.n580 0.103337
R3367 VPWR VPWR.n5 0.103337
R3368 VPWR VPWR.n14 0.103337
R3369 VPWR VPWR.n23 0.103337
R3370 VPWR.n144 VPWR.n142 0.103002
R3371 VPWR.n369 VPWR.n367 0.103002
R3372 VPWR.n52 VPWR.n26 0.10175
R3373 VPWR.n134 VPWR.n93 0.10175
R3374 VPWR.n150 VPWR.n149 0.10175
R3375 VPWR.n187 VPWR.n186 0.10175
R3376 VPWR.n262 VPWR.n261 0.10175
R3377 VPWR.n283 VPWR.n250 0.10175
R3378 VPWR.n334 VPWR.n312 0.10175
R3379 VPWR.n375 VPWR.n374 0.10175
R3380 VPWR.n396 VPWR.n363 0.10175
R3381 VPWR.n510 VPWR.n488 0.10175
R3382 VPWR.n526 VPWR.n525 0.10175
R3383 VPWR.n1 VPWR.n0 0.10175
R3384 VPWR.n159 VPWR.n158 0.100789
R3385 VPWR.n196 VPWR.n195 0.100789
R3386 VPWR.n294 VPWR.n286 0.100789
R3387 VPWR.n324 VPWR.n323 0.100789
R3388 VPWR.n345 VPWR.n337 0.100789
R3389 VPWR.n500 VPWR.n499 0.100789
R3390 VPWR.n535 VPWR.n534 0.100789
R3391 VPWR.n68 VPWR.n67 0.1005
R3392 VPWR.n111 VPWR.n110 0.1005
R3393 VPWR.n225 VPWR.n224 0.1005
R3394 VPWR.n413 VPWR.n412 0.1005
R3395 VPWR.n462 VPWR.n461 0.1005
R3396 VPWR.n564 VPWR.n563 0.1005
R3397 VPWR.n144 VPWR.n143 0.09925
R3398 VPWR.n181 VPWR.n180 0.09925
R3399 VPWR.n256 VPWR.n255 0.09925
R3400 VPWR.n369 VPWR.n368 0.09925
R3401 VPWR.n520 VPWR.n519 0.09925
R3402 VPWR.n157 VPWR.n156 0.095789
R3403 VPWR.n194 VPWR.n193 0.095789
R3404 VPWR.n290 VPWR.n289 0.095789
R3405 VPWR.n317 VPWR.n316 0.095789
R3406 VPWR.n341 VPWR.n340 0.095789
R3407 VPWR.n493 VPWR.n492 0.095789
R3408 VPWR.n533 VPWR.n532 0.095789
R3409 VPWR.n120 VPWR.n119 0.0955
R3410 VPWR.n132 VPWR.n131 0.0955
R3411 VPWR.n475 VPWR.n474 0.0955
R3412 VPWR VPWR.n98 0.0908945
R3413 VPWR.n32 VPWR.n28 0.0892512
R3414 VPWR.n61 VPWR.n57 0.0892512
R3415 VPWR.n218 VPWR.n214 0.0892512
R3416 VPWR.n304 VPWR.n299 0.0892512
R3417 VPWR.n355 VPWR.n350 0.0892512
R3418 VPWR.n406 VPWR.n402 0.0892512
R3419 VPWR.n557 VPWR.n553 0.0892512
R3420 VPWR.n6 VPWR.n2 0.0892512
R3421 VPWR.n96 VPWR.n95 0.08675
R3422 VPWR.n442 VPWR.n441 0.08675
R3423 VPWR.n115 VPWR.n114 0.0855
R3424 VPWR.n149 VPWR.n148 0.0855
R3425 VPWR.n186 VPWR.n185 0.0855
R3426 VPWR.n261 VPWR.n260 0.0855
R3427 VPWR.n374 VPWR.n373 0.0855
R3428 VPWR.n460 VPWR.n459 0.0855
R3429 VPWR.n466 VPWR.n465 0.0855
R3430 VPWR.n525 VPWR.n524 0.0855
R3431 VPWR.n456 VPWR.n455 0.08175
R3432 VPWR.n314 VPWR 0.0813395
R3433 VPWR.n490 VPWR 0.0813395
R3434 VPWR.n143 VPWR.n141 0.080789
R3435 VPWR.n154 VPWR.n153 0.080789
R3436 VPWR.n180 VPWR.n178 0.080789
R3437 VPWR.n191 VPWR.n190 0.080789
R3438 VPWR.n255 VPWR.n253 0.080789
R3439 VPWR.n288 VPWR.n287 0.080789
R3440 VPWR.n339 VPWR.n338 0.080789
R3441 VPWR.n368 VPWR.n366 0.080789
R3442 VPWR.n455 VPWR.n440 0.080789
R3443 VPWR.n519 VPWR.n517 0.080789
R3444 VPWR.n530 VPWR.n529 0.080789
R3445 VPWR.n96 VPWR 0.0807397
R3446 VPWR.n442 VPWR 0.0807397
R3447 VPWR.n116 VPWR.n115 0.0805
R3448 VPWR.n125 VPWR.n124 0.0805
R3449 VPWR.n471 VPWR.n470 0.0805
R3450 VPWR.n105 VPWR.n104 0.07925
R3451 VPWR.n53 VPWR.n52 0.0705
R3452 VPWR.n109 VPWR.n108 0.0705
R3453 VPWR.n119 VPWR.n118 0.0705
R3454 VPWR.n284 VPWR.n283 0.0705
R3455 VPWR.n335 VPWR.n334 0.0705
R3456 VPWR.n397 VPWR.n396 0.0705
R3457 VPWR.n464 VPWR.n463 0.0705
R3458 VPWR.n470 VPWR.n469 0.0705
R3459 VPWR.n511 VPWR.n510 0.0705
R3460 VPWR.n589 VPWR.n1 0.0705
R3461 VPWR.n33 VPWR.n32 0.065789
R3462 VPWR.n62 VPWR.n61 0.065789
R3463 VPWR.n77 VPWR.n76 0.065789
R3464 VPWR.n219 VPWR.n218 0.065789
R3465 VPWR.n234 VPWR.n233 0.065789
R3466 VPWR.n272 VPWR.n271 0.065789
R3467 VPWR.n305 VPWR.n304 0.065789
R3468 VPWR.n356 VPWR.n355 0.065789
R3469 VPWR.n385 VPWR.n384 0.065789
R3470 VPWR.n407 VPWR.n406 0.065789
R3471 VPWR.n422 VPWR.n421 0.065789
R3472 VPWR.n449 VPWR.n440 0.065789
R3473 VPWR.n558 VPWR.n557 0.065789
R3474 VPWR.n573 VPWR.n572 0.065789
R3475 VPWR.n7 VPWR.n6 0.065789
R3476 VPWR.n112 VPWR.n111 0.0655
R3477 VPWR.n267 VPWR.n266 0.0655
R3478 VPWR.n380 VPWR.n379 0.0655
R3479 VPWR.n467 VPWR.n466 0.0655
R3480 VPWR.n473 VPWR.n472 0.0655
R3481 VPWR.n480 VPWR.n478 0.06425
R3482 VPWR.n41 VPWR.n37 0.062039
R3483 VPWR.n15 VPWR.n11 0.062039
R3484 VPWR VPWR.n35 0.0605
R3485 VPWR.n36 VPWR 0.0605
R3486 VPWR VPWR.n44 0.0605
R3487 VPWR.n45 VPWR 0.0605
R3488 VPWR.n27 VPWR 0.0605
R3489 VPWR VPWR.n64 0.0605
R3490 VPWR.n65 VPWR 0.0605
R3491 VPWR VPWR.n80 0.0605
R3492 VPWR.n81 VPWR 0.0605
R3493 VPWR.n88 VPWR 0.0605
R3494 VPWR.n56 VPWR 0.0605
R3495 VPWR VPWR.n106 0.0605
R3496 VPWR.n107 VPWR 0.0605
R3497 VPWR VPWR.n121 0.0605
R3498 VPWR VPWR.n134 0.0605
R3499 VPWR.n94 VPWR 0.0605
R3500 VPWR VPWR.n162 0.0605
R3501 VPWR.n163 VPWR 0.0605
R3502 VPWR.n170 VPWR 0.0605
R3503 VPWR.n139 VPWR 0.0605
R3504 VPWR VPWR.n199 0.0605
R3505 VPWR.n200 VPWR 0.0605
R3506 VPWR.n207 VPWR 0.0605
R3507 VPWR.n176 VPWR 0.0605
R3508 VPWR VPWR.n221 0.0605
R3509 VPWR.n222 VPWR 0.0605
R3510 VPWR VPWR.n237 0.0605
R3511 VPWR.n238 VPWR 0.0605
R3512 VPWR.n245 VPWR 0.0605
R3513 VPWR.n213 VPWR 0.0605
R3514 VPWR.n265 VPWR 0.0605
R3515 VPWR VPWR.n275 0.0605
R3516 VPWR.n276 VPWR 0.0605
R3517 VPWR.n251 VPWR 0.0605
R3518 VPWR.n298 VPWR 0.0605
R3519 VPWR.n307 VPWR 0.0605
R3520 VPWR.n297 VPWR 0.0605
R3521 VPWR.n297 VPWR 0.0605
R3522 VPWR VPWR.n326 0.0605
R3523 VPWR.n327 VPWR 0.0605
R3524 VPWR.n313 VPWR 0.0605
R3525 VPWR.n349 VPWR 0.0605
R3526 VPWR.n358 VPWR 0.0605
R3527 VPWR.n348 VPWR 0.0605
R3528 VPWR.n348 VPWR 0.0605
R3529 VPWR.n378 VPWR 0.0605
R3530 VPWR VPWR.n388 0.0605
R3531 VPWR.n389 VPWR 0.0605
R3532 VPWR.n364 VPWR 0.0605
R3533 VPWR VPWR.n409 0.0605
R3534 VPWR.n410 VPWR 0.0605
R3535 VPWR VPWR.n425 0.0605
R3536 VPWR.n426 VPWR 0.0605
R3537 VPWR.n433 VPWR 0.0605
R3538 VPWR.n401 VPWR 0.0605
R3539 VPWR VPWR.n457 0.0605
R3540 VPWR.n458 VPWR 0.0605
R3541 VPWR VPWR.n476 0.0605
R3542 VPWR.n483 VPWR 0.0605
R3543 VPWR.n439 VPWR 0.0605
R3544 VPWR VPWR.n502 0.0605
R3545 VPWR.n503 VPWR 0.0605
R3546 VPWR.n489 VPWR 0.0605
R3547 VPWR VPWR.n538 0.0605
R3548 VPWR.n539 VPWR 0.0605
R3549 VPWR.n546 VPWR 0.0605
R3550 VPWR.n515 VPWR 0.0605
R3551 VPWR VPWR.n560 0.0605
R3552 VPWR.n561 VPWR 0.0605
R3553 VPWR VPWR.n576 0.0605
R3554 VPWR.n577 VPWR 0.0605
R3555 VPWR.n584 VPWR 0.0605
R3556 VPWR.n552 VPWR 0.0605
R3557 VPWR VPWR.n9 0.0605
R3558 VPWR.n10 VPWR 0.0605
R3559 VPWR VPWR.n18 0.0605
R3560 VPWR.n19 VPWR 0.0605
R3561 VPWR VPWR.n592 0.0605
R3562 VPWR.n481 VPWR.n480 0.05675
R3563 VPWR.n268 VPWR.n267 0.056625
R3564 VPWR.n381 VPWR.n380 0.056625
R3565 VPWR.n113 VPWR.n112 0.0555
R3566 VPWR.n123 VPWR.n122 0.0555
R3567 VPWR.n468 VPWR.n467 0.0555
R3568 VPWR.n474 VPWR.n473 0.0555
R3569 VPWR.n83 VPWR.n82 0.05425
R3570 VPWR.n165 VPWR.n164 0.05425
R3571 VPWR.n202 VPWR.n201 0.05425
R3572 VPWR.n240 VPWR.n239 0.05425
R3573 VPWR.n428 VPWR.n427 0.05425
R3574 VPWR.n438 VPWR 0.05425
R3575 VPWR.n541 VPWR.n540 0.05425
R3576 VPWR.n579 VPWR.n578 0.05425
R3577 VPWR.n76 VPWR 0.0536485
R3578 VPWR.n233 VPWR 0.0536485
R3579 VPWR.n421 VPWR 0.0536485
R3580 VPWR.n449 VPWR 0.0536485
R3581 VPWR.n572 VPWR 0.0536485
R3582 VPWR.n79 VPWR.n78 0.05175
R3583 VPWR.n236 VPWR.n235 0.05175
R3584 VPWR.n424 VPWR.n423 0.05175
R3585 VPWR.n575 VPWR.n574 0.05175
R3586 VPWR.n53 VPWR.n25 0.0505
R3587 VPWR.n90 VPWR.n54 0.0505
R3588 VPWR.n108 VPWR.n107 0.0505
R3589 VPWR.n118 VPWR.n117 0.0505
R3590 VPWR.n135 VPWR.n92 0.0505
R3591 VPWR.n152 VPWR.n151 0.0505
R3592 VPWR.n172 VPWR.n137 0.0505
R3593 VPWR.n189 VPWR.n188 0.0505
R3594 VPWR.n209 VPWR.n174 0.0505
R3595 VPWR.n247 VPWR.n211 0.0505
R3596 VPWR.n264 VPWR.n263 0.0505
R3597 VPWR.n284 VPWR.n249 0.0505
R3598 VPWR.n335 VPWR.n311 0.0505
R3599 VPWR.n377 VPWR.n376 0.0505
R3600 VPWR.n397 VPWR.n362 0.0505
R3601 VPWR.n435 VPWR.n399 0.0505
R3602 VPWR.n463 VPWR.n462 0.0505
R3603 VPWR.n469 VPWR.n468 0.0505
R3604 VPWR.n511 VPWR.n487 0.0505
R3605 VPWR.n528 VPWR.n527 0.0505
R3606 VPWR.n548 VPWR.n513 0.0505
R3607 VPWR.n586 VPWR.n550 0.0505
R3608 VPWR.n590 VPWR.n589 0.0505
R3609 VPWR VPWR.n140 0.04925
R3610 VPWR VPWR.n177 0.04925
R3611 VPWR VPWR.n252 0.04925
R3612 VPWR VPWR.n365 0.04925
R3613 VPWR VPWR.n516 0.04925
R3614 VPWR.n90 VPWR.n89 0.0455
R3615 VPWR.n155 VPWR.n154 0.0455
R3616 VPWR.n158 VPWR.n157 0.0455
R3617 VPWR.n161 VPWR.n160 0.0455
R3618 VPWR.n172 VPWR.n171 0.0455
R3619 VPWR.n192 VPWR.n191 0.0455
R3620 VPWR.n195 VPWR.n194 0.0455
R3621 VPWR.n198 VPWR.n197 0.0455
R3622 VPWR.n209 VPWR.n208 0.0455
R3623 VPWR.n247 VPWR.n246 0.0455
R3624 VPWR.n309 VPWR.n308 0.0455
R3625 VPWR.n360 VPWR.n359 0.0455
R3626 VPWR.n435 VPWR.n434 0.0455
R3627 VPWR.n485 VPWR.n484 0.0455
R3628 VPWR.n531 VPWR.n530 0.0455
R3629 VPWR.n534 VPWR.n533 0.0455
R3630 VPWR.n537 VPWR.n536 0.0455
R3631 VPWR.n548 VPWR.n547 0.0455
R3632 VPWR.n586 VPWR.n585 0.0455
R3633 VPWR.n42 VPWR.n41 0.0448003
R3634 VPWR.n16 VPWR.n15 0.0448003
R3635 VPWR.n50 VPWR.n49 0.0423097
R3636 VPWR.n86 VPWR.n85 0.0423097
R3637 VPWR.n168 VPWR.n167 0.0423097
R3638 VPWR.n205 VPWR.n204 0.0423097
R3639 VPWR.n243 VPWR.n242 0.0423097
R3640 VPWR.n281 VPWR.n280 0.0423097
R3641 VPWR.n332 VPWR.n331 0.0423097
R3642 VPWR.n394 VPWR.n393 0.0423097
R3643 VPWR.n431 VPWR.n430 0.0423097
R3644 VPWR.n508 VPWR.n507 0.0423097
R3645 VPWR.n544 VPWR.n543 0.0423097
R3646 VPWR.n582 VPWR.n581 0.0423097
R3647 VPWR.n24 VPWR.n20 0.0423097
R3648 VPWR.n55 VPWR 0.04175
R3649 VPWR.n138 VPWR 0.04175
R3650 VPWR.n175 VPWR 0.04175
R3651 VPWR.n212 VPWR 0.04175
R3652 VPWR.n400 VPWR 0.04175
R3653 VPWR.n514 VPWR 0.04175
R3654 VPWR.n551 VPWR 0.04175
R3655 VPWR.n117 VPWR.n116 0.0405
R3656 VPWR.n126 VPWR.n125 0.0405
R3657 VPWR.n472 VPWR.n471 0.0405
R3658 VPWR.n478 VPWR.n477 0.0405
R3659 VPWR.n104 VPWR.n95 0.0355
R3660 VPWR.n114 VPWR.n113 0.0355
R3661 VPWR.n148 VPWR.n147 0.0355
R3662 VPWR.n185 VPWR.n184 0.0355
R3663 VPWR.n260 VPWR.n259 0.0355
R3664 VPWR.n373 VPWR.n372 0.0355
R3665 VPWR.n459 VPWR.n458 0.0355
R3666 VPWR.n465 VPWR.n464 0.0355
R3667 VPWR.n524 VPWR.n523 0.0355
R3668 VPWR.n481 VPWR.n437 0.03425
R3669 VPWR.n99 VPWR 0.033
R3670 VPWR.n98 VPWR 0.031
R3671 VPWR.n447 VPWR.n446 0.030637
R3672 VPWR.n101 VPWR.n100 0.028
R3673 VPWR.n32 VPWR 0.0263824
R3674 VPWR.n41 VPWR 0.0263824
R3675 VPWR.n49 VPWR 0.0263824
R3676 VPWR.n61 VPWR 0.0263824
R3677 VPWR.n85 VPWR 0.0263824
R3678 VPWR.n167 VPWR 0.0263824
R3679 VPWR.n204 VPWR 0.0263824
R3680 VPWR.n218 VPWR 0.0263824
R3681 VPWR.n242 VPWR 0.0263824
R3682 VPWR.n271 VPWR 0.0263824
R3683 VPWR.n280 VPWR 0.0263824
R3684 VPWR.n304 VPWR 0.0263824
R3685 VPWR.n331 VPWR 0.0263824
R3686 VPWR.n355 VPWR 0.0263824
R3687 VPWR.n384 VPWR 0.0263824
R3688 VPWR.n393 VPWR 0.0263824
R3689 VPWR.n406 VPWR 0.0263824
R3690 VPWR.n430 VPWR 0.0263824
R3691 VPWR.n507 VPWR 0.0263824
R3692 VPWR.n543 VPWR 0.0263824
R3693 VPWR.n557 VPWR 0.0263824
R3694 VPWR.n581 VPWR 0.0263824
R3695 VPWR.n6 VPWR 0.0263824
R3696 VPWR.n15 VPWR 0.0263824
R3697 VPWR.n24 VPWR 0.0263824
R3698 VPWR.n89 VPWR.n88 0.0255
R3699 VPWR.n121 VPWR.n120 0.0255
R3700 VPWR.n131 VPWR.n92 0.0255
R3701 VPWR.n162 VPWR.n161 0.0255
R3702 VPWR.n171 VPWR.n170 0.0255
R3703 VPWR.n199 VPWR.n198 0.0255
R3704 VPWR.n208 VPWR.n207 0.0255
R3705 VPWR.n246 VPWR.n245 0.0255
R3706 VPWR.n308 VPWR.n307 0.0255
R3707 VPWR.n326 VPWR.n325 0.0255
R3708 VPWR.n359 VPWR.n358 0.0255
R3709 VPWR.n434 VPWR.n433 0.0255
R3710 VPWR.n476 VPWR.n475 0.0255
R3711 VPWR.n484 VPWR.n483 0.0255
R3712 VPWR.n502 VPWR.n501 0.0255
R3713 VPWR.n538 VPWR.n537 0.0255
R3714 VPWR.n547 VPWR.n546 0.0255
R3715 VPWR.n585 VPWR.n584 0.0255
R3716 VPWR.n67 VPWR.n66 0.0205
R3717 VPWR.n110 VPWR.n109 0.0205
R3718 VPWR.n224 VPWR.n223 0.0205
R3719 VPWR.n412 VPWR.n411 0.0205
R3720 VPWR.n461 VPWR.n460 0.0205
R3721 VPWR.n477 VPWR 0.0205
R3722 VPWR.n563 VPWR.n562 0.0205
R3723 VPWR.n35 VPWR.n34 0.01925
R3724 VPWR.n44 VPWR.n43 0.01925
R3725 VPWR.n27 VPWR.n26 0.01925
R3726 VPWR.n64 VPWR.n63 0.01925
R3727 VPWR.n80 VPWR.n79 0.01925
R3728 VPWR.n56 VPWR.n55 0.01925
R3729 VPWR.n94 VPWR.n93 0.01925
R3730 VPWR.n151 VPWR.n150 0.01925
R3731 VPWR.n139 VPWR.n138 0.01925
R3732 VPWR.n188 VPWR.n187 0.01925
R3733 VPWR.n176 VPWR.n175 0.01925
R3734 VPWR.n221 VPWR.n220 0.01925
R3735 VPWR.n237 VPWR.n236 0.01925
R3736 VPWR.n213 VPWR.n212 0.01925
R3737 VPWR.n263 VPWR.n262 0.01925
R3738 VPWR.n275 VPWR.n274 0.01925
R3739 VPWR.n251 VPWR.n250 0.01925
R3740 VPWR.n300 VPWR.n298 0.01925
R3741 VPWR.n313 VPWR.n312 0.01925
R3742 VPWR.n351 VPWR.n349 0.01925
R3743 VPWR.n376 VPWR.n375 0.01925
R3744 VPWR.n388 VPWR.n387 0.01925
R3745 VPWR.n364 VPWR.n363 0.01925
R3746 VPWR.n409 VPWR.n408 0.01925
R3747 VPWR.n425 VPWR.n424 0.01925
R3748 VPWR.n401 VPWR.n400 0.01925
R3749 VPWR.n457 VPWR.n456 0.01925
R3750 VPWR.n489 VPWR.n488 0.01925
R3751 VPWR.n527 VPWR.n526 0.01925
R3752 VPWR.n515 VPWR.n514 0.01925
R3753 VPWR.n560 VPWR.n559 0.01925
R3754 VPWR.n576 VPWR.n575 0.01925
R3755 VPWR.n552 VPWR.n551 0.01925
R3756 VPWR.n9 VPWR.n8 0.01925
R3757 VPWR.n18 VPWR.n17 0.01925
R3758 VPWR.n592 VPWR.n0 0.01925
R3759 VPWR.n485 VPWR.n437 0.01675
R3760 VPWR.n74 VPWR.n73 0.0131337
R3761 VPWR.n231 VPWR.n230 0.0131337
R3762 VPWR.n419 VPWR.n418 0.0131337
R3763 VPWR.n570 VPWR.n569 0.0131337
R3764 VPWR.n452 VPWR.n451 0.012698
R3765 VPWR.n39 VPWR.n36 0.01175
R3766 VPWR.n46 VPWR.n45 0.01175
R3767 VPWR.n72 VPWR.n65 0.01175
R3768 VPWR.n83 VPWR.n81 0.01175
R3769 VPWR.n127 VPWR.n123 0.01175
R3770 VPWR.n165 VPWR.n163 0.01175
R3771 VPWR.n202 VPWR.n200 0.01175
R3772 VPWR.n229 VPWR.n222 0.01175
R3773 VPWR.n240 VPWR.n238 0.01175
R3774 VPWR.n269 VPWR.n265 0.01175
R3775 VPWR.n277 VPWR.n276 0.01175
R3776 VPWR.n328 VPWR.n327 0.01175
R3777 VPWR.n382 VPWR.n378 0.01175
R3778 VPWR.n390 VPWR.n389 0.01175
R3779 VPWR.n417 VPWR.n410 0.01175
R3780 VPWR.n428 VPWR.n426 0.01175
R3781 VPWR.n504 VPWR.n503 0.01175
R3782 VPWR.n541 VPWR.n539 0.01175
R3783 VPWR.n568 VPWR.n561 0.01175
R3784 VPWR.n579 VPWR.n577 0.01175
R3785 VPWR.n13 VPWR.n10 0.01175
R3786 VPWR.n22 VPWR.n19 0.01175
R3787 VPWR.n454 VPWR 0.0109554
R3788 VPWR.n97 VPWR.n96 0.0106712
R3789 VPWR.n443 VPWR.n442 0.0106712
R3790 VPWR.n135 VPWR 0.0105
R3791 VPWR VPWR.n152 0.0105
R3792 VPWR VPWR.n189 0.0105
R3793 VPWR VPWR.n264 0.0105
R3794 VPWR VPWR.n377 0.0105
R3795 VPWR VPWR.n528 0.0105
R3796 VPWR.n103 VPWR.n99 0.00878767
R3797 VPWR.n74 VPWR.n71 0.00790594
R3798 VPWR.n231 VPWR.n228 0.00790594
R3799 VPWR.n419 VPWR.n416 0.00790594
R3800 VPWR.n452 VPWR.n450 0.00790594
R3801 VPWR.n570 VPWR.n567 0.00790594
R3802 VPWR.n75 VPWR.n70 0.0074703
R3803 VPWR.n76 VPWR.n75 0.0074703
R3804 VPWR.n232 VPWR.n227 0.0074703
R3805 VPWR.n233 VPWR.n232 0.0074703
R3806 VPWR.n420 VPWR.n415 0.0074703
R3807 VPWR.n421 VPWR.n420 0.0074703
R3808 VPWR.n453 VPWR.n449 0.0074703
R3809 VPWR.n571 VPWR.n566 0.0074703
R3810 VPWR.n572 VPWR.n571 0.0074703
R3811 VPWR.n106 VPWR.n105 0.00675
R3812 VPWR.n274 VPWR.n273 0.00675
R3813 VPWR.n387 VPWR.n386 0.00675
R3814 VPWR.n439 VPWR.n438 0.00675
R3815 VPWR.n70 VPWR.n69 0.00659901
R3816 VPWR.n227 VPWR.n226 0.00659901
R3817 VPWR.n415 VPWR.n414 0.00659901
R3818 VPWR.n566 VPWR.n565 0.00659901
R3819 VPWR.n49 VPWR.n25 0.0055
R3820 VPWR.n85 VPWR.n54 0.0055
R3821 VPWR.n122 VPWR 0.0055
R3822 VPWR.n147 VPWR.n146 0.0055
R3823 VPWR.n167 VPWR.n137 0.0055
R3824 VPWR.n184 VPWR.n183 0.0055
R3825 VPWR.n204 VPWR.n174 0.0055
R3826 VPWR.n242 VPWR.n211 0.0055
R3827 VPWR.n259 VPWR.n258 0.0055
R3828 VPWR.n280 VPWR.n249 0.0055
R3829 VPWR.n331 VPWR.n311 0.0055
R3830 VPWR.n372 VPWR.n371 0.0055
R3831 VPWR.n393 VPWR.n362 0.0055
R3832 VPWR.n430 VPWR.n399 0.0055
R3833 VPWR.n507 VPWR.n487 0.0055
R3834 VPWR.n523 VPWR.n522 0.0055
R3835 VPWR.n543 VPWR.n513 0.0055
R3836 VPWR.n581 VPWR.n550 0.0055
R3837 VPWR.n590 VPWR.n24 0.0055
R3838 VPWR.n102 VPWR.n101 0.00426712
R3839 VPWR.n100 VPWR.n97 0.00313699
R3840 VPWR.n446 VPWR.n443 0.00313699
R3841 VPWR VPWR.n453 0.00311386
R3842 VPWR.n103 VPWR.n102 0.00276027
R3843 VPWR.n445 VPWR.n444 0.00276027
R3844 VPWR.n71 VPWR.n68 0.00175
R3845 VPWR.n129 VPWR.n126 0.00175
R3846 VPWR.n132 VPWR.n130 0.00175
R3847 VPWR.n145 VPWR.n144 0.00175
R3848 VPWR.n182 VPWR.n181 0.00175
R3849 VPWR.n228 VPWR.n225 0.00175
R3850 VPWR.n257 VPWR.n256 0.00175
R3851 VPWR.n370 VPWR.n369 0.00175
R3852 VPWR.n416 VPWR.n413 0.00175
R3853 VPWR.n450 VPWR.n441 0.00175
R3854 VPWR.n521 VPWR.n520 0.00175
R3855 VPWR.n567 VPWR.n564 0.00175
R3856 VPWR.n447 VPWR.n445 0.00163014
R3857 VPWR.n271 VPWR.n268 0.00162498
R3858 VPWR.n384 VPWR.n381 0.00162498
R3859 VPWR.n73 VPWR.n69 0.00115347
R3860 VPWR.n230 VPWR.n226 0.00115347
R3861 VPWR.n418 VPWR.n414 0.00115347
R3862 VPWR.n454 VPWR.n448 0.00115347
R3863 VPWR.n569 VPWR.n565 0.00115347
R3864 VPWR.n451 VPWR.n448 0.000935644
R3865 dr[1].n0 dr[1] 32.8039
R3866 dr[1].n0 dr[1].t0 4.95768
R3867 dr[1] dr[1].n0 0.148317
R3868 db[3].n0 db[3] 29.5303
R3869 db[3].n0 db[3].t0 4.95768
R3870 db[3] db[3].n0 0.148317
R3871 dr[4].n0 dr[4] 30.6127
R3872 dr[4].n0 dr[4].t0 4.95768
R3873 dr[4] dr[4].n0 0.148317
R3874 db[5].n0 db[5] 32.2759
R3875 db[5].n0 db[5].t0 4.95768
R3876 db[5] db[5].n0 0.148317
R3877 dr[6].n0 dr[6] 10.1791
R3878 dr[6].n0 dr[6].t0 4.95768
R3879 dr[6] dr[6].n0 0.148317
R3880 r[6].t0 r[6] 17.1634
R3881 r[6].n3 r[6].t0 17.0005
R3882 r[6].n10 r[6] 11.9744
R3883 r[6].n5 r[6].t3 8.52233
R3884 r[6].n7 r[6].t1 8.5005
R3885 r[6].n11 r[6].t2 8.5005
R3886 r[6].n0 r[6].t7 6.31247
R3887 r[6].n2 r[6].t5 5.79041
R3888 r[6].n0 r[6].t6 5.78997
R3889 r[6].n1 r[6].t4 5.78997
R3890 r[6].n6 r[6] 1.48874
R3891 r[6].n9 r[6] 0.828735
R3892 r[6].n1 r[6].n0 0.523
R3893 r[6].n2 r[6].n1 0.523
R3894 r[6].n5 r[6] 0.514393
R3895 r[6].n12 r[6].n4 0.492265
R3896 r[6].n6 r[6].n5 0.492265
R3897 r[6].n9 r[6].n8 0.492265
R3898 r[6].n4 r[6].n2 0.396077
R3899 r[6].n8 r[6] 0.3405
R3900 r[6] r[6].n12 0.171798
R3901 r[6].n4 r[6] 0.168735
R3902 r[6].n12 r[6].n11 0.0223321
R3903 r[6].n7 r[6].n6 0.0221667
R3904 r[6].n8 r[6].n7 0.0221667
R3905 r[6].n10 r[6].n9 0.0214924
R3906 r[6].n3 r[6] 0.0195385
R3907 r[6].n4 r[6].n3 0.0174231
R3908 r[6].n11 r[6].n10 0.00133969
R3909 b[3].n9 b[3] 12.1214
R3910 b[3].n7 b[3].t0 8.56366
R3911 b[3].n0 b[3].t2 8.52233
R3912 b[3].n2 b[3].t1 8.5005
R3913 b[3].n5 b[3].t3 8.5005
R3914 b[3].n8 b[3].t6 6.31291
R3915 b[3].n8 b[3].t7 5.79041
R3916 b[3].n11 b[3].t4 5.79041
R3917 b[3].n9 b[3].t5 5.60428
R3918 b[3].n1 b[3] 1.48874
R3919 b[3].n4 b[3] 0.828735
R3920 b[3].n11 b[3].n10 0.523
R3921 b[3].n10 b[3].n8 0.523
R3922 b[3].n0 b[3] 0.514393
R3923 b[3].n1 b[3].n0 0.492265
R3924 b[3].n4 b[3].n3 0.492265
R3925 b[3].n7 b[3].n6 0.492265
R3926 b[3] b[3].n11 0.360115
R3927 b[3].n3 b[3] 0.3405
R3928 b[3].n10 b[3].n9 0.186974
R3929 b[3].n6 b[3] 0.171798
R3930 b[3].n7 b[3] 0.168735
R3931 b[3] b[3].n7 0.0364615
R3932 b[3].n5 b[3].n4 0.0223321
R3933 b[3].n6 b[3].n5 0.0223321
R3934 b[3].n2 b[3].n1 0.0221667
R3935 b[3].n3 b[3].n2 0.0221667
R3936 r[5].n9 r[5] 10.8542
R3937 r[5].n7 r[5].t0 8.56366
R3938 r[5].n0 r[5].t2 8.52233
R3939 r[5].n2 r[5].t1 8.5005
R3940 r[5].n5 r[5].t3 8.5005
R3941 r[5].n8 r[5].t6 6.31291
R3942 r[5].n8 r[5].t5 5.79041
R3943 r[5].n11 r[5].t4 5.79041
R3944 r[5].n9 r[5].t7 5.60428
R3945 r[5].n1 r[5] 1.48874
R3946 r[5].n4 r[5] 0.828735
R3947 r[5].n11 r[5].n10 0.523
R3948 r[5].n10 r[5].n8 0.523
R3949 r[5].n0 r[5] 0.514393
R3950 r[5].n1 r[5].n0 0.492265
R3951 r[5].n4 r[5].n3 0.492265
R3952 r[5].n7 r[5].n6 0.492265
R3953 r[5] r[5].n11 0.360115
R3954 r[5].n3 r[5] 0.3405
R3955 r[5].n10 r[5].n9 0.186974
R3956 r[5].n6 r[5] 0.171798
R3957 r[5].n7 r[5] 0.168735
R3958 r[5] r[5].n7 0.0364615
R3959 r[5].n5 r[5].n4 0.0223321
R3960 r[5].n6 r[5].n5 0.0223321
R3961 r[5].n2 r[5].n1 0.0221667
R3962 r[5].n3 r[5].n2 0.0221667
R3963 r[1].n9 r[1] 11.0654
R3964 r[1].n7 r[1].t1 8.56366
R3965 r[1].n0 r[1].t2 8.52233
R3966 r[1].n2 r[1].t0 8.5005
R3967 r[1].n5 r[1].t3 8.5005
R3968 r[1].n8 r[1].t5 6.31291
R3969 r[1].n8 r[1].t7 5.79041
R3970 r[1].n11 r[1].t6 5.79041
R3971 r[1].n9 r[1].t4 5.60428
R3972 r[1].n1 r[1] 1.48874
R3973 r[1].n4 r[1] 0.828735
R3974 r[1].n11 r[1].n10 0.523
R3975 r[1].n10 r[1].n8 0.523
R3976 r[1].n0 r[1] 0.514393
R3977 r[1].n1 r[1].n0 0.492265
R3978 r[1].n4 r[1].n3 0.492265
R3979 r[1].n7 r[1].n6 0.492265
R3980 r[1] r[1].n11 0.360115
R3981 r[1].n3 r[1] 0.3405
R3982 r[1].n10 r[1].n9 0.186974
R3983 r[1].n6 r[1] 0.171798
R3984 r[1].n7 r[1] 0.168735
R3985 r[1] r[1].n7 0.0364615
R3986 r[1].n5 r[1].n4 0.0223321
R3987 r[1].n6 r[1].n5 0.0223321
R3988 r[1].n2 r[1].n1 0.0221667
R3989 r[1].n3 r[1].n2 0.0221667
R3990 b[1].n9 b[1] 11.4878
R3991 b[1].n7 b[1].t0 8.56366
R3992 b[1].n0 b[1].t2 8.52233
R3993 b[1].n2 b[1].t1 8.5005
R3994 b[1].n5 b[1].t3 8.5005
R3995 b[1].n8 b[1].t5 6.31291
R3996 b[1].n8 b[1].t4 5.79041
R3997 b[1].n11 b[1].t6 5.79041
R3998 b[1].n9 b[1].t7 5.60428
R3999 b[1].n1 b[1] 1.48874
R4000 b[1].n4 b[1] 0.828735
R4001 b[1].n11 b[1].n10 0.523
R4002 b[1].n10 b[1].n8 0.523
R4003 b[1].n0 b[1] 0.514393
R4004 b[1].n1 b[1].n0 0.492265
R4005 b[1].n4 b[1].n3 0.492265
R4006 b[1].n7 b[1].n6 0.492265
R4007 b[1] b[1].n11 0.360115
R4008 b[1].n3 b[1] 0.3405
R4009 b[1].n10 b[1].n9 0.186974
R4010 b[1].n6 b[1] 0.171798
R4011 b[1].n7 b[1] 0.168735
R4012 b[1] b[1].n7 0.0364615
R4013 b[1].n5 b[1].n4 0.0223321
R4014 b[1].n6 b[1].n5 0.0223321
R4015 b[1].n2 b[1].n1 0.0221667
R4016 b[1].n3 b[1].n2 0.0221667
R4017 g[6].t3 g[6] 17.1634
R4018 g[6].n3 g[6].t3 17.0005
R4019 g[6].n10 g[6] 10.7072
R4020 g[6].n5 g[6].t0 8.52233
R4021 g[6].n7 g[6].t2 8.5005
R4022 g[6].n11 g[6].t1 8.5005
R4023 g[6].n0 g[6].t4 6.31247
R4024 g[6].n2 g[6].t7 5.79041
R4025 g[6].n0 g[6].t6 5.78997
R4026 g[6].n1 g[6].t5 5.78997
R4027 g[6].n6 g[6] 1.48874
R4028 g[6].n9 g[6] 0.828735
R4029 g[6].n1 g[6].n0 0.523
R4030 g[6].n2 g[6].n1 0.523
R4031 g[6].n5 g[6] 0.514393
R4032 g[6].n12 g[6].n4 0.492265
R4033 g[6].n6 g[6].n5 0.492265
R4034 g[6].n9 g[6].n8 0.492265
R4035 g[6].n4 g[6].n2 0.396077
R4036 g[6].n8 g[6] 0.3405
R4037 g[6] g[6].n12 0.171798
R4038 g[6].n4 g[6] 0.168735
R4039 g[6].n12 g[6].n11 0.0223321
R4040 g[6].n7 g[6].n6 0.0221667
R4041 g[6].n8 g[6].n7 0.0221667
R4042 g[6].n10 g[6].n9 0.0214924
R4043 g[6].n3 g[6] 0.0195385
R4044 g[6].n4 g[6].n3 0.0174231
R4045 g[6].n11 g[6].n10 0.00133969
R4046 g[1].n9 g[1] 10.8542
R4047 g[1].n7 g[1].t1 8.56366
R4048 g[1].n0 g[1].t0 8.52233
R4049 g[1].n2 g[1].t3 8.5005
R4050 g[1].n5 g[1].t2 8.5005
R4051 g[1].n8 g[1].t4 6.31291
R4052 g[1].n8 g[1].t6 5.79041
R4053 g[1].n11 g[1].t7 5.79041
R4054 g[1].n9 g[1].t5 5.60428
R4055 g[1].n1 g[1] 1.48874
R4056 g[1].n4 g[1] 0.828735
R4057 g[1].n11 g[1].n10 0.523
R4058 g[1].n10 g[1].n8 0.523
R4059 g[1].n0 g[1] 0.514393
R4060 g[1].n1 g[1].n0 0.492265
R4061 g[1].n4 g[1].n3 0.492265
R4062 g[1].n7 g[1].n6 0.492265
R4063 g[1] g[1].n11 0.360115
R4064 g[1].n3 g[1] 0.3405
R4065 g[1].n10 g[1].n9 0.186974
R4066 g[1].n6 g[1] 0.171798
R4067 g[1].n7 g[1] 0.168735
R4068 g[1] g[1].n7 0.0364615
R4069 g[1].n5 g[1].n4 0.0223321
R4070 g[1].n6 g[1].n5 0.0223321
R4071 g[1].n2 g[1].n1 0.0221667
R4072 g[1].n3 g[1].n2 0.0221667
R4073 g[2].t2 g[2] 17.1634
R4074 g[2].n3 g[2].t2 17.0005
R4075 g[2].n10 g[2] 10.7072
R4076 g[2].n5 g[2].t1 8.52233
R4077 g[2].n7 g[2].t0 8.5005
R4078 g[2].n11 g[2].t3 8.5005
R4079 g[2].n0 g[2].t4 6.31247
R4080 g[2].n2 g[2].t5 5.79041
R4081 g[2].n0 g[2].t7 5.78997
R4082 g[2].n1 g[2].t6 5.78997
R4083 g[2].n6 g[2] 1.48874
R4084 g[2].n9 g[2] 0.828735
R4085 g[2].n1 g[2].n0 0.523
R4086 g[2].n2 g[2].n1 0.523
R4087 g[2].n5 g[2] 0.514393
R4088 g[2].n12 g[2].n4 0.492265
R4089 g[2].n6 g[2].n5 0.492265
R4090 g[2].n9 g[2].n8 0.492265
R4091 g[2].n4 g[2].n2 0.396077
R4092 g[2].n8 g[2] 0.3405
R4093 g[2] g[2].n12 0.171798
R4094 g[2].n4 g[2] 0.168735
R4095 g[2].n12 g[2].n11 0.0223321
R4096 g[2].n7 g[2].n6 0.0221667
R4097 g[2].n8 g[2].n7 0.0221667
R4098 g[2].n10 g[2].n9 0.0214924
R4099 g[2].n3 g[2] 0.0195385
R4100 g[2].n4 g[2].n3 0.0174231
R4101 g[2].n11 g[2].n10 0.00133969
R4102 b[2].t0 b[2] 17.1634
R4103 b[2].n3 b[2].t0 17.0005
R4104 b[2].n10 b[2] 10.7072
R4105 b[2].n5 b[2].t3 8.52233
R4106 b[2].n7 b[2].t1 8.5005
R4107 b[2].n11 b[2].t2 8.5005
R4108 b[2].n0 b[2].t7 6.31247
R4109 b[2].n2 b[2].t4 5.79041
R4110 b[2].n0 b[2].t5 5.78997
R4111 b[2].n1 b[2].t6 5.78997
R4112 b[2].n6 b[2] 1.48874
R4113 b[2].n9 b[2] 0.828735
R4114 b[2].n1 b[2].n0 0.523
R4115 b[2].n2 b[2].n1 0.523
R4116 b[2].n5 b[2] 0.514393
R4117 b[2].n12 b[2].n4 0.492265
R4118 b[2].n6 b[2].n5 0.492265
R4119 b[2].n9 b[2].n8 0.492265
R4120 b[2].n4 b[2].n2 0.396077
R4121 b[2].n8 b[2] 0.3405
R4122 b[2] b[2].n12 0.171798
R4123 b[2].n4 b[2] 0.168735
R4124 b[2].n12 b[2].n11 0.0223321
R4125 b[2].n7 b[2].n6 0.0221667
R4126 b[2].n8 b[2].n7 0.0221667
R4127 b[2].n10 b[2].n9 0.0214924
R4128 b[2].n3 b[2] 0.0195385
R4129 b[2].n4 b[2].n3 0.0174231
R4130 b[2].n11 b[2].n10 0.00133969
R4131 r[0].t1 r[0] 17.1634
R4132 r[0].n3 r[0].t1 17.0005
R4133 r[0].n10 r[0] 10.7072
R4134 r[0].n5 r[0].t2 8.52233
R4135 r[0].n7 r[0].t0 8.5005
R4136 r[0].n11 r[0].t3 8.5005
R4137 r[0].n0 r[0].t6 6.31247
R4138 r[0].n2 r[0].t4 5.79041
R4139 r[0].n0 r[0].t5 5.78997
R4140 r[0].n1 r[0].t7 5.78997
R4141 r[0].n6 r[0] 1.48874
R4142 r[0].n9 r[0] 0.828735
R4143 r[0].n1 r[0].n0 0.523
R4144 r[0].n2 r[0].n1 0.523
R4145 r[0].n5 r[0] 0.514393
R4146 r[0].n12 r[0].n4 0.492265
R4147 r[0].n6 r[0].n5 0.492265
R4148 r[0].n9 r[0].n8 0.492265
R4149 r[0].n4 r[0].n2 0.396077
R4150 r[0].n8 r[0] 0.3405
R4151 r[0] r[0].n12 0.171798
R4152 r[0].n4 r[0] 0.168735
R4153 r[0].n12 r[0].n11 0.0223321
R4154 r[0].n7 r[0].n6 0.0221667
R4155 r[0].n8 r[0].n7 0.0221667
R4156 r[0].n10 r[0].n9 0.0214924
R4157 r[0].n3 r[0] 0.0195385
R4158 r[0].n4 r[0].n3 0.0174231
R4159 r[0].n11 r[0].n10 0.00133969
R4160 r[7].n9 r[7] 10.8542
R4161 r[7].n7 r[7].t1 8.56366
R4162 r[7].n0 r[7].t2 8.52233
R4163 r[7].n2 r[7].t0 8.5005
R4164 r[7].n5 r[7].t3 8.5005
R4165 r[7].n8 r[7].t6 6.31291
R4166 r[7].n8 r[7].t4 5.79041
R4167 r[7].n11 r[7].t5 5.79041
R4168 r[7].n9 r[7].t7 5.60428
R4169 r[7].n1 r[7] 1.48874
R4170 r[7].n4 r[7] 0.828735
R4171 r[7].n11 r[7].n10 0.523
R4172 r[7].n10 r[7].n8 0.523
R4173 r[7].n0 r[7] 0.514393
R4174 r[7].n1 r[7].n0 0.492265
R4175 r[7].n4 r[7].n3 0.492265
R4176 r[7].n7 r[7].n6 0.492265
R4177 r[7] r[7].n11 0.360115
R4178 r[7].n3 r[7] 0.3405
R4179 r[7].n10 r[7].n9 0.186974
R4180 r[7].n6 r[7] 0.171798
R4181 r[7].n7 r[7] 0.168735
R4182 r[7] r[7].n7 0.0364615
R4183 r[7].n5 r[7].n4 0.0223321
R4184 r[7].n6 r[7].n5 0.0223321
R4185 r[7].n2 r[7].n1 0.0221667
R4186 r[7].n3 r[7].n2 0.0221667
R4187 dr[5].n0 dr[5] 11.9703
R4188 dr[5].n0 dr[5].t0 4.95768
R4189 dr[5] dr[5].n0 0.148317
R4190 db[7].n0 db[7] 33.7543
R4191 db[7].n0 db[7].t0 4.95768
R4192 db[7] db[7].n0 0.148317
R4193 b[6].t0 b[6] 17.1634
R4194 b[6].n3 b[6].t0 17.0005
R4195 b[6].n10 b[6] 11.9744
R4196 b[6].n5 b[6].t2 8.52233
R4197 b[6].n7 b[6].t3 8.5005
R4198 b[6].n11 b[6].t1 8.5005
R4199 b[6].n0 b[6].t6 6.31247
R4200 b[6].n2 b[6].t4 5.79041
R4201 b[6].n0 b[6].t5 5.78997
R4202 b[6].n1 b[6].t7 5.78997
R4203 b[6].n6 b[6] 1.48874
R4204 b[6].n9 b[6] 0.828735
R4205 b[6].n1 b[6].n0 0.523
R4206 b[6].n2 b[6].n1 0.523
R4207 b[6].n5 b[6] 0.514393
R4208 b[6].n12 b[6].n4 0.492265
R4209 b[6].n6 b[6].n5 0.492265
R4210 b[6].n9 b[6].n8 0.492265
R4211 b[6].n4 b[6].n2 0.396077
R4212 b[6].n8 b[6] 0.3405
R4213 b[6] b[6].n12 0.171798
R4214 b[6].n4 b[6] 0.168735
R4215 b[6].n12 b[6].n11 0.0223321
R4216 b[6].n7 b[6].n6 0.0221667
R4217 b[6].n8 b[6].n7 0.0221667
R4218 b[6].n10 b[6].n9 0.0214924
R4219 b[6].n3 b[6] 0.0195385
R4220 b[6].n4 b[6].n3 0.0174231
R4221 b[6].n11 b[6].n10 0.00133969
R4222 r[4].t2 r[4] 17.1634
R4223 r[4].n3 r[4].t2 17.0005
R4224 r[4].n10 r[4] 10.7072
R4225 r[4].n5 r[4].t3 8.52233
R4226 r[4].n7 r[4].t1 8.5005
R4227 r[4].n11 r[4].t0 8.5005
R4228 r[4].n0 r[4].t6 6.31247
R4229 r[4].n2 r[4].t4 5.79041
R4230 r[4].n0 r[4].t5 5.78997
R4231 r[4].n1 r[4].t7 5.78997
R4232 r[4].n6 r[4] 1.48874
R4233 r[4].n9 r[4] 0.828735
R4234 r[4].n1 r[4].n0 0.523
R4235 r[4].n2 r[4].n1 0.523
R4236 r[4].n5 r[4] 0.514393
R4237 r[4].n12 r[4].n4 0.492265
R4238 r[4].n6 r[4].n5 0.492265
R4239 r[4].n9 r[4].n8 0.492265
R4240 r[4].n4 r[4].n2 0.396077
R4241 r[4].n8 r[4] 0.3405
R4242 r[4] r[4].n12 0.171798
R4243 r[4].n4 r[4] 0.168735
R4244 r[4].n12 r[4].n11 0.0223321
R4245 r[4].n7 r[4].n6 0.0221667
R4246 r[4].n8 r[4].n7 0.0221667
R4247 r[4].n10 r[4].n9 0.0214924
R4248 r[4].n3 r[4] 0.0195385
R4249 r[4].n4 r[4].n3 0.0174231
R4250 r[4].n11 r[4].n10 0.00133969
R4251 dg[0].n0 dg[0] 30.4543
R4252 dg[0].n0 dg[0].t0 4.95768
R4253 dg[0] dg[0].n0 0.148317
R4254 b[7].n9 b[7] 10.8542
R4255 b[7].n7 b[7].t0 8.56366
R4256 b[7].n0 b[7].t3 8.52233
R4257 b[7].n2 b[7].t1 8.5005
R4258 b[7].n5 b[7].t2 8.5005
R4259 b[7].n8 b[7].t5 6.31291
R4260 b[7].n8 b[7].t7 5.79041
R4261 b[7].n11 b[7].t6 5.79041
R4262 b[7].n9 b[7].t4 5.60428
R4263 b[7].n1 b[7] 1.48874
R4264 b[7].n4 b[7] 0.828735
R4265 b[7].n11 b[7].n10 0.523
R4266 b[7].n10 b[7].n8 0.523
R4267 b[7].n0 b[7] 0.514393
R4268 b[7].n1 b[7].n0 0.492265
R4269 b[7].n4 b[7].n3 0.492265
R4270 b[7].n7 b[7].n6 0.492265
R4271 b[7] b[7].n11 0.360115
R4272 b[7].n3 b[7] 0.3405
R4273 b[7].n10 b[7].n9 0.186974
R4274 b[7].n6 b[7] 0.171798
R4275 b[7].n7 b[7] 0.168735
R4276 b[7] b[7].n7 0.0364615
R4277 b[7].n5 b[7].n4 0.0223321
R4278 b[7].n6 b[7].n5 0.0223321
R4279 b[7].n2 b[7].n1 0.0221667
R4280 b[7].n3 b[7].n2 0.0221667
R4281 db[6].n0 db[6] 31.9327
R4282 db[6].n0 db[6].t0 4.95768
R4283 db[6] db[6].n0 0.148317
R4284 db[0].n0 db[0] 11.8159
R4285 db[0].n0 db[0].t0 4.95768
R4286 db[0] db[0].n0 0.148317
R4287 g[0].t0 g[0] 17.1634
R4288 g[0].n3 g[0].t0 17.0005
R4289 g[0].n10 g[0] 11.9744
R4290 g[0].n5 g[0].t3 8.52233
R4291 g[0].n7 g[0].t1 8.5005
R4292 g[0].n11 g[0].t2 8.5005
R4293 g[0].n0 g[0].t7 6.31247
R4294 g[0].n2 g[0].t4 5.79041
R4295 g[0].n0 g[0].t5 5.78997
R4296 g[0].n1 g[0].t6 5.78997
R4297 g[0].n6 g[0] 1.48874
R4298 g[0].n9 g[0] 0.828735
R4299 g[0].n1 g[0].n0 0.523
R4300 g[0].n2 g[0].n1 0.523
R4301 g[0].n5 g[0] 0.514393
R4302 g[0].n12 g[0].n4 0.492265
R4303 g[0].n6 g[0].n5 0.492265
R4304 g[0].n9 g[0].n8 0.492265
R4305 g[0].n4 g[0].n2 0.396077
R4306 g[0].n8 g[0] 0.3405
R4307 g[0] g[0].n12 0.171798
R4308 g[0].n4 g[0] 0.168735
R4309 g[0].n12 g[0].n11 0.0223321
R4310 g[0].n7 g[0].n6 0.0221667
R4311 g[0].n8 g[0].n7 0.0221667
R4312 g[0].n10 g[0].n9 0.0214924
R4313 g[0].n3 g[0] 0.0195385
R4314 g[0].n4 g[0].n3 0.0174231
R4315 g[0].n11 g[0].n10 0.00133969
R4316 b[0].t2 b[0] 17.1634
R4317 b[0].n3 b[0].t2 17.0005
R4318 b[0].n10 b[0] 10.7072
R4319 b[0].n5 b[0].t1 8.52233
R4320 b[0].n7 b[0].t3 8.5005
R4321 b[0].n11 b[0].t0 8.5005
R4322 b[0].n0 b[0].t5 6.31247
R4323 b[0].n2 b[0].t6 5.79041
R4324 b[0].n0 b[0].t7 5.78997
R4325 b[0].n1 b[0].t4 5.78997
R4326 b[0].n6 b[0] 1.48874
R4327 b[0].n9 b[0] 0.828735
R4328 b[0].n1 b[0].n0 0.523
R4329 b[0].n2 b[0].n1 0.523
R4330 b[0].n5 b[0] 0.514393
R4331 b[0].n12 b[0].n4 0.492265
R4332 b[0].n6 b[0].n5 0.492265
R4333 b[0].n9 b[0].n8 0.492265
R4334 b[0].n4 b[0].n2 0.396077
R4335 b[0].n8 b[0] 0.3405
R4336 b[0] b[0].n12 0.171798
R4337 b[0].n4 b[0] 0.168735
R4338 b[0].n12 b[0].n11 0.0223321
R4339 b[0].n7 b[0].n6 0.0221667
R4340 b[0].n8 b[0].n7 0.0221667
R4341 b[0].n10 b[0].n9 0.0214924
R4342 b[0].n3 b[0] 0.0195385
R4343 b[0].n4 b[0].n3 0.0174231
R4344 b[0].n11 b[0].n10 0.00133969
R4345 g[5].n9 g[5] 10.8542
R4346 g[5].n7 g[5].t3 8.56366
R4347 g[5].n0 g[5].t0 8.52233
R4348 g[5].n2 g[5].t2 8.5005
R4349 g[5].n5 g[5].t1 8.5005
R4350 g[5].n8 g[5].t6 6.31291
R4351 g[5].n8 g[5].t4 5.79041
R4352 g[5].n11 g[5].t5 5.79041
R4353 g[5].n9 g[5].t7 5.60428
R4354 g[5].n1 g[5] 1.48874
R4355 g[5].n4 g[5] 0.828735
R4356 g[5].n11 g[5].n10 0.523
R4357 g[5].n10 g[5].n8 0.523
R4358 g[5].n0 g[5] 0.514393
R4359 g[5].n1 g[5].n0 0.492265
R4360 g[5].n4 g[5].n3 0.492265
R4361 g[5].n7 g[5].n6 0.492265
R4362 g[5] g[5].n11 0.360115
R4363 g[5].n3 g[5] 0.3405
R4364 g[5].n10 g[5].n9 0.186974
R4365 g[5].n6 g[5] 0.171798
R4366 g[5].n7 g[5] 0.168735
R4367 g[5] g[5].n7 0.0364615
R4368 g[5].n5 g[5].n4 0.0223321
R4369 g[5].n6 g[5].n5 0.0223321
R4370 g[5].n2 g[5].n1 0.0221667
R4371 g[5].n3 g[5].n2 0.0221667
R4372 g[3].n9 g[3] 12.1214
R4373 g[3].n7 g[3].t2 8.56366
R4374 g[3].n0 g[3].t1 8.52233
R4375 g[3].n2 g[3].t3 8.5005
R4376 g[3].n5 g[3].t0 8.5005
R4377 g[3].n8 g[3].t7 6.31291
R4378 g[3].n8 g[3].t6 5.79041
R4379 g[3].n11 g[3].t5 5.79041
R4380 g[3].n9 g[3].t4 5.60428
R4381 g[3].n1 g[3] 1.48874
R4382 g[3].n4 g[3] 0.828735
R4383 g[3].n11 g[3].n10 0.523
R4384 g[3].n10 g[3].n8 0.523
R4385 g[3].n0 g[3] 0.514393
R4386 g[3].n1 g[3].n0 0.492265
R4387 g[3].n4 g[3].n3 0.492265
R4388 g[3].n7 g[3].n6 0.492265
R4389 g[3] g[3].n11 0.360115
R4390 g[3].n3 g[3] 0.3405
R4391 g[3].n10 g[3].n9 0.186974
R4392 g[3].n6 g[3] 0.171798
R4393 g[3].n7 g[3] 0.168735
R4394 g[3] g[3].n7 0.0364615
R4395 g[3].n5 g[3].n4 0.0223321
R4396 g[3].n6 g[3].n5 0.0223321
R4397 g[3].n2 g[3].n1 0.0221667
R4398 g[3].n3 g[3].n2 0.0221667
R4399 db[4].n0 db[4] 30.4543
R4400 db[4].n0 db[4].t0 4.95768
R4401 db[4] db[4].n0 0.148317
R4402 b[4].t0 b[4] 17.1634
R4403 b[4].n3 b[4].t0 17.0005
R4404 b[4].n10 b[4] 11.9744
R4405 b[4].n5 b[4].t2 8.52233
R4406 b[4].n7 b[4].t1 8.5005
R4407 b[4].n11 b[4].t3 8.5005
R4408 b[4].n0 b[4].t6 6.31247
R4409 b[4].n2 b[4].t5 5.79041
R4410 b[4].n0 b[4].t4 5.78997
R4411 b[4].n1 b[4].t7 5.78997
R4412 b[4].n6 b[4] 1.48874
R4413 b[4].n9 b[4] 0.828735
R4414 b[4].n1 b[4].n0 0.523
R4415 b[4].n2 b[4].n1 0.523
R4416 b[4].n5 b[4] 0.514393
R4417 b[4].n12 b[4].n4 0.492265
R4418 b[4].n6 b[4].n5 0.492265
R4419 b[4].n9 b[4].n8 0.492265
R4420 b[4].n4 b[4].n2 0.396077
R4421 b[4].n8 b[4] 0.3405
R4422 b[4] b[4].n12 0.171798
R4423 b[4].n4 b[4] 0.168735
R4424 b[4].n12 b[4].n11 0.0223321
R4425 b[4].n7 b[4].n6 0.0221667
R4426 b[4].n8 b[4].n7 0.0221667
R4427 b[4].n10 b[4].n9 0.0214924
R4428 b[4].n3 b[4] 0.0195385
R4429 b[4].n4 b[4].n3 0.0174231
R4430 b[4].n11 b[4].n10 0.00133969
R4431 dg[2].n0 dg[2] 12.0975
R4432 dg[2].n0 dg[2].t0 4.95768
R4433 dg[2] dg[2].n0 0.148317
R4434 dr[7].n0 dr[7] 11.9703
R4435 dr[7].n0 dr[7].t0 4.95768
R4436 dr[7] dr[7].n0 0.148317
R4437 dg[4].n0 dg[4] 10.5487
R4438 dg[4].n0 dg[4].t0 4.95768
R4439 dg[4] dg[4].n0 0.148317
R4440 g[4].t2 g[4] 17.1634
R4441 g[4].n3 g[4].t2 17.0005
R4442 g[4].n10 g[4] 11.9744
R4443 g[4].n5 g[4].t1 8.52233
R4444 g[4].n7 g[4].t3 8.5005
R4445 g[4].n11 g[4].t0 8.5005
R4446 g[4].n0 g[4].t7 6.31247
R4447 g[4].n2 g[4].t4 5.79041
R4448 g[4].n0 g[4].t5 5.78997
R4449 g[4].n1 g[4].t6 5.78997
R4450 g[4].n6 g[4] 1.48874
R4451 g[4].n9 g[4] 0.828735
R4452 g[4].n1 g[4].n0 0.523
R4453 g[4].n2 g[4].n1 0.523
R4454 g[4].n5 g[4] 0.514393
R4455 g[4].n12 g[4].n4 0.492265
R4456 g[4].n6 g[4].n5 0.492265
R4457 g[4].n9 g[4].n8 0.492265
R4458 g[4].n4 g[4].n2 0.396077
R4459 g[4].n8 g[4] 0.3405
R4460 g[4] g[4].n12 0.171798
R4461 g[4].n4 g[4] 0.168735
R4462 g[4].n12 g[4].n11 0.0223321
R4463 g[4].n7 g[4].n6 0.0221667
R4464 g[4].n8 g[4].n7 0.0221667
R4465 g[4].n10 g[4].n9 0.0214924
R4466 g[4].n3 g[4] 0.0195385
R4467 g[4].n4 g[4].n3 0.0174231
R4468 g[4].n11 g[4].n10 0.00133969
R4469 dr[3].n0 dr[3] 30.2695
R4470 dr[3].n0 dr[3].t0 4.95768
R4471 dr[3] dr[3].n0 0.148317
R4472 r[3].n9 r[3] 12.1214
R4473 r[3].n7 r[3].t0 8.56366
R4474 r[3].n0 r[3].t3 8.52233
R4475 r[3].n2 r[3].t1 8.5005
R4476 r[3].n5 r[3].t2 8.5005
R4477 r[3].n8 r[3].t5 6.31291
R4478 r[3].n8 r[3].t7 5.79041
R4479 r[3].n11 r[3].t6 5.79041
R4480 r[3].n9 r[3].t4 5.60428
R4481 r[3].n1 r[3] 1.48874
R4482 r[3].n4 r[3] 0.828735
R4483 r[3].n11 r[3].n10 0.523
R4484 r[3].n10 r[3].n8 0.523
R4485 r[3].n0 r[3] 0.514393
R4486 r[3].n1 r[3].n0 0.492265
R4487 r[3].n4 r[3].n3 0.492265
R4488 r[3].n7 r[3].n6 0.492265
R4489 r[3] r[3].n11 0.360115
R4490 r[3].n3 r[3] 0.3405
R4491 r[3].n10 r[3].n9 0.186974
R4492 r[3].n6 r[3] 0.171798
R4493 r[3].n7 r[3] 0.168735
R4494 r[3] r[3].n7 0.0364615
R4495 r[3].n5 r[3].n4 0.0223321
R4496 r[3].n6 r[3].n5 0.0223321
R4497 r[3].n2 r[3].n1 0.0221667
R4498 r[3].n3 r[3].n2 0.0221667
R4499 db[1].n0 db[1] 10.6855
R4500 db[1].n0 db[1].t0 4.95768
R4501 db[1] db[1].n0 0.148317
R4502 dr[0].n0 dr[0] 33.5695
R4503 dr[0].n0 dr[0].t0 4.95768
R4504 dr[0] dr[0].n0 0.148317
R4505 dg[1].n0 dg[1] 31.1671
R4506 dg[1].n0 dg[1].t0 4.95768
R4507 dg[1] dg[1].n0 0.148317
R4508 dr[2].n0 dr[2] 30.8239
R4509 dr[2].n0 dr[2].t0 4.95768
R4510 dr[2] dr[2].n0 0.148317
R4511 dg[3].n0 dg[3] 10.3639
R4512 dg[3].n0 dg[3].t0 4.95768
R4513 dg[3] dg[3].n0 0.148317
R4514 r[2].t0 r[2] 17.1634
R4515 r[2].n3 r[2].t0 17.0005
R4516 r[2].n10 r[2] 11.9744
R4517 r[2].n5 r[2].t3 8.52233
R4518 r[2].n7 r[2].t1 8.5005
R4519 r[2].n11 r[2].t2 8.5005
R4520 r[2].n0 r[2].t7 6.31247
R4521 r[2].n2 r[2].t4 5.79041
R4522 r[2].n0 r[2].t5 5.78997
R4523 r[2].n1 r[2].t6 5.78997
R4524 r[2].n6 r[2] 1.48874
R4525 r[2].n9 r[2] 0.828735
R4526 r[2].n1 r[2].n0 0.523
R4527 r[2].n2 r[2].n1 0.523
R4528 r[2].n5 r[2] 0.514393
R4529 r[2].n12 r[2].n4 0.492265
R4530 r[2].n6 r[2].n5 0.492265
R4531 r[2].n9 r[2].n8 0.492265
R4532 r[2].n4 r[2].n2 0.396077
R4533 r[2].n8 r[2] 0.3405
R4534 r[2] r[2].n12 0.171798
R4535 r[2].n4 r[2] 0.168735
R4536 r[2].n12 r[2].n11 0.0223321
R4537 r[2].n7 r[2].n6 0.0221667
R4538 r[2].n8 r[2].n7 0.0221667
R4539 r[2].n10 r[2].n9 0.0214924
R4540 r[2].n3 r[2] 0.0195385
R4541 r[2].n4 r[2].n3 0.0174231
R4542 r[2].n11 r[2].n10 0.00133969
R4543 dg[5].n0 dg[5] 30.4279
R4544 dg[5].n0 dg[5].t0 4.95768
R4545 dg[5] dg[5].n0 0.148317
R4546 g[7].n9 g[7] 12.1214
R4547 g[7].n7 g[7].t2 8.56366
R4548 g[7].n0 g[7].t1 8.52233
R4549 g[7].n2 g[7].t3 8.5005
R4550 g[7].n5 g[7].t0 8.5005
R4551 g[7].n8 g[7].t5 6.31291
R4552 g[7].n8 g[7].t6 5.79041
R4553 g[7].n11 g[7].t7 5.79041
R4554 g[7].n9 g[7].t4 5.60428
R4555 g[7].n1 g[7] 1.48874
R4556 g[7].n4 g[7] 0.828735
R4557 g[7].n11 g[7].n10 0.523
R4558 g[7].n10 g[7].n8 0.523
R4559 g[7].n0 g[7] 0.514393
R4560 g[7].n1 g[7].n0 0.492265
R4561 g[7].n4 g[7].n3 0.492265
R4562 g[7].n7 g[7].n6 0.492265
R4563 g[7] g[7].n11 0.360115
R4564 g[7].n3 g[7] 0.3405
R4565 g[7].n10 g[7].n9 0.186974
R4566 g[7].n6 g[7] 0.171798
R4567 g[7].n7 g[7] 0.168735
R4568 g[7] g[7].n7 0.0364615
R4569 g[7].n5 g[7].n4 0.0223321
R4570 g[7].n6 g[7].n5 0.0223321
R4571 g[7].n2 g[7].n1 0.0221667
R4572 g[7].n3 g[7].n2 0.0221667
R4573 dg[7].n0 dg[7] 30.6391
R4574 dg[7].n0 dg[7].t0 4.95768
R4575 dg[7] dg[7].n0 0.148317
R4576 db[2].n0 db[2] 30.2431
R4577 db[2].n0 db[2].t0 4.95768
R4578 db[2] db[2].n0 0.148317
R4579 dg[6].n0 dg[6] 31.3519
R4580 dg[6].n0 dg[6].t0 4.95768
R4581 dg[6] dg[6].n0 0.148317
C0 b[6] db[7] 0.02006f
C1 VPWR a_320_4330# 0.0021f
C2 db[1] b[1] 0.00213f
C3 a_490_22762# r[1] 0.00183f
C4 dg[2] g[3] 0.002f
C5 a_1066_5376# a_1066_4618# 0.02326f
C6 a_1066_12178# dg[6] 0.00301f
C7 VPWR r[0] 1.3325f
C8 VPWR r[7] 1.8358f
C9 dr[4] dr[5] 0.08395f
C10 r[3] r[5] 0.00163f
C11 dr[4] a_490_18984# 0.00483f
C12 dr[6] a_1066_18226# 0.65532f
C13 VPWR b[6] 1.3707f
C14 dg[6] dg[7] 0.10089f
C15 VPWR g[2] 1.3431f
C16 VPWR db[1] 0.27457f
C17 VPWR a_320_10620# 0.00167f
C18 db[6] a_2240_4782# 0.00195f
C19 dr[1] r[1] 0.00217f
C20 dr[0] r[2] 0.01652f
C21 dg[0] g[0] 0.00828f
C22 a_1066_21250# dr[3] 0.00164f
C23 a_490_14448# a_490_13690# 0.02326f
C24 a_1066_12936# g[3] 1.15042f
C25 a_2152_22474# dr[1] 0.00251f
C26 a_490_10666# g[5] 0.00414f
C27 a_1066_4618# b[3] 0.00897f
C28 VPWR a_320_19902# 0.07562f
C29 dg[1] g[2] 0.00517f
C30 r[5] a_320_19106# 0.00425f
C31 db[7] b[7] 0.00444f
C32 db[6] db[3] 0.00961f
C33 b[1] db[2] 0.00201f
C34 dg[3] g[3] 0.00586f
C35 a_778_6888# db[0] 0.00754f
C36 a_328_22130# r[0] 0.00467f
C37 VPWR r[1] 1.84546f
C38 VPWR g[0] 1.3748f
C39 a_2240_20618# dr[0] 0.00171f
C40 VPWR a_2152_22474# 0.00121f
C41 r[4] r[5] 0.05597f
C42 r[3] a_1066_21250# 0.00135f
C43 a_2240_5498# db[3] 0.01808f
C44 a_1066_5376# db[1] 0.0013f
C45 dr[7] a_1066_18226# 0.01326f
C46 dr[5] a_490_18984# 0.64976f
C47 a_490_19738# a_320_19902# 0.01277f
C48 VPWR b[7] 1.8358f
C49 VPWR db[2] 0.52754f
C50 VPWR g[3] 2.00084f
C51 VPWR a_320_13644# 0.00167f
C52 dr[1] r[2] 0.00241f
C53 VPWR a_320_11890# 0.0021f
C54 g[0] dg[1] 0.00363f
C55 a_320_13854# g[2] 0.00406f
C56 a_1066_12936# g[4] 0.00126f
C57 a_586_22008# dr[0] 0.01859f
C58 a_490_7642# db[0] 0.67355f
C59 a_490_10666# g[6] 1.15206f
C60 a_1066_20496# dr[0] 0.01316f
C61 a_490_11424# g[4] 0.02529f
C62 a_1066_4618# b[4] 1.15154f
C63 r[4] a_320_19450# 0.00117f
C64 a_1066_3106# b[4] 0.00157f
C65 db[7] db[3] 0.00474f
C66 b[5] b[4] 0.06698f
C67 db[6] db[4] 0.0911f
C68 VPWR a_2240_4782# 0.0641f
C69 g[7] g[6] 0.04801f
C70 db[2] b[2] 0.00957f
C71 a_490_22762# a_586_22008# 0.02155f
C72 a_1066_5376# a_2240_5842# 0.0017f
C73 a_778_6888# db[1] 0.64255f
C74 a_328_22130# r[1] 0.013f
C75 a_490_13690# dg[2] 0.66099f
C76 a_320_3986# b[4] 0.00128f
C77 VPWR r[2] 1.37586f
C78 a_2240_20618# dr[1] 0.0064f
C79 dr[4] dr[0] 0.00147f
C80 dr[5] dr[6] 0.06337f
C81 a_1066_21250# a_2240_21204# 0.0017f
C82 a_2240_5498# db[4] 0.00165f
C83 a_1066_5376# db[2] 0.00861f
C84 a_490_3864# b[4] 0.02529f
C85 VPWR db[3] 0.26027f
C86 dg[0] a_2240_15366# 0.01778f
C87 VPWR g[4] 1.36503f
C88 a_1066_3106# a_2240_3060# 0.0017f
C89 dr[2] r[2] 0.00223f
C90 a_320_4330# b[4] 0.00117f
C91 a_586_22008# dr[1] 0.64209f
C92 a_320_14570# g[1] 0.00425f
C93 a_490_11424# g[5] 1.15098f
C94 a_490_13690# a_1066_12936# 0.0063f
C95 a_1066_20496# dr[1] 0.02158f
C96 a_1066_9912# a_2240_10034# 0.0073f
C97 VPWR a_2240_20618# 0.06455f
C98 db[7] a_490_2352# 0.64766f
C99 a_490_6130# db[2] 0.66955f
C100 VPWR a_1066_18226# 1.01815f
C101 db[6] db[5] 0.86735f
C102 b[6] b[4] 0.01758f
C103 db[7] db[4] 0.09382f
C104 a_320_10830# g[6] 0.00406f
C105 VPWR a_2240_15366# 0.06525f
C106 dg[4] g[4] 0.00781f
C107 db[2] b[3] 0.00287f
C108 b[2] db[3] 0.00213f
C109 VPWR a_320_2474# 0.07622f
C110 a_778_6888# db[2] 0.02325f
C111 a_328_22474# r[0] 0.0041f
C112 a_2240_20618# dr[2] 0.00165f
C113 dr[5] dr[7] 0.00806f
C114 r[5] r[6] 0.02576f
C115 VPWR a_586_22008# 1.10011f
C116 a_2240_5498# db[5] 0.00507f
C117 VPWR a_490_2352# 1.1249f
C118 a_1066_5376# db[3] 0.66185f
C119 a_490_10666# g[7] 0.00439f
C120 VPWR a_1066_20496# 1.00693f
C121 VPWR db[4] 0.23403f
C122 VPWR g[5] 1.82849f
C123 VPWR a_320_2818# 0.0021f
C124 VPWR a_490_13690# 1.12103f
C125 a_1066_18226# a_2240_18390# 0.0073f
C126 VPWR a_2240_12342# 0.06422f
C127 a_490_11424# g[6] 0.00126f
C128 a_1066_20496# dr[2] 0.00305f
C129 VPWR dr[4] 0.34867f
C130 r[4] a_320_19902# 0.00406f
C131 a_1066_20496# a_490_19738# 0.00532f
C132 a_490_10666# a_1066_9912# 0.0063f
C133 a_490_6130# db[3] 0.00438f
C134 g[0] a_1066_15202# 1.15166f
C135 dg[1] a_490_13690# 0.01355f
C136 r[6] a_490_17472# 0.02529f
C137 db[7] db[5] 0.07748f
C138 db[3] b[3] 0.00751f
C139 g[4] dg[5] 0.0105f
C140 db[6] a_2240_3270# 0.01809f
C141 a_328_22474# r[1] 0.002f
C142 a_586_22008# a_328_22130# 0.01205f
C143 a_2240_12342# dg[4] 0.02153f
C144 a_2240_20618# dr[3] 0.01725f
C145 a_1066_9912# g[7] 1.15042f
C146 r[3] r[2] 0.08922f
C147 dr[6] dr[7] 0.0645f
C148 a_2240_13058# dg[2] 0.00171f
C149 a_1066_5376# db[4] 0.00873f
C150 a_490_10666# a_320_10830# 0.01277f
C151 dr[4] a_490_19738# 0.64761f
C152 a_1066_20496# a_2240_20962# 0.0017f
C153 a_1066_4618# a_1066_3106# 0.00243f
C154 VPWR db[5] 0.39582f
C155 g[0] a_320_14570# 0.00128f
C156 VPWR g[6] 1.34345f
C157 VPWR a_2240_10034# 0.06525f
C158 a_490_13690# a_320_13854# 0.01277f
C159 a_1066_20496# dr[3] 0.6657f
C160 a_1066_12178# g[3] 0.00897f
C161 a_2240_21414# dr[1] 0.00165f
C162 b[5] a_320_3986# 0.00425f
C163 a_1066_4618# a_490_3864# 0.0063f
C164 a_1066_12936# a_2240_13058# 0.0073f
C165 g[0] a_320_14914# 0.00117f
C166 VPWR dr[5] 0.47656f
C167 dg[0] a_490_14448# 0.00422f
C168 r[7] a_490_17472# 1.15098f
C169 VPWR a_490_18984# 1.11142f
C170 a_490_3864# a_1066_3106# 0.00532f
C171 b[5] a_490_3864# 1.15098f
C172 a_490_11424# a_490_10666# 0.02326f
C173 VPWR a_320_17594# 0.07622f
C174 dg[5] g[5] 0.0034f
C175 g[4] dg[6] 0.00184f
C176 b[3] db[4] 0.00221f
C177 a_320_22926# r[0] 0.00406f
C178 a_490_3864# a_320_3986# 0.01277f
C179 dr[4] dr[3] 0.24848f
C180 a_2240_12342# dg[5] 0.0024f
C181 a_2240_13058# dg[3] 0.02318f
C182 r[6] r[7] 0.06698f
C183 VPWR a_320_22716# 0.00167f
C184 a_1066_5376# db[5] 0.01683f
C185 VPWR a_2240_21414# 0.06364f
C186 r[3] a_1066_20496# 1.15042f
C187 a_490_19738# a_490_18984# 0.02591f
C188 VPWR a_2240_3270# 0.06515f
C189 VPWR a_490_14448# 1.12096f
C190 b[6] a_1066_3106# 1.15166f
C191 b[5] b[6] 0.02576f
C192 VPWR a_2240_13058# 0.06422f
C193 a_490_22762# dr[0] 0.64761f
C194 db[0] db[1] 0.07594f
C195 g[1] g[2] 0.02795f
C196 a_1066_12178# g[4] 1.15154f
C197 VPWR a_490_10666# 1.12103f
C198 a_1066_15202# a_2240_15366# 0.0073f
C199 a_2152_22130# dr[0] 0.00224f
C200 a_2240_21414# dr[2] 0.02098f
C201 VPWR dr[6] 0.23226f
C202 r[3] dr[4] 0.00596f
C203 dg[1] a_490_14448# 0.65445f
C204 b[6] a_490_3864# 0.00436f
C205 b[3] db[5] 0.00452f
C206 db[4] b[4] 0.00199f
C207 g[5] dg[6] 0.01042f
C208 VPWR g[7] 2.02f
C209 dr[0] dr[1] 0.46489f
C210 a_1066_12936# dg[2] 0.02091f
C211 g[0] g[1] 0.06698f
C212 dr[6] a_2240_18390# 0.02264f
C213 db[6] db[7] 1.18306f
C214 VPWR a_1066_9912# 1.01188f
C215 b[0] b[1] 0.04703f
C216 db[0] db[2] 0.00207f
C217 dg[2] dg[3] 0.07094f
C218 a_2152_22130# dr[1] 0.01286f
C219 VPWR dr[0] 0.42298f
C220 VPWR dr[7] 0.34015f
C221 dr[4] r[4] 0.00466f
C222 a_1066_12178# a_2240_12342# 0.0073f
C223 VPWR a_320_19692# 0.00167f
C224 r[3] a_490_18984# 0.00297f
C225 a_1066_4618# a_2240_4782# 0.0073f
C226 VPWR db[6] 0.31727f
C227 VPWR a_320_10830# 0.07532f
C228 b[4] db[5] 0.00414f
C229 dg[6] g[6] 0.00957f
C230 g[5] dg[7] 0.00129f
C231 VPWR b[0] 1.34042f
C232 VPWR dg[2] 0.26735f
C233 VPWR a_320_17938# 0.0021f
C234 dr[0] dr[2] 0.072f
C235 r[0] r[1] 0.05203f
C236 a_1066_12936# dg[3] 0.67444f
C237 a_1066_21250# r[2] 1.15166f
C238 VPWR a_490_22762# 1.10943f
C239 VPWR a_2240_5498# 0.06421f
C240 a_490_10666# dg[5] 0.00119f
C241 VPWR a_2152_22130# 0.15108f
C242 a_1066_4618# db[3] 0.00114f
C243 g[0] g[2] 0.00164f
C244 dg[1] dg[2] 0.46545f
C245 a_490_18984# a_320_19106# 0.01277f
C246 b[6] b[7] 0.06698f
C247 VPWR a_1066_12936# 1.00776f
C248 db[1] db[2] 0.09781f
C249 g[2] g[3] 0.04801f
C250 a_1066_18226# a_490_17472# 0.0063f
C251 db[7] a_2240_4572# 0.00202f
C252 VPWR a_490_11424# 1.12097f
C253 a_2152_22130# dr[2] 0.00183f
C254 a_320_13644# g[2] 0.00243f
C255 VPWR dr[1] 0.3574f
C256 a_320_11546# g[4] 0.00128f
C257 a_2240_20962# dr[0] 0.00203f
C258 VPWR dg[0] 0.35563f
C259 dr[4] r[5] 0.00199f
C260 db[6] a_1066_5376# 0.0026f
C261 r[6] a_1066_18226# 1.15166f
C262 r[4] a_490_18984# 0.00943f
C263 VPWR db[7] 0.42772f
C264 VPWR b[1] 1.92816f
C265 g[6] dg[7] 0.00213f
C266 VPWR dg[3] 0.24318f
C267 a_1066_5376# a_2240_5498# 0.0073f
C268 dr[1] dr[2] 0.80225f
C269 dr[0] dr[3] 0.03854f
C270 a_2240_10034# dg[7] 0.01774f
C271 a_1066_15202# a_490_14448# 0.0063f
C272 dg[0] dg[1] 0.11715f
C273 a_1066_12936# dg[4] 0.00171f
C274 a_586_22008# a_1066_21250# 0.00713f
C275 a_490_10666# dg[6] 0.66522f
C276 a_1066_21250# a_1066_20496# 0.02591f
C277 a_1066_4618# db[4] 0.64051f
C278 a_1066_3106# a_490_2352# 0.0063f
C279 dg[0] a_2240_15156# 0.00101f
C280 g[7] dg[6] 0.00287f
C281 b[1] b[2] 0.03406f
C282 dg[2] dg[5] 0.00336f
C283 dg[3] dg[4] 0.06652f
C284 a_778_6888# b[0] 0.00191f
C285 a_490_14448# a_320_14570# 0.01277f
C286 a_490_13690# g[1] 0.00414f
C287 a_320_11546# g[5] 0.00425f
C288 VPWR dr[2] 0.25226f
C289 a_2240_20962# dr[1] 0.00112f
C290 VPWR dg[1] 0.45075f
C291 dr[5] r[5] 0.00895f
C292 a_490_3864# a_490_2352# 0.00188f
C293 a_320_7596# b[0] 0.00243f
C294 VPWR a_490_19738# 1.1119f
C295 r[5] a_490_18984# 1.15098f
C296 VPWR b[2] 1.34342f
C297 VPWR a_2240_18390# 0.06525f
C298 VPWR dg[4] 0.26497f
C299 a_320_7806# b[0] 0.00406f
C300 r[1] r[2] 0.0313f
C301 dr[1] dr[3] 0.18994f
C302 a_1066_9912# dg[6] 0.00816f
C303 a_586_22008# r[0] 0.00649f
C304 b[6] a_320_2474# 0.00128f
C305 VPWR a_1066_5376# 1.00736f
C306 a_490_10666# dg[7] 0.00535f
C307 a_490_7642# b[0] 1.15184f
C308 a_490_11424# dg[5] 0.64029f
C309 VPWR a_328_22130# 0.14967f
C310 a_1066_4618# db[5] 0.01394f
C311 a_2240_5842# db[3] 0.00141f
C312 b[6] a_490_2352# 0.02529f
C313 a_490_6130# b[1] 0.01153f
C314 VPWR a_320_6084# 0.00167f
C315 a_1066_3106# db[5] 0.01158f
C316 db[6] b[4] 0.01058f
C317 b[5] db[5] 0.00213f
C318 b[1] b[3] 0.00814f
C319 VPWR a_320_13854# 0.07532f
C320 g[7] dg[7] 0.00751f
C321 db[2] db[3] 0.07209f
C322 g[3] g[4] 0.06684f
C323 a_490_18984# a_490_17472# 0.00188f
C324 a_1066_18226# a_2240_18180# 0.0017f
C325 b[6] a_320_2818# 0.00117f
C326 VPWR a_320_6294# 0.07626f
C327 a_778_6888# b[1] 1.15043f
C328 a_490_13690# g[2] 1.15206f
C329 a_490_17472# a_320_17594# 0.01277f
C330 VPWR dr[3] 0.32417f
C331 r[3] dr[1] 0.00554f
C332 a_320_11890# g[4] 0.00117f
C333 dr[5] r[6] 0.00379f
C334 a_2240_21204# dr[0] 0.00117f
C335 VPWR a_490_6130# 1.1286f
C336 r[4] a_320_19692# 0.00243f
C337 r[6] a_490_18984# 0.00436f
C338 a_490_3864# db[5] 0.64209f
C339 VPWR b[3] 2.00047f
C340 VPWR dg[5] 0.30967f
C341 r[6] a_320_17594# 0.00128f
C342 VPWR a_778_6888# 1.09781f
C343 a_320_6084# b[2] 0.00243f
C344 dr[2] dr[3] 0.15884f
C345 a_1066_9912# dg[7] 0.66117f
C346 a_586_22008# r[1] 1.15098f
C347 b[7] a_320_2474# 0.00425f
C348 a_320_6294# b[2] 0.00406f
C349 VPWR a_320_7596# 0.00167f
C350 a_490_7642# b[1] 0.00311f
C351 a_490_11424# dg[6] 0.04561f
C352 a_490_19738# dr[3] 0.00671f
C353 a_1066_21250# a_2240_21414# 0.0073f
C354 a_2240_5842# db[4] 0.00111f
C355 VPWR r[3] 1.99159f
C356 b[7] a_490_2352# 1.15098f
C357 VPWR a_320_7806# 0.07622f
C358 a_490_6130# b[2] 1.15206f
C359 dg[0] a_1066_15202# 0.66113f
C360 g[0] a_490_13690# 0.00294f
C361 b[6] db[5] 0.00379f
C362 db[7] b[4] 0.00709f
C363 b[2] b[3] 0.04801f
C364 dg[4] dg[5] 0.08036f
C365 a_1066_3106# a_2240_3270# 0.0073f
C366 VPWR a_490_7642# 1.11542f
C367 a_320_10620# g[6] 0.00243f
C368 a_490_13690# g[3] 0.00439f
C369 a_490_14448# g[1] 1.15098f
C370 a_490_6130# a_1066_5376# 0.0063f
C371 dr[6] r[6] 0.00371f
C372 a_1066_9912# a_2240_10378# 0.0017f
C373 a_1066_5376# b[3] 1.15042f
C374 a_1066_12936# a_1066_12178# 0.02326f
C375 r[3] a_490_19738# 0.01905f
C376 VPWR b[4] 1.36578f
C377 a_1066_12178# a_490_11424# 0.0063f
C378 VPWR dg[6] 0.39096f
C379 VPWR a_320_19106# 0.07551f
C380 r[7] a_320_17594# 0.00425f
C381 VPWR a_1066_15202# 1.01184f
C382 a_490_6130# a_320_6294# 0.01277f
C383 a_2240_4782# db[4] 0.02175f
C384 a_586_22008# r[2] 0.00419f
C385 a_320_22716# r[0] 0.00243f
C386 a_1066_20496# r[2] 0.00943f
C387 a_2240_12132# dg[5] 0.00249f
C388 VPWR a_328_22474# 0.00734f
C389 VPWR r[4] 1.32853f
C390 a_490_6130# b[3] 0.00439f
C391 dg[1] a_1066_15202# 0.00646f
C392 dr[7] a_490_17472# 0.64642f
C393 a_778_6888# a_490_6130# 0.01178f
C394 dg[4] dg[6] 0.00112f
C395 g[4] g[5] 0.06698f
C396 VPWR a_320_14570# 0.07533f
C397 db[3] db[4] 0.13267f
C398 VPWR a_1066_12178# 1.00772f
C399 a_490_14448# g[2] 0.00126f
C400 r[3] dr[3] 0.01032f
C401 a_2240_21204# dr[2] 0.00191f
C402 a_1066_15202# a_2240_15156# 0.0017f
C403 a_1066_21250# dr[0] 0.04045f
C404 r[6] dr[7] 0.00363f
C405 a_1066_5376# b[4] 0.00126f
C406 a_1066_20496# a_2240_20618# 0.0073f
C407 r[4] a_490_19738# 1.15206f
C408 db[6] a_1066_4618# 0.04761f
C409 VPWR a_320_14914# 0.0021f
C410 VPWR dg[7] 0.37476f
C411 r[6] a_320_17938# 0.00117f
C412 a_490_2352# a_320_2474# 0.01277f
C413 db[6] a_1066_3106# 0.65369f
C414 a_490_22762# a_320_22926# 0.01277f
C415 a_490_7642# a_490_6130# 0.00185f
C416 a_2240_4782# db[5] 0.00165f
C417 db[0] b[0] 0.01316f
C418 a_1066_12178# dg[4] 0.68543f
C419 a_2240_13402# dg[2] 0.00217f
C420 a_490_7642# a_778_6888# 0.01399f
C421 VPWR r[5] 1.83028f
C422 g[0] a_490_14448# 0.02529f
C423 dr[6] a_2240_18180# 0.001f
C424 b[3] b[4] 0.06684f
C425 db[3] db[5] 0.0087f
C426 g[4] g[6] 0.00164f
C427 dg[5] dg[6] 0.72227f
C428 a_490_7642# a_320_7806# 0.01277f
C429 dr[0] r[0] 0.00466f
C430 r[4] dr[3] 0.00432f
C431 a_1066_21250# dr[1] 0.01975f
C432 dr[7] r[7] 0.00358f
C433 a_1066_12936# a_2240_13402# 0.0017f
C434 dr[4] a_1066_20496# 0.01041f
C435 r[5] a_490_19738# 0.00135f
C436 db[7] a_1066_4618# 0.02952f
C437 a_1066_12178# a_2240_12132# 0.0017f
C438 dg[0] g[1] 0.00204f
C439 VPWR a_320_19450# 0.0021f
C440 a_1066_4618# a_2240_4572# 0.0017f
C441 a_490_11424# a_320_11546# 0.01277f
C442 VPWR a_490_17472# 1.1249f
C443 db[7] a_1066_3106# 0.04045f
C444 db[6] b[6] 0.00215f
C445 b[5] db[7] 0.00575f
C446 a_490_22762# r[0] 1.15206f
C447 dg[2] g[2] 0.0087f
C448 a_1066_12178# dg[5] 0.03739f
C449 VPWR a_320_22926# 0.0758f
C450 VPWR a_1066_4618# 1.00725f
C451 VPWR r[6] 1.3707f
C452 VPWR a_1066_21250# 1.00882f
C453 r[3] r[4] 0.03875f
C454 dr[7] a_2240_18180# 0.00131f
C455 dr[5] a_1066_18226# 0.01707f
C456 db[7] a_490_3864# 0.01366f
C457 VPWR a_1066_3106# 1.01769f
C458 VPWR b[5] 1.83283f
C459 db[4] db[5] 0.65184f
C460 dg[5] dg[7] 0.00283f
C461 g[5] g[6] 0.02795f
C462 VPWR g[1] 1.82867f
C463 VPWR db[0] 0.28315f
C464 a_490_18984# a_1066_18226# 0.00532f
C465 VPWR a_320_3986# 0.07625f
C466 dr[0] r[1] 0.00672f
C467 VPWR a_320_11546# 0.07533f
C468 a_1066_21250# dr[2] 0.64284f
C469 a_2152_22474# dr[0] 0.00244f
C470 a_490_10666# g[4] 0.00294f
C471 VPWR a_490_3864# 1.12917f
C472 dg[1] g[1] 0.00776f
C473 r[4] a_320_19106# 0.00134f
C474 b[7] VGND 0.95169f
C475 db[7] VGND 1.61374f
C476 b[6] VGND 1.30075f
C477 db[6] VGND 1.02917f
C478 b[5] VGND 0.924f
C479 db[5] VGND 1.21713f
C480 b[4] VGND 1.26821f
C481 db[4] VGND 1.01911f
C482 b[3] VGND 0.79436f
C483 db[3] VGND 1.07501f
C484 b[2] VGND 1.06941f
C485 db[2] VGND 1.07414f
C486 b[1] VGND 0.95311f
C487 db[1] VGND 0.90922f
C488 b[0] VGND 1.09565f
C489 db[0] VGND 1.6139f
C490 g[7] VGND 0.87541f
C491 dg[7] VGND 1.26226f
C492 g[6] VGND 1.06833f
C493 dg[6] VGND 1.27247f
C494 g[5] VGND 0.91524f
C495 dg[5] VGND 1.1662f
C496 g[4] VGND 1.28865f
C497 dg[4] VGND 0.82346f
C498 g[3] VGND 0.80492f
C499 dg[3] VGND 0.80967f
C500 g[2] VGND 1.06311f
C501 dg[2] VGND 1.23607f
C502 g[1] VGND 0.91685f
C503 dg[1] VGND 1.20506f
C504 g[0] VGND 1.35238f
C505 dg[0] VGND 1.2299f
C506 r[7] VGND 0.95169f
C507 dr[7] VGND 1.28669f
C508 r[6] VGND 1.32279f
C509 dr[6] VGND 0.80329f
C510 r[5] VGND 0.91887f
C511 dr[5] VGND 1.05116f
C512 r[4] VGND 1.05902f
C513 dr[4] VGND 1.29389f
C514 r[3] VGND 1.02807f
C515 dr[3] VGND 1.05765f
C516 r[2] VGND 1.31214f
C517 dr[2] VGND 1.05883f
C518 r[1] VGND 0.934f
C519 dr[1] VGND 1.19729f
C520 r[0] VGND 1.0886f
C521 dr[0] VGND 1.61666f
C522 VPWR VGND 89.44511f
C523 a_320_2474# VGND 0.08041f $ **FLOATING
C524 a_490_2352# VGND 2.34771f
C525 a_320_2818# VGND 0.00719f $ **FLOATING
C526 a_2240_3060# VGND 0.00521f $ **FLOATING
C527 a_2240_3270# VGND 0.08013f $ **FLOATING
C528 a_1066_3106# VGND 2.36735f
C529 a_320_3986# VGND 0.08039f $ **FLOATING
C530 a_490_3864# VGND 2.33953f
C531 a_320_4330# VGND 0.00719f $ **FLOATING
C532 a_2240_4572# VGND 0.00513f $ **FLOATING
C533 a_2240_4782# VGND 0.07916f $ **FLOATING
C534 a_1066_4618# VGND 2.35547f
C535 a_2240_5498# VGND 0.07954f $ **FLOATING
C536 a_2240_5842# VGND 0.00521f $ **FLOATING
C537 a_1066_5376# VGND 2.35695f
C538 a_320_6084# VGND 0.00719f $ **FLOATING
C539 a_320_6294# VGND 0.08039f $ **FLOATING
C540 a_490_6130# VGND 2.32929f
C541 a_778_6888# VGND 2.35993f
C542 a_320_7596# VGND 0.00719f $ **FLOATING
C543 a_320_7806# VGND 0.08042f $ **FLOATING
C544 a_490_7642# VGND 2.34585f
C545 a_2240_10034# VGND 0.08052f $ **FLOATING
C546 a_2240_10378# VGND 0.00521f $ **FLOATING
C547 a_1066_9912# VGND 2.38495f
C548 a_320_10620# VGND 0.00719f $ **FLOATING
C549 a_320_10830# VGND 0.07989f $ **FLOATING
C550 a_490_10666# VGND 2.32325f
C551 a_320_11546# VGND 0.07989f $ **FLOATING
C552 a_490_11424# VGND 2.32128f
C553 a_320_11890# VGND 0.00719f $ **FLOATING
C554 a_2240_12132# VGND 0.00513f $ **FLOATING
C555 a_2240_12342# VGND 0.07962f $ **FLOATING
C556 a_1066_12178# VGND 2.35882f
C557 a_2240_13058# VGND 0.07954f $ **FLOATING
C558 a_2240_13402# VGND 0.00513f $ **FLOATING
C559 a_1066_12936# VGND 2.35921f
C560 a_320_13644# VGND 0.00719f $ **FLOATING
C561 a_320_13854# VGND 0.07989f $ **FLOATING
C562 a_490_13690# VGND 2.32388f
C563 a_320_14570# VGND 0.07989f $ **FLOATING
C564 a_490_14448# VGND 2.32557f
C565 a_320_14914# VGND 0.00719f $ **FLOATING
C566 a_2240_15156# VGND 0.00521f $ **FLOATING
C567 a_2240_15366# VGND 0.08052f $ **FLOATING
C568 a_1066_15202# VGND 2.3849f
C569 a_320_17594# VGND 0.08041f $ **FLOATING
C570 a_490_17472# VGND 2.34771f
C571 a_320_17938# VGND 0.00719f $ **FLOATING
C572 a_2240_18180# VGND 0.00521f $ **FLOATING
C573 a_2240_18390# VGND 0.08043f $ **FLOATING
C574 a_1066_18226# VGND 2.37104f
C575 a_320_19106# VGND 0.07955f $ **FLOATING
C576 a_490_18984# VGND 2.33124f
C577 a_320_19450# VGND 0.00719f $ **FLOATING
C578 a_320_19692# VGND 0.00719f $ **FLOATING
C579 a_320_19902# VGND 0.07995f $ **FLOATING
C580 a_490_19738# VGND 2.33364f
C581 a_2240_20618# VGND 0.07958f $ **FLOATING
C582 a_2240_20962# VGND 0.00513f $ **FLOATING
C583 a_1066_20496# VGND 2.35889f
C584 a_2240_21204# VGND 0.00521f $ **FLOATING
C585 a_2240_21414# VGND 0.07889f $ **FLOATING
C586 a_1066_21250# VGND 2.35321f
C587 a_2152_22130# VGND 0.12627f $ **FLOATING
C588 a_2152_22474# VGND 0.02388f $ **FLOATING
C589 a_328_22130# VGND 0.12215f $ **FLOATING
C590 a_586_22008# VGND 2.34335f
C591 a_328_22474# VGND 0.0226f $ **FLOATING
C592 a_320_22716# VGND 0.00719f $ **FLOATING
C593 a_320_22926# VGND 0.08008f $ **FLOATING
C594 a_490_22762# VGND 2.34603f
C595 g[7].t1 VGND 0.07912f
C596 g[7].n0 VGND 0.34756f
C597 g[7].n1 VGND 0.08515f
C598 g[7].t3 VGND 0.07903f
C599 g[7].n2 VGND 0.02411f
C600 g[7].n3 VGND 0.2194f
C601 g[7].n4 VGND 0.0607f
C602 g[7].t0 VGND 0.07903f
C603 g[7].n5 VGND 0.02393f
C604 g[7].n6 VGND 0.124f
C605 g[7].t2 VGND 0.07935f
C606 g[7].n7 VGND 0.06844f
C607 g[7].t7 VGND 0.12115f
C608 g[7].t5 VGND 0.12879f
C609 g[7].t6 VGND 0.12117f
C610 g[7].n8 VGND 0.19433f
C611 g[7].t4 VGND 0.11963f
C612 g[7].n9 VGND 0.09718f
C613 g[7].n10 VGND 0.0634f
C614 g[7].n11 VGND 0.11747f
C615 g[3].t1 VGND 0.07912f
C616 g[3].n0 VGND 0.34756f
C617 g[3].n1 VGND 0.08515f
C618 g[3].t3 VGND 0.07903f
C619 g[3].n2 VGND 0.02411f
C620 g[3].n3 VGND 0.2194f
C621 g[3].n4 VGND 0.0607f
C622 g[3].t0 VGND 0.07903f
C623 g[3].n5 VGND 0.02393f
C624 g[3].n6 VGND 0.124f
C625 g[3].t2 VGND 0.07935f
C626 g[3].n7 VGND 0.06844f
C627 g[3].t5 VGND 0.12115f
C628 g[3].t7 VGND 0.12879f
C629 g[3].t6 VGND 0.12117f
C630 g[3].n8 VGND 0.19433f
C631 g[3].t4 VGND 0.11963f
C632 g[3].n9 VGND 0.09718f
C633 g[3].n10 VGND 0.0634f
C634 g[3].n11 VGND 0.11747f
C635 b[3].t2 VGND 0.07912f
C636 b[3].n0 VGND 0.34756f
C637 b[3].n1 VGND 0.08515f
C638 b[3].t1 VGND 0.07903f
C639 b[3].n2 VGND 0.02411f
C640 b[3].n3 VGND 0.2194f
C641 b[3].n4 VGND 0.0607f
C642 b[3].t3 VGND 0.07903f
C643 b[3].n5 VGND 0.02393f
C644 b[3].n6 VGND 0.124f
C645 b[3].t0 VGND 0.07935f
C646 b[3].n7 VGND 0.06844f
C647 b[3].t4 VGND 0.12115f
C648 b[3].t6 VGND 0.12879f
C649 b[3].t7 VGND 0.12117f
C650 b[3].n8 VGND 0.19433f
C651 b[3].t5 VGND 0.11963f
C652 b[3].n9 VGND 0.09718f
C653 b[3].n10 VGND 0.0634f
C654 b[3].n11 VGND 0.11747f
C655 VPWR.t203 VGND 0.00138f
C656 VPWR.t178 VGND 0.00139f
C657 VPWR.n0 VGND 0.00306f
C658 VPWR.t489 VGND 0.00511f
C659 VPWR.n3 VGND 0.00626f
C660 VPWR.t183 VGND 0.00287f
C661 VPWR.n4 VGND 0.00384f
C662 VPWR.t156 VGND 0.00287f
C663 VPWR.t448 VGND 0.00511f
C664 VPWR.n5 VGND 0.00583f
C665 VPWR.n6 VGND 0.00545f
C666 VPWR.t184 VGND 0.00138f
C667 VPWR.t157 VGND 0.00139f
C668 VPWR.n8 VGND 0.00334f
C669 VPWR.t488 VGND 0.00511f
C670 VPWR.n12 VGND 0.00626f
C671 VPWR.t190 VGND 0.00287f
C672 VPWR.n13 VGND 0.00333f
C673 VPWR.t160 VGND 0.00287f
C674 VPWR.t449 VGND 0.00511f
C675 VPWR.n14 VGND 0.00583f
C676 VPWR.n15 VGND 0.00521f
C677 VPWR.t191 VGND 0.00138f
C678 VPWR.t161 VGND 0.00139f
C679 VPWR.n17 VGND 0.00341f
C680 VPWR.t497 VGND 0.00511f
C681 VPWR.n21 VGND 0.00626f
C682 VPWR.t202 VGND 0.00287f
C683 VPWR.n22 VGND 0.00339f
C684 VPWR.t177 VGND 0.00287f
C685 VPWR.t496 VGND 0.00511f
C686 VPWR.n23 VGND 0.00583f
C687 VPWR.n24 VGND 0.00481f
C688 VPWR.t167 VGND 0.00138f
C689 VPWR.t154 VGND 0.00139f
C690 VPWR.n26 VGND 0.00306f
C691 VPWR.t478 VGND 0.00511f
C692 VPWR.n29 VGND 0.00626f
C693 VPWR.t152 VGND 0.00287f
C694 VPWR.n30 VGND 0.00384f
C695 VPWR.t141 VGND 0.00287f
C696 VPWR.t456 VGND 0.00511f
C697 VPWR.n31 VGND 0.00583f
C698 VPWR.n32 VGND 0.00545f
C699 VPWR.t243 VGND 0.00138f
C700 VPWR.t225 VGND 0.00139f
C701 VPWR.n34 VGND 0.00334f
C702 VPWR.t460 VGND 0.00511f
C703 VPWR.n38 VGND 0.00626f
C704 VPWR.t158 VGND 0.00287f
C705 VPWR.n39 VGND 0.00333f
C706 VPWR.t150 VGND 0.00287f
C707 VPWR.t473 VGND 0.00511f
C708 VPWR.n40 VGND 0.00583f
C709 VPWR.n41 VGND 0.00521f
C710 VPWR.t159 VGND 0.00138f
C711 VPWR.t151 VGND 0.00139f
C712 VPWR.n43 VGND 0.00341f
C713 VPWR.n46 VGND 0.00339f
C714 VPWR.t466 VGND 0.00511f
C715 VPWR.t166 VGND 0.00287f
C716 VPWR.n47 VGND 0.00626f
C717 VPWR.t153 VGND 0.00287f
C718 VPWR.t444 VGND 0.00511f
C719 VPWR.n48 VGND 0.00583f
C720 VPWR.n49 VGND 0.00481f
C721 VPWR.t140 VGND 0.16772f
C722 VPWR.n51 VGND 0.01183f
C723 VPWR.n53 VGND 0.00577f
C724 VPWR.t83 VGND 0.00157f
C725 VPWR.t145 VGND 0.00138f
C726 VPWR.n55 VGND 0.00153f
C727 VPWR.t465 VGND 0.00511f
C728 VPWR.n58 VGND 0.00626f
C729 VPWR.t217 VGND 0.00287f
C730 VPWR.n59 VGND 0.00384f
C731 VPWR.t198 VGND 0.00287f
C732 VPWR.t468 VGND 0.00511f
C733 VPWR.n60 VGND 0.00583f
C734 VPWR.n61 VGND 0.00545f
C735 VPWR.t218 VGND 0.00138f
C736 VPWR.t199 VGND 0.00139f
C737 VPWR.n63 VGND 0.00334f
C738 VPWR.t399 VGND 0.00169f
C739 VPWR.n67 VGND 0.00139f
C740 VPWR.t82 VGND 0.00169f
C741 VPWR.n70 VGND 0.00246f
C742 VPWR.n71 VGND 0.0027f
C743 VPWR.n72 VGND 0.00173f
C744 VPWR.t194 VGND 0.00287f
C745 VPWR.n73 VGND 0.00151f
C746 VPWR.n74 VGND 0.00227f
C747 VPWR.t482 VGND 0.00507f
C748 VPWR.n75 VGND 0.00158f
C749 VPWR.n76 VGND 0.00723f
C750 VPWR.t301 VGND 0.00138f
C751 VPWR.t85 VGND 0.00169f
C752 VPWR.n78 VGND 0.00179f
C753 VPWR.n79 VGND 0.00156f
C754 VPWR.t81 VGND 0.00169f
C755 VPWR.n82 VGND 0.00186f
C756 VPWR.t457 VGND 0.00511f
C757 VPWR.n83 VGND 0.00154f
C758 VPWR.t144 VGND 0.00287f
C759 VPWR.n84 VGND 0.00626f
C760 VPWR.t80 VGND 0.00169f
C761 VPWR.n85 VGND 0.00439f
C762 VPWR.t79 VGND 0.16772f
C763 VPWR.n87 VGND 0.01183f
C764 VPWR.n89 VGND 0.00164f
C765 VPWR.n90 VGND 0.00288f
C766 VPWR.n91 VGND 0.13433f
C767 VPWR.t263 VGND 0.00139f
C768 VPWR.n93 VGND 0.00174f
C769 VPWR.n96 VGND 0.00372f
C770 VPWR.n99 VGND 0.00197f
C771 VPWR.t286 VGND 0.00133f
C772 VPWR.t15 VGND 0.00169f
C773 VPWR.t464 VGND 0.00252f
C774 VPWR.n100 VGND 0.00255f
C775 VPWR.n101 VGND 0.00217f
C776 VPWR.t287 VGND 0.00135f
C777 VPWR.t14 VGND 0.00169f
C778 VPWR.n104 VGND 0.00137f
C779 VPWR.n105 VGND 0.00135f
C780 VPWR.t102 VGND 0.00169f
C781 VPWR.n108 VGND 0.00154f
C782 VPWR.t412 VGND 0.00169f
C783 VPWR.n110 VGND 0.00139f
C784 VPWR.t99 VGND 0.00169f
C785 VPWR.n112 VGND 0.00154f
C786 VPWR.t386 VGND 0.00169f
C787 VPWR.n114 VGND 0.00139f
C788 VPWR.t103 VGND 0.00169f
C789 VPWR.n116 VGND 0.00155f
C790 VPWR.t380 VGND 0.00169f
C791 VPWR.n118 VGND 0.00154f
C792 VPWR.t98 VGND 0.00157f
C793 VPWR.n120 VGND 0.00182f
C794 VPWR.t379 VGND 0.00169f
C795 VPWR.n122 VGND 0.00133f
C796 VPWR.t381 VGND 0.00169f
C797 VPWR.n125 VGND 0.00155f
C798 VPWR.n127 VGND 0.00173f
C799 VPWR.t196 VGND 0.00287f
C800 VPWR.t474 VGND 0.00511f
C801 VPWR.n128 VGND 0.00583f
C802 VPWR.n129 VGND 0.00144f
C803 VPWR.n130 VGND 0.00217f
C804 VPWR.t384 VGND 0.00157f
C805 VPWR.n131 VGND 0.00182f
C806 VPWR.t13 VGND 0.16772f
C807 VPWR.n133 VGND 0.01183f
C808 VPWR.n135 VGND 0.00276f
C809 VPWR.n136 VGND 0.06762f
C810 VPWR.t393 VGND 0.00157f
C811 VPWR.t249 VGND 0.00138f
C812 VPWR.n138 VGND 0.00153f
C813 VPWR.n140 VGND 0.00198f
C814 VPWR.t447 VGND 0.00511f
C815 VPWR.t169 VGND 0.00287f
C816 VPWR.n142 VGND 0.00583f
C817 VPWR.t133 VGND 0.00169f
C818 VPWR.n143 VGND 0.00175f
C819 VPWR.n144 VGND 0.0021f
C820 VPWR.n146 VGND 0.00146f
C821 VPWR.t2 VGND 0.00169f
C822 VPWR.n148 VGND 0.00139f
C823 VPWR.t266 VGND 0.00139f
C824 VPWR.n150 VGND 0.00174f
C825 VPWR.t3 VGND 0.00169f
C826 VPWR.n152 VGND 0.00133f
C827 VPWR.t1 VGND 0.00169f
C828 VPWR.t431 VGND 0.00169f
C829 VPWR.n154 VGND 0.00157f
C830 VPWR.n155 VGND 0.00178f
C831 VPWR.t4 VGND 0.00169f
C832 VPWR.t392 VGND 0.00169f
C833 VPWR.n157 VGND 0.00159f
C834 VPWR.n158 VGND 0.00176f
C835 VPWR.t7 VGND 0.00157f
C836 VPWR.t395 VGND 0.00169f
C837 VPWR.n160 VGND 0.00177f
C838 VPWR.n161 VGND 0.00164f
C839 VPWR.t391 VGND 0.00169f
C840 VPWR.n164 VGND 0.00186f
C841 VPWR.t451 VGND 0.00511f
C842 VPWR.n165 VGND 0.00154f
C843 VPWR.t188 VGND 0.00287f
C844 VPWR.n166 VGND 0.00626f
C845 VPWR.t390 VGND 0.00169f
C846 VPWR.n167 VGND 0.00439f
C847 VPWR.t0 VGND 0.16772f
C848 VPWR.n169 VGND 0.01183f
C849 VPWR.n171 VGND 0.00164f
C850 VPWR.n172 VGND 0.00288f
C851 VPWR.n173 VGND 0.06762f
C852 VPWR.t118 VGND 0.00157f
C853 VPWR.t247 VGND 0.00139f
C854 VPWR.n175 VGND 0.00153f
C855 VPWR.n177 VGND 0.00198f
C856 VPWR.t173 VGND 0.00287f
C857 VPWR.t470 VGND 0.00511f
C858 VPWR.n179 VGND 0.00583f
C859 VPWR.t130 VGND 0.00169f
C860 VPWR.n180 VGND 0.00175f
C861 VPWR.n181 VGND 0.0021f
C862 VPWR.n183 VGND 0.00146f
C863 VPWR.t24 VGND 0.00169f
C864 VPWR.n185 VGND 0.00139f
C865 VPWR.t270 VGND 0.00138f
C866 VPWR.n187 VGND 0.00174f
C867 VPWR.t20 VGND 0.00169f
C868 VPWR.n189 VGND 0.00133f
C869 VPWR.t22 VGND 0.00169f
C870 VPWR.t88 VGND 0.00169f
C871 VPWR.n191 VGND 0.00157f
C872 VPWR.n192 VGND 0.00178f
C873 VPWR.t18 VGND 0.00169f
C874 VPWR.t90 VGND 0.00169f
C875 VPWR.n194 VGND 0.00159f
C876 VPWR.n195 VGND 0.00176f
C877 VPWR.t21 VGND 0.00157f
C878 VPWR.t120 VGND 0.00169f
C879 VPWR.n197 VGND 0.00177f
C880 VPWR.n198 VGND 0.00164f
C881 VPWR.t116 VGND 0.00169f
C882 VPWR.n201 VGND 0.00186f
C883 VPWR.t115 VGND 0.0017f
C884 VPWR.n202 VGND 0.00154f
C885 VPWR.t185 VGND 0.00287f
C886 VPWR.t458 VGND 0.00511f
C887 VPWR.n203 VGND 0.00583f
C888 VPWR.n204 VGND 0.0042f
C889 VPWR.t17 VGND 0.16772f
C890 VPWR.n206 VGND 0.01183f
C891 VPWR.n208 VGND 0.00164f
C892 VPWR.n209 VGND 0.00288f
C893 VPWR.n210 VGND 0.06762f
C894 VPWR.t322 VGND 0.00157f
C895 VPWR.t272 VGND 0.00139f
C896 VPWR.n212 VGND 0.00153f
C897 VPWR.t484 VGND 0.00511f
C898 VPWR.n215 VGND 0.00626f
C899 VPWR.t149 VGND 0.00287f
C900 VPWR.n216 VGND 0.00384f
C901 VPWR.t175 VGND 0.00287f
C902 VPWR.t479 VGND 0.00511f
C903 VPWR.n217 VGND 0.00583f
C904 VPWR.n218 VGND 0.00545f
C905 VPWR.t228 VGND 0.00138f
C906 VPWR.t176 VGND 0.00139f
C907 VPWR.n220 VGND 0.00334f
C908 VPWR.t441 VGND 0.00169f
C909 VPWR.n224 VGND 0.00139f
C910 VPWR.t321 VGND 0.00169f
C911 VPWR.n227 VGND 0.00246f
C912 VPWR.n228 VGND 0.0027f
C913 VPWR.n229 VGND 0.00173f
C914 VPWR.t148 VGND 0.00287f
C915 VPWR.n230 VGND 0.00151f
C916 VPWR.n231 VGND 0.00227f
C917 VPWR.t445 VGND 0.00507f
C918 VPWR.n232 VGND 0.00158f
C919 VPWR.n233 VGND 0.00723f
C920 VPWR.t257 VGND 0.00139f
C921 VPWR.t318 VGND 0.00169f
C922 VPWR.n235 VGND 0.00179f
C923 VPWR.n236 VGND 0.00156f
C924 VPWR.t320 VGND 0.00169f
C925 VPWR.n239 VGND 0.00186f
C926 VPWR.t319 VGND 0.0017f
C927 VPWR.n240 VGND 0.00154f
C928 VPWR.t201 VGND 0.00287f
C929 VPWR.t471 VGND 0.00511f
C930 VPWR.n241 VGND 0.00583f
C931 VPWR.n242 VGND 0.0042f
C932 VPWR.t147 VGND 0.16772f
C933 VPWR.n244 VGND 0.01183f
C934 VPWR.n246 VGND 0.00164f
C935 VPWR.n247 VGND 0.00288f
C936 VPWR.n248 VGND 0.06762f
C937 VPWR.t268 VGND 0.00138f
C938 VPWR.t234 VGND 0.00139f
C939 VPWR.n250 VGND 0.00306f
C940 VPWR.n252 VGND 0.00198f
C941 VPWR.t171 VGND 0.00287f
C942 VPWR.t476 VGND 0.00511f
C943 VPWR.n254 VGND 0.00583f
C944 VPWR.t435 VGND 0.00169f
C945 VPWR.n255 VGND 0.00175f
C946 VPWR.n256 VGND 0.0021f
C947 VPWR.n258 VGND 0.00146f
C948 VPWR.t74 VGND 0.00169f
C949 VPWR.n260 VGND 0.00139f
C950 VPWR.t172 VGND 0.00138f
C951 VPWR.n262 VGND 0.00174f
C952 VPWR.t75 VGND 0.00169f
C953 VPWR.n264 VGND 0.00133f
C954 VPWR.t72 VGND 0.00169f
C955 VPWR.n267 VGND 0.00154f
C956 VPWR.n269 VGND 0.00173f
C957 VPWR.t143 VGND 0.00287f
C958 VPWR.t454 VGND 0.00511f
C959 VPWR.n270 VGND 0.00626f
C960 VPWR.t76 VGND 0.00169f
C961 VPWR.n271 VGND 0.0048f
C962 VPWR.t254 VGND 0.00138f
C963 VPWR.t71 VGND 0.00157f
C964 VPWR.n273 VGND 0.00204f
C965 VPWR.n274 VGND 0.00141f
C966 VPWR.n277 VGND 0.00339f
C967 VPWR.t462 VGND 0.00511f
C968 VPWR.t197 VGND 0.00287f
C969 VPWR.n278 VGND 0.00626f
C970 VPWR.t168 VGND 0.00287f
C971 VPWR.t487 VGND 0.00511f
C972 VPWR.n279 VGND 0.00583f
C973 VPWR.n280 VGND 0.00481f
C974 VPWR.t70 VGND 0.16772f
C975 VPWR.n282 VGND 0.01183f
C976 VPWR.n284 VGND 0.00297f
C977 VPWR.n285 VGND 0.06762f
C978 VPWR.t59 VGND 0.00157f
C979 VPWR.t416 VGND 0.00157f
C980 VPWR.t95 VGND 0.00169f
C981 VPWR.t437 VGND 0.00169f
C982 VPWR.n288 VGND 0.00302f
C983 VPWR.t58 VGND 0.00169f
C984 VPWR.t415 VGND 0.00169f
C985 VPWR.n290 VGND 0.003f
C986 VPWR.t53 VGND 0.00169f
C987 VPWR.t418 VGND 0.00169f
C988 VPWR.n292 VGND 0.00328f
C989 VPWR.t54 VGND 0.00169f
C990 VPWR.t419 VGND 0.00169f
C991 VPWR.n294 VGND 0.0033f
C992 VPWR.t57 VGND 0.00169f
C993 VPWR.t417 VGND 0.00169f
C994 VPWR.n295 VGND 0.00328f
C995 VPWR.t137 VGND 0.00138f
C996 VPWR.t282 VGND 0.00139f
C997 VPWR.n300 VGND 0.00334f
C998 VPWR.t450 VGND 0.00511f
C999 VPWR.n301 VGND 0.00626f
C1000 VPWR.t136 VGND 0.00287f
C1001 VPWR.n302 VGND 0.00384f
C1002 VPWR.t193 VGND 0.00287f
C1003 VPWR.t486 VGND 0.00511f
C1004 VPWR.n303 VGND 0.00583f
C1005 VPWR.n304 VGND 0.00545f
C1006 VPWR.t52 VGND 0.16772f
C1007 VPWR.n306 VGND 0.01183f
C1008 VPWR.n308 VGND 0.00305f
C1009 VPWR.n309 VGND 0.0032f
C1010 VPWR.n310 VGND 0.06762f
C1011 VPWR.t206 VGND 0.00138f
C1012 VPWR.t182 VGND 0.00139f
C1013 VPWR.n312 VGND 0.00306f
C1014 VPWR.t370 VGND 0.00169f
C1015 VPWR.t388 VGND 0.00169f
C1016 VPWR.n315 VGND 0.00317f
C1017 VPWR.t332 VGND 0.00169f
C1018 VPWR.t387 VGND 0.00169f
C1019 VPWR.n317 VGND 0.003f
C1020 VPWR.t328 VGND 0.00169f
C1021 VPWR.t408 VGND 0.00169f
C1022 VPWR.n319 VGND 0.00328f
C1023 VPWR.t330 VGND 0.00169f
C1024 VPWR.t405 VGND 0.00169f
C1025 VPWR.n321 VGND 0.00328f
C1026 VPWR.t326 VGND 0.00169f
C1027 VPWR.t409 VGND 0.00169f
C1028 VPWR.n323 VGND 0.0033f
C1029 VPWR.t329 VGND 0.00157f
C1030 VPWR.t404 VGND 0.00157f
C1031 VPWR.n325 VGND 0.00351f
C1032 VPWR.n328 VGND 0.00339f
C1033 VPWR.t480 VGND 0.00511f
C1034 VPWR.t205 VGND 0.00287f
C1035 VPWR.n329 VGND 0.00626f
C1036 VPWR.t181 VGND 0.00287f
C1037 VPWR.t490 VGND 0.00511f
C1038 VPWR.n330 VGND 0.00583f
C1039 VPWR.n331 VGND 0.00481f
C1040 VPWR.t180 VGND 0.16772f
C1041 VPWR.n333 VGND 0.01183f
C1042 VPWR.n335 VGND 0.00297f
C1043 VPWR.n336 VGND 0.06762f
C1044 VPWR.t344 VGND 0.00157f
C1045 VPWR.t50 VGND 0.00157f
C1046 VPWR.t338 VGND 0.00169f
C1047 VPWR.t10 VGND 0.00169f
C1048 VPWR.n339 VGND 0.00302f
C1049 VPWR.t337 VGND 0.00169f
C1050 VPWR.t12 VGND 0.00169f
C1051 VPWR.n341 VGND 0.003f
C1052 VPWR.t340 VGND 0.00169f
C1053 VPWR.t44 VGND 0.00169f
C1054 VPWR.n343 VGND 0.00328f
C1055 VPWR.t341 VGND 0.00169f
C1056 VPWR.t45 VGND 0.00169f
C1057 VPWR.n345 VGND 0.0033f
C1058 VPWR.t342 VGND 0.00169f
C1059 VPWR.t48 VGND 0.00169f
C1060 VPWR.n346 VGND 0.00328f
C1061 VPWR.t289 VGND 0.00138f
C1062 VPWR.t220 VGND 0.00139f
C1063 VPWR.n351 VGND 0.00334f
C1064 VPWR.t455 VGND 0.00511f
C1065 VPWR.n352 VGND 0.00626f
C1066 VPWR.t204 VGND 0.00287f
C1067 VPWR.n353 VGND 0.00384f
C1068 VPWR.t219 VGND 0.00287f
C1069 VPWR.t469 VGND 0.00511f
C1070 VPWR.n354 VGND 0.00583f
C1071 VPWR.n355 VGND 0.00545f
C1072 VPWR.t9 VGND 0.16772f
C1073 VPWR.n357 VGND 0.01183f
C1074 VPWR.n359 VGND 0.00305f
C1075 VPWR.n360 VGND 0.0032f
C1076 VPWR.n361 VGND 0.06762f
C1077 VPWR.t261 VGND 0.00138f
C1078 VPWR.t230 VGND 0.00139f
C1079 VPWR.n363 VGND 0.00306f
C1080 VPWR.n365 VGND 0.00198f
C1081 VPWR.t446 VGND 0.00511f
C1082 VPWR.t138 VGND 0.00287f
C1083 VPWR.n367 VGND 0.00583f
C1084 VPWR.t401 VGND 0.00169f
C1085 VPWR.n368 VGND 0.00175f
C1086 VPWR.n369 VGND 0.0021f
C1087 VPWR.n371 VGND 0.00146f
C1088 VPWR.t112 VGND 0.00169f
C1089 VPWR.n373 VGND 0.00139f
C1090 VPWR.t139 VGND 0.00139f
C1091 VPWR.n375 VGND 0.00174f
C1092 VPWR.t108 VGND 0.00169f
C1093 VPWR.n377 VGND 0.00133f
C1094 VPWR.t111 VGND 0.00169f
C1095 VPWR.n380 VGND 0.00154f
C1096 VPWR.t107 VGND 0.0017f
C1097 VPWR.n382 VGND 0.00173f
C1098 VPWR.t146 VGND 0.00287f
C1099 VPWR.t452 VGND 0.00511f
C1100 VPWR.n383 VGND 0.00583f
C1101 VPWR.n384 VGND 0.00461f
C1102 VPWR.t251 VGND 0.00139f
C1103 VPWR.t113 VGND 0.00157f
C1104 VPWR.n386 VGND 0.00204f
C1105 VPWR.n387 VGND 0.00141f
C1106 VPWR.n390 VGND 0.00339f
C1107 VPWR.t461 VGND 0.00511f
C1108 VPWR.t260 VGND 0.00287f
C1109 VPWR.n391 VGND 0.00626f
C1110 VPWR.t229 VGND 0.00287f
C1111 VPWR.t475 VGND 0.00511f
C1112 VPWR.n392 VGND 0.00583f
C1113 VPWR.n393 VGND 0.00481f
C1114 VPWR.t106 VGND 0.16772f
C1115 VPWR.n395 VGND 0.01183f
C1116 VPWR.n397 VGND 0.00297f
C1117 VPWR.n398 VGND 0.06762f
C1118 VPWR.t31 VGND 0.00157f
C1119 VPWR.t223 VGND 0.00138f
C1120 VPWR.n400 VGND 0.00153f
C1121 VPWR.t492 VGND 0.00511f
C1122 VPWR.n403 VGND 0.00626f
C1123 VPWR.t290 VGND 0.00287f
C1124 VPWR.n404 VGND 0.00384f
C1125 VPWR.t231 VGND 0.00287f
C1126 VPWR.t481 VGND 0.00511f
C1127 VPWR.n405 VGND 0.00583f
C1128 VPWR.n406 VGND 0.00545f
C1129 VPWR.t291 VGND 0.00138f
C1130 VPWR.t232 VGND 0.00139f
C1131 VPWR.n408 VGND 0.00334f
C1132 VPWR.t127 VGND 0.00169f
C1133 VPWR.n412 VGND 0.00139f
C1134 VPWR.t34 VGND 0.00169f
C1135 VPWR.n415 VGND 0.00246f
C1136 VPWR.n416 VGND 0.0027f
C1137 VPWR.n417 VGND 0.00173f
C1138 VPWR.t235 VGND 0.00287f
C1139 VPWR.n418 VGND 0.00151f
C1140 VPWR.n419 VGND 0.00227f
C1141 VPWR.t491 VGND 0.00507f
C1142 VPWR.n420 VGND 0.00158f
C1143 VPWR.n421 VGND 0.00723f
C1144 VPWR.t236 VGND 0.00138f
C1145 VPWR.t28 VGND 0.00169f
C1146 VPWR.n423 VGND 0.00179f
C1147 VPWR.n424 VGND 0.00156f
C1148 VPWR.t32 VGND 0.00169f
C1149 VPWR.n427 VGND 0.00186f
C1150 VPWR.t443 VGND 0.00511f
C1151 VPWR.n428 VGND 0.00154f
C1152 VPWR.t222 VGND 0.00287f
C1153 VPWR.n429 VGND 0.00626f
C1154 VPWR.t27 VGND 0.00169f
C1155 VPWR.n430 VGND 0.00439f
C1156 VPWR.t26 VGND 0.16772f
C1157 VPWR.n432 VGND 0.01183f
C1158 VPWR.n434 VGND 0.00164f
C1159 VPWR.n435 VGND 0.00288f
C1160 VPWR.n436 VGND 0.06762f
C1161 VPWR.t38 VGND 0.00157f
C1162 VPWR.t259 VGND 0.00135f
C1163 VPWR.n438 VGND 0.00127f
C1164 VPWR.n442 VGND 0.00372f
C1165 VPWR.n444 VGND 0.00244f
C1166 VPWR.t296 VGND 0.00133f
C1167 VPWR.t463 VGND 0.00252f
C1168 VPWR.n446 VGND 0.00265f
C1169 VPWR.n447 VGND 0.0025f
C1170 VPWR.t208 VGND 0.00287f
C1171 VPWR.n449 VGND 0.00723f
C1172 VPWR.n450 VGND 0.00146f
C1173 VPWR.t297 VGND 0.00135f
C1174 VPWR.n451 VGND 0.00249f
C1175 VPWR.n452 VGND 0.00222f
C1176 VPWR.t472 VGND 0.00507f
C1177 VPWR.n453 VGND 0.00109f
C1178 VPWR.n454 VGND 0.00126f
C1179 VPWR.t209 VGND 0.00139f
C1180 VPWR.t352 VGND 0.00169f
C1181 VPWR.n455 VGND 0.00169f
C1182 VPWR.n456 VGND 0.00167f
C1183 VPWR.t312 VGND 0.00169f
C1184 VPWR.n459 VGND 0.00139f
C1185 VPWR.t376 VGND 0.00169f
C1186 VPWR.n461 VGND 0.00139f
C1187 VPWR.t310 VGND 0.00169f
C1188 VPWR.n463 VGND 0.00154f
C1189 VPWR.t41 VGND 0.00169f
C1190 VPWR.n465 VGND 0.00139f
C1191 VPWR.t311 VGND 0.00169f
C1192 VPWR.n467 VGND 0.00154f
C1193 VPWR.t37 VGND 0.00169f
C1194 VPWR.n469 VGND 0.00154f
C1195 VPWR.t316 VGND 0.00169f
C1196 VPWR.n471 VGND 0.00155f
C1197 VPWR.t39 VGND 0.00169f
C1198 VPWR.n473 VGND 0.00154f
C1199 VPWR.t313 VGND 0.00157f
C1200 VPWR.n475 VGND 0.00182f
C1201 VPWR.t36 VGND 0.00169f
C1202 VPWR.n477 VGND 0.00134f
C1203 VPWR.t485 VGND 0.00252f
C1204 VPWR.t258 VGND 0.00133f
C1205 VPWR.n479 VGND 0.00322f
C1206 VPWR.n480 VGND 0.00149f
C1207 VPWR.t35 VGND 0.16772f
C1208 VPWR.n482 VGND 0.01183f
C1209 VPWR.n484 VGND 0.00164f
C1210 VPWR.n485 VGND 0.00276f
C1211 VPWR.n486 VGND 0.06762f
C1212 VPWR.t163 VGND 0.00138f
C1213 VPWR.t279 VGND 0.00139f
C1214 VPWR.n488 VGND 0.00306f
C1215 VPWR.t348 VGND 0.00169f
C1216 VPWR.t374 VGND 0.00169f
C1217 VPWR.n491 VGND 0.00317f
C1218 VPWR.t349 VGND 0.00169f
C1219 VPWR.t65 VGND 0.00169f
C1220 VPWR.n493 VGND 0.003f
C1221 VPWR.t357 VGND 0.00169f
C1222 VPWR.t62 VGND 0.00169f
C1223 VPWR.n495 VGND 0.00328f
C1224 VPWR.t355 VGND 0.00169f
C1225 VPWR.t64 VGND 0.00169f
C1226 VPWR.n497 VGND 0.00328f
C1227 VPWR.t356 VGND 0.00169f
C1228 VPWR.t63 VGND 0.00169f
C1229 VPWR.n499 VGND 0.0033f
C1230 VPWR.t354 VGND 0.00157f
C1231 VPWR.t66 VGND 0.00157f
C1232 VPWR.n501 VGND 0.00351f
C1233 VPWR.n504 VGND 0.00339f
C1234 VPWR.t477 VGND 0.00511f
C1235 VPWR.t162 VGND 0.00287f
C1236 VPWR.n505 VGND 0.00626f
C1237 VPWR.t278 VGND 0.00287f
C1238 VPWR.t493 VGND 0.00511f
C1239 VPWR.n506 VGND 0.00583f
C1240 VPWR.n507 VGND 0.00481f
C1241 VPWR.t61 VGND 0.16772f
C1242 VPWR.n509 VGND 0.01183f
C1243 VPWR.n511 VGND 0.00297f
C1244 VPWR.n512 VGND 0.06762f
C1245 VPWR.t368 VGND 0.00157f
C1246 VPWR.t240 VGND 0.00139f
C1247 VPWR.n514 VGND 0.00153f
C1248 VPWR.n516 VGND 0.00198f
C1249 VPWR.t214 VGND 0.00287f
C1250 VPWR.t467 VGND 0.00511f
C1251 VPWR.n518 VGND 0.00583f
C1252 VPWR.t334 VGND 0.00169f
C1253 VPWR.n519 VGND 0.00175f
C1254 VPWR.n520 VGND 0.0021f
C1255 VPWR.n522 VGND 0.00146f
C1256 VPWR.t304 VGND 0.00169f
C1257 VPWR.n524 VGND 0.00139f
C1258 VPWR.t215 VGND 0.00138f
C1259 VPWR.n526 VGND 0.00174f
C1260 VPWR.t308 VGND 0.00169f
C1261 VPWR.n528 VGND 0.00133f
C1262 VPWR.t303 VGND 0.00169f
C1263 VPWR.t124 VGND 0.00169f
C1264 VPWR.n530 VGND 0.00157f
C1265 VPWR.n531 VGND 0.00178f
C1266 VPWR.t302 VGND 0.00169f
C1267 VPWR.t126 VGND 0.00169f
C1268 VPWR.n533 VGND 0.00159f
C1269 VPWR.n534 VGND 0.00176f
C1270 VPWR.t305 VGND 0.00157f
C1271 VPWR.t365 VGND 0.00169f
C1272 VPWR.n536 VGND 0.00177f
C1273 VPWR.n537 VGND 0.00164f
C1274 VPWR.t362 VGND 0.00169f
C1275 VPWR.n540 VGND 0.00186f
C1276 VPWR.t364 VGND 0.0017f
C1277 VPWR.n541 VGND 0.00154f
C1278 VPWR.t239 VGND 0.00287f
C1279 VPWR.t453 VGND 0.00511f
C1280 VPWR.n542 VGND 0.00583f
C1281 VPWR.n543 VGND 0.0042f
C1282 VPWR.t123 VGND 0.16772f
C1283 VPWR.n545 VGND 0.01183f
C1284 VPWR.n547 VGND 0.00164f
C1285 VPWR.n548 VGND 0.00288f
C1286 VPWR.n549 VGND 0.06762f
C1287 VPWR.t429 VGND 0.00157f
C1288 VPWR.t274 VGND 0.00139f
C1289 VPWR.n551 VGND 0.00153f
C1290 VPWR.t483 VGND 0.00511f
C1291 VPWR.n554 VGND 0.00626f
C1292 VPWR.t186 VGND 0.00287f
C1293 VPWR.n555 VGND 0.00384f
C1294 VPWR.t164 VGND 0.00287f
C1295 VPWR.t495 VGND 0.00511f
C1296 VPWR.n556 VGND 0.00583f
C1297 VPWR.n557 VGND 0.00545f
C1298 VPWR.t187 VGND 0.00138f
C1299 VPWR.t165 VGND 0.00139f
C1300 VPWR.n559 VGND 0.00334f
C1301 VPWR.t92 VGND 0.00169f
C1302 VPWR.n563 VGND 0.00139f
C1303 VPWR.t94 VGND 0.00169f
C1304 VPWR.n566 VGND 0.00246f
C1305 VPWR.n567 VGND 0.0027f
C1306 VPWR.n568 VGND 0.00173f
C1307 VPWR.t179 VGND 0.00287f
C1308 VPWR.n569 VGND 0.00151f
C1309 VPWR.n570 VGND 0.00227f
C1310 VPWR.t494 VGND 0.00507f
C1311 VPWR.n571 VGND 0.00158f
C1312 VPWR.n572 VGND 0.00723f
C1313 VPWR.t284 VGND 0.00139f
C1314 VPWR.t426 VGND 0.00169f
C1315 VPWR.n574 VGND 0.00179f
C1316 VPWR.n575 VGND 0.00156f
C1317 VPWR.t423 VGND 0.00169f
C1318 VPWR.n578 VGND 0.00186f
C1319 VPWR.t425 VGND 0.0017f
C1320 VPWR.n579 VGND 0.00154f
C1321 VPWR.t273 VGND 0.00287f
C1322 VPWR.t459 VGND 0.00511f
C1323 VPWR.n580 VGND 0.00583f
C1324 VPWR.n581 VGND 0.0042f
C1325 VPWR.t91 VGND 0.16772f
C1326 VPWR.n583 VGND 0.01183f
C1327 VPWR.n585 VGND 0.00164f
C1328 VPWR.n586 VGND 0.00288f
C1329 VPWR.n587 VGND 0.06762f
C1330 VPWR.n588 VGND 0.0523f
C1331 VPWR.n589 VGND 0.00297f
C1332 VPWR.t155 VGND 0.16772f
C1333 VPWR.n591 VGND 0.01183f
.ends

