magic
tech ihp-sg13g2
magscale 1 2
timestamp 1746816402
<< nwell >>
rect -48 350 816 834
<< pwell >>
rect 32 292 324 314
rect 32 56 745 292
rect -26 -56 794 56
<< nmos >>
rect 129 160 155 288
rect 204 160 230 288
rect 409 118 435 266
rect 523 118 549 266
rect 625 118 651 266
<< pmos >>
rect 166 429 192 597
rect 268 429 294 597
rect 409 412 435 636
rect 486 412 512 636
rect 598 412 624 636
<< ndiff >>
rect 58 274 129 288
rect 58 242 75 274
rect 107 242 129 274
rect 58 206 129 242
rect 58 174 75 206
rect 107 174 129 206
rect 58 160 129 174
rect 155 160 204 288
rect 230 274 298 288
rect 230 242 252 274
rect 284 242 298 274
rect 230 206 298 242
rect 230 174 252 206
rect 284 174 298 206
rect 230 160 298 174
rect 341 195 409 266
rect 341 163 355 195
rect 387 163 409 195
rect 341 118 409 163
rect 435 128 523 266
rect 435 118 463 128
rect 449 96 463 118
rect 495 118 523 128
rect 549 195 625 266
rect 549 163 571 195
rect 603 163 625 195
rect 549 118 625 163
rect 651 249 719 266
rect 651 217 673 249
rect 705 217 719 249
rect 651 165 719 217
rect 651 133 673 165
rect 705 133 719 165
rect 651 118 719 133
rect 495 96 509 118
rect 449 82 509 96
<< pdiff >>
rect 341 622 409 636
rect 341 597 355 622
rect 58 574 166 597
rect 58 542 74 574
rect 106 542 166 574
rect 58 482 166 542
rect 58 450 74 482
rect 106 450 166 482
rect 58 429 166 450
rect 192 574 268 597
rect 192 542 214 574
rect 246 542 268 574
rect 192 506 268 542
rect 192 474 214 506
rect 246 474 268 506
rect 192 429 268 474
rect 294 590 355 597
rect 387 590 409 622
rect 294 543 409 590
rect 294 511 355 543
rect 387 511 409 543
rect 294 429 409 511
rect 341 412 409 429
rect 435 412 486 636
rect 512 622 598 636
rect 512 590 544 622
rect 576 590 598 622
rect 512 543 598 590
rect 512 511 544 543
rect 576 511 598 543
rect 512 463 598 511
rect 512 431 544 463
rect 576 431 598 463
rect 512 412 598 431
rect 624 622 692 636
rect 624 590 646 622
rect 678 590 692 622
rect 624 520 692 590
rect 624 488 646 520
rect 678 488 692 520
rect 624 412 692 488
<< ndiffc >>
rect 75 242 107 274
rect 75 174 107 206
rect 252 242 284 274
rect 252 174 284 206
rect 355 163 387 195
rect 463 96 495 128
rect 571 163 603 195
rect 673 217 705 249
rect 673 133 705 165
<< pdiffc >>
rect 74 542 106 574
rect 74 450 106 482
rect 214 542 246 574
rect 214 474 246 506
rect 355 590 387 622
rect 355 511 387 543
rect 544 590 576 622
rect 544 511 576 543
rect 544 431 576 463
rect 646 590 678 622
rect 646 488 678 520
<< psubdiff >>
rect 0 16 768 30
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 608 16
rect 640 -16 704 16
rect 736 -16 768 16
rect 0 -30 768 -16
<< nsubdiff >>
rect 0 772 768 786
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 608 772
rect 640 740 704 772
rect 736 740 768 772
rect 0 726 768 740
<< psubdiffcont >>
rect 32 -16 64 16
rect 128 -16 160 16
rect 224 -16 256 16
rect 320 -16 352 16
rect 416 -16 448 16
rect 512 -16 544 16
rect 608 -16 640 16
rect 704 -16 736 16
<< nsubdiffcont >>
rect 32 740 64 772
rect 128 740 160 772
rect 224 740 256 772
rect 320 740 352 772
rect 416 740 448 772
rect 512 740 544 772
rect 608 740 640 772
rect 704 740 736 772
<< poly >>
rect 409 636 435 672
rect 486 636 512 672
rect 598 636 624 672
rect 166 597 192 633
rect 268 597 294 633
rect 166 414 192 429
rect 129 382 192 414
rect 268 397 294 429
rect 129 288 155 382
rect 248 380 314 397
rect 409 380 435 412
rect 486 380 512 412
rect 248 348 265 380
rect 297 348 314 380
rect 248 336 314 348
rect 204 306 314 336
rect 362 363 435 380
rect 362 331 379 363
rect 411 331 435 363
rect 362 314 435 331
rect 471 363 549 380
rect 598 370 624 412
rect 471 331 503 363
rect 535 331 549 363
rect 471 314 549 331
rect 204 288 230 306
rect 409 266 435 314
rect 523 266 549 314
rect 594 353 660 370
rect 594 321 611 353
rect 643 321 660 353
rect 594 304 660 321
rect 625 266 651 304
rect 129 88 155 160
rect 204 124 230 160
rect 409 88 435 118
rect 129 62 435 88
rect 523 82 549 118
rect 625 82 651 118
<< polycont >>
rect 265 348 297 380
rect 379 331 411 363
rect 503 331 535 363
rect 611 321 643 353
<< metal1 >>
rect 0 772 768 800
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 608 772
rect 640 740 704 772
rect 736 740 768 772
rect 0 712 768 740
rect 64 574 112 712
rect 345 622 399 712
rect 345 590 355 622
rect 387 590 399 622
rect 64 542 74 574
rect 106 542 112 574
rect 64 482 112 542
rect 194 574 248 586
rect 194 542 214 574
rect 246 542 248 574
rect 194 522 248 542
rect 64 450 74 482
rect 106 450 112 482
rect 64 440 112 450
rect 148 506 248 522
rect 345 543 399 590
rect 345 511 355 543
rect 387 511 399 543
rect 345 508 399 511
rect 468 622 596 626
rect 468 590 544 622
rect 576 590 596 622
rect 468 543 596 590
rect 468 511 544 543
rect 576 511 596 543
rect 468 508 596 511
rect 148 474 214 506
rect 246 474 248 506
rect 148 461 248 474
rect 64 274 112 288
rect 64 242 75 274
rect 107 242 112 274
rect 64 206 112 242
rect 64 174 75 206
rect 107 174 112 206
rect 64 44 112 174
rect 148 199 180 461
rect 284 434 496 468
rect 284 392 316 434
rect 248 380 316 392
rect 248 348 265 380
rect 297 348 316 380
rect 248 314 316 348
rect 352 363 415 392
rect 352 331 379 363
rect 411 331 415 363
rect 352 305 415 331
rect 451 380 496 434
rect 534 463 596 508
rect 636 622 688 712
rect 636 590 646 622
rect 678 590 688 622
rect 636 520 688 590
rect 636 488 646 520
rect 678 488 688 520
rect 636 484 688 488
rect 534 431 544 463
rect 576 448 596 463
rect 576 431 714 448
rect 534 416 714 431
rect 451 363 539 380
rect 451 331 503 363
rect 535 331 539 363
rect 451 305 539 331
rect 586 353 646 370
rect 586 321 611 353
rect 643 321 646 353
rect 586 304 646 321
rect 242 274 294 278
rect 242 242 252 274
rect 284 268 294 274
rect 586 268 620 304
rect 284 242 620 268
rect 682 263 714 416
rect 242 236 620 242
rect 663 249 714 263
rect 242 206 294 236
rect 242 199 252 206
rect 148 174 252 199
rect 284 174 294 206
rect 663 217 673 249
rect 705 217 714 249
rect 148 167 294 174
rect 345 195 613 200
rect 345 163 355 195
rect 387 166 571 195
rect 387 163 405 166
rect 345 160 405 163
rect 554 163 571 166
rect 603 163 613 195
rect 554 158 613 163
rect 663 165 714 217
rect 663 133 673 165
rect 705 133 714 165
rect 453 128 505 130
rect 453 96 463 128
rect 495 96 505 128
rect 663 121 714 133
rect 453 44 505 96
rect 0 16 768 44
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 608 16
rect 640 -16 704 16
rect 736 -16 768 16
rect 0 -44 768 -16
<< labels >>
flabel metal1 s 534 416 596 626 0 FreeSans 400 0 0 0 Y
port 2 nsew
flabel metal1 s 248 314 316 392 0 FreeSans 400 0 0 0 B
port 3 nsew
flabel metal1 s 0 712 768 800 0 FreeSans 400 0 0 0 VDD
port 4 nsew
flabel metal1 s 352 305 415 392 0 FreeSans 400 0 0 0 A
port 5 nsew
flabel metal1 s 0 -44 768 44 0 FreeSans 400 0 0 0 VSS
port 6 nsew
<< properties >>
string FIXED_BBOX 0 0 768 756
string GDS_END 72138
string GDS_FILE ../gds/controller.gds
string GDS_START 65828
<< end >>
