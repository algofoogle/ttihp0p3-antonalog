magic
tech ihp-sg13g2
magscale 1 2
timestamp 1746816402
<< nwell >>
rect -48 350 1296 834
<< pwell >>
rect 1 56 1236 292
rect -26 -56 1274 56
<< nmos >>
rect 96 118 122 266
rect 198 118 224 266
rect 300 118 326 266
rect 402 118 428 266
rect 504 118 530 266
rect 606 118 632 266
rect 708 118 734 266
rect 810 118 836 266
rect 912 118 938 266
rect 1014 118 1040 266
rect 1116 118 1142 266
<< pmos >>
rect 96 412 122 636
rect 198 412 224 636
rect 300 412 326 636
rect 402 412 428 636
rect 504 412 530 636
rect 606 412 632 636
rect 708 412 734 636
rect 810 412 836 636
rect 912 412 938 636
rect 1014 412 1040 636
rect 1116 412 1142 636
<< ndiff >>
rect 27 251 96 266
rect 27 219 42 251
rect 74 219 96 251
rect 27 165 96 219
rect 27 133 42 165
rect 74 133 96 165
rect 27 118 96 133
rect 122 195 198 266
rect 122 163 144 195
rect 176 163 198 195
rect 122 118 198 163
rect 224 251 300 266
rect 224 219 246 251
rect 278 219 300 251
rect 224 165 300 219
rect 224 133 246 165
rect 278 133 300 165
rect 224 118 300 133
rect 326 195 402 266
rect 326 163 348 195
rect 380 163 402 195
rect 326 118 402 163
rect 428 251 504 266
rect 428 219 450 251
rect 482 219 504 251
rect 428 165 504 219
rect 428 133 450 165
rect 482 133 504 165
rect 428 118 504 133
rect 530 185 606 266
rect 530 153 552 185
rect 584 153 606 185
rect 530 118 606 153
rect 632 251 708 266
rect 632 219 654 251
rect 686 219 708 251
rect 632 165 708 219
rect 632 133 654 165
rect 686 133 708 165
rect 632 118 708 133
rect 734 185 810 266
rect 734 153 756 185
rect 788 153 810 185
rect 734 118 810 153
rect 836 251 912 266
rect 836 219 858 251
rect 890 219 912 251
rect 836 165 912 219
rect 836 133 858 165
rect 890 133 912 165
rect 836 118 912 133
rect 938 185 1014 266
rect 938 153 960 185
rect 992 153 1014 185
rect 938 118 1014 153
rect 1040 251 1116 266
rect 1040 219 1062 251
rect 1094 219 1116 251
rect 1040 165 1116 219
rect 1040 133 1062 165
rect 1094 133 1116 165
rect 1040 118 1116 133
rect 1142 251 1210 266
rect 1142 219 1164 251
rect 1196 219 1210 251
rect 1142 165 1210 219
rect 1142 133 1164 165
rect 1196 133 1210 165
rect 1142 118 1210 133
<< pdiff >>
rect 28 621 96 636
rect 28 589 42 621
rect 74 589 96 621
rect 28 551 96 589
rect 28 519 42 551
rect 74 519 96 551
rect 28 481 96 519
rect 28 449 42 481
rect 74 449 96 481
rect 28 412 96 449
rect 122 621 198 636
rect 122 589 144 621
rect 176 589 198 621
rect 122 551 198 589
rect 122 519 144 551
rect 176 519 198 551
rect 122 412 198 519
rect 224 621 300 636
rect 224 589 246 621
rect 278 589 300 621
rect 224 551 300 589
rect 224 519 246 551
rect 278 519 300 551
rect 224 481 300 519
rect 224 449 246 481
rect 278 449 300 481
rect 224 412 300 449
rect 326 621 402 636
rect 326 589 348 621
rect 380 589 402 621
rect 326 550 402 589
rect 326 518 348 550
rect 380 518 402 550
rect 326 412 402 518
rect 428 621 504 636
rect 428 589 450 621
rect 482 589 504 621
rect 428 540 504 589
rect 428 508 450 540
rect 482 508 504 540
rect 428 459 504 508
rect 428 427 450 459
rect 482 427 504 459
rect 428 412 504 427
rect 530 621 606 636
rect 530 589 552 621
rect 584 589 606 621
rect 530 521 606 589
rect 530 489 552 521
rect 584 489 606 521
rect 530 412 606 489
rect 632 621 708 636
rect 632 589 654 621
rect 686 589 708 621
rect 632 540 708 589
rect 632 508 654 540
rect 686 508 708 540
rect 632 459 708 508
rect 632 427 654 459
rect 686 427 708 459
rect 632 412 708 427
rect 734 621 810 636
rect 734 589 756 621
rect 788 589 810 621
rect 734 521 810 589
rect 734 489 756 521
rect 788 489 810 521
rect 734 412 810 489
rect 836 621 912 636
rect 836 589 858 621
rect 890 589 912 621
rect 836 540 912 589
rect 836 508 858 540
rect 890 508 912 540
rect 836 459 912 508
rect 836 427 858 459
rect 890 427 912 459
rect 836 412 912 427
rect 938 621 1014 636
rect 938 589 960 621
rect 992 589 1014 621
rect 938 521 1014 589
rect 938 489 960 521
rect 992 489 1014 521
rect 938 412 1014 489
rect 1040 621 1116 636
rect 1040 589 1062 621
rect 1094 589 1116 621
rect 1040 540 1116 589
rect 1040 508 1062 540
rect 1094 508 1116 540
rect 1040 459 1116 508
rect 1040 427 1062 459
rect 1094 427 1116 459
rect 1040 412 1116 427
rect 1142 621 1211 636
rect 1142 589 1164 621
rect 1196 589 1211 621
rect 1142 540 1211 589
rect 1142 508 1164 540
rect 1196 508 1211 540
rect 1142 459 1211 508
rect 1142 427 1164 459
rect 1196 427 1211 459
rect 1142 412 1211 427
<< ndiffc >>
rect 42 219 74 251
rect 42 133 74 165
rect 144 163 176 195
rect 246 219 278 251
rect 246 133 278 165
rect 348 163 380 195
rect 450 219 482 251
rect 450 133 482 165
rect 552 153 584 185
rect 654 219 686 251
rect 654 133 686 165
rect 756 153 788 185
rect 858 219 890 251
rect 858 133 890 165
rect 960 153 992 185
rect 1062 219 1094 251
rect 1062 133 1094 165
rect 1164 219 1196 251
rect 1164 133 1196 165
<< pdiffc >>
rect 42 589 74 621
rect 42 519 74 551
rect 42 449 74 481
rect 144 589 176 621
rect 144 519 176 551
rect 246 589 278 621
rect 246 519 278 551
rect 246 449 278 481
rect 348 589 380 621
rect 348 518 380 550
rect 450 589 482 621
rect 450 508 482 540
rect 450 427 482 459
rect 552 589 584 621
rect 552 489 584 521
rect 654 589 686 621
rect 654 508 686 540
rect 654 427 686 459
rect 756 589 788 621
rect 756 489 788 521
rect 858 589 890 621
rect 858 508 890 540
rect 858 427 890 459
rect 960 589 992 621
rect 960 489 992 521
rect 1062 589 1094 621
rect 1062 508 1094 540
rect 1062 427 1094 459
rect 1164 589 1196 621
rect 1164 508 1196 540
rect 1164 427 1196 459
<< psubdiff >>
rect 0 16 1248 30
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 608 16
rect 640 -16 704 16
rect 736 -16 800 16
rect 832 -16 896 16
rect 928 -16 992 16
rect 1024 -16 1088 16
rect 1120 -16 1184 16
rect 1216 -16 1248 16
rect 0 -30 1248 -16
<< nsubdiff >>
rect 0 772 1248 786
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 608 772
rect 640 740 704 772
rect 736 740 800 772
rect 832 740 896 772
rect 928 740 992 772
rect 1024 740 1088 772
rect 1120 740 1184 772
rect 1216 740 1248 772
rect 0 726 1248 740
<< psubdiffcont >>
rect 32 -16 64 16
rect 128 -16 160 16
rect 224 -16 256 16
rect 320 -16 352 16
rect 416 -16 448 16
rect 512 -16 544 16
rect 608 -16 640 16
rect 704 -16 736 16
rect 800 -16 832 16
rect 896 -16 928 16
rect 992 -16 1024 16
rect 1088 -16 1120 16
rect 1184 -16 1216 16
<< nsubdiffcont >>
rect 32 740 64 772
rect 128 740 160 772
rect 224 740 256 772
rect 320 740 352 772
rect 416 740 448 772
rect 512 740 544 772
rect 608 740 640 772
rect 704 740 736 772
rect 800 740 832 772
rect 896 740 928 772
rect 992 740 1024 772
rect 1088 740 1120 772
rect 1184 740 1216 772
<< poly >>
rect 96 636 122 672
rect 198 636 224 672
rect 300 636 326 672
rect 402 636 428 672
rect 504 636 530 672
rect 606 636 632 672
rect 708 636 734 672
rect 810 636 836 672
rect 912 636 938 672
rect 1014 636 1040 672
rect 1116 636 1142 672
rect 96 380 122 412
rect 198 380 224 412
rect 300 380 326 412
rect 96 363 326 380
rect 402 370 428 412
rect 504 370 530 412
rect 606 370 632 412
rect 708 370 734 412
rect 810 370 836 412
rect 912 370 938 412
rect 1014 370 1040 412
rect 1116 370 1142 412
rect 96 331 124 363
rect 156 331 192 363
rect 224 331 260 363
rect 292 331 326 363
rect 96 314 326 331
rect 96 266 122 314
rect 198 266 224 314
rect 300 266 326 314
rect 385 353 1142 370
rect 385 321 402 353
rect 434 321 470 353
rect 502 321 538 353
rect 570 321 606 353
rect 638 321 674 353
rect 706 321 742 353
rect 774 321 810 353
rect 842 321 878 353
rect 910 321 946 353
rect 978 321 1142 353
rect 385 304 1142 321
rect 385 298 428 304
rect 402 266 428 298
rect 504 266 530 304
rect 606 266 632 304
rect 708 266 734 304
rect 810 266 836 304
rect 912 266 938 304
rect 1014 266 1040 304
rect 1116 266 1142 304
rect 96 82 122 118
rect 198 82 224 118
rect 300 82 326 118
rect 402 82 428 118
rect 504 82 530 118
rect 606 82 632 118
rect 708 82 734 118
rect 810 82 836 118
rect 912 82 938 118
rect 1014 82 1040 118
rect 1116 82 1142 118
<< polycont >>
rect 124 331 156 363
rect 192 331 224 363
rect 260 331 292 363
rect 402 321 434 353
rect 470 321 502 353
rect 538 321 570 353
rect 606 321 638 353
rect 674 321 706 353
rect 742 321 774 353
rect 810 321 842 353
rect 878 321 910 353
rect 946 321 978 353
<< metal1 >>
rect 0 772 1248 800
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 608 772
rect 640 740 704 772
rect 736 740 800 772
rect 832 740 896 772
rect 928 740 992 772
rect 1024 740 1088 772
rect 1120 740 1184 772
rect 1216 740 1248 772
rect 0 712 1248 740
rect 32 621 84 625
rect 32 589 42 621
rect 74 589 84 621
rect 32 551 84 589
rect 32 519 42 551
rect 74 519 84 551
rect 32 481 84 519
rect 134 621 186 712
rect 134 589 144 621
rect 176 589 186 621
rect 134 551 186 589
rect 134 519 144 551
rect 176 519 186 551
rect 134 515 186 519
rect 236 621 288 625
rect 236 589 246 621
rect 278 589 288 621
rect 236 551 288 589
rect 236 519 246 551
rect 278 519 288 551
rect 32 449 42 481
rect 74 468 84 481
rect 236 481 288 519
rect 338 621 390 712
rect 338 589 348 621
rect 380 589 390 621
rect 338 550 390 589
rect 338 518 348 550
rect 380 518 390 550
rect 338 515 390 518
rect 440 621 492 624
rect 440 589 450 621
rect 482 589 492 621
rect 440 540 492 589
rect 236 468 246 481
rect 74 449 246 468
rect 278 468 288 481
rect 440 508 450 540
rect 482 508 492 540
rect 278 449 388 468
rect 32 434 388 449
rect 59 363 310 390
rect 59 331 124 363
rect 156 331 192 363
rect 224 331 260 363
rect 292 331 310 363
rect 59 314 310 331
rect 354 363 388 434
rect 440 459 492 508
rect 542 621 594 712
rect 542 589 552 621
rect 584 589 594 621
rect 542 521 594 589
rect 542 489 552 521
rect 584 489 594 521
rect 542 486 594 489
rect 644 621 696 625
rect 644 589 654 621
rect 686 589 696 621
rect 644 540 696 589
rect 644 508 654 540
rect 686 508 696 540
rect 440 427 450 459
rect 482 446 492 459
rect 644 459 696 508
rect 746 621 798 712
rect 746 589 756 621
rect 788 589 798 621
rect 746 521 798 589
rect 746 489 756 521
rect 788 489 798 521
rect 746 486 798 489
rect 848 621 900 626
rect 848 589 858 621
rect 890 589 900 621
rect 848 540 900 589
rect 848 508 858 540
rect 890 508 900 540
rect 644 446 654 459
rect 482 427 654 446
rect 686 446 696 459
rect 848 459 900 508
rect 950 621 1002 712
rect 950 589 960 621
rect 992 589 1002 621
rect 950 521 1002 589
rect 950 489 960 521
rect 992 489 1002 521
rect 950 484 1002 489
rect 1052 621 1104 624
rect 1052 589 1062 621
rect 1094 589 1104 621
rect 1052 540 1104 589
rect 1052 508 1062 540
rect 1094 508 1104 540
rect 848 446 858 459
rect 686 427 858 446
rect 890 446 900 459
rect 1052 459 1104 508
rect 1052 446 1062 459
rect 890 427 1062 446
rect 1094 427 1104 459
rect 440 414 1104 427
rect 1154 621 1206 712
rect 1154 589 1164 621
rect 1196 589 1206 621
rect 1154 540 1206 589
rect 1154 508 1164 540
rect 1196 508 1206 540
rect 1154 459 1206 508
rect 1154 427 1164 459
rect 1196 427 1206 459
rect 1154 424 1206 427
rect 354 353 995 363
rect 354 321 402 353
rect 434 321 470 353
rect 502 321 538 353
rect 570 321 606 353
rect 638 321 674 353
rect 706 321 742 353
rect 774 321 810 353
rect 842 321 878 353
rect 910 321 946 353
rect 978 321 995 353
rect 354 311 995 321
rect 354 270 388 311
rect 32 251 388 270
rect 1052 260 1104 414
rect 32 219 42 251
rect 74 236 246 251
rect 74 219 84 236
rect 32 165 84 219
rect 236 219 246 236
rect 278 236 388 251
rect 440 251 1104 260
rect 278 219 288 236
rect 32 133 42 165
rect 74 133 84 165
rect 32 128 84 133
rect 134 195 186 199
rect 134 163 144 195
rect 176 163 186 195
rect 134 44 186 163
rect 236 165 288 219
rect 440 219 450 251
rect 482 226 654 251
rect 482 219 492 226
rect 236 133 246 165
rect 278 133 288 165
rect 236 129 288 133
rect 338 195 390 198
rect 338 163 348 195
rect 380 163 390 195
rect 338 44 390 163
rect 440 165 492 219
rect 644 219 654 226
rect 686 226 858 251
rect 686 219 696 226
rect 440 133 450 165
rect 482 133 492 165
rect 440 129 492 133
rect 542 185 594 190
rect 542 153 552 185
rect 584 153 594 185
rect 542 44 594 153
rect 644 165 696 219
rect 848 219 858 226
rect 890 226 1062 251
rect 890 219 900 226
rect 644 133 654 165
rect 686 133 696 165
rect 644 128 696 133
rect 746 185 798 190
rect 746 153 756 185
rect 788 153 798 185
rect 746 44 798 153
rect 848 165 900 219
rect 1052 219 1062 226
rect 1094 219 1104 251
rect 848 133 858 165
rect 890 133 900 165
rect 848 129 900 133
rect 950 185 1002 189
rect 950 153 960 185
rect 992 153 1002 185
rect 950 44 1002 153
rect 1052 165 1104 219
rect 1052 133 1062 165
rect 1094 133 1104 165
rect 1052 130 1104 133
rect 1154 251 1206 255
rect 1154 219 1164 251
rect 1196 219 1206 251
rect 1154 165 1206 219
rect 1154 133 1164 165
rect 1196 133 1206 165
rect 1154 44 1206 133
rect 0 16 1248 44
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 608 16
rect 640 -16 704 16
rect 736 -16 800 16
rect 832 -16 896 16
rect 928 -16 992 16
rect 1024 -16 1088 16
rect 1120 -16 1184 16
rect 1216 -16 1248 16
rect 0 -44 1248 -16
<< labels >>
flabel metal1 s 440 226 1104 260 0 FreeSans 400 0 0 0 X
port 2 nsew
flabel metal1 s 0 712 1248 800 0 FreeSans 400 0 0 0 VDD
port 3 nsew
flabel metal1 s 59 314 310 390 0 FreeSans 400 0 0 0 A
port 4 nsew
flabel metal1 s 0 -44 1248 44 0 FreeSans 400 0 0 0 VSS
port 5 nsew
<< properties >>
string FIXED_BBOX 0 0 1248 756
string GDS_END 247864
string GDS_FILE ../gds/controller.gds
string GDS_START 237696
<< end >>
