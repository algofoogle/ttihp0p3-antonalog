magic
tech ihp-sg13g2
magscale 1 2
timestamp 1746816402
<< nwell >>
rect -48 350 432 834
<< pwell >>
rect 33 56 343 298
rect -26 -56 410 56
<< nmos >>
rect 127 195 153 272
rect 223 96 249 272
<< pmos >>
rect 127 494 153 554
rect 223 451 249 660
<< ndiff >>
rect 59 250 127 272
rect 59 218 73 250
rect 105 218 127 250
rect 59 195 127 218
rect 153 195 223 272
rect 167 141 223 195
rect 59 103 223 141
rect 59 71 114 103
rect 146 96 223 103
rect 249 238 317 272
rect 249 206 271 238
rect 303 206 317 238
rect 249 142 317 206
rect 249 110 271 142
rect 303 110 317 142
rect 249 96 317 110
rect 146 71 203 96
rect 59 36 203 71
<< pdiff >>
rect 59 676 203 720
rect 59 644 108 676
rect 140 660 203 676
rect 140 644 223 660
rect 59 608 223 644
rect 171 554 223 608
rect 59 540 127 554
rect 59 508 73 540
rect 105 508 127 540
rect 59 494 127 508
rect 153 494 223 554
rect 177 451 223 494
rect 249 565 317 660
rect 249 533 271 565
rect 303 533 317 565
rect 249 497 317 533
rect 249 465 271 497
rect 303 465 317 497
rect 249 451 317 465
<< ndiffc >>
rect 73 218 105 250
rect 114 71 146 103
rect 271 206 303 238
rect 271 110 303 142
<< pdiffc >>
rect 108 644 140 676
rect 73 508 105 540
rect 271 533 303 565
rect 271 465 303 497
<< psubdiff >>
rect 59 30 203 36
rect 0 16 384 30
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 384 16
rect 0 -30 384 -16
<< nsubdiff >>
rect 0 772 384 786
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 384 772
rect 0 726 384 740
rect 59 720 203 726
<< psubdiffcont >>
rect 32 -16 64 16
rect 128 -16 160 16
rect 224 -16 256 16
rect 320 -16 352 16
<< nsubdiffcont >>
rect 32 740 64 772
rect 128 740 160 772
rect 224 740 256 772
rect 320 740 352 772
<< poly >>
rect 223 660 249 698
rect 127 554 153 592
rect 127 478 153 494
rect 59 464 153 478
rect 59 432 73 464
rect 105 452 153 464
rect 105 432 135 452
rect 59 418 135 432
rect 109 314 135 418
rect 223 416 249 451
rect 171 402 249 416
rect 171 370 185 402
rect 217 387 249 402
rect 217 370 231 387
rect 171 363 231 370
rect 171 362 230 363
rect 171 361 229 362
rect 171 360 228 361
rect 171 359 227 360
rect 171 358 226 359
rect 171 357 225 358
rect 171 356 224 357
rect 267 347 320 348
rect 266 346 320 347
rect 265 345 320 346
rect 264 344 320 345
rect 263 343 320 344
rect 262 342 320 343
rect 261 341 320 342
rect 260 334 320 341
rect 260 314 274 334
rect 109 288 153 314
rect 127 272 153 288
rect 223 302 274 314
rect 306 302 320 334
rect 223 288 320 302
rect 223 272 249 288
rect 127 157 153 195
rect 223 58 249 96
<< polycont >>
rect 73 432 105 464
rect 185 370 217 402
rect 274 302 306 334
<< metal1 >>
rect 0 772 384 800
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 384 772
rect 0 712 384 740
rect 91 676 156 712
rect 91 644 108 676
rect 140 644 156 676
rect 91 633 156 644
rect 261 565 316 575
rect 63 540 115 552
rect 63 508 73 540
rect 105 508 115 540
rect 63 464 115 508
rect 63 432 73 464
rect 105 432 115 464
rect 63 422 115 432
rect 261 533 271 565
rect 303 533 316 565
rect 261 497 316 533
rect 261 465 271 497
rect 303 465 316 497
rect 175 402 223 412
rect 175 370 185 402
rect 217 370 223 402
rect 175 258 223 370
rect 261 334 316 465
rect 261 302 274 334
rect 306 302 316 334
rect 261 292 316 302
rect 63 250 223 258
rect 63 218 73 250
rect 105 218 223 250
rect 63 206 223 218
rect 259 238 317 246
rect 259 206 271 238
rect 303 206 317 238
rect 259 155 317 206
rect 219 142 317 155
rect 93 103 163 121
rect 93 71 114 103
rect 146 71 163 103
rect 219 110 271 142
rect 303 110 317 142
rect 219 97 317 110
rect 93 44 163 71
rect 0 16 384 44
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 384 16
rect 0 -44 384 -16
<< labels >>
flabel metal1 s 259 97 317 246 0 FreeSans 400 0 0 0 L_LO
port 2 nsew
flabel metal1 s 0 712 384 800 0 FreeSans 400 0 0 0 VDD
port 3 nsew
flabel metal1 s 0 -44 384 44 0 FreeSans 400 0 0 0 VSS
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 384 756
string GDS_END 257808
string GDS_FILE ../gds/controller.gds
string GDS_START 254068
<< end >>
