magic
tech ihp-sg13g2
magscale 1 2
timestamp 1747056038
<< nwell >>
rect -48 350 720 834
<< pwell >>
rect 50 56 672 314
rect -26 -56 698 56
<< nmos >>
rect 144 160 170 288
rect 246 160 272 288
rect 348 160 374 288
rect 450 140 476 288
rect 552 140 578 288
<< pmos >>
rect 144 471 170 639
rect 246 471 272 639
rect 348 471 374 639
rect 450 434 476 658
rect 552 434 578 658
<< ndiff >>
rect 76 253 144 288
rect 76 221 90 253
rect 122 221 144 253
rect 76 160 144 221
rect 170 160 246 288
rect 272 160 348 288
rect 374 210 450 288
rect 374 178 396 210
rect 428 178 450 210
rect 374 160 450 178
rect 388 140 450 160
rect 476 263 552 288
rect 476 231 498 263
rect 530 231 552 263
rect 476 195 552 231
rect 476 163 498 195
rect 530 163 552 195
rect 476 140 552 163
rect 578 195 646 288
rect 578 163 600 195
rect 632 163 646 195
rect 578 140 646 163
<< pdiff >>
rect 388 639 450 658
rect 76 618 144 639
rect 76 586 90 618
rect 122 586 144 618
rect 76 527 144 586
rect 76 495 90 527
rect 122 495 144 527
rect 76 471 144 495
rect 170 580 246 639
rect 170 548 192 580
rect 224 548 246 580
rect 170 471 246 548
rect 272 613 348 639
rect 272 581 294 613
rect 326 581 348 613
rect 272 534 348 581
rect 272 502 294 534
rect 326 502 348 534
rect 272 471 348 502
rect 374 626 450 639
rect 374 594 396 626
rect 428 594 450 626
rect 374 558 450 594
rect 374 526 396 558
rect 428 526 450 558
rect 374 471 450 526
rect 404 434 450 471
rect 476 644 552 658
rect 476 612 498 644
rect 530 612 552 644
rect 476 572 552 612
rect 476 540 498 572
rect 530 540 552 572
rect 476 434 552 540
rect 578 644 648 658
rect 578 612 602 644
rect 634 612 648 644
rect 578 434 648 612
<< ndiffc >>
rect 90 221 122 253
rect 396 178 428 210
rect 498 231 530 263
rect 498 163 530 195
rect 600 163 632 195
<< pdiffc >>
rect 90 586 122 618
rect 90 495 122 527
rect 192 548 224 580
rect 294 581 326 613
rect 294 502 326 534
rect 396 594 428 626
rect 396 526 428 558
rect 498 612 530 644
rect 498 540 530 572
rect 602 612 634 644
<< psubdiff >>
rect 0 16 672 30
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 608 16
rect 640 -16 672 16
rect 0 -30 672 -16
<< nsubdiff >>
rect 0 772 672 786
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 608 772
rect 640 740 672 772
rect 0 726 672 740
<< psubdiffcont >>
rect 32 -16 64 16
rect 128 -16 160 16
rect 224 -16 256 16
rect 320 -16 352 16
rect 416 -16 448 16
rect 512 -16 544 16
rect 608 -16 640 16
<< nsubdiffcont >>
rect 32 740 64 772
rect 128 740 160 772
rect 224 740 256 772
rect 320 740 352 772
rect 416 740 448 772
rect 512 740 544 772
rect 608 740 640 772
<< poly >>
rect 144 639 170 675
rect 246 639 272 675
rect 348 639 374 675
rect 450 658 476 701
rect 552 658 578 700
rect 144 288 170 471
rect 246 396 272 471
rect 348 400 374 471
rect 450 413 476 434
rect 552 413 578 434
rect 218 379 284 396
rect 218 347 235 379
rect 267 347 284 379
rect 218 330 284 347
rect 346 383 412 400
rect 346 351 363 383
rect 395 351 412 383
rect 346 334 412 351
rect 450 396 578 413
rect 450 364 480 396
rect 512 364 578 396
rect 450 347 578 364
rect 246 288 272 330
rect 348 288 374 334
rect 450 288 476 347
rect 552 288 578 347
rect 144 146 170 160
rect 70 132 204 146
rect 70 100 87 132
rect 119 100 155 132
rect 187 100 204 132
rect 246 108 272 160
rect 348 109 374 160
rect 450 104 476 140
rect 552 103 578 140
rect 70 78 204 100
<< polycont >>
rect 235 347 267 379
rect 363 351 395 383
rect 480 364 512 396
rect 87 100 119 132
rect 155 100 187 132
<< metal1 >>
rect 0 772 672 800
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 608 772
rect 640 740 672 772
rect 0 712 672 740
rect 80 618 132 623
rect 80 586 90 618
rect 122 586 132 618
rect 80 527 132 586
rect 182 580 234 712
rect 386 626 438 712
rect 182 548 192 580
rect 224 548 234 580
rect 182 546 234 548
rect 284 613 336 617
rect 284 581 294 613
rect 326 581 336 613
rect 80 495 90 527
rect 122 495 132 527
rect 80 464 132 495
rect 284 534 336 581
rect 284 502 294 534
rect 326 502 336 534
rect 386 594 396 626
rect 428 594 438 626
rect 386 558 438 594
rect 386 526 396 558
rect 428 526 438 558
rect 386 523 438 526
rect 487 644 541 672
rect 487 612 498 644
rect 530 612 541 644
rect 487 572 541 612
rect 591 644 645 712
rect 591 612 602 644
rect 634 612 645 644
rect 591 575 645 612
rect 487 540 498 572
rect 530 540 541 572
rect 487 538 541 540
rect 487 502 613 538
rect 284 464 336 502
rect 80 432 481 464
rect 80 253 132 432
rect 449 413 481 432
rect 449 396 529 413
rect 218 379 308 396
rect 218 347 235 379
rect 267 347 308 379
rect 218 280 308 347
rect 346 383 412 390
rect 346 351 363 383
rect 395 351 412 383
rect 346 280 412 351
rect 449 364 480 396
rect 512 364 529 396
rect 449 347 529 364
rect 567 310 613 502
rect 80 221 90 253
rect 122 221 132 253
rect 488 263 613 310
rect 488 231 498 263
rect 530 258 613 263
rect 530 231 540 258
rect 80 218 132 221
rect 245 158 318 218
rect 70 132 318 158
rect 70 100 87 132
rect 119 100 155 132
rect 187 100 318 132
rect 70 95 318 100
rect 386 210 438 228
rect 386 178 396 210
rect 428 178 438 210
rect 386 44 438 178
rect 488 195 540 231
rect 488 163 498 195
rect 530 163 540 195
rect 488 154 540 163
rect 590 195 642 218
rect 590 163 600 195
rect 632 163 642 195
rect 590 44 642 163
rect 0 16 672 44
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 608 16
rect 640 -16 672 16
rect 0 -44 672 -16
<< labels >>
flabel metal1 s 488 258 613 310 0 FreeSans 400 0 0 0 X
port 2 nsew
flabel metal1 s 218 280 308 396 0 FreeSans 400 0 0 0 B
port 3 nsew
flabel metal1 s 0 712 672 800 0 FreeSans 400 0 0 0 VDD
port 4 nsew
flabel metal1 s 0 -44 672 44 0 FreeSans 400 0 0 0 VSS
port 5 nsew
flabel metal1 s 346 280 412 390 0 FreeSans 400 0 0 0 C
port 6 nsew
flabel metal1 s 245 95 318 218 0 FreeSans 400 0 0 0 A
port 7 nsew
<< properties >>
string FIXED_BBOX 0 0 672 756
string GDS_END 206726
string GDS_FILE ../gds/controller.gds
string GDS_START 200978
<< end >>
