* NGSPICE file created from r2r_dac_parax.ext - technology: ihp-sg13g2

.subckt r2r_dac_parax IN[0] IN[1] IN[2] IN[3] IN[4] IN[5] IN[6] IN[7] OUT GND
X0 IN[3].t0 wi3 rhigh l=6u w=1u
X1 wJ5 wi5 rhigh l=6u w=1u
X2 wJ1 wJ0 rhigh l=6u w=1u
X3 wJ5 wJ6 rhigh l=6u w=1u
X4 wg0 GND.t0 rhigh l=6u w=1u
X5 wi0 wJ0 rhigh l=6u w=1u
X6 wi4 IN[4].t0 rhigh l=6u w=1u
X7 OUT.t0 wi7 rhigh l=6u w=1u
X8 wi2 wJ2 rhigh l=6u w=1u
X9 wJ3 wJ2 rhigh l=6u w=1u
X10 IN[1].t0 wi1 rhigh l=6u w=1u
X11 wi0 IN[0].t0 rhigh l=6u w=1u
X12 wJ3 wi3 rhigh l=6u w=1u
X13 wJ3 wJ4 rhigh l=6u w=1u
X14 wJ5 wJ4 rhigh l=6u w=1u
X15 IN[5].t0 wi5 rhigh l=6u w=1u
X16 wJ1 wJ2 rhigh l=6u w=1u
X17 wJ1 wi1 rhigh l=6u w=1u
X18 wi6 wJ6 rhigh l=6u w=1u
X19 OUT.t1 wJ6 rhigh l=6u w=1u
X20 wg0 wJ0 rhigh l=6u w=1u
X21 IN[7].t0 wi7 rhigh l=6u w=1u
X22 wi2 IN[2].t0 rhigh l=6u w=1u
X23 wi4 wJ4 rhigh l=6u w=1u
X24 wi6 IN[6].t0 rhigh l=6u w=1u
R0 IN[3] IN[3].t0 5.05324
R1 GND GND.t0 5.03325
R2 IN[4] IN[4].t0 5.05324
R3 OUT.n0 OUT.t0 5.19036
R4 OUT.n0 OUT.t1 5.0005
R5 OUT OUT.n0 0.0532397
R6 IN[1] IN[1].t0 5.05324
R7 IN[0] IN[0].t0 5.05324
R8 IN[5] IN[5].t0 5.05324
R9 IN[7] IN[7].t0 5.05324
R10 IN[2] IN[2].t0 5.05324
R11 IN[6] IN[6].t0 5.05324
C0 a_n1828_n720# wi0 0.0454f
C1 a_n1828_n720# wJ0 0.13277f
C2 IN[3] wJ3 0.21494f
C3 a_1952_n720# wJ6 0.00468f
C4 wJ1 a_n1576_n720# 0.06789f
C5 a_3212_n720# wi7 0.04606f
C6 wJ3 a_440_n720# 0.13277f
C7 a_1448_n720# a_1196_n720# 0.29305f
C8 wJ2 wJ1 0.00581f
C9 wJ2 IN[2] 0.21494f
C10 wJ3 a_n316_n720# 0.00468f
C11 wi6 a_2708_n720# 0.0454f
C12 wi6 a_2456_n720# 0.0454f
C13 wi4 a_1196_n720# 0.0454f
C14 wJ6 IN[6] 0.21494f
C15 a_n1324_n720# wJ1 0.12652f
C16 wJ4 a_440_n720# 0.00468f
C17 wg0 a_n2332_n720# 0.04606f
C18 a_2204_n720# wJ5 0.12652f
C19 wJ2 a_188_n720# 0.02248f
C20 wi5 a_1700_n720# 0.0454f
C21 a_1952_n720# IN[5] 0.02298f
C22 wi5 wJ5 0.01312f
C23 a_n568_n720# a_n316_n720# 0.29305f
C24 IN[4] IN[2] 0.00132f
C25 a_440_n720# wi3 0.0454f
C26 wJ0 wi0 0.01312f
C27 wg0 a_n2584_n720# 0.04606f
C28 a_n1828_n720# a_n2080_n720# 0.29305f
C29 wJ2 a_n1072_n720# 0.00468f
C30 wi2 a_n316_n720# 0.0454f
C31 wJ3 wJ5 0.0072f
C32 OUT wi7 0.00483f
C33 wJ0 wi1 0.07984f
C34 a_3464_n720# wJ6 0.00468f
C35 a_2204_n720# wJ6 0.06789f
C36 a_n1072_n720# a_n1324_n720# 0.29305f
C37 wJ5 a_2708_n720# 0.00468f
C38 wJ5 a_2456_n720# 0.02248f
C39 wJ4 a_1700_n720# 0.02248f
C40 wJ3 wJ1 0.0072f
C41 wJ4 wJ5 0.00581f
C42 wi5 wJ6 0.07984f
C43 a_n64_n720# a_n316_n720# 0.29305f
C44 a_n1324_n720# a_n1576_n720# 0.29305f
C45 a_3212_n720# a_2960_n720# 0.29305f
C46 a_692_n720# a_440_n720# 0.29305f
C47 a_2204_n720# a_1952_n720# 0.29305f
C48 wJ2 a_n1324_n720# 0.00183f
C49 wJ3 a_188_n720# 0.12652f
C50 a_2708_n720# wJ6 0.13277f
C51 a_n568_n720# wJ1 0.02248f
C52 wJ6 a_2456_n720# 0.12652f
C53 wi5 a_1952_n720# 0.0454f
C54 wi0 a_n2080_n720# 0.0454f
C55 IN[0] IN[2] 0.00132f
C56 IN[4] IN[6] 0.00132f
C57 wJ4 wJ6 0.0072f
C58 wJ0 a_n2080_n720# 0.12652f
C59 wi2 wJ1 0.07984f
C60 IN[3] IN[1] 0.00132f
C61 wJ1 a_n820_n720# 0.12652f
C62 wJ4 a_188_n720# 0.00183f
C63 OUT a_3212_n720# 0.04606f
C64 a_n1828_n720# wJ1 0.00468f
C65 a_1196_n720# wJ5 0.00468f
C66 wJ3 a_944_n720# 0.02248f
C67 OUT a_2960_n720# 0.0454f
C68 wJ4 a_1952_n720# 0.00468f
C69 IN[7] a_3464_n720# 0.04606f
C70 a_188_n720# wi3 0.0454f
C71 a_n64_n720# wJ1 0.00183f
C72 wJ6 wi7 0.07984f
C73 wJ2 wJ3 0.00581f
C74 a_1448_n720# a_1700_n720# 0.29305f
C75 a_1448_n720# wJ5 0.06789f
C76 wJ4 a_944_n720# 0.12652f
C77 wg0 wi0 0.07984f
C78 a_2708_n720# IN[6] 0.02298f
C79 a_n1072_n720# a_n820_n720# 0.29305f
C80 wg0 wJ0 0.00483f
C81 a_n64_n720# a_188_n720# 0.29305f
C82 IN[3] a_440_n720# 0.02298f
C83 wi4 wJ5 0.07984f
C84 wJ2 wJ4 0.0072f
C85 wJ2 a_n568_n720# 0.12652f
C86 wi6 OUT 0.07984f
C87 wJ1 wi0 0.07984f
C88 a_n1828_n720# a_n1576_n720# 0.29305f
C89 wJ2 wi2 0.01312f
C90 wJ2 a_n820_n720# 0.06789f
C91 wJ5 a_2960_n720# 0.00183f
C92 wJ1 wJ0 0.00581f
C93 wJ2 wi3 0.07984f
C94 wJ1 wi1 0.01312f
C95 IN[1] wJ1 0.21494f
C96 a_n2584_n720# a_n2332_n720# 0.29305f
C97 a_2204_n720# a_2456_n720# 0.29305f
C98 wJ4 IN[4] 0.21494f
C99 a_2204_n720# wJ4 0.00183f
C100 a_1196_n720# a_944_n720# 0.29305f
C101 wJ6 a_3212_n720# 0.02248f
C102 wJ2 a_n64_n720# 0.12652f
C103 a_692_n720# a_944_n720# 0.29305f
C104 wJ4 wi5 0.07984f
C105 IN[7] wi7 0.00483f
C106 wJ6 a_2960_n720# 0.12652f
C107 wi6 wJ5 0.07984f
C108 a_n1072_n720# wJ0 0.00468f
C109 wJ4 wJ3 0.00581f
C110 a_3464_n720# wi7 0.04606f
C111 a_n1072_n720# wi1 0.0454f
C112 wJ2 a_692_n720# 0.00183f
C113 a_n1072_n720# IN[1] 0.02298f
C114 a_2708_n720# a_2456_n720# 0.29305f
C115 wJ3 a_n568_n720# 0.00183f
C116 wi4 a_944_n720# 0.0454f
C117 wJ1 a_n2080_n720# 0.00183f
C118 wJ0 a_n1576_n720# 0.12652f
C119 wJ3 wi2 0.07984f
C120 IN[4] a_1196_n720# 0.02298f
C121 wJ3 wi3 0.01312f
C122 wJ1 a_n316_n720# 0.00468f
C123 wJ2 wJ0 0.0072f
C124 a_n316_n720# IN[2] 0.02298f
C125 wi6 wJ6 0.01312f
C126 wJ2 wi1 0.07984f
C127 a_188_n720# a_440_n720# 0.29305f
C128 OUT wJ6 0.00581f
C129 a_n1324_n720# wJ0 0.02248f
C130 a_n1324_n720# wi1 0.0454f
C131 a_1700_n720# wJ5 0.12652f
C132 a_n64_n720# wJ3 0.06789f
C133 wJ4 wi3 0.07984f
C134 wi2 a_n568_n720# 0.0454f
C135 a_n568_n720# a_n820_n720# 0.29305f
C136 wJ3 a_1196_n720# 0.00468f
C137 a_n1828_n720# IN[0] 0.02298f
C138 IN[3] IN[5] 0.00132f
C139 a_3464_n720# a_3212_n720# 0.29305f
C140 a_692_n720# wJ3 0.12652f
C141 wJ0 a_n2332_n720# 0.06854f
C142 OUT IN[5] 0.00216f
C143 a_1448_n720# wJ3 0.00183f
C144 wJ4 a_1196_n720# 0.13277f
C145 a_1700_n720# wJ6 0.00183f
C146 wJ5 wJ6 0.00581f
C147 wJ2 a_440_n720# 0.00468f
C148 a_692_n720# wJ4 0.06789f
C149 wi4 wJ3 0.07984f
C150 a_n2584_n720# wJ0 0.00468f
C151 a_1448_n720# wJ4 0.12652f
C152 wJ2 a_n316_n720# 0.13277f
C153 a_1700_n720# a_1952_n720# 0.29305f
C154 wJ5 a_1952_n720# 0.13277f
C155 IN[7] OUT 0.12089f
C156 wJ4 wi4 0.01312f
C157 a_944_n720# wJ5 0.00183f
C158 IN[0] wJ0 0.21494f
C159 wJ5 IN[5] 0.21494f
C160 a_2708_n720# a_2960_n720# 0.29305f
C161 a_n2332_n720# a_n2080_n720# 0.29305f
C162 a_n1072_n720# wJ1 0.13277f
C163 wJ0 a_n820_n720# 0.00183f
C164 IN[7] GND 0.22507f
C165 OUT GND 0.39088f
C166 IN[6] GND 0.19677f
C167 IN[5] GND 0.19457f
C168 IN[4] GND 0.19552f
C169 IN[3] GND 0.19552f
C170 IN[2] GND 0.19552f
C171 IN[1] GND 0.19688f
C172 IN[0] GND 0.19671f
C173 a_3464_n720# GND 0.87154f $ **FLOATING
C174 wi7 GND 0.35118f
C175 a_3212_n720# GND 0.66978f $ **FLOATING
C176 a_2960_n720# GND 0.66978f $ **FLOATING
C177 a_2708_n720# GND 0.66978f $ **FLOATING
C178 a_2456_n720# GND 0.66978f $ **FLOATING
C179 wi6 GND 0.31577f
C180 wJ6 GND 0.54599f
C181 a_2204_n720# GND 0.66978f $ **FLOATING
C182 a_1952_n720# GND 0.66978f $ **FLOATING
C183 wi5 GND 0.31577f
C184 a_1700_n720# GND 0.66978f $ **FLOATING
C185 a_1448_n720# GND 0.66978f $ **FLOATING
C186 wJ5 GND 0.54102f
C187 a_1196_n720# GND 0.66978f $ **FLOATING
C188 a_944_n720# GND 0.66978f $ **FLOATING
C189 wi4 GND 0.31577f
C190 wJ4 GND 0.536f
C191 a_692_n720# GND 0.66978f $ **FLOATING
C192 a_440_n720# GND 0.66978f $ **FLOATING
C193 wi3 GND 0.31577f
C194 a_188_n720# GND 0.66978f $ **FLOATING
C195 a_n64_n720# GND 0.66978f $ **FLOATING
C196 wJ3 GND 0.536f
C197 a_n316_n720# GND 0.66978f $ **FLOATING
C198 a_n568_n720# GND 0.66978f $ **FLOATING
C199 wi2 GND 0.31577f
C200 wJ2 GND 0.536f
C201 a_n820_n720# GND 0.66978f $ **FLOATING
C202 a_n1072_n720# GND 0.6701f $ **FLOATING
C203 wi1 GND 0.31577f
C204 a_n1324_n720# GND 0.67141f $ **FLOATING
C205 a_n1576_n720# GND 0.67281f $ **FLOATING
C206 wJ1 GND 0.54094f
C207 a_n1828_n720# GND 0.67474f $ **FLOATING
C208 a_n2080_n720# GND 0.67932f $ **FLOATING
C209 wi0 GND 0.31577f
C210 wJ0 GND 0.62584f
C211 a_n2332_n720# GND 0.69982f $ **FLOATING
C212 a_n2584_n720# GND 1.12317f $ **FLOATING
C213 wg0 GND 0.42845f
.ends

