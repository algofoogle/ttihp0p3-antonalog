magic
tech ihp-sg13g2
timestamp 1747537721
<< nwell >>
rect -24 175 312 417
<< pwell >>
rect 15 120 269 146
rect 15 28 275 120
rect -13 -28 301 28
<< nmos >>
rect 62 59 75 133
rect 113 59 126 133
rect 164 59 177 133
rect 215 59 228 133
<< pmos >>
rect 62 206 75 318
rect 104 206 117 318
rect 161 206 174 318
rect 218 206 231 318
<< ndiff >>
rect 28 120 62 133
rect 28 104 35 120
rect 51 104 62 120
rect 28 82 62 104
rect 28 66 35 82
rect 51 66 62 82
rect 28 59 62 66
rect 75 125 113 133
rect 75 109 86 125
rect 102 109 113 125
rect 75 82 113 109
rect 75 66 86 82
rect 102 66 113 82
rect 75 59 113 66
rect 126 97 164 133
rect 126 81 137 97
rect 153 81 164 97
rect 126 59 164 81
rect 177 125 215 133
rect 177 109 188 125
rect 204 109 215 125
rect 177 82 215 109
rect 177 66 188 82
rect 204 66 215 82
rect 177 59 215 66
rect 228 107 256 133
rect 228 93 262 107
rect 228 77 239 93
rect 255 77 262 93
rect 228 59 262 77
<< pdiff >>
rect 28 310 62 318
rect 28 294 35 310
rect 51 294 62 310
rect 28 270 62 294
rect 28 254 35 270
rect 51 254 62 270
rect 28 229 62 254
rect 28 213 35 229
rect 51 213 62 229
rect 28 206 62 213
rect 75 206 104 318
rect 117 206 161 318
rect 174 206 218 318
rect 231 310 267 318
rect 231 294 244 310
rect 260 294 267 310
rect 231 276 267 294
rect 231 260 244 276
rect 260 260 267 276
rect 231 241 267 260
rect 231 225 244 241
rect 260 225 267 241
rect 231 206 267 225
<< ndiffc >>
rect 35 104 51 120
rect 35 66 51 82
rect 86 109 102 125
rect 86 66 102 82
rect 137 81 153 97
rect 188 109 204 125
rect 188 66 204 82
rect 239 77 255 93
<< pdiffc >>
rect 35 294 51 310
rect 35 254 51 270
rect 35 213 51 229
rect 244 294 260 310
rect 244 260 260 276
rect 244 225 260 241
<< psubdiff >>
rect 0 8 288 15
rect 0 -8 16 8
rect 32 -8 64 8
rect 80 -8 112 8
rect 128 -8 160 8
rect 176 -8 208 8
rect 224 -8 256 8
rect 272 -8 288 8
rect 0 -15 288 -8
<< nsubdiff >>
rect 0 386 288 393
rect 0 370 16 386
rect 32 370 64 386
rect 80 370 112 386
rect 128 370 160 386
rect 176 370 208 386
rect 224 370 256 386
rect 272 370 288 386
rect 0 363 288 370
<< psubdiffcont >>
rect 16 -8 32 8
rect 64 -8 80 8
rect 112 -8 128 8
rect 160 -8 176 8
rect 208 -8 224 8
rect 256 -8 272 8
<< nsubdiffcont >>
rect 16 370 32 386
rect 64 370 80 386
rect 112 370 128 386
rect 160 370 176 386
rect 208 370 224 386
rect 256 370 272 386
<< poly >>
rect 62 318 75 336
rect 104 318 117 336
rect 161 318 174 336
rect 218 318 231 336
rect 62 198 75 206
rect 104 198 117 206
rect 161 198 174 206
rect 218 198 231 206
rect 60 177 75 198
rect 26 168 75 177
rect 26 152 34 168
rect 50 152 75 168
rect 93 190 120 198
rect 93 181 126 190
rect 93 165 102 181
rect 118 165 126 181
rect 93 157 126 165
rect 144 181 177 198
rect 144 165 152 181
rect 168 165 177 181
rect 144 157 177 165
rect 195 181 234 198
rect 195 165 208 181
rect 224 165 234 181
rect 195 157 234 165
rect 26 144 75 152
rect 62 133 75 144
rect 113 133 126 157
rect 164 133 177 157
rect 215 133 228 157
rect 62 41 75 59
rect 113 41 126 59
rect 164 41 177 59
rect 215 41 228 59
<< polycont >>
rect 34 152 50 168
rect 102 165 118 181
rect 152 165 168 181
rect 208 165 224 181
<< metal1 >>
rect 0 386 288 400
rect 0 370 16 386
rect 32 370 64 386
rect 80 370 112 386
rect 128 370 160 386
rect 176 370 208 386
rect 224 370 256 386
rect 272 370 288 386
rect 0 356 288 370
rect 30 310 56 356
rect 30 294 35 310
rect 51 294 56 310
rect 30 270 56 294
rect 30 254 35 270
rect 51 254 56 270
rect 30 229 56 254
rect 30 213 35 229
rect 51 213 56 229
rect 30 212 56 213
rect 19 168 63 183
rect 19 152 34 168
rect 50 152 63 168
rect 83 181 126 311
rect 222 310 270 320
rect 222 294 244 310
rect 260 294 270 310
rect 222 276 270 294
rect 222 260 244 276
rect 260 260 270 276
rect 222 241 270 260
rect 83 165 102 181
rect 118 165 126 181
rect 83 157 126 165
rect 144 181 174 237
rect 222 225 244 241
rect 260 225 270 241
rect 222 217 270 225
rect 144 165 152 181
rect 168 165 174 181
rect 144 157 174 165
rect 195 181 232 198
rect 195 165 208 181
rect 224 165 232 181
rect 195 157 232 165
rect 19 141 63 152
rect 250 139 270 217
rect 81 125 270 139
rect 29 120 56 123
rect 29 104 35 120
rect 51 104 56 120
rect 29 82 56 104
rect 29 66 35 82
rect 51 66 56 82
rect 29 22 56 66
rect 81 109 86 125
rect 102 117 188 125
rect 102 109 107 117
rect 81 82 107 109
rect 183 109 188 117
rect 204 117 270 125
rect 204 109 209 117
rect 81 66 86 82
rect 102 66 107 82
rect 81 64 107 66
rect 132 97 158 99
rect 132 81 137 97
rect 153 81 158 97
rect 132 22 158 81
rect 183 82 209 109
rect 183 66 188 82
rect 204 66 209 82
rect 183 64 209 66
rect 234 93 260 96
rect 234 77 239 93
rect 255 77 260 93
rect 234 22 260 77
rect 0 8 288 22
rect 0 -8 16 8
rect 32 -8 64 8
rect 80 -8 112 8
rect 128 -8 160 8
rect 176 -8 208 8
rect 224 -8 256 8
rect 272 -8 288 8
rect 0 -22 288 -8
<< labels >>
flabel metal1 s 0 -22 288 22 0 FreeSans 200 0 0 0 VSS
port 2 nsew
flabel metal1 s 0 356 288 400 0 FreeSans 200 0 0 0 VDD
port 3 nsew
flabel metal1 s 83 157 126 311 0 FreeSans 200 0 0 0 B
port 4 nsew
flabel metal1 s 144 157 174 237 0 FreeSans 200 0 0 0 C
port 5 nsew
flabel metal1 s 222 217 270 320 0 FreeSans 200 0 0 0 Y
port 6 nsew
flabel metal1 s 19 141 63 183 0 FreeSans 200 0 0 0 A
port 7 nsew
flabel metal1 s 195 157 232 198 0 FreeSans 200 0 0 0 D
port 8 nsew
<< properties >>
string FIXED_BBOX 0 0 288 378
string GDS_END 204846
string GDS_FILE ../gds/controller.gds
string GDS_START 199404
<< end >>
