magic
tech ihp-sg13g2
magscale 1 2
timestamp 1747056038
<< nwell >>
rect -48 350 624 834
<< pwell >>
rect 19 56 547 314
rect -26 -56 602 56
<< nmos >>
rect 113 160 139 288
rect 215 160 241 288
rect 317 140 343 288
rect 419 140 445 288
<< pmos >>
rect 113 468 139 636
rect 215 468 241 636
rect 317 412 343 636
rect 419 412 445 636
<< ndiff >>
rect 45 268 113 288
rect 45 236 59 268
rect 91 236 113 268
rect 45 160 113 236
rect 139 160 215 288
rect 241 229 317 288
rect 241 197 263 229
rect 295 197 317 229
rect 241 160 317 197
rect 271 140 317 160
rect 343 269 419 288
rect 343 237 365 269
rect 397 237 419 269
rect 343 191 419 237
rect 343 159 365 191
rect 397 159 419 191
rect 343 140 419 159
rect 445 229 521 288
rect 445 197 467 229
rect 499 197 521 229
rect 445 140 521 197
<< pdiff >>
rect 45 620 113 636
rect 45 588 59 620
rect 91 588 113 620
rect 45 519 113 588
rect 45 487 59 519
rect 91 487 113 519
rect 45 468 113 487
rect 139 620 215 636
rect 139 588 161 620
rect 193 588 215 620
rect 139 519 215 588
rect 139 487 161 519
rect 193 487 215 519
rect 139 468 215 487
rect 241 620 317 636
rect 241 588 263 620
rect 295 588 317 620
rect 241 531 317 588
rect 241 499 263 531
rect 295 499 317 531
rect 241 468 317 499
rect 271 412 317 468
rect 343 620 419 636
rect 343 588 365 620
rect 397 588 419 620
rect 343 543 419 588
rect 343 511 365 543
rect 397 511 419 543
rect 343 463 419 511
rect 343 431 365 463
rect 397 431 419 463
rect 343 412 419 431
rect 445 620 521 636
rect 445 588 467 620
rect 499 588 521 620
rect 445 531 521 588
rect 445 499 467 531
rect 499 499 521 531
rect 445 412 521 499
<< ndiffc >>
rect 59 236 91 268
rect 263 197 295 229
rect 365 237 397 269
rect 365 159 397 191
rect 467 197 499 229
<< pdiffc >>
rect 59 588 91 620
rect 59 487 91 519
rect 161 588 193 620
rect 161 487 193 519
rect 263 588 295 620
rect 263 499 295 531
rect 365 588 397 620
rect 365 511 397 543
rect 365 431 397 463
rect 467 588 499 620
rect 467 499 499 531
<< psubdiff >>
rect 0 16 576 30
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 576 16
rect 0 -30 576 -16
<< nsubdiff >>
rect 0 772 576 786
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 576 772
rect 0 726 576 740
<< psubdiffcont >>
rect 32 -16 64 16
rect 128 -16 160 16
rect 224 -16 256 16
rect 320 -16 352 16
rect 416 -16 448 16
rect 512 -16 544 16
<< nsubdiffcont >>
rect 32 740 64 772
rect 128 740 160 772
rect 224 740 256 772
rect 320 740 352 772
rect 416 740 448 772
rect 512 740 544 772
<< poly >>
rect 113 636 139 672
rect 215 636 241 672
rect 317 636 343 672
rect 419 636 445 672
rect 113 288 139 468
rect 215 380 241 468
rect 317 380 343 412
rect 419 380 445 412
rect 175 363 241 380
rect 175 331 192 363
rect 224 331 241 363
rect 175 314 241 331
rect 277 363 445 380
rect 277 331 306 363
rect 338 331 445 363
rect 277 314 445 331
rect 215 288 241 314
rect 317 288 343 314
rect 419 288 445 314
rect 113 146 139 160
rect 21 128 155 146
rect 21 96 38 128
rect 70 96 106 128
rect 138 96 155 128
rect 215 124 241 160
rect 317 104 343 140
rect 419 104 445 140
rect 21 82 155 96
<< polycont >>
rect 192 331 224 363
rect 306 331 338 363
rect 38 96 70 128
rect 106 96 138 128
<< metal1 >>
rect 0 772 576 800
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 576 772
rect 0 712 576 740
rect 49 620 101 712
rect 49 588 59 620
rect 91 588 101 620
rect 49 519 101 588
rect 49 487 59 519
rect 91 487 101 519
rect 49 485 101 487
rect 151 620 203 622
rect 151 588 161 620
rect 193 588 203 620
rect 151 519 203 588
rect 151 487 161 519
rect 193 487 203 519
rect 253 620 305 712
rect 253 588 263 620
rect 295 588 305 620
rect 253 531 305 588
rect 253 499 263 531
rect 295 499 305 531
rect 253 497 305 499
rect 355 620 421 622
rect 355 588 365 620
rect 397 588 421 620
rect 355 543 421 588
rect 355 511 365 543
rect 397 511 421 543
rect 151 448 203 487
rect 355 463 421 511
rect 457 620 509 712
rect 457 588 467 620
rect 499 588 509 620
rect 457 531 509 588
rect 457 499 467 531
rect 499 499 509 531
rect 457 497 509 499
rect 49 410 312 448
rect 355 431 365 463
rect 397 431 421 463
rect 355 428 421 431
rect 49 268 101 410
rect 280 380 312 410
rect 156 363 234 374
rect 156 331 192 363
rect 224 331 234 363
rect 156 287 234 331
rect 280 363 348 380
rect 280 331 306 363
rect 338 331 348 363
rect 280 314 348 331
rect 384 272 421 428
rect 49 236 59 268
rect 91 236 101 268
rect 49 228 101 236
rect 355 269 421 272
rect 355 237 365 269
rect 397 237 421 269
rect 253 229 305 231
rect 253 197 263 229
rect 295 197 305 229
rect 21 128 156 192
rect 21 96 38 128
rect 70 96 106 128
rect 138 96 156 128
rect 21 81 156 96
rect 253 44 305 197
rect 355 191 421 237
rect 355 159 365 191
rect 397 159 421 191
rect 355 156 421 159
rect 457 229 509 231
rect 457 197 467 229
rect 499 197 509 229
rect 457 44 509 197
rect 0 16 576 44
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 576 16
rect 0 -44 576 -16
<< labels >>
flabel metal1 s 355 428 421 622 0 FreeSans 400 0 0 0 X
port 2 nsew
flabel metal1 s 0 -44 576 44 0 FreeSans 400 0 0 0 VSS
port 3 nsew
flabel metal1 s 0 712 576 800 0 FreeSans 400 0 0 0 VDD
port 4 nsew
flabel metal1 s 156 287 234 374 0 FreeSans 400 0 0 0 B
port 5 nsew
flabel metal1 s 21 81 156 192 0 FreeSans 400 0 0 0 A
port 6 nsew
<< properties >>
string FIXED_BBOX 0 0 576 756
string GDS_END 234828
string GDS_FILE ../gds/controller.gds
string GDS_START 230118
<< end >>
