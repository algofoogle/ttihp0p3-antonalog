magic
tech ihp-sg13g2
timestamp 1747537721
<< nwell >>
rect -24 175 312 417
<< pwell >>
rect 9 28 273 157
rect -13 -28 301 28
<< nmos >>
rect 56 80 69 144
rect 107 80 120 144
rect 158 70 171 144
rect 209 70 222 144
<< pmos >>
rect 56 234 69 318
rect 107 234 120 318
rect 158 206 171 318
rect 209 206 222 318
<< ndiff >>
rect 22 134 56 144
rect 22 118 29 134
rect 45 118 56 134
rect 22 80 56 118
rect 69 80 107 144
rect 120 114 158 144
rect 120 98 131 114
rect 147 98 158 114
rect 120 80 158 98
rect 135 70 158 80
rect 171 134 209 144
rect 171 118 182 134
rect 198 118 209 134
rect 171 95 209 118
rect 171 79 182 95
rect 198 79 209 95
rect 171 70 209 79
rect 222 114 260 144
rect 222 98 233 114
rect 249 98 260 114
rect 222 70 260 98
<< pdiff >>
rect 22 310 56 318
rect 22 294 29 310
rect 45 294 56 310
rect 22 259 56 294
rect 22 243 29 259
rect 45 243 56 259
rect 22 234 56 243
rect 69 310 107 318
rect 69 294 80 310
rect 96 294 107 310
rect 69 259 107 294
rect 69 243 80 259
rect 96 243 107 259
rect 69 234 107 243
rect 120 310 158 318
rect 120 294 131 310
rect 147 294 158 310
rect 120 265 158 294
rect 120 249 131 265
rect 147 249 158 265
rect 120 234 158 249
rect 135 206 158 234
rect 171 310 209 318
rect 171 294 182 310
rect 198 294 209 310
rect 171 271 209 294
rect 171 255 182 271
rect 198 255 209 271
rect 171 231 209 255
rect 171 215 182 231
rect 198 215 209 231
rect 171 206 209 215
rect 222 310 260 318
rect 222 294 233 310
rect 249 294 260 310
rect 222 265 260 294
rect 222 249 233 265
rect 249 249 260 265
rect 222 206 260 249
<< ndiffc >>
rect 29 118 45 134
rect 131 98 147 114
rect 182 118 198 134
rect 182 79 198 95
rect 233 98 249 114
<< pdiffc >>
rect 29 294 45 310
rect 29 243 45 259
rect 80 294 96 310
rect 80 243 96 259
rect 131 294 147 310
rect 131 249 147 265
rect 182 294 198 310
rect 182 255 198 271
rect 182 215 198 231
rect 233 294 249 310
rect 233 249 249 265
<< psubdiff >>
rect 0 8 288 15
rect 0 -8 16 8
rect 32 -8 64 8
rect 80 -8 112 8
rect 128 -8 160 8
rect 176 -8 208 8
rect 224 -8 256 8
rect 272 -8 288 8
rect 0 -15 288 -8
<< nsubdiff >>
rect 0 386 288 393
rect 0 370 16 386
rect 32 370 64 386
rect 80 370 112 386
rect 128 370 160 386
rect 176 370 208 386
rect 224 370 256 386
rect 272 370 288 386
rect 0 363 288 370
<< psubdiffcont >>
rect 16 -8 32 8
rect 64 -8 80 8
rect 112 -8 128 8
rect 160 -8 176 8
rect 208 -8 224 8
rect 256 -8 272 8
<< nsubdiffcont >>
rect 16 370 32 386
rect 64 370 80 386
rect 112 370 128 386
rect 160 370 176 386
rect 208 370 224 386
rect 256 370 272 386
<< poly >>
rect 56 318 69 336
rect 107 318 120 336
rect 158 318 171 336
rect 209 318 222 336
rect 56 144 69 234
rect 107 190 120 234
rect 158 190 171 206
rect 209 190 222 206
rect 87 181 120 190
rect 87 165 96 181
rect 112 165 120 181
rect 87 157 120 165
rect 138 181 222 190
rect 138 165 153 181
rect 169 165 222 181
rect 138 157 222 165
rect 107 144 120 157
rect 158 144 171 157
rect 209 144 222 157
rect 56 73 69 80
rect 10 64 77 73
rect 10 48 19 64
rect 35 48 53 64
rect 69 48 77 64
rect 107 62 120 80
rect 158 52 171 70
rect 209 52 222 70
rect 10 41 77 48
<< polycont >>
rect 96 165 112 181
rect 153 165 169 181
rect 19 48 35 64
rect 53 48 69 64
<< metal1 >>
rect 0 386 288 400
rect 0 370 16 386
rect 32 370 64 386
rect 80 370 112 386
rect 128 370 160 386
rect 176 370 208 386
rect 224 370 256 386
rect 272 370 288 386
rect 0 356 288 370
rect 24 310 50 356
rect 24 294 29 310
rect 45 294 50 310
rect 24 259 50 294
rect 24 243 29 259
rect 45 243 50 259
rect 24 242 50 243
rect 75 310 101 311
rect 75 294 80 310
rect 96 294 101 310
rect 75 259 101 294
rect 75 243 80 259
rect 96 243 101 259
rect 126 310 152 356
rect 126 294 131 310
rect 147 294 152 310
rect 126 265 152 294
rect 126 249 131 265
rect 147 249 152 265
rect 126 248 152 249
rect 177 310 210 311
rect 177 294 182 310
rect 198 294 210 310
rect 177 271 210 294
rect 177 255 182 271
rect 198 255 210 271
rect 75 224 101 243
rect 177 231 210 255
rect 228 310 254 356
rect 228 294 233 310
rect 249 294 254 310
rect 228 265 254 294
rect 228 249 233 265
rect 249 249 254 265
rect 228 248 254 249
rect 24 205 156 224
rect 177 215 182 231
rect 198 215 210 231
rect 177 214 210 215
rect 24 134 50 205
rect 140 190 156 205
rect 78 181 117 187
rect 78 165 96 181
rect 112 165 117 181
rect 78 143 117 165
rect 140 181 174 190
rect 140 165 153 181
rect 169 165 174 181
rect 140 157 174 165
rect 192 136 210 214
rect 24 118 29 134
rect 45 118 50 134
rect 24 114 50 118
rect 177 134 210 136
rect 177 118 182 134
rect 198 118 210 134
rect 126 114 152 115
rect 126 98 131 114
rect 147 98 152 114
rect 10 64 78 96
rect 10 48 19 64
rect 35 48 53 64
rect 69 48 78 64
rect 10 40 78 48
rect 126 22 152 98
rect 177 95 210 118
rect 177 79 182 95
rect 198 79 210 95
rect 177 78 210 79
rect 228 114 254 115
rect 228 98 233 114
rect 249 98 254 114
rect 228 22 254 98
rect 0 8 288 22
rect 0 -8 16 8
rect 32 -8 64 8
rect 80 -8 112 8
rect 128 -8 160 8
rect 176 -8 208 8
rect 224 -8 256 8
rect 272 -8 288 8
rect 0 -22 288 -8
<< labels >>
flabel metal1 s 177 214 210 311 0 FreeSans 200 0 0 0 X
port 2 nsew
flabel metal1 s 0 -22 288 22 0 FreeSans 200 0 0 0 VSS
port 3 nsew
flabel metal1 s 0 356 288 400 0 FreeSans 200 0 0 0 VDD
port 4 nsew
flabel metal1 s 78 143 117 187 0 FreeSans 200 0 0 0 B
port 5 nsew
flabel metal1 s 10 40 78 96 0 FreeSans 200 0 0 0 A
port 6 nsew
<< properties >>
string FIXED_BBOX 0 0 288 378
string GDS_END 236660
string GDS_FILE ../gds/controller.gds
string GDS_START 231950
<< end >>
