magic
tech ihp-sg13g2
timestamp 1747537721
<< nwell >>
rect -24 175 1032 417
rect 74 161 456 175
<< pwell >>
rect 638 151 786 157
rect 638 136 999 151
rect 22 28 999 136
rect -13 -28 1021 28
<< nmos >>
rect 69 59 82 123
rect 141 59 154 123
rect 178 59 191 123
rect 237 59 250 123
rect 322 59 335 123
rect 392 59 405 123
rect 430 59 443 123
rect 498 59 511 123
rect 535 59 548 123
rect 675 80 688 144
rect 726 80 739 144
rect 882 74 895 138
rect 939 64 952 138
<< pmos >>
rect 79 206 92 306
rect 134 192 147 292
rect 230 192 243 292
rect 281 192 294 292
rect 326 192 339 292
rect 389 192 402 292
rect 440 215 453 315
rect 541 215 554 315
rect 581 215 594 315
rect 683 218 696 318
rect 741 218 754 318
rect 863 215 876 315
rect 941 206 954 318
<< ndiff >>
rect 35 116 69 123
rect 35 100 42 116
rect 58 100 69 116
rect 35 82 69 100
rect 35 66 42 82
rect 58 66 69 82
rect 35 59 69 66
rect 82 82 141 123
rect 82 66 103 82
rect 119 66 141 82
rect 82 59 141 66
rect 154 59 178 123
rect 191 111 237 123
rect 191 95 210 111
rect 226 95 237 111
rect 191 59 237 95
rect 250 59 322 123
rect 335 82 392 123
rect 335 66 356 82
rect 372 66 392 82
rect 335 59 392 66
rect 405 59 430 123
rect 443 82 498 123
rect 443 66 462 82
rect 478 66 498 82
rect 443 59 498 66
rect 511 59 535 123
rect 548 91 582 123
rect 651 114 675 144
rect 548 75 559 91
rect 575 75 582 91
rect 548 59 582 75
rect 609 107 675 114
rect 609 91 616 107
rect 632 91 675 107
rect 609 80 675 91
rect 688 137 726 144
rect 688 121 699 137
rect 715 121 726 137
rect 688 80 726 121
rect 739 103 773 144
rect 739 87 750 103
rect 766 87 773 103
rect 739 80 773 87
rect 846 131 882 138
rect 846 115 853 131
rect 869 115 882 131
rect 846 97 882 115
rect 846 81 853 97
rect 869 81 882 97
rect 609 62 668 80
rect 609 46 616 62
rect 632 46 668 62
rect 609 39 668 46
rect 846 74 882 81
rect 895 131 939 138
rect 895 115 908 131
rect 924 115 939 131
rect 895 97 939 115
rect 895 81 908 97
rect 924 81 939 97
rect 895 74 939 81
rect 912 64 939 74
rect 952 131 986 138
rect 952 115 963 131
rect 979 115 986 131
rect 952 88 986 115
rect 952 72 963 88
rect 979 72 986 88
rect 952 64 986 72
<< pdiff >>
rect 45 297 79 306
rect 45 281 52 297
rect 68 281 79 297
rect 45 263 79 281
rect 45 247 52 263
rect 68 247 79 263
rect 45 229 79 247
rect 45 213 52 229
rect 68 213 79 229
rect 45 206 79 213
rect 92 297 127 306
rect 92 281 103 297
rect 119 292 127 297
rect 350 314 380 321
rect 350 298 357 314
rect 373 298 380 314
rect 350 292 380 298
rect 412 292 440 315
rect 119 281 134 292
rect 92 263 134 281
rect 92 247 103 263
rect 119 247 134 263
rect 92 229 134 247
rect 92 213 103 229
rect 119 213 134 229
rect 92 206 134 213
rect 108 192 134 206
rect 147 192 230 292
rect 243 284 281 292
rect 243 268 254 284
rect 270 268 281 284
rect 243 250 281 268
rect 243 234 254 250
rect 270 234 281 250
rect 243 216 281 234
rect 243 200 254 216
rect 270 200 281 216
rect 243 192 281 200
rect 294 192 326 292
rect 339 192 389 292
rect 402 215 440 292
rect 453 287 541 315
rect 453 271 464 287
rect 480 271 514 287
rect 530 271 541 287
rect 453 239 541 271
rect 453 223 464 239
rect 480 223 514 239
rect 530 223 541 239
rect 453 215 541 223
rect 554 215 581 315
rect 594 307 628 315
rect 594 291 605 307
rect 621 291 628 307
rect 594 215 628 291
rect 649 311 683 318
rect 649 295 656 311
rect 672 295 683 311
rect 649 276 683 295
rect 649 260 656 276
rect 672 260 683 276
rect 649 241 683 260
rect 649 225 656 241
rect 672 225 683 241
rect 649 218 683 225
rect 696 310 741 318
rect 696 294 709 310
rect 725 294 741 310
rect 696 276 741 294
rect 696 260 709 276
rect 725 260 741 276
rect 696 241 741 260
rect 696 225 709 241
rect 725 225 741 241
rect 696 218 741 225
rect 754 287 788 318
rect 909 315 941 318
rect 754 271 765 287
rect 781 271 788 287
rect 754 241 788 271
rect 754 225 765 241
rect 781 225 788 241
rect 754 218 788 225
rect 829 287 863 315
rect 829 271 836 287
rect 852 271 863 287
rect 829 241 863 271
rect 829 225 836 241
rect 852 225 863 241
rect 402 192 430 215
rect 829 215 863 225
rect 876 309 941 315
rect 876 293 914 309
rect 930 293 941 309
rect 876 275 941 293
rect 876 259 914 275
rect 930 259 941 275
rect 876 215 941 259
rect 916 206 941 215
rect 954 302 988 318
rect 954 286 965 302
rect 981 286 988 302
rect 954 206 988 286
<< ndiffc >>
rect 42 100 58 116
rect 42 66 58 82
rect 103 66 119 82
rect 210 95 226 111
rect 356 66 372 82
rect 462 66 478 82
rect 559 75 575 91
rect 616 91 632 107
rect 699 121 715 137
rect 750 87 766 103
rect 853 115 869 131
rect 853 81 869 97
rect 616 46 632 62
rect 908 115 924 131
rect 908 81 924 97
rect 963 115 979 131
rect 963 72 979 88
<< pdiffc >>
rect 52 281 68 297
rect 52 247 68 263
rect 52 213 68 229
rect 103 281 119 297
rect 357 298 373 314
rect 103 247 119 263
rect 103 213 119 229
rect 254 268 270 284
rect 254 234 270 250
rect 254 200 270 216
rect 464 271 480 287
rect 514 271 530 287
rect 464 223 480 239
rect 514 223 530 239
rect 605 291 621 307
rect 656 295 672 311
rect 656 260 672 276
rect 656 225 672 241
rect 709 294 725 310
rect 709 260 725 276
rect 709 225 725 241
rect 765 271 781 287
rect 765 225 781 241
rect 836 271 852 287
rect 836 225 852 241
rect 914 293 930 309
rect 914 259 930 275
rect 965 286 981 302
<< psubdiff >>
rect 0 8 1008 15
rect 0 -8 16 8
rect 32 -8 64 8
rect 80 -8 112 8
rect 128 -8 160 8
rect 176 -8 208 8
rect 224 -8 256 8
rect 272 -8 304 8
rect 320 -8 352 8
rect 368 -8 400 8
rect 416 -8 448 8
rect 464 -8 496 8
rect 512 -8 544 8
rect 560 -8 592 8
rect 608 -8 640 8
rect 656 -8 688 8
rect 704 -8 736 8
rect 752 -8 784 8
rect 800 -8 832 8
rect 848 -8 880 8
rect 896 -8 928 8
rect 944 -8 976 8
rect 992 -8 1008 8
rect 0 -15 1008 -8
<< nsubdiff >>
rect 0 386 1008 393
rect 0 370 16 386
rect 32 370 64 386
rect 80 370 112 386
rect 128 370 160 386
rect 176 370 208 386
rect 224 370 256 386
rect 272 370 304 386
rect 320 370 352 386
rect 368 370 400 386
rect 416 370 448 386
rect 464 370 496 386
rect 512 370 544 386
rect 560 370 592 386
rect 608 370 640 386
rect 656 370 688 386
rect 704 370 736 386
rect 752 370 784 386
rect 800 370 832 386
rect 848 370 880 386
rect 896 370 928 386
rect 944 370 976 386
rect 992 370 1008 386
rect 0 363 1008 370
<< psubdiffcont >>
rect 16 -8 32 8
rect 64 -8 80 8
rect 112 -8 128 8
rect 160 -8 176 8
rect 208 -8 224 8
rect 256 -8 272 8
rect 304 -8 320 8
rect 352 -8 368 8
rect 400 -8 416 8
rect 448 -8 464 8
rect 496 -8 512 8
rect 544 -8 560 8
rect 592 -8 608 8
rect 640 -8 656 8
rect 688 -8 704 8
rect 736 -8 752 8
rect 784 -8 800 8
rect 832 -8 848 8
rect 880 -8 896 8
rect 928 -8 944 8
rect 976 -8 992 8
<< nsubdiffcont >>
rect 16 370 32 386
rect 64 370 80 386
rect 112 370 128 386
rect 160 370 176 386
rect 208 370 224 386
rect 256 370 272 386
rect 304 370 320 386
rect 352 370 368 386
rect 400 370 416 386
rect 448 370 464 386
rect 496 370 512 386
rect 544 370 560 386
rect 592 370 608 386
rect 640 370 656 386
rect 688 370 704 386
rect 736 370 752 386
rect 784 370 800 386
rect 832 370 848 386
rect 880 370 896 386
rect 928 370 944 386
rect 976 370 992 386
<< poly >>
rect 79 328 453 342
rect 79 306 92 328
rect 134 292 147 310
rect 230 292 243 328
rect 440 315 453 328
rect 541 315 554 333
rect 581 315 594 333
rect 683 318 696 336
rect 741 318 754 336
rect 281 292 294 310
rect 326 292 339 310
rect 389 292 402 310
rect 79 176 92 206
rect 863 315 876 333
rect 941 318 954 336
rect 440 206 453 215
rect 134 176 147 192
rect 230 185 243 192
rect 68 168 102 176
rect 68 152 78 168
rect 94 152 102 168
rect 68 143 102 152
rect 124 168 157 176
rect 124 152 132 168
rect 148 152 157 168
rect 124 143 157 152
rect 175 166 208 175
rect 175 150 183 166
rect 199 150 208 166
rect 69 123 82 143
rect 141 123 154 143
rect 175 142 208 150
rect 178 123 191 142
rect 230 130 250 185
rect 281 167 294 192
rect 326 176 339 192
rect 389 176 402 192
rect 440 191 502 206
rect 541 199 554 215
rect 322 168 355 176
rect 268 158 301 167
rect 268 142 276 158
rect 292 142 301 158
rect 268 134 301 142
rect 322 152 330 168
rect 346 152 355 168
rect 322 143 355 152
rect 376 168 409 176
rect 376 152 384 168
rect 400 152 409 168
rect 376 143 409 152
rect 430 158 463 167
rect 237 123 250 130
rect 322 123 335 143
rect 392 123 405 143
rect 430 142 438 158
rect 454 142 463 158
rect 430 134 463 142
rect 487 145 502 191
rect 523 191 554 199
rect 523 175 531 191
rect 547 175 554 191
rect 523 166 554 175
rect 581 199 594 215
rect 581 191 640 199
rect 581 175 615 191
rect 631 175 640 191
rect 581 145 640 175
rect 683 171 696 218
rect 741 181 754 218
rect 785 191 818 199
rect 785 181 793 191
rect 430 123 443 134
rect 487 130 511 145
rect 498 123 511 130
rect 535 130 640 145
rect 675 156 696 171
rect 726 175 793 181
rect 809 175 818 191
rect 726 166 818 175
rect 863 190 876 215
rect 941 190 954 206
rect 863 181 895 190
rect 675 144 688 156
rect 726 144 739 166
rect 863 165 871 181
rect 887 165 895 181
rect 863 157 895 165
rect 916 181 954 190
rect 916 165 925 181
rect 941 165 954 181
rect 916 157 954 165
rect 535 123 548 130
rect 882 138 895 157
rect 939 138 952 157
rect 69 41 82 59
rect 141 41 154 59
rect 178 41 191 59
rect 237 41 250 59
rect 322 41 335 59
rect 392 41 405 59
rect 430 41 443 59
rect 498 41 511 59
rect 535 41 548 59
rect 675 44 688 80
rect 726 62 739 80
rect 882 44 895 74
rect 939 46 952 64
rect 675 31 895 44
<< polycont >>
rect 78 152 94 168
rect 132 152 148 168
rect 183 150 199 166
rect 276 142 292 158
rect 330 152 346 168
rect 384 152 400 168
rect 438 142 454 158
rect 531 175 547 191
rect 615 175 631 191
rect 793 175 809 191
rect 871 165 887 181
rect 925 165 941 181
<< metal1 >>
rect 0 386 1008 400
rect 0 370 16 386
rect 32 370 64 386
rect 80 370 112 386
rect 128 370 160 386
rect 176 370 208 386
rect 224 370 256 386
rect 272 370 304 386
rect 320 370 352 386
rect 368 370 400 386
rect 416 370 448 386
rect 464 370 496 386
rect 512 370 544 386
rect 560 370 592 386
rect 608 370 640 386
rect 656 370 688 386
rect 704 370 736 386
rect 752 370 784 386
rect 800 370 832 386
rect 848 370 880 386
rect 896 370 928 386
rect 944 370 976 386
rect 992 370 1008 386
rect 0 356 1008 370
rect 33 297 74 298
rect 33 281 52 297
rect 68 281 74 297
rect 33 263 74 281
rect 33 247 52 263
rect 68 247 74 263
rect 33 229 74 247
rect 33 213 52 229
rect 68 213 74 229
rect 33 212 74 213
rect 98 297 124 356
rect 352 314 378 356
rect 352 298 357 314
rect 373 298 378 314
rect 352 297 378 298
rect 401 312 577 329
rect 98 281 103 297
rect 119 281 124 297
rect 98 263 124 281
rect 98 247 103 263
rect 119 247 124 263
rect 98 229 124 247
rect 98 213 103 229
rect 119 213 124 229
rect 98 212 124 213
rect 226 284 277 290
rect 226 268 254 284
rect 270 272 277 284
rect 401 272 424 312
rect 270 268 424 272
rect 226 255 424 268
rect 452 287 538 294
rect 452 271 464 287
rect 480 271 514 287
rect 530 271 538 287
rect 226 250 277 255
rect 226 234 254 250
rect 270 234 277 250
rect 452 239 538 271
rect 557 272 577 312
rect 595 307 628 356
rect 595 291 605 307
rect 621 291 628 307
rect 595 290 628 291
rect 651 311 678 320
rect 651 295 656 311
rect 672 295 678 311
rect 651 276 678 295
rect 651 272 656 276
rect 557 260 656 272
rect 672 260 678 276
rect 557 255 678 260
rect 226 216 277 234
rect 33 120 50 212
rect 226 200 254 216
rect 270 200 277 216
rect 226 195 277 200
rect 70 168 104 192
rect 70 152 78 168
rect 94 152 104 168
rect 70 143 104 152
rect 124 168 157 192
rect 124 152 132 168
rect 148 152 157 168
rect 124 143 157 152
rect 175 166 208 175
rect 175 150 183 166
rect 199 150 208 166
rect 175 142 208 150
rect 175 120 191 142
rect 226 120 242 195
rect 322 168 354 237
rect 33 116 191 120
rect 33 100 42 116
rect 58 102 191 116
rect 58 100 64 102
rect 33 82 64 100
rect 33 66 42 82
rect 58 66 64 82
rect 33 59 64 66
rect 98 82 124 84
rect 98 66 103 82
rect 119 66 124 82
rect 98 22 124 66
rect 175 64 191 102
rect 209 111 242 120
rect 209 95 210 111
rect 226 95 242 111
rect 209 87 242 95
rect 268 158 301 167
rect 268 142 276 158
rect 292 142 301 158
rect 322 152 330 168
rect 346 152 354 168
rect 322 143 354 152
rect 372 168 409 237
rect 452 223 464 239
rect 480 223 514 239
rect 530 237 538 239
rect 651 241 678 255
rect 530 223 588 237
rect 452 220 588 223
rect 372 152 384 168
rect 400 152 409 168
rect 480 191 553 197
rect 480 175 531 191
rect 547 175 553 191
rect 372 143 409 152
rect 430 158 461 167
rect 268 121 301 142
rect 430 142 438 158
rect 454 142 461 158
rect 430 121 461 142
rect 480 166 553 175
rect 480 121 497 166
rect 571 138 588 220
rect 651 225 656 241
rect 672 225 678 241
rect 651 217 678 225
rect 607 191 640 200
rect 607 175 615 191
rect 631 175 640 191
rect 607 156 640 175
rect 268 105 497 121
rect 515 121 637 138
rect 268 64 285 105
rect 515 87 532 121
rect 611 107 637 121
rect 175 47 285 64
rect 349 82 377 83
rect 349 66 356 82
rect 372 66 377 82
rect 349 22 377 66
rect 455 82 532 87
rect 455 66 462 82
rect 478 66 532 82
rect 455 59 532 66
rect 554 91 580 101
rect 554 75 559 91
rect 575 75 580 91
rect 554 22 580 75
rect 611 91 616 107
rect 632 91 637 107
rect 611 62 637 91
rect 658 98 678 217
rect 701 312 891 329
rect 701 310 730 312
rect 701 294 709 310
rect 725 294 730 310
rect 701 276 730 294
rect 701 260 709 276
rect 725 260 730 276
rect 701 241 730 260
rect 701 225 709 241
rect 725 225 730 241
rect 701 150 730 225
rect 696 137 730 150
rect 696 121 699 137
rect 715 133 730 137
rect 751 287 786 292
rect 751 271 765 287
rect 781 271 786 287
rect 751 241 786 271
rect 751 225 765 241
rect 781 225 786 241
rect 751 222 786 225
rect 819 287 857 292
rect 819 271 836 287
rect 852 271 857 287
rect 819 241 857 271
rect 819 225 836 241
rect 852 225 857 241
rect 751 148 767 222
rect 819 217 857 225
rect 875 240 891 312
rect 909 309 935 356
rect 909 293 914 309
rect 930 293 935 309
rect 909 275 935 293
rect 964 302 990 307
rect 964 286 965 302
rect 981 286 990 302
rect 964 278 990 286
rect 909 259 914 275
rect 930 259 935 275
rect 909 258 935 259
rect 875 223 946 240
rect 819 199 835 217
rect 785 191 835 199
rect 785 175 793 191
rect 809 175 835 191
rect 785 166 835 175
rect 715 121 721 133
rect 751 132 801 148
rect 696 116 721 121
rect 745 103 767 108
rect 745 98 750 103
rect 658 87 750 98
rect 766 87 767 103
rect 658 82 767 87
rect 611 46 616 62
rect 632 60 637 62
rect 785 60 801 132
rect 819 138 835 166
rect 853 181 895 198
rect 853 165 871 181
rect 887 165 895 181
rect 853 156 895 165
rect 919 181 946 223
rect 919 165 925 181
rect 941 165 946 181
rect 919 157 946 165
rect 819 131 874 138
rect 966 136 990 278
rect 819 115 853 131
rect 869 115 874 131
rect 819 97 874 115
rect 819 81 853 97
rect 869 81 874 97
rect 819 75 874 81
rect 903 131 929 132
rect 903 115 908 131
rect 924 115 929 131
rect 903 97 929 115
rect 903 81 908 97
rect 924 81 929 97
rect 632 46 801 60
rect 611 44 801 46
rect 903 22 929 81
rect 947 131 990 136
rect 947 115 963 131
rect 979 115 990 131
rect 947 88 990 115
rect 947 72 963 88
rect 979 72 990 88
rect 947 62 990 72
rect 0 8 1008 22
rect 0 -8 16 8
rect 32 -8 64 8
rect 80 -8 112 8
rect 128 -8 160 8
rect 176 -8 208 8
rect 224 -8 256 8
rect 272 -8 304 8
rect 320 -8 352 8
rect 368 -8 400 8
rect 416 -8 448 8
rect 464 -8 496 8
rect 512 -8 544 8
rect 560 -8 592 8
rect 608 -8 640 8
rect 656 -8 688 8
rect 704 -8 736 8
rect 752 -8 784 8
rect 800 -8 832 8
rect 848 -8 880 8
rect 896 -8 928 8
rect 944 -8 976 8
rect 992 -8 1008 8
rect 0 -22 1008 -8
<< labels >>
flabel metal1 s 947 62 990 136 0 FreeSans 200 0 0 0 X
port 2 nsew
flabel metal1 s 322 143 354 237 0 FreeSans 200 0 0 0 A1
port 3 nsew
flabel metal1 s 372 143 409 237 0 FreeSans 200 0 0 0 A2
port 4 nsew
flabel metal1 s 70 143 104 192 0 FreeSans 200 0 0 0 S0
port 5 nsew
flabel metal1 s 0 356 1008 400 0 FreeSans 200 0 0 0 VDD
port 6 nsew
flabel metal1 s 0 -22 1008 22 0 FreeSans 200 0 0 0 VSS
port 7 nsew
flabel metal1 s 853 156 895 198 0 FreeSans 200 0 0 0 S1
port 8 nsew
flabel metal1 s 124 143 157 192 0 FreeSans 200 0 0 0 A0
port 9 nsew
flabel metal1 s 607 156 640 200 0 FreeSans 200 0 0 0 A3
port 10 nsew
<< properties >>
string FIXED_BBOX 0 0 1008 378
string GDS_END 171634
string GDS_FILE ../gds/controller.gds
string GDS_START 159636
<< end >>
