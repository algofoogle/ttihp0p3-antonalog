magic
tech ihp-sg13g2
magscale 1 2
timestamp 1746839692
<< pwell >>
rect 830 1624 1338 1740
rect 834 446 1046 630
rect 538 330 1046 446
rect 834 322 1046 330
rect 1126 180 1342 446
<< metal1 >>
rect -94 444 98 2036
rect 238 1630 746 1752
rect 830 1624 1338 1740
rect 1420 1738 1928 1744
rect 1420 1618 1930 1738
rect 2016 1642 2224 1892
rect 1730 1478 1930 1618
rect 2314 1478 2514 1734
rect 2608 1626 3120 1740
rect 3186 1736 3714 1742
rect 3186 1614 3720 1736
rect 3790 1644 4004 1894
rect 1730 1278 2514 1478
rect 3510 1482 3720 1614
rect 4091 1482 4301 1731
rect 4376 1620 4896 1744
rect 4976 1728 5484 1736
rect 4976 1624 5490 1728
rect 5572 1642 5786 1900
rect 6772 1732 7222 1900
rect 3510 1272 4301 1482
rect 5282 1470 5490 1624
rect 5862 1470 6070 1730
rect 6154 1622 6670 1732
rect 6750 1620 7260 1732
rect 7346 1620 7556 1900
rect 5282 1262 6070 1470
rect 834 550 1636 762
rect 834 446 1046 550
rect -100 24 460 444
rect 538 330 1046 446
rect 834 322 1046 330
rect 1126 180 1342 446
rect 1424 340 1636 550
rect 2612 544 3414 760
rect 2612 460 2828 544
rect 1716 324 2232 426
rect 2308 324 2828 460
rect 2308 316 2822 324
rect 2902 174 3114 454
rect 3198 330 3414 544
rect 4394 548 5187 762
rect 3482 336 4010 464
rect 4394 458 4608 548
rect 4080 340 4608 458
rect 4080 334 4600 340
rect 4670 166 4894 460
rect 4973 345 5187 548
rect 6170 548 6965 762
rect 5270 340 5778 452
rect 6170 444 6384 548
rect 5858 340 6384 444
rect 5858 334 6374 340
rect 6446 170 6670 442
rect 6751 341 6965 548
rect 7044 332 7554 444
use resistors  resistors_0
timestamp 1746839677
transform 1 0 2660 0 1 1006
box -2802 -1024 5262 1056
<< labels >>
flabel metal1 250 160 424 296 0 FreeSans 320 0 0 0 GND
port 0 nsew
flabel metal1 1166 220 1302 300 0 FreeSans 320 0 0 0 IN[0]
port 1 nsew
flabel metal1 2058 1776 2186 1868 0 FreeSans 320 0 0 0 IN[1]
port 2 nsew
flabel metal1 2950 218 3068 302 0 FreeSans 320 0 0 0 IN[2]
port 3 nsew
flabel metal1 3834 1780 3964 1860 0 FreeSans 320 0 0 0 IN[3]
port 4 nsew
flabel metal1 4722 218 4850 306 0 FreeSans 320 0 0 0 IN[4]
port 5 nsew
flabel metal1 5612 1764 5744 1860 0 FreeSans 320 0 0 0 IN[5]
port 6 nsew
flabel metal1 6484 212 6632 302 0 FreeSans 320 0 0 0 IN[6]
port 7 nsew
flabel metal1 7386 1768 7520 1858 0 FreeSans 320 0 0 0 IN[7]
port 8 nsew
flabel metal1 6856 1772 7158 1864 0 FreeSans 320 0 0 0 OUT
port 9 nsew
<< end >>
