magic
tech ihp-sg13g2
timestamp 1747537721
<< nwell >>
rect -27 175 360 417
<< pwell >>
rect 12 28 326 157
rect -13 -28 349 28
<< nmos >>
rect 59 80 72 144
rect 113 72 126 144
rect 164 72 177 144
rect 215 72 228 144
rect 266 72 279 144
<< pmos >>
rect 59 206 72 306
rect 113 206 126 318
rect 164 206 177 318
rect 215 206 228 318
rect 266 206 279 318
<< ndiff >>
rect 25 137 59 144
rect 25 121 32 137
rect 48 121 59 137
rect 25 80 59 121
rect 72 137 113 144
rect 72 121 86 137
rect 102 121 113 137
rect 72 95 113 121
rect 72 80 86 95
rect 79 79 86 80
rect 102 79 113 95
rect 79 72 113 79
rect 126 131 164 144
rect 126 115 137 131
rect 153 115 164 131
rect 126 95 164 115
rect 126 79 137 95
rect 153 79 164 95
rect 126 72 164 79
rect 177 95 215 144
rect 177 79 188 95
rect 204 79 215 95
rect 177 72 215 79
rect 228 131 266 144
rect 228 115 239 131
rect 255 115 266 131
rect 228 95 266 115
rect 228 79 239 95
rect 255 79 266 95
rect 228 72 266 79
rect 279 131 313 144
rect 279 115 290 131
rect 306 115 313 131
rect 279 95 313 115
rect 279 79 290 95
rect 306 79 313 95
rect 279 72 313 79
<< pdiff >>
rect 79 311 113 318
rect 79 306 86 311
rect 25 299 59 306
rect 25 283 32 299
rect 48 283 59 299
rect 25 264 59 283
rect 25 248 32 264
rect 48 248 59 264
rect 25 229 59 248
rect 25 213 32 229
rect 48 213 59 229
rect 25 206 59 213
rect 72 295 86 306
rect 102 295 113 311
rect 72 271 113 295
rect 72 255 86 271
rect 102 255 113 271
rect 72 229 113 255
rect 72 213 86 229
rect 102 213 113 229
rect 72 206 113 213
rect 126 311 164 318
rect 126 295 137 311
rect 153 295 164 311
rect 126 271 164 295
rect 126 255 137 271
rect 153 255 164 271
rect 126 206 164 255
rect 177 263 215 318
rect 177 247 188 263
rect 204 247 215 263
rect 177 229 215 247
rect 177 213 188 229
rect 204 213 215 229
rect 177 206 215 213
rect 228 311 266 318
rect 228 295 239 311
rect 255 295 266 311
rect 228 271 266 295
rect 228 255 239 271
rect 255 255 266 271
rect 228 229 266 255
rect 228 213 239 229
rect 255 213 266 229
rect 228 206 266 213
rect 279 311 313 318
rect 279 295 290 311
rect 306 295 313 311
rect 279 271 313 295
rect 279 255 290 271
rect 306 255 313 271
rect 279 229 313 255
rect 279 213 290 229
rect 306 213 313 229
rect 279 206 313 213
<< ndiffc >>
rect 32 121 48 137
rect 86 121 102 137
rect 86 79 102 95
rect 137 115 153 131
rect 137 79 153 95
rect 188 79 204 95
rect 239 115 255 131
rect 239 79 255 95
rect 290 115 306 131
rect 290 79 306 95
<< pdiffc >>
rect 32 283 48 299
rect 32 248 48 264
rect 32 213 48 229
rect 86 295 102 311
rect 86 255 102 271
rect 86 213 102 229
rect 137 295 153 311
rect 137 255 153 271
rect 188 247 204 263
rect 188 213 204 229
rect 239 295 255 311
rect 239 255 255 271
rect 239 213 255 229
rect 290 295 306 311
rect 290 255 306 271
rect 290 213 306 229
<< psubdiff >>
rect 0 8 336 15
rect 0 -8 16 8
rect 32 -8 64 8
rect 80 -8 112 8
rect 128 -8 160 8
rect 176 -8 208 8
rect 224 -8 256 8
rect 272 -8 304 8
rect 320 -8 336 8
rect 0 -15 336 -8
<< nsubdiff >>
rect 0 386 336 393
rect 0 370 16 386
rect 32 370 64 386
rect 80 370 112 386
rect 128 370 160 386
rect 176 370 208 386
rect 224 370 256 386
rect 272 370 304 386
rect 320 370 336 386
rect 0 363 336 370
<< psubdiffcont >>
rect 16 -8 32 8
rect 64 -8 80 8
rect 112 -8 128 8
rect 160 -8 176 8
rect 208 -8 224 8
rect 256 -8 272 8
rect 304 -8 320 8
<< nsubdiffcont >>
rect 16 370 32 386
rect 64 370 80 386
rect 112 370 128 386
rect 160 370 176 386
rect 208 370 224 386
rect 256 370 272 386
rect 304 370 320 386
<< poly >>
rect 59 306 72 324
rect 113 318 126 336
rect 164 318 177 336
rect 215 318 228 336
rect 266 318 279 336
rect 59 144 72 206
rect 113 193 126 206
rect 90 186 126 193
rect 90 170 97 186
rect 113 170 126 186
rect 90 163 126 170
rect 113 144 126 163
rect 164 189 177 206
rect 215 189 228 206
rect 164 182 248 189
rect 164 166 225 182
rect 241 166 248 182
rect 164 159 248 166
rect 164 144 177 159
rect 215 144 228 159
rect 266 144 279 206
rect 59 70 72 80
rect 35 63 72 70
rect 35 47 42 63
rect 58 47 72 63
rect 35 40 72 47
rect 113 35 126 72
rect 164 54 177 72
rect 215 54 228 72
rect 266 35 279 72
rect 113 22 279 35
<< polycont >>
rect 97 170 113 186
rect 225 166 241 182
rect 42 47 58 63
<< metal1 >>
rect 0 386 336 400
rect 0 370 16 386
rect 32 370 64 386
rect 80 370 112 386
rect 128 370 160 386
rect 176 370 208 386
rect 224 370 256 386
rect 272 370 304 386
rect 320 370 336 386
rect 0 356 336 370
rect 81 311 107 356
rect 27 299 53 304
rect 27 283 32 299
rect 48 283 53 299
rect 27 264 53 283
rect 27 248 32 264
rect 48 248 53 264
rect 27 229 53 248
rect 27 213 32 229
rect 48 213 53 229
rect 27 186 53 213
rect 81 295 86 311
rect 102 295 107 311
rect 81 271 107 295
rect 81 255 86 271
rect 102 255 107 271
rect 81 229 107 255
rect 132 311 260 326
rect 132 295 137 311
rect 153 308 239 311
rect 153 295 158 308
rect 132 271 158 295
rect 234 295 239 308
rect 255 295 260 311
rect 132 255 137 271
rect 153 255 158 271
rect 132 247 158 255
rect 183 263 209 290
rect 183 247 188 263
rect 204 247 209 263
rect 81 213 86 229
rect 102 213 107 229
rect 183 229 209 247
rect 183 220 188 229
rect 81 208 107 213
rect 136 213 188 220
rect 204 213 209 229
rect 136 200 209 213
rect 234 271 260 295
rect 234 255 239 271
rect 255 255 260 271
rect 234 229 260 255
rect 234 213 239 229
rect 255 213 260 229
rect 234 208 260 213
rect 285 311 311 356
rect 285 295 290 311
rect 306 295 311 311
rect 285 271 311 295
rect 285 255 290 271
rect 306 255 311 271
rect 285 229 311 255
rect 285 213 290 229
rect 306 213 311 229
rect 285 208 311 213
rect 27 170 97 186
rect 113 170 118 186
rect 27 137 53 170
rect 27 121 32 137
rect 48 121 53 137
rect 27 116 53 121
rect 81 137 107 142
rect 81 121 86 137
rect 102 121 107 137
rect 136 136 158 200
rect 217 166 225 182
rect 241 166 296 182
rect 217 154 296 166
rect 37 63 63 96
rect 37 47 42 63
rect 58 47 63 63
rect 37 40 63 47
rect 81 95 107 121
rect 81 79 86 95
rect 102 79 107 95
rect 81 22 107 79
rect 132 131 260 136
rect 132 115 137 131
rect 153 116 239 131
rect 153 115 158 116
rect 132 95 158 115
rect 234 115 239 116
rect 255 115 260 131
rect 132 79 137 95
rect 153 79 158 95
rect 132 72 158 79
rect 183 95 209 98
rect 183 79 188 95
rect 204 79 209 95
rect 183 22 209 79
rect 234 95 260 115
rect 234 79 239 95
rect 255 79 260 95
rect 234 72 260 79
rect 285 131 311 136
rect 285 115 290 131
rect 306 115 311 131
rect 285 95 311 115
rect 285 79 290 95
rect 306 79 311 95
rect 285 22 311 79
rect 0 8 336 22
rect 0 -8 16 8
rect 32 -8 64 8
rect 80 -8 112 8
rect 128 -8 160 8
rect 176 -8 208 8
rect 224 -8 256 8
rect 272 -8 304 8
rect 320 -8 336 8
rect 0 -22 336 -8
<< labels >>
flabel metal1 s 217 154 296 182 0 FreeSans 200 0 0 0 A
port 2 nsew
flabel metal1 s 37 40 63 96 0 FreeSans 200 0 0 0 B_N
port 3 nsew
flabel metal1 s 0 356 336 400 0 FreeSans 200 0 0 0 VDD
port 4 nsew
flabel metal1 s 132 116 260 136 0 FreeSans 200 0 0 0 Y
port 5 nsew
flabel metal1 s 0 -22 336 22 0 FreeSans 200 0 0 0 VSS
port 6 nsew
<< properties >>
string FIXED_BBOX 0 0 336 378
string GDS_END 231904
string GDS_FILE ../gds/controller.gds
string GDS_START 226776
<< end >>
