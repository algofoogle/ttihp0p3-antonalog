magic
tech ihp-sg13g2
magscale 1 2
timestamp 1747056097
<< nwell >>
rect -48 350 720 834
<< pwell >>
rect 5 56 669 240
rect -26 -56 698 56
<< nmos >>
rect 99 130 299 214
rect 375 130 575 214
<< pmos >>
rect 101 437 301 637
rect 377 437 577 637
<< ndiff >>
rect 31 188 99 214
rect 31 156 45 188
rect 77 156 99 188
rect 31 130 99 156
rect 299 188 375 214
rect 299 156 321 188
rect 353 156 375 188
rect 299 130 375 156
rect 575 188 643 214
rect 575 156 597 188
rect 629 156 643 188
rect 575 130 643 156
<< pdiff >>
rect 33 623 101 637
rect 33 591 47 623
rect 79 591 101 623
rect 33 552 101 591
rect 33 520 47 552
rect 79 520 101 552
rect 33 484 101 520
rect 33 452 47 484
rect 79 452 101 484
rect 33 437 101 452
rect 301 623 377 637
rect 301 591 323 623
rect 355 591 377 623
rect 301 555 377 591
rect 301 523 323 555
rect 355 523 377 555
rect 301 487 377 523
rect 301 455 323 487
rect 355 455 377 487
rect 301 437 377 455
rect 577 623 645 637
rect 577 591 599 623
rect 631 591 645 623
rect 577 552 645 591
rect 577 520 599 552
rect 631 520 645 552
rect 577 484 645 520
rect 577 452 599 484
rect 631 452 645 484
rect 577 437 645 452
<< ndiffc >>
rect 45 156 77 188
rect 321 156 353 188
rect 597 156 629 188
<< pdiffc >>
rect 47 591 79 623
rect 47 520 79 552
rect 47 452 79 484
rect 323 591 355 623
rect 323 523 355 555
rect 323 455 355 487
rect 599 591 631 623
rect 599 520 631 552
rect 599 452 631 484
<< psubdiff >>
rect 0 16 672 30
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 608 16
rect 640 -16 672 16
rect 0 -30 672 -16
<< nsubdiff >>
rect 0 772 672 786
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 608 772
rect 640 740 672 772
rect 0 726 672 740
<< psubdiffcont >>
rect 32 -16 64 16
rect 128 -16 160 16
rect 224 -16 256 16
rect 320 -16 352 16
rect 416 -16 448 16
rect 512 -16 544 16
rect 608 -16 640 16
<< nsubdiffcont >>
rect 32 740 64 772
rect 128 740 160 772
rect 224 740 256 772
rect 320 740 352 772
rect 416 740 448 772
rect 512 740 544 772
rect 608 740 640 772
<< poly >>
rect 101 637 301 673
rect 377 637 577 673
rect 101 401 301 437
rect 377 401 577 437
rect 101 344 167 401
rect 101 312 118 344
rect 150 312 167 344
rect 101 296 167 312
rect 244 343 431 361
rect 244 311 260 343
rect 292 311 381 343
rect 413 311 431 343
rect 244 283 431 311
rect 511 344 577 401
rect 511 312 526 344
rect 558 312 577 344
rect 511 296 577 312
rect 244 250 299 283
rect 99 214 299 250
rect 375 250 431 283
rect 375 214 575 250
rect 99 94 299 130
rect 375 94 575 130
<< polycont >>
rect 118 312 150 344
rect 260 311 292 343
rect 381 311 413 343
rect 526 312 558 344
<< metal1 >>
rect 0 772 672 800
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 608 772
rect 640 740 672 772
rect 0 712 672 740
rect 37 623 89 712
rect 37 591 47 623
rect 79 591 89 623
rect 37 552 89 591
rect 37 520 47 552
rect 79 520 89 552
rect 37 484 89 520
rect 37 452 47 484
rect 79 452 89 484
rect 37 441 89 452
rect 244 623 431 712
rect 244 591 323 623
rect 355 591 431 623
rect 244 555 431 591
rect 244 523 323 555
rect 355 523 431 555
rect 244 487 431 523
rect 244 455 323 487
rect 355 455 431 487
rect 104 344 162 362
rect 104 312 118 344
rect 150 312 162 344
rect 104 198 162 312
rect 244 343 431 455
rect 589 623 641 712
rect 589 591 599 623
rect 631 591 641 623
rect 589 552 641 591
rect 589 520 599 552
rect 631 520 641 552
rect 589 484 641 520
rect 589 452 599 484
rect 631 452 641 484
rect 589 442 641 452
rect 244 311 260 343
rect 292 311 381 343
rect 413 311 431 343
rect 244 295 431 311
rect 517 344 567 362
rect 517 312 526 344
rect 558 312 567 344
rect 35 188 162 198
rect 35 156 45 188
rect 77 156 162 188
rect 35 44 162 156
rect 306 188 367 206
rect 306 156 321 188
rect 353 156 367 188
rect 306 44 367 156
rect 517 198 567 312
rect 517 188 639 198
rect 517 156 597 188
rect 629 156 639 188
rect 517 44 639 156
rect 0 16 672 44
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 608 16
rect 640 -16 672 16
rect 0 -44 672 -16
<< labels >>
flabel metal1 s 0 712 672 800 0 FreeSans 400 0 0 0 VDD
port 2 nsew
flabel metal1 s 0 -44 672 44 0 FreeSans 400 0 0 0 VSS
port 3 nsew
<< properties >>
string FIXED_BBOX 0 0 672 756
string GDS_END 3472
string GDS_FILE ../gds/rgb_buffers.gds
string GDS_START 116
<< end >>
