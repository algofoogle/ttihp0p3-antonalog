magic
tech ihp-sg13g2
magscale 1 2
timestamp 1747056038
<< nwell >>
rect -48 350 1008 834
<< pwell >>
rect 33 56 945 292
rect -26 -56 986 56
<< nmos >>
rect 127 156 153 266
rect 259 118 285 266
rect 356 118 382 266
rect 470 118 496 266
rect 678 118 704 266
rect 784 118 810 266
<< pmos >>
rect 127 412 153 580
rect 259 412 285 612
rect 418 412 444 612
rect 533 412 559 612
rect 678 412 704 612
rect 784 412 810 636
<< ndiff >>
rect 59 226 127 266
rect 59 194 73 226
rect 105 194 127 226
rect 59 156 127 194
rect 153 252 259 266
rect 153 220 181 252
rect 213 220 259 252
rect 153 164 259 220
rect 153 156 181 164
rect 167 132 181 156
rect 213 132 259 164
rect 167 118 259 132
rect 285 118 356 266
rect 382 164 470 266
rect 382 132 412 164
rect 444 132 470 164
rect 382 118 470 132
rect 496 118 678 266
rect 704 165 784 266
rect 704 133 730 165
rect 762 133 784 165
rect 704 118 784 133
rect 810 248 919 266
rect 810 216 866 248
rect 898 216 919 248
rect 810 167 919 216
rect 810 135 866 167
rect 898 135 919 167
rect 810 118 919 135
<< pdiff >>
rect 718 612 784 636
rect 183 580 259 612
rect 59 566 127 580
rect 59 534 73 566
rect 105 534 127 566
rect 59 471 127 534
rect 59 439 73 471
rect 105 439 127 471
rect 59 412 127 439
rect 153 561 259 580
rect 153 529 205 561
rect 237 529 259 561
rect 153 412 259 529
rect 285 412 418 612
rect 444 573 533 612
rect 444 541 470 573
rect 502 541 533 573
rect 444 458 533 541
rect 444 426 470 458
rect 502 426 533 458
rect 444 412 533 426
rect 559 412 678 612
rect 704 596 784 612
rect 704 564 730 596
rect 762 564 784 596
rect 704 526 784 564
rect 704 494 730 526
rect 762 494 784 526
rect 704 458 784 494
rect 704 426 730 458
rect 762 426 784 458
rect 704 412 784 426
rect 810 622 918 636
rect 810 590 866 622
rect 898 590 918 622
rect 810 539 918 590
rect 810 507 866 539
rect 898 507 918 539
rect 810 458 918 507
rect 810 426 866 458
rect 898 426 918 458
rect 810 412 918 426
<< ndiffc >>
rect 73 194 105 226
rect 181 220 213 252
rect 181 132 213 164
rect 412 132 444 164
rect 730 133 762 165
rect 866 216 898 248
rect 866 135 898 167
<< pdiffc >>
rect 73 534 105 566
rect 73 439 105 471
rect 205 529 237 561
rect 470 541 502 573
rect 470 426 502 458
rect 730 564 762 596
rect 730 494 762 526
rect 730 426 762 458
rect 866 590 898 622
rect 866 507 898 539
rect 866 426 898 458
<< psubdiff >>
rect 0 16 960 30
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 608 16
rect 640 -16 704 16
rect 736 -16 800 16
rect 832 -16 896 16
rect 928 -16 960 16
rect 0 -30 960 -16
<< nsubdiff >>
rect 0 772 960 786
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 608 772
rect 640 740 704 772
rect 736 740 800 772
rect 832 740 896 772
rect 928 740 960 772
rect 0 726 960 740
<< psubdiffcont >>
rect 32 -16 64 16
rect 128 -16 160 16
rect 224 -16 256 16
rect 320 -16 352 16
rect 416 -16 448 16
rect 512 -16 544 16
rect 608 -16 640 16
rect 704 -16 736 16
rect 800 -16 832 16
rect 896 -16 928 16
<< nsubdiffcont >>
rect 32 740 64 772
rect 128 740 160 772
rect 224 740 256 772
rect 320 740 352 772
rect 416 740 448 772
rect 512 740 544 772
rect 608 740 640 772
rect 704 740 736 772
rect 800 740 832 772
rect 896 740 928 772
<< poly >>
rect 127 580 153 616
rect 259 612 285 648
rect 418 612 444 648
rect 533 612 559 648
rect 678 612 704 648
rect 784 636 810 672
rect 127 380 153 412
rect 259 380 285 412
rect 127 362 285 380
rect 127 330 141 362
rect 173 330 285 362
rect 418 354 444 412
rect 533 354 559 412
rect 678 374 704 412
rect 678 356 744 374
rect 127 314 285 330
rect 127 266 153 314
rect 259 266 285 314
rect 322 336 382 350
rect 322 304 336 336
rect 368 304 382 336
rect 322 290 382 304
rect 356 266 382 290
rect 418 336 496 354
rect 418 304 434 336
rect 466 304 496 336
rect 418 288 496 304
rect 533 336 599 354
rect 533 304 549 336
rect 581 304 599 336
rect 533 288 599 304
rect 678 324 694 356
rect 726 324 744 356
rect 678 308 744 324
rect 784 370 810 412
rect 784 352 850 370
rect 784 320 802 352
rect 834 320 850 352
rect 470 266 496 288
rect 678 266 704 308
rect 784 304 850 320
rect 784 266 810 304
rect 127 120 153 156
rect 259 82 285 118
rect 356 82 382 118
rect 470 82 496 118
rect 678 82 704 118
rect 784 82 810 118
<< polycont >>
rect 141 330 173 362
rect 336 304 368 336
rect 434 304 466 336
rect 549 304 581 336
rect 694 324 726 356
rect 802 320 834 352
<< metal1 >>
rect 0 772 960 800
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 608 772
rect 640 740 704 772
rect 736 740 800 772
rect 832 740 896 772
rect 928 740 960 772
rect 0 712 960 740
rect 29 566 115 569
rect 29 534 73 566
rect 105 534 115 566
rect 29 492 115 534
rect 195 561 247 712
rect 195 529 205 561
rect 237 529 247 561
rect 195 528 247 529
rect 296 625 685 659
rect 296 492 328 625
rect 29 471 328 492
rect 29 439 73 471
rect 105 460 328 471
rect 460 573 512 575
rect 460 541 470 573
rect 502 541 512 573
rect 105 439 115 460
rect 29 434 115 439
rect 460 458 512 541
rect 29 236 70 434
rect 460 429 470 458
rect 364 426 470 429
rect 502 426 512 458
rect 364 424 512 426
rect 254 393 512 424
rect 254 391 378 393
rect 120 362 218 381
rect 120 330 141 362
rect 173 330 218 362
rect 120 300 218 330
rect 171 252 218 262
rect 29 226 115 236
rect 29 194 73 226
rect 105 194 115 226
rect 29 184 115 194
rect 171 220 181 252
rect 213 220 218 252
rect 171 164 218 220
rect 171 132 181 164
rect 213 132 218 164
rect 171 44 218 132
rect 254 166 286 391
rect 650 374 685 625
rect 726 596 766 712
rect 726 564 730 596
rect 762 564 766 596
rect 726 526 766 564
rect 726 494 730 526
rect 762 494 766 526
rect 726 458 766 494
rect 726 426 730 458
rect 762 426 766 458
rect 726 416 766 426
rect 827 622 937 640
rect 827 590 866 622
rect 898 590 937 622
rect 827 539 937 590
rect 827 507 866 539
rect 898 507 937 539
rect 827 458 937 507
rect 827 426 866 458
rect 898 426 937 458
rect 827 408 937 426
rect 322 336 378 351
rect 322 304 336 336
rect 368 304 378 336
rect 322 288 378 304
rect 342 240 378 288
rect 418 336 496 357
rect 418 304 434 336
rect 466 304 496 336
rect 418 280 496 304
rect 539 336 598 357
rect 539 304 549 336
rect 581 304 598 336
rect 650 356 744 374
rect 650 324 694 356
rect 726 324 744 356
rect 650 308 744 324
rect 789 352 849 370
rect 789 320 802 352
rect 834 320 849 352
rect 539 240 598 304
rect 789 304 849 320
rect 789 240 827 304
rect 903 263 937 408
rect 342 206 598 240
rect 639 206 827 240
rect 863 248 937 263
rect 863 216 866 248
rect 898 216 937 248
rect 639 166 673 206
rect 254 164 673 166
rect 254 132 412 164
rect 444 132 673 164
rect 254 122 673 132
rect 720 165 772 169
rect 720 133 730 165
rect 762 133 772 165
rect 720 44 772 133
rect 863 167 937 216
rect 863 135 866 167
rect 898 135 937 167
rect 863 114 937 135
rect 0 16 960 44
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 608 16
rect 640 -16 704 16
rect 736 -16 800 16
rect 832 -16 896 16
rect 928 -16 960 16
rect 0 -44 960 -16
<< labels >>
flabel metal1 s 539 206 598 357 0 FreeSans 400 0 0 0 A1
port 2 nsew
flabel metal1 s 827 408 937 640 0 FreeSans 400 0 0 0 X
port 3 nsew
flabel metal1 s 120 300 218 381 0 FreeSans 400 0 0 0 S
port 4 nsew
flabel metal1 s 0 712 960 800 0 FreeSans 400 0 0 0 VDD
port 5 nsew
flabel metal1 s 0 -44 960 44 0 FreeSans 400 0 0 0 VSS
port 6 nsew
flabel metal1 s 418 280 496 357 0 FreeSans 400 0 0 0 A0
port 7 nsew
<< properties >>
string FIXED_BBOX 0 0 960 756
string GDS_END 179930
string GDS_FILE ../gds/controller.gds
string GDS_START 172918
<< end >>
