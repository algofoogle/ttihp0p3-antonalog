magic
tech ihp-sg13g2
magscale 1 2
timestamp 1747056038
<< nwell >>
rect -48 350 528 834
<< pwell >>
rect 31 56 449 314
rect -26 -56 506 56
<< nmos >>
rect 125 140 151 288
rect 227 140 253 288
rect 329 140 355 288
<< pmos >>
rect 125 412 151 636
rect 227 412 253 636
rect 329 412 355 636
<< ndiff >>
rect 57 186 125 288
rect 57 154 71 186
rect 103 154 125 186
rect 57 140 125 154
rect 151 274 227 288
rect 151 242 173 274
rect 205 242 227 274
rect 151 186 227 242
rect 151 154 173 186
rect 205 154 227 186
rect 151 140 227 154
rect 253 140 329 288
rect 355 274 423 288
rect 355 242 377 274
rect 409 242 423 274
rect 355 186 423 242
rect 355 154 377 186
rect 409 154 423 186
rect 355 140 423 154
<< pdiff >>
rect 57 622 125 636
rect 57 590 71 622
rect 103 590 125 622
rect 57 543 125 590
rect 57 511 71 543
rect 103 511 125 543
rect 57 458 125 511
rect 57 426 71 458
rect 103 426 125 458
rect 57 412 125 426
rect 151 622 227 636
rect 151 590 173 622
rect 205 590 227 622
rect 151 543 227 590
rect 151 511 173 543
rect 205 511 227 543
rect 151 412 227 511
rect 253 622 329 636
rect 253 590 275 622
rect 307 590 329 622
rect 253 412 329 590
rect 355 622 423 636
rect 355 590 377 622
rect 409 590 423 622
rect 355 543 423 590
rect 355 511 377 543
rect 409 511 423 543
rect 355 458 423 511
rect 355 426 377 458
rect 409 426 423 458
rect 355 412 423 426
<< ndiffc >>
rect 71 154 103 186
rect 173 242 205 274
rect 173 154 205 186
rect 377 242 409 274
rect 377 154 409 186
<< pdiffc >>
rect 71 590 103 622
rect 71 511 103 543
rect 71 426 103 458
rect 173 590 205 622
rect 173 511 205 543
rect 275 590 307 622
rect 377 590 409 622
rect 377 511 409 543
rect 377 426 409 458
<< psubdiff >>
rect 0 16 480 30
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 480 16
rect 0 -30 480 -16
<< nsubdiff >>
rect 0 772 480 786
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 480 772
rect 0 726 480 740
<< psubdiffcont >>
rect 32 -16 64 16
rect 128 -16 160 16
rect 224 -16 256 16
rect 320 -16 352 16
rect 416 -16 448 16
<< nsubdiffcont >>
rect 32 740 64 772
rect 128 740 160 772
rect 224 740 256 772
rect 320 740 352 772
rect 416 740 448 772
<< poly >>
rect 125 636 151 672
rect 227 636 253 672
rect 329 636 355 672
rect 125 380 151 412
rect 227 380 253 412
rect 329 380 355 412
rect 57 366 151 380
rect 57 334 71 366
rect 103 334 151 366
rect 57 320 151 334
rect 210 366 270 380
rect 210 334 224 366
rect 256 334 270 366
rect 210 320 270 334
rect 329 366 423 380
rect 329 334 377 366
rect 409 334 423 366
rect 329 320 423 334
rect 125 288 151 320
rect 227 288 253 320
rect 329 288 355 320
rect 125 104 151 140
rect 227 104 253 140
rect 329 104 355 140
<< polycont >>
rect 71 334 103 366
rect 224 334 256 366
rect 377 334 409 366
<< metal1 >>
rect 0 772 480 800
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 480 772
rect 0 712 480 740
rect 265 622 317 712
rect 61 590 71 622
rect 103 590 113 622
rect 61 543 113 590
rect 61 511 71 543
rect 103 511 113 543
rect 163 590 173 622
rect 205 590 215 622
rect 163 543 215 590
rect 265 590 275 622
rect 307 590 317 622
rect 265 580 317 590
rect 367 590 377 622
rect 409 590 419 622
rect 367 543 419 590
rect 163 511 173 543
rect 205 511 377 543
rect 409 511 419 543
rect 61 458 113 511
rect 215 458 419 511
rect 61 426 71 458
rect 103 426 178 458
rect 215 426 377 458
rect 409 426 419 458
rect 61 366 106 380
rect 61 334 71 366
rect 103 334 106 366
rect 61 231 106 334
rect 143 274 178 426
rect 353 366 419 390
rect 214 334 224 366
rect 256 334 317 366
rect 214 324 317 334
rect 143 242 173 274
rect 205 242 215 274
rect 163 186 215 242
rect 61 154 71 186
rect 103 154 113 186
rect 163 154 173 186
rect 205 154 215 186
rect 265 154 317 324
rect 353 334 377 366
rect 409 334 419 366
rect 353 310 419 334
rect 367 242 377 274
rect 409 242 419 274
rect 367 186 419 242
rect 367 154 377 186
rect 409 154 419 186
rect 61 44 113 154
rect 367 44 419 154
rect 0 16 480 44
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 480 16
rect 0 -44 480 -16
<< labels >>
flabel metal1 s 0 712 480 800 0 FreeSans 400 0 0 0 VDD
port 2 nsew
flabel metal1 s 0 -44 480 44 0 FreeSans 400 0 0 0 VSS
port 3 nsew
flabel metal1 s 362 310 394 390 0 FreeSans 400 0 0 0 A2
port 4 nsew
flabel metal1 s 266 154 298 366 0 FreeSans 400 0 0 0 A1
port 5 nsew
flabel metal1 s 74 231 106 380 0 FreeSans 400 0 0 0 B1
port 6 nsew
flabel metal1 s 74 426 106 622 0 FreeSans 400 0 0 0 Y
port 7 nsew
<< properties >>
string FIXED_BBOX 0 0 480 756
string GDS_END 45568
string GDS_FILE ../gds/controller.gds
string GDS_START 41548
<< end >>
