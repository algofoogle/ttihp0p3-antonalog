magic
tech ihp-sg13g2
magscale 1 2
timestamp 1746816402
<< nwell >>
rect -48 350 912 834
<< pwell >>
rect 495 272 855 292
rect 109 56 855 272
rect -26 -56 890 56
<< nmos >>
rect 203 118 229 246
rect 281 118 307 246
rect 359 118 385 246
rect 473 118 499 246
rect 575 118 601 266
rect 705 118 731 266
<< pmos >>
rect 149 468 175 636
rect 251 468 277 636
rect 353 468 379 636
rect 467 468 493 636
rect 575 412 601 636
rect 705 412 731 636
<< ndiff >>
rect 521 246 575 266
rect 135 232 203 246
rect 135 200 149 232
rect 181 200 203 232
rect 135 164 203 200
rect 135 132 149 164
rect 181 132 203 164
rect 135 118 203 132
rect 229 118 281 246
rect 307 118 359 246
rect 385 118 473 246
rect 499 232 575 246
rect 499 200 521 232
rect 553 200 575 232
rect 499 164 575 200
rect 499 132 521 164
rect 553 132 575 164
rect 499 118 575 132
rect 601 252 705 266
rect 601 220 651 252
rect 683 220 705 252
rect 601 164 705 220
rect 601 132 651 164
rect 683 132 705 164
rect 601 118 705 132
rect 731 252 829 266
rect 731 220 783 252
rect 815 220 829 252
rect 731 164 829 220
rect 731 132 783 164
rect 815 132 829 164
rect 731 118 829 132
<< pdiff >>
rect 81 622 149 636
rect 81 590 95 622
rect 127 590 149 622
rect 81 546 149 590
rect 81 514 95 546
rect 127 514 149 546
rect 81 468 149 514
rect 175 622 251 636
rect 175 590 197 622
rect 229 590 251 622
rect 175 515 251 590
rect 175 483 197 515
rect 229 483 251 515
rect 175 468 251 483
rect 277 622 353 636
rect 277 590 299 622
rect 331 590 353 622
rect 277 546 353 590
rect 277 514 299 546
rect 331 514 353 546
rect 277 468 353 514
rect 379 622 467 636
rect 379 590 407 622
rect 439 590 467 622
rect 379 515 467 590
rect 379 483 407 515
rect 439 483 467 515
rect 379 468 467 483
rect 493 622 575 636
rect 493 590 518 622
rect 550 590 575 622
rect 493 552 575 590
rect 493 520 518 552
rect 550 520 575 552
rect 493 468 575 520
rect 529 412 575 468
rect 601 622 705 636
rect 601 590 651 622
rect 683 590 705 622
rect 601 543 705 590
rect 601 511 651 543
rect 683 511 705 543
rect 601 458 705 511
rect 601 426 651 458
rect 683 426 705 458
rect 601 412 705 426
rect 731 622 829 636
rect 731 590 783 622
rect 815 590 829 622
rect 731 543 829 590
rect 731 511 783 543
rect 815 511 829 543
rect 731 458 829 511
rect 731 426 783 458
rect 815 426 829 458
rect 731 412 829 426
<< ndiffc >>
rect 149 200 181 232
rect 149 132 181 164
rect 521 200 553 232
rect 521 132 553 164
rect 651 220 683 252
rect 651 132 683 164
rect 783 220 815 252
rect 783 132 815 164
<< pdiffc >>
rect 95 590 127 622
rect 95 514 127 546
rect 197 590 229 622
rect 197 483 229 515
rect 299 590 331 622
rect 299 514 331 546
rect 407 590 439 622
rect 407 483 439 515
rect 518 590 550 622
rect 518 520 550 552
rect 651 590 683 622
rect 651 511 683 543
rect 651 426 683 458
rect 783 590 815 622
rect 783 511 815 543
rect 783 426 815 458
<< psubdiff >>
rect 0 16 864 30
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 608 16
rect 640 -16 704 16
rect 736 -16 800 16
rect 832 -16 864 16
rect 0 -30 864 -16
<< nsubdiff >>
rect 0 772 864 786
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 608 772
rect 640 740 704 772
rect 736 740 800 772
rect 832 740 864 772
rect 0 726 864 740
<< psubdiffcont >>
rect 32 -16 64 16
rect 128 -16 160 16
rect 224 -16 256 16
rect 320 -16 352 16
rect 416 -16 448 16
rect 512 -16 544 16
rect 608 -16 640 16
rect 704 -16 736 16
rect 800 -16 832 16
<< nsubdiffcont >>
rect 32 740 64 772
rect 128 740 160 772
rect 224 740 256 772
rect 320 740 352 772
rect 416 740 448 772
rect 512 740 544 772
rect 608 740 640 772
rect 704 740 736 772
rect 800 740 832 772
<< poly >>
rect 149 636 175 672
rect 251 636 277 672
rect 353 636 379 672
rect 467 636 493 672
rect 575 636 601 672
rect 705 636 731 672
rect 149 453 175 468
rect 251 453 277 468
rect 147 402 183 453
rect 247 405 283 453
rect 353 426 379 468
rect 139 384 205 402
rect 139 352 155 384
rect 187 352 205 384
rect 139 316 205 352
rect 247 387 317 405
rect 353 402 425 426
rect 247 355 267 387
rect 299 355 317 387
rect 247 339 317 355
rect 359 384 425 402
rect 359 352 375 384
rect 407 352 425 384
rect 139 284 155 316
rect 187 291 205 316
rect 187 284 229 291
rect 139 261 229 284
rect 203 246 229 261
rect 281 246 307 339
rect 359 316 425 352
rect 359 284 375 316
rect 407 284 425 316
rect 467 380 493 468
rect 575 380 601 412
rect 705 380 731 412
rect 467 362 533 380
rect 467 330 483 362
rect 515 330 533 362
rect 467 314 533 330
rect 575 356 731 380
rect 575 324 591 356
rect 623 324 731 356
rect 359 268 425 284
rect 359 246 385 268
rect 473 246 499 314
rect 575 308 731 324
rect 575 266 601 308
rect 705 266 731 308
rect 203 82 229 118
rect 281 82 307 118
rect 359 82 385 118
rect 473 82 499 118
rect 575 82 601 118
rect 705 82 731 118
<< polycont >>
rect 155 352 187 384
rect 267 355 299 387
rect 375 352 407 384
rect 155 284 187 316
rect 375 284 407 316
rect 483 330 515 362
rect 591 324 623 356
<< metal1 >>
rect 0 772 864 800
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 608 772
rect 640 740 704 772
rect 736 740 800 772
rect 832 740 864 772
rect 0 712 864 740
rect 85 622 137 712
rect 85 590 95 622
rect 127 590 137 622
rect 85 546 137 590
rect 85 514 95 546
rect 127 514 137 546
rect 85 512 137 514
rect 187 622 239 625
rect 187 590 197 622
rect 229 590 239 622
rect 187 515 239 590
rect 187 483 197 515
rect 229 483 239 515
rect 289 622 341 712
rect 289 590 299 622
rect 331 590 341 622
rect 289 546 341 590
rect 289 514 299 546
rect 331 514 341 546
rect 289 512 341 514
rect 397 622 449 624
rect 397 590 407 622
rect 439 590 449 622
rect 397 515 449 590
rect 508 622 560 712
rect 508 590 518 622
rect 550 590 560 622
rect 508 552 560 590
rect 508 520 518 552
rect 550 520 560 552
rect 508 517 560 520
rect 641 622 737 624
rect 641 590 651 622
rect 683 590 737 622
rect 641 543 737 590
rect 187 476 239 483
rect 397 483 407 515
rect 439 483 449 515
rect 397 476 449 483
rect 641 511 651 543
rect 683 511 737 543
rect 71 444 602 476
rect 71 234 105 444
rect 141 384 214 402
rect 141 352 155 384
rect 187 352 214 384
rect 141 316 214 352
rect 141 284 155 316
rect 187 284 214 316
rect 141 270 214 284
rect 251 387 313 405
rect 251 355 267 387
rect 299 355 313 387
rect 71 232 199 234
rect 71 200 149 232
rect 181 200 199 232
rect 71 164 199 200
rect 71 132 149 164
rect 181 132 199 164
rect 251 132 313 355
rect 359 384 425 402
rect 359 352 375 384
rect 407 352 425 384
rect 359 316 425 352
rect 359 284 375 316
rect 407 284 425 316
rect 463 362 533 400
rect 463 330 483 362
rect 515 330 533 362
rect 463 314 533 330
rect 570 374 602 444
rect 641 458 737 511
rect 641 426 651 458
rect 683 426 737 458
rect 773 622 825 712
rect 773 590 783 622
rect 815 590 825 622
rect 773 543 825 590
rect 773 511 783 543
rect 815 511 825 543
rect 773 458 825 511
rect 773 426 783 458
rect 815 426 825 458
rect 641 414 737 426
rect 570 356 641 374
rect 570 324 591 356
rect 623 324 641 356
rect 570 308 641 324
rect 359 132 425 284
rect 705 252 737 414
rect 510 232 563 242
rect 510 200 521 232
rect 553 200 563 232
rect 510 164 563 200
rect 510 132 521 164
rect 553 132 563 164
rect 71 129 199 132
rect 510 44 563 132
rect 641 220 651 252
rect 683 220 737 252
rect 641 164 737 220
rect 641 132 651 164
rect 683 132 737 164
rect 641 128 737 132
rect 773 220 783 252
rect 815 220 825 252
rect 773 164 825 220
rect 773 132 783 164
rect 815 132 825 164
rect 773 44 825 132
rect 0 16 864 44
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 608 16
rect 640 -16 704 16
rect 736 -16 800 16
rect 832 -16 864 16
rect 0 -44 864 -16
<< labels >>
flabel metal1 s 641 414 737 624 0 FreeSans 400 0 0 0 X
port 2 nsew
flabel metal1 s 251 132 313 405 0 FreeSans 400 0 0 0 B
port 3 nsew
flabel metal1 s 141 270 214 402 0 FreeSans 400 0 0 0 A
port 4 nsew
flabel metal1 s 0 712 864 800 0 FreeSans 400 0 0 0 VDD
port 5 nsew
flabel metal1 s 0 -44 864 44 0 FreeSans 400 0 0 0 VSS
port 6 nsew
flabel metal1 s 359 132 425 402 0 FreeSans 400 0 0 0 C
port 7 nsew
flabel metal1 s 463 314 533 400 0 FreeSans 400 0 0 0 D
port 8 nsew
<< properties >>
string FIXED_BBOX 0 0 864 756
string GDS_END 254024
string GDS_FILE ../gds/controller.gds
string GDS_START 247910
<< end >>
