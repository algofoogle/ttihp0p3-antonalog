magic
tech ihp-sg13g2
magscale 1 2
timestamp 1747056038
<< nwell >>
rect -48 350 720 834
<< pwell >>
rect 50 56 570 314
rect -26 -56 698 56
<< nmos >>
rect 144 160 170 288
rect 246 160 272 288
rect 348 160 374 288
rect 450 140 476 288
<< pmos >>
rect 144 471 170 639
rect 246 471 272 639
rect 348 471 374 639
rect 518 434 544 658
<< ndiff >>
rect 76 253 144 288
rect 76 221 90 253
rect 122 221 144 253
rect 76 160 144 221
rect 170 160 246 288
rect 272 160 348 288
rect 374 210 450 288
rect 374 178 396 210
rect 428 178 450 210
rect 374 160 450 178
rect 388 140 450 160
rect 476 263 544 288
rect 476 231 498 263
rect 530 231 544 263
rect 476 195 544 231
rect 476 163 498 195
rect 530 163 544 195
rect 476 140 544 163
<< pdiff >>
rect 388 639 518 658
rect 76 618 144 639
rect 76 586 90 618
rect 122 586 144 618
rect 76 527 144 586
rect 76 495 90 527
rect 122 495 144 527
rect 76 471 144 495
rect 170 580 246 639
rect 170 548 192 580
rect 224 548 246 580
rect 170 471 246 548
rect 272 613 348 639
rect 272 581 294 613
rect 326 581 348 613
rect 272 534 348 581
rect 272 502 294 534
rect 326 502 348 534
rect 272 471 348 502
rect 374 626 518 639
rect 374 594 396 626
rect 428 594 464 626
rect 496 594 518 626
rect 374 558 518 594
rect 374 526 396 558
rect 428 526 464 558
rect 496 526 518 558
rect 374 471 518 526
rect 456 434 518 471
rect 544 644 612 658
rect 544 612 566 644
rect 598 612 612 644
rect 544 572 612 612
rect 544 540 566 572
rect 598 540 612 572
rect 544 492 612 540
rect 544 460 566 492
rect 598 460 612 492
rect 544 434 612 460
<< ndiffc >>
rect 90 221 122 253
rect 396 178 428 210
rect 498 231 530 263
rect 498 163 530 195
<< pdiffc >>
rect 90 586 122 618
rect 90 495 122 527
rect 192 548 224 580
rect 294 581 326 613
rect 294 502 326 534
rect 396 594 428 626
rect 464 594 496 626
rect 396 526 428 558
rect 464 526 496 558
rect 566 612 598 644
rect 566 540 598 572
rect 566 460 598 492
<< psubdiff >>
rect 0 16 672 30
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 608 16
rect 640 -16 672 16
rect 0 -30 672 -16
<< nsubdiff >>
rect 0 772 672 786
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 608 772
rect 640 740 672 772
rect 0 726 672 740
<< psubdiffcont >>
rect 32 -16 64 16
rect 128 -16 160 16
rect 224 -16 256 16
rect 320 -16 352 16
rect 416 -16 448 16
rect 512 -16 544 16
rect 608 -16 640 16
<< nsubdiffcont >>
rect 32 740 64 772
rect 128 740 160 772
rect 224 740 256 772
rect 320 740 352 772
rect 416 740 448 772
rect 512 740 544 772
rect 608 740 640 772
<< poly >>
rect 144 639 170 675
rect 246 639 272 675
rect 348 639 374 675
rect 518 658 544 701
rect 144 288 170 471
rect 246 396 272 471
rect 348 400 374 471
rect 218 379 284 396
rect 218 347 235 379
rect 267 347 284 379
rect 218 330 284 347
rect 346 383 412 400
rect 346 351 363 383
rect 395 351 412 383
rect 518 380 544 434
rect 346 334 412 351
rect 450 363 544 380
rect 246 288 272 330
rect 348 288 374 334
rect 450 331 480 363
rect 512 331 544 363
rect 450 314 544 331
rect 450 288 476 314
rect 144 146 170 160
rect 70 132 204 146
rect 70 100 87 132
rect 119 100 155 132
rect 187 100 204 132
rect 246 108 272 160
rect 348 109 374 160
rect 450 104 476 140
rect 70 78 204 100
<< polycont >>
rect 235 347 267 379
rect 363 351 395 383
rect 480 331 512 363
rect 87 100 119 132
rect 155 100 187 132
<< metal1 >>
rect 0 772 672 800
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 608 772
rect 640 740 672 772
rect 0 712 672 740
rect 80 618 132 623
rect 80 586 90 618
rect 122 586 132 618
rect 80 527 132 586
rect 182 580 234 712
rect 386 626 506 712
rect 182 548 192 580
rect 224 548 234 580
rect 182 546 234 548
rect 284 613 336 617
rect 284 581 294 613
rect 326 581 336 613
rect 80 495 90 527
rect 122 495 132 527
rect 80 464 132 495
rect 284 534 336 581
rect 284 502 294 534
rect 326 502 336 534
rect 386 594 396 626
rect 428 594 464 626
rect 496 594 506 626
rect 386 558 506 594
rect 386 526 396 558
rect 428 526 464 558
rect 496 526 506 558
rect 386 523 506 526
rect 556 644 613 654
rect 556 612 566 644
rect 598 612 613 644
rect 556 572 613 612
rect 556 540 566 572
rect 598 540 613 572
rect 284 464 336 502
rect 556 492 613 540
rect 80 432 481 464
rect 556 460 566 492
rect 598 460 613 492
rect 556 434 613 460
rect 80 253 132 432
rect 218 379 308 396
rect 218 347 235 379
rect 267 347 308 379
rect 218 280 308 347
rect 346 383 412 390
rect 346 351 363 383
rect 395 351 412 383
rect 346 280 412 351
rect 449 380 481 432
rect 449 363 529 380
rect 449 331 480 363
rect 512 331 529 363
rect 449 314 529 331
rect 579 277 613 434
rect 80 221 90 253
rect 122 221 132 253
rect 488 263 613 277
rect 488 231 498 263
rect 530 231 613 263
rect 80 218 132 221
rect 245 158 318 218
rect 70 132 318 158
rect 70 100 87 132
rect 119 100 155 132
rect 187 100 318 132
rect 70 95 318 100
rect 386 210 438 228
rect 386 178 396 210
rect 428 178 438 210
rect 386 44 438 178
rect 488 225 613 231
rect 488 195 540 225
rect 488 163 498 195
rect 530 163 540 195
rect 488 154 540 163
rect 0 16 672 44
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 608 16
rect 640 -16 672 16
rect 0 -44 672 -16
<< labels >>
flabel metal1 s 488 225 613 277 0 FreeSans 400 0 0 0 X
port 2 nsew
flabel metal1 s 218 280 308 396 0 FreeSans 400 0 0 0 B
port 3 nsew
flabel metal1 s 0 712 672 800 0 FreeSans 400 0 0 0 VDD
port 4 nsew
flabel metal1 s 0 -44 672 44 0 FreeSans 400 0 0 0 VSS
port 5 nsew
flabel metal1 s 346 280 412 390 0 FreeSans 400 0 0 0 C
port 6 nsew
flabel metal1 s 245 95 318 218 0 FreeSans 400 0 0 0 A
port 7 nsew
<< properties >>
string FIXED_BBOX 0 0 672 756
string GDS_END 108634
string GDS_FILE ../gds/controller.gds
string GDS_START 102998
<< end >>
