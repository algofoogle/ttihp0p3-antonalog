magic
tech ihp-sg13g2
timestamp 1747537721
<< nwell >>
rect -24 175 408 417
<< pwell >>
rect -2 28 363 142
rect -13 -28 397 28
<< nmos >>
rect 45 74 58 129
rect 149 57 162 129
rect 200 57 213 129
rect 252 57 265 129
rect 303 57 316 129
<< pmos >>
rect 45 206 58 290
rect 149 206 162 318
rect 200 206 213 318
rect 252 206 265 318
rect 303 206 316 318
<< ndiff >>
rect 11 122 45 129
rect 11 106 18 122
rect 34 106 45 122
rect 11 74 45 106
rect 58 122 92 129
rect 58 106 69 122
rect 85 106 92 122
rect 58 74 92 106
rect 113 115 149 129
rect 113 99 120 115
rect 136 99 149 115
rect 113 81 149 99
rect 113 65 121 81
rect 137 65 149 81
rect 113 57 149 65
rect 162 80 200 129
rect 162 64 173 80
rect 189 64 200 80
rect 162 57 200 64
rect 213 116 252 129
rect 213 100 224 116
rect 240 100 252 116
rect 213 82 252 100
rect 213 66 224 82
rect 240 66 252 82
rect 213 57 252 66
rect 265 121 303 129
rect 265 105 276 121
rect 292 105 303 121
rect 265 57 303 105
rect 316 115 350 129
rect 316 99 327 115
rect 343 99 350 115
rect 316 81 350 99
rect 316 65 327 81
rect 343 65 350 81
rect 316 57 350 65
<< pdiff >>
rect 113 311 149 318
rect 113 295 120 311
rect 136 295 149 311
rect 11 283 45 290
rect 11 267 18 283
rect 34 267 45 283
rect 11 229 45 267
rect 11 213 18 229
rect 34 213 45 229
rect 11 206 45 213
rect 58 283 92 290
rect 58 267 69 283
rect 85 267 92 283
rect 58 229 92 267
rect 58 213 69 229
rect 85 213 92 229
rect 58 206 92 213
rect 113 270 149 295
rect 113 254 120 270
rect 136 254 149 270
rect 113 230 149 254
rect 113 214 120 230
rect 136 214 149 230
rect 113 206 149 214
rect 162 311 200 318
rect 162 295 173 311
rect 189 295 200 311
rect 162 271 200 295
rect 162 255 173 271
rect 189 255 200 271
rect 162 231 200 255
rect 162 215 173 231
rect 189 215 200 231
rect 162 206 200 215
rect 213 311 252 318
rect 213 295 224 311
rect 240 295 252 311
rect 213 206 252 295
rect 265 311 303 318
rect 265 295 276 311
rect 292 295 303 311
rect 265 271 303 295
rect 265 255 276 271
rect 292 255 303 271
rect 265 237 303 255
rect 265 221 276 237
rect 292 221 303 237
rect 265 206 303 221
rect 316 311 351 318
rect 316 295 327 311
rect 343 295 351 311
rect 316 270 351 295
rect 316 254 327 270
rect 343 254 351 270
rect 316 233 351 254
rect 316 217 327 233
rect 343 217 351 233
rect 316 206 351 217
<< ndiffc >>
rect 18 106 34 122
rect 69 106 85 122
rect 120 99 136 115
rect 121 65 137 81
rect 173 64 189 80
rect 224 100 240 116
rect 224 66 240 82
rect 276 105 292 121
rect 327 99 343 115
rect 327 65 343 81
<< pdiffc >>
rect 120 295 136 311
rect 18 267 34 283
rect 18 213 34 229
rect 69 267 85 283
rect 69 213 85 229
rect 120 254 136 270
rect 120 214 136 230
rect 173 295 189 311
rect 173 255 189 271
rect 173 215 189 231
rect 224 295 240 311
rect 276 295 292 311
rect 276 255 292 271
rect 276 221 292 237
rect 327 295 343 311
rect 327 254 343 270
rect 327 217 343 233
<< psubdiff >>
rect 0 8 384 15
rect 0 -8 16 8
rect 32 -8 64 8
rect 80 -8 112 8
rect 128 -8 160 8
rect 176 -8 208 8
rect 224 -8 256 8
rect 272 -8 304 8
rect 320 -8 352 8
rect 368 -8 384 8
rect 0 -15 384 -8
<< nsubdiff >>
rect 0 386 384 393
rect 0 370 16 386
rect 32 370 64 386
rect 80 370 112 386
rect 128 370 160 386
rect 176 370 208 386
rect 224 370 256 386
rect 272 370 304 386
rect 320 370 352 386
rect 368 370 384 386
rect 0 363 384 370
<< psubdiffcont >>
rect 16 -8 32 8
rect 64 -8 80 8
rect 112 -8 128 8
rect 160 -8 176 8
rect 208 -8 224 8
rect 256 -8 272 8
rect 304 -8 320 8
rect 352 -8 368 8
<< nsubdiffcont >>
rect 16 370 32 386
rect 64 370 80 386
rect 112 370 128 386
rect 160 370 176 386
rect 208 370 224 386
rect 256 370 272 386
rect 304 370 320 386
rect 352 370 368 386
<< poly >>
rect 149 318 162 336
rect 200 318 213 336
rect 252 318 265 336
rect 303 318 316 336
rect 45 290 58 308
rect 45 183 58 206
rect 149 187 162 206
rect 200 187 213 206
rect 149 186 213 187
rect 252 199 265 206
rect 303 199 316 206
rect 252 186 316 199
rect 33 176 63 183
rect 33 160 40 176
rect 56 160 63 176
rect 33 153 63 160
rect 119 179 213 186
rect 119 163 126 179
rect 142 163 213 179
rect 119 156 213 163
rect 231 179 316 186
rect 231 163 238 179
rect 254 168 316 179
rect 254 163 265 168
rect 231 156 265 163
rect 45 129 58 153
rect 149 129 162 156
rect 200 129 213 156
rect 252 129 265 156
rect 303 129 316 168
rect 45 56 58 74
rect 149 39 162 57
rect 200 39 213 57
rect 252 39 265 57
rect 303 39 316 57
<< polycont >>
rect 40 160 56 176
rect 126 163 142 179
rect 238 163 254 179
<< metal1 >>
rect 0 386 384 400
rect 0 370 16 386
rect 32 370 64 386
rect 80 370 112 386
rect 128 370 160 386
rect 176 370 208 386
rect 224 370 256 386
rect 272 370 304 386
rect 320 370 352 386
rect 368 370 384 386
rect 0 356 384 370
rect 13 283 39 356
rect 115 311 141 356
rect 115 295 120 311
rect 136 295 141 311
rect 13 267 18 283
rect 34 267 39 283
rect 13 229 39 267
rect 13 213 18 229
rect 34 213 39 229
rect 13 208 39 213
rect 64 283 90 288
rect 64 267 69 283
rect 85 267 90 283
rect 64 234 90 267
rect 115 270 141 295
rect 115 254 120 270
rect 136 254 141 270
rect 64 229 96 234
rect 64 213 69 229
rect 85 213 96 229
rect 64 208 96 213
rect 115 230 141 254
rect 115 214 120 230
rect 136 214 141 230
rect 167 311 193 318
rect 167 295 173 311
rect 189 295 193 311
rect 167 271 193 295
rect 218 311 244 356
rect 218 295 224 311
rect 240 295 244 311
rect 218 290 244 295
rect 272 311 298 318
rect 272 295 276 311
rect 292 295 298 311
rect 167 255 173 271
rect 189 255 193 271
rect 167 236 193 255
rect 272 271 298 295
rect 272 255 276 271
rect 292 255 298 271
rect 272 237 298 255
rect 272 236 276 237
rect 167 231 276 236
rect 167 215 173 231
rect 189 221 276 231
rect 292 221 298 237
rect 189 215 298 221
rect 167 214 298 215
rect 115 212 141 214
rect 15 176 61 186
rect 15 160 40 176
rect 56 160 61 176
rect 15 147 61 160
rect 80 184 96 208
rect 80 179 147 184
rect 80 163 126 179
rect 142 163 147 179
rect 80 158 147 163
rect 184 179 259 192
rect 184 163 238 179
rect 254 163 259 179
rect 80 127 96 158
rect 184 157 259 163
rect 277 139 298 214
rect 322 311 348 356
rect 322 295 327 311
rect 343 295 348 311
rect 322 270 348 295
rect 322 254 327 270
rect 343 254 348 270
rect 322 233 348 254
rect 322 217 327 233
rect 343 217 348 233
rect 322 212 348 217
rect 13 122 39 127
rect 13 106 18 122
rect 34 106 39 122
rect 13 22 39 106
rect 64 122 96 127
rect 64 106 69 122
rect 85 106 96 122
rect 271 121 298 139
rect 64 101 96 106
rect 115 116 245 120
rect 115 115 224 116
rect 115 99 120 115
rect 136 103 224 115
rect 136 99 141 103
rect 115 81 141 99
rect 218 100 224 103
rect 240 100 245 116
rect 271 105 276 121
rect 292 105 298 121
rect 271 100 298 105
rect 320 115 348 120
rect 115 65 121 81
rect 137 65 141 81
rect 115 50 141 65
rect 168 80 194 85
rect 168 64 173 80
rect 189 64 194 80
rect 168 22 194 64
rect 218 82 245 100
rect 218 66 224 82
rect 240 76 245 82
rect 320 99 327 115
rect 343 99 348 115
rect 320 81 348 99
rect 320 76 327 81
rect 240 66 327 76
rect 218 65 327 66
rect 343 65 348 81
rect 218 53 348 65
rect 0 8 384 22
rect 0 -8 16 8
rect 32 -8 64 8
rect 80 -8 112 8
rect 128 -8 160 8
rect 176 -8 208 8
rect 224 -8 256 8
rect 272 -8 304 8
rect 320 -8 352 8
rect 368 -8 384 8
rect 0 -22 384 -8
<< labels >>
flabel metal1 s 15 147 61 186 0 FreeSans 200 0 0 0 A_N
port 2 nsew
flabel metal1 s 276 214 298 318 0 FreeSans 200 0 0 0 Y
port 3 nsew
flabel metal1 s 0 356 384 400 0 FreeSans 200 0 0 0 VDD
port 4 nsew
flabel metal1 s 0 -22 384 22 0 FreeSans 200 0 0 0 VSS
port 5 nsew
flabel metal1 s 184 157 259 192 0 FreeSans 200 0 0 0 B
port 6 nsew
<< properties >>
string FIXED_BBOX 0 0 384 378
string GDS_END 220936
string GDS_FILE ../gds/controller.gds
string GDS_START 215392
<< end >>
