magic
tech ihp-sg13g2
magscale 1 2
timestamp 1747537721
<< nwell >>
rect -48 350 528 834
<< pwell >>
rect 206 232 421 270
rect -4 56 421 232
rect -26 -56 506 56
<< nmos >>
rect 90 96 116 206
rect 192 96 218 206
rect 301 96 327 244
<< pmos >>
rect 90 492 116 660
rect 192 492 218 660
rect 301 436 327 660
<< ndiff >>
rect 232 210 301 244
rect 232 206 247 210
rect 22 192 90 206
rect 22 160 36 192
rect 68 160 90 192
rect 22 96 90 160
rect 116 192 192 206
rect 116 160 138 192
rect 170 160 192 192
rect 116 96 192 160
rect 218 178 247 206
rect 279 178 301 210
rect 218 142 301 178
rect 218 110 244 142
rect 276 110 301 142
rect 218 96 301 110
rect 327 230 395 244
rect 327 198 349 230
rect 381 198 395 230
rect 327 142 395 198
rect 327 110 349 142
rect 381 110 395 142
rect 327 96 395 110
<< pdiff >>
rect 22 646 90 660
rect 22 614 36 646
rect 68 614 90 646
rect 22 538 90 614
rect 22 506 36 538
rect 68 506 90 538
rect 22 492 90 506
rect 116 492 192 660
rect 218 646 301 660
rect 218 614 244 646
rect 276 614 301 646
rect 218 567 301 614
rect 218 535 244 567
rect 276 535 301 567
rect 218 499 301 535
rect 218 492 246 499
rect 232 467 246 492
rect 278 467 301 499
rect 232 436 301 467
rect 327 646 398 660
rect 327 614 350 646
rect 382 614 398 646
rect 327 567 398 614
rect 327 535 350 567
rect 382 535 398 567
rect 327 482 398 535
rect 327 450 350 482
rect 382 450 398 482
rect 327 436 398 450
<< ndiffc >>
rect 36 160 68 192
rect 138 160 170 192
rect 247 178 279 210
rect 244 110 276 142
rect 349 198 381 230
rect 349 110 381 142
<< pdiffc >>
rect 36 614 68 646
rect 36 506 68 538
rect 244 614 276 646
rect 244 535 276 567
rect 246 467 278 499
rect 350 614 382 646
rect 350 535 382 567
rect 350 450 382 482
<< psubdiff >>
rect 0 16 480 30
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 480 16
rect 0 -30 480 -16
<< nsubdiff >>
rect 0 772 480 786
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 480 772
rect 0 726 480 740
<< psubdiffcont >>
rect 32 -16 64 16
rect 128 -16 160 16
rect 224 -16 256 16
rect 320 -16 352 16
rect 416 -16 448 16
<< nsubdiffcont >>
rect 32 740 64 772
rect 128 740 160 772
rect 224 740 256 772
rect 320 740 352 772
rect 416 740 448 772
<< poly >>
rect 90 660 116 704
rect 192 660 218 705
rect 301 660 327 706
rect 90 478 116 492
rect 90 464 156 478
rect 90 432 109 464
rect 141 432 156 464
rect 90 418 156 432
rect 90 206 116 418
rect 192 383 218 492
rect 169 369 229 383
rect 169 337 183 369
rect 215 337 229 369
rect 169 323 229 337
rect 192 206 218 323
rect 301 320 327 436
rect 271 306 334 320
rect 271 274 286 306
rect 318 274 334 306
rect 271 258 334 274
rect 301 244 327 258
rect 90 44 116 96
rect 192 44 218 96
rect 301 44 327 96
<< polycont >>
rect 109 432 141 464
rect 183 337 215 369
rect 286 274 318 306
<< metal1 >>
rect 0 772 480 800
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 480 772
rect 0 712 480 740
rect 236 646 288 712
rect 26 614 36 646
rect 68 614 78 646
rect 26 538 78 614
rect 26 506 36 538
rect 68 506 78 538
rect 234 614 244 646
rect 276 614 288 646
rect 234 567 288 614
rect 234 535 244 567
rect 276 535 288 567
rect 26 279 63 506
rect 130 470 181 530
rect 99 464 181 470
rect 99 432 109 464
rect 141 432 181 464
rect 234 499 288 535
rect 234 467 246 499
rect 278 467 288 499
rect 234 450 288 467
rect 340 614 350 646
rect 382 614 392 646
rect 340 567 392 614
rect 340 535 350 567
rect 382 535 392 567
rect 340 482 392 535
rect 340 450 350 482
rect 382 450 392 482
rect 99 426 181 432
rect 143 369 227 389
rect 143 337 183 369
rect 215 337 227 369
rect 143 315 227 337
rect 271 306 323 316
rect 271 279 286 306
rect 26 274 286 279
rect 318 274 323 306
rect 26 263 323 274
rect 26 246 304 263
rect 26 232 180 246
rect 128 192 180 232
rect 359 230 391 450
rect 26 160 36 192
rect 68 160 78 192
rect 128 160 138 192
rect 170 160 180 192
rect 237 178 247 210
rect 279 178 289 210
rect 26 44 78 160
rect 237 142 289 178
rect 237 110 244 142
rect 276 110 289 142
rect 339 198 349 230
rect 381 198 391 230
rect 339 142 391 198
rect 339 110 349 142
rect 381 110 391 142
rect 237 44 289 110
rect 0 16 480 44
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 480 16
rect 0 -44 480 -16
<< labels >>
flabel metal1 s 143 315 227 389 0 FreeSans 400 0 0 0 A
port 2 nsew
flabel metal1 s 0 -44 480 44 0 FreeSans 400 0 0 0 VSS
port 3 nsew
flabel metal1 s 130 426 181 530 0 FreeSans 400 0 0 0 B
port 4 nsew
flabel metal1 s 359 230 391 450 0 FreeSans 400 0 0 0 X
port 5 nsew
flabel metal1 s 0 712 480 800 0 FreeSans 400 0 0 0 VDD
port 6 nsew
<< properties >>
string FIXED_BBOX 0 0 480 756
string GDS_END 65488
string GDS_FILE ../gds/controller.gds
string GDS_START 61194
<< end >>
