magic
tech ihp-sg13g2
magscale 1 2
timestamp 1746816402
<< nwell >>
rect -60 374 2556 834
rect -60 350 319 374
rect 669 368 2556 374
rect 1153 350 2556 368
rect 1153 329 1551 350
<< pwell >>
rect 353 272 669 327
rect 1193 272 1322 293
rect 353 271 1322 272
rect 353 232 1408 271
rect 50 227 1408 232
rect 1879 227 2441 292
rect 50 56 2441 227
rect -26 -56 2522 56
<< nmos >>
rect 144 122 170 206
rect 218 122 244 206
rect 447 153 473 301
rect 549 153 575 301
rect 800 162 826 246
rect 902 162 928 246
rect 980 162 1006 246
rect 1052 162 1078 246
rect 1176 117 1202 245
rect 1310 117 1336 245
rect 1504 117 1530 201
rect 1582 117 1608 201
rect 1694 117 1720 201
rect 1765 117 1791 201
rect 1973 118 1999 266
rect 2213 118 2239 228
rect 2321 118 2347 266
<< pmos >>
rect 135 552 161 636
rect 237 552 263 636
rect 441 436 467 636
rect 543 436 569 636
rect 775 507 801 591
rect 877 507 903 591
rect 952 507 978 591
rect 1067 507 1093 591
rect 1303 391 1329 591
rect 1405 391 1431 591
rect 1535 515 1561 599
rect 1602 515 1628 599
rect 1704 515 1730 599
rect 1806 515 1832 599
rect 1918 412 1944 636
rect 2213 468 2239 636
rect 2315 412 2341 636
<< ndiff >>
rect 379 232 447 301
rect 76 179 144 206
rect 76 147 90 179
rect 122 147 144 179
rect 76 122 144 147
rect 170 122 218 206
rect 244 179 312 206
rect 244 147 266 179
rect 298 147 312 179
rect 379 200 393 232
rect 425 200 447 232
rect 379 153 447 200
rect 473 197 549 301
rect 473 165 495 197
rect 527 165 549 197
rect 473 153 549 165
rect 575 199 643 301
rect 575 167 597 199
rect 629 167 643 199
rect 575 153 643 167
rect 732 221 800 246
rect 732 189 746 221
rect 778 189 800 221
rect 732 162 800 189
rect 826 221 902 246
rect 826 189 848 221
rect 880 189 902 221
rect 826 162 902 189
rect 928 162 980 246
rect 1006 162 1052 246
rect 1078 245 1142 246
rect 1219 245 1296 267
rect 1078 162 1176 245
rect 244 122 312 147
rect 487 130 535 153
rect 1092 126 1176 162
rect 1092 94 1106 126
rect 1138 117 1176 126
rect 1202 218 1310 245
rect 1202 186 1256 218
rect 1288 186 1310 218
rect 1202 117 1310 186
rect 1336 201 1382 245
rect 1336 172 1504 201
rect 1336 140 1442 172
rect 1474 140 1504 172
rect 1336 117 1504 140
rect 1530 117 1582 201
rect 1608 170 1694 201
rect 1608 138 1636 170
rect 1668 138 1694 170
rect 1608 117 1694 138
rect 1720 117 1765 201
rect 1791 175 1859 201
rect 1791 143 1813 175
rect 1845 143 1859 175
rect 1791 117 1859 143
rect 1905 164 1973 266
rect 1905 132 1919 164
rect 1951 132 1973 164
rect 1905 118 1973 132
rect 1999 252 2074 266
rect 1999 220 2028 252
rect 2060 220 2074 252
rect 2253 252 2321 266
rect 2253 228 2267 252
rect 1999 164 2074 220
rect 1999 132 2028 164
rect 2060 132 2074 164
rect 1999 118 2074 132
rect 2145 187 2213 228
rect 2145 155 2159 187
rect 2191 155 2213 187
rect 2145 118 2213 155
rect 2239 220 2267 228
rect 2299 220 2321 252
rect 2239 165 2321 220
rect 2239 133 2267 165
rect 2299 133 2321 165
rect 2239 118 2321 133
rect 2347 252 2415 266
rect 2347 220 2369 252
rect 2401 220 2415 252
rect 2347 164 2415 220
rect 2347 132 2369 164
rect 2401 132 2415 164
rect 2347 118 2415 132
rect 1138 94 1161 117
rect 1092 79 1161 94
<< pdiff >>
rect 67 609 135 636
rect 67 577 81 609
rect 113 577 135 609
rect 67 552 135 577
rect 161 609 237 636
rect 161 577 183 609
rect 215 577 237 609
rect 161 552 237 577
rect 263 622 331 636
rect 263 590 285 622
rect 317 590 331 622
rect 263 552 331 590
rect 373 482 441 636
rect 373 450 387 482
rect 419 450 441 482
rect 373 436 441 450
rect 467 620 543 636
rect 467 588 489 620
rect 521 588 543 620
rect 467 436 543 588
rect 569 482 637 636
rect 569 450 591 482
rect 623 450 637 482
rect 569 436 637 450
rect 992 609 1053 623
rect 992 591 1006 609
rect 707 564 775 591
rect 707 532 721 564
rect 753 532 775 564
rect 707 507 775 532
rect 801 577 877 591
rect 801 545 823 577
rect 855 545 877 577
rect 801 507 877 545
rect 903 507 952 591
rect 978 577 1006 591
rect 1038 591 1053 609
rect 1846 609 1918 636
rect 1846 599 1860 609
rect 1482 591 1535 599
rect 1038 577 1067 591
rect 978 507 1067 577
rect 1093 562 1166 591
rect 1093 530 1119 562
rect 1151 530 1166 562
rect 1093 507 1166 530
rect 1235 577 1303 591
rect 1235 545 1249 577
rect 1281 545 1303 577
rect 1235 508 1303 545
rect 1235 476 1249 508
rect 1281 476 1303 508
rect 1235 440 1303 476
rect 1235 408 1249 440
rect 1281 408 1303 440
rect 1235 391 1303 408
rect 1329 577 1405 591
rect 1329 545 1351 577
rect 1383 545 1405 577
rect 1329 506 1405 545
rect 1329 474 1351 506
rect 1383 474 1405 506
rect 1329 437 1405 474
rect 1329 405 1351 437
rect 1383 405 1405 437
rect 1329 391 1405 405
rect 1431 565 1535 591
rect 1431 533 1461 565
rect 1493 533 1535 565
rect 1431 515 1535 533
rect 1561 515 1602 599
rect 1628 572 1704 599
rect 1628 540 1650 572
rect 1682 540 1704 572
rect 1628 515 1704 540
rect 1730 572 1806 599
rect 1730 540 1752 572
rect 1784 540 1806 572
rect 1730 515 1806 540
rect 1832 577 1860 599
rect 1892 577 1918 609
rect 1832 515 1918 577
rect 1431 391 1478 515
rect 1846 513 1918 515
rect 1846 481 1860 513
rect 1892 481 1918 513
rect 1846 412 1918 481
rect 1944 622 2080 636
rect 1944 590 1966 622
rect 1998 590 2034 622
rect 2066 590 2080 622
rect 1944 539 2080 590
rect 1944 507 1966 539
rect 1998 507 2034 539
rect 2066 507 2080 539
rect 1944 458 2080 507
rect 2145 621 2213 636
rect 2145 589 2159 621
rect 2191 589 2213 621
rect 2145 514 2213 589
rect 2145 482 2159 514
rect 2191 482 2213 514
rect 2145 468 2213 482
rect 2239 622 2315 636
rect 2239 590 2261 622
rect 2293 590 2315 622
rect 2239 539 2315 590
rect 2239 507 2261 539
rect 2293 507 2315 539
rect 2239 468 2315 507
rect 1944 426 1966 458
rect 1998 426 2034 458
rect 2066 426 2080 458
rect 1944 412 2080 426
rect 2255 412 2315 468
rect 2341 622 2409 636
rect 2341 590 2363 622
rect 2395 590 2409 622
rect 2341 539 2409 590
rect 2341 507 2363 539
rect 2395 507 2409 539
rect 2341 458 2409 507
rect 2341 426 2363 458
rect 2395 426 2409 458
rect 2341 412 2409 426
<< ndiffc >>
rect 90 147 122 179
rect 266 147 298 179
rect 393 200 425 232
rect 495 165 527 197
rect 597 167 629 199
rect 746 189 778 221
rect 848 189 880 221
rect 1106 94 1138 126
rect 1256 186 1288 218
rect 1442 140 1474 172
rect 1636 138 1668 170
rect 1813 143 1845 175
rect 1919 132 1951 164
rect 2028 220 2060 252
rect 2028 132 2060 164
rect 2159 155 2191 187
rect 2267 220 2299 252
rect 2267 133 2299 165
rect 2369 220 2401 252
rect 2369 132 2401 164
<< pdiffc >>
rect 81 577 113 609
rect 183 577 215 609
rect 285 590 317 622
rect 387 450 419 482
rect 489 588 521 620
rect 591 450 623 482
rect 721 532 753 564
rect 823 545 855 577
rect 1006 577 1038 609
rect 1119 530 1151 562
rect 1249 545 1281 577
rect 1249 476 1281 508
rect 1249 408 1281 440
rect 1351 545 1383 577
rect 1351 474 1383 506
rect 1351 405 1383 437
rect 1461 533 1493 565
rect 1650 540 1682 572
rect 1752 540 1784 572
rect 1860 577 1892 609
rect 1860 481 1892 513
rect 1966 590 1998 622
rect 2034 590 2066 622
rect 1966 507 1998 539
rect 2034 507 2066 539
rect 2159 589 2191 621
rect 2159 482 2191 514
rect 2261 590 2293 622
rect 2261 507 2293 539
rect 1966 426 1998 458
rect 2034 426 2066 458
rect 2363 590 2395 622
rect 2363 507 2395 539
rect 2363 426 2395 458
<< psubdiff >>
rect 0 16 2496 30
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 608 16
rect 640 -16 704 16
rect 736 -16 800 16
rect 832 -16 896 16
rect 928 -16 992 16
rect 1024 -16 1088 16
rect 1120 -16 1184 16
rect 1216 -16 1280 16
rect 1312 -16 1376 16
rect 1408 -16 1472 16
rect 1504 -16 1568 16
rect 1600 -16 1664 16
rect 1696 -16 1760 16
rect 1792 -16 1856 16
rect 1888 -16 1952 16
rect 1984 -16 2048 16
rect 2080 -16 2144 16
rect 2176 -16 2240 16
rect 2272 -16 2336 16
rect 2368 -16 2432 16
rect 2464 -16 2496 16
rect 0 -30 2496 -16
<< nsubdiff >>
rect 0 772 2496 786
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 608 772
rect 640 740 704 772
rect 736 740 800 772
rect 832 740 896 772
rect 928 740 992 772
rect 1024 740 1088 772
rect 1120 740 1184 772
rect 1216 740 1280 772
rect 1312 740 1376 772
rect 1408 740 1472 772
rect 1504 740 1568 772
rect 1600 740 1664 772
rect 1696 740 1760 772
rect 1792 740 1856 772
rect 1888 740 1952 772
rect 1984 740 2048 772
rect 2080 740 2144 772
rect 2176 740 2240 772
rect 2272 740 2336 772
rect 2368 740 2432 772
rect 2464 740 2496 772
rect 0 726 2496 740
<< psubdiffcont >>
rect 32 -16 64 16
rect 128 -16 160 16
rect 224 -16 256 16
rect 320 -16 352 16
rect 416 -16 448 16
rect 512 -16 544 16
rect 608 -16 640 16
rect 704 -16 736 16
rect 800 -16 832 16
rect 896 -16 928 16
rect 992 -16 1024 16
rect 1088 -16 1120 16
rect 1184 -16 1216 16
rect 1280 -16 1312 16
rect 1376 -16 1408 16
rect 1472 -16 1504 16
rect 1568 -16 1600 16
rect 1664 -16 1696 16
rect 1760 -16 1792 16
rect 1856 -16 1888 16
rect 1952 -16 1984 16
rect 2048 -16 2080 16
rect 2144 -16 2176 16
rect 2240 -16 2272 16
rect 2336 -16 2368 16
rect 2432 -16 2464 16
<< nsubdiffcont >>
rect 32 740 64 772
rect 128 740 160 772
rect 224 740 256 772
rect 320 740 352 772
rect 416 740 448 772
rect 512 740 544 772
rect 608 740 640 772
rect 704 740 736 772
rect 800 740 832 772
rect 896 740 928 772
rect 992 740 1024 772
rect 1088 740 1120 772
rect 1184 740 1216 772
rect 1280 740 1312 772
rect 1376 740 1408 772
rect 1472 740 1504 772
rect 1568 740 1600 772
rect 1664 740 1696 772
rect 1760 740 1792 772
rect 1856 740 1888 772
rect 1952 740 1984 772
rect 2048 740 2080 772
rect 2144 740 2176 772
rect 2240 740 2272 772
rect 2336 740 2368 772
rect 2432 740 2464 772
<< poly >>
rect 135 636 161 672
rect 237 636 263 672
rect 441 636 467 672
rect 543 636 569 672
rect 651 663 1431 689
rect 135 537 161 552
rect 237 537 263 552
rect 128 514 164 537
rect 89 428 170 514
rect 89 396 105 428
rect 137 396 170 428
rect 89 360 170 396
rect 89 328 105 360
rect 137 328 170 360
rect 89 292 170 328
rect 89 260 105 292
rect 137 260 170 292
rect 89 244 170 260
rect 144 206 170 244
rect 218 472 270 537
rect 218 454 311 472
rect 218 422 261 454
rect 293 422 311 454
rect 218 386 311 422
rect 441 399 467 436
rect 543 399 569 436
rect 651 399 677 663
rect 775 591 801 627
rect 877 591 903 663
rect 1390 645 1431 663
rect 952 591 978 627
rect 1067 591 1093 627
rect 1303 591 1329 627
rect 1405 591 1431 645
rect 1918 636 1944 672
rect 2213 636 2239 672
rect 2315 636 2341 672
rect 1535 599 1561 635
rect 1602 599 1628 635
rect 1704 599 1730 635
rect 1806 599 1832 635
rect 775 486 801 507
rect 775 441 810 486
rect 877 471 903 507
rect 952 475 978 507
rect 1067 492 1093 507
rect 1062 475 1098 492
rect 952 457 1026 475
rect 952 445 976 457
rect 218 354 261 386
rect 293 354 311 386
rect 218 318 311 354
rect 425 381 496 399
rect 425 349 446 381
rect 478 349 496 381
rect 425 326 496 349
rect 543 371 677 399
rect 744 423 810 441
rect 744 391 760 423
rect 792 391 810 423
rect 744 386 810 391
rect 960 425 976 445
rect 1008 425 1026 457
rect 960 389 1026 425
rect 744 381 918 386
rect 746 379 918 381
rect 748 377 918 379
rect 750 375 918 377
rect 752 373 918 375
rect 754 371 918 373
rect 543 339 579 371
rect 611 358 677 371
rect 756 369 918 371
rect 758 367 918 369
rect 760 365 918 367
rect 762 363 918 365
rect 764 361 918 363
rect 766 359 918 361
rect 611 356 706 358
rect 768 356 918 359
rect 611 354 708 356
rect 611 352 710 354
rect 611 350 712 352
rect 611 348 714 350
rect 611 346 716 348
rect 611 344 718 346
rect 611 342 720 344
rect 611 340 722 342
rect 611 339 724 340
rect 543 338 724 339
rect 543 336 726 338
rect 543 326 729 336
rect 218 286 261 318
rect 293 286 311 318
rect 447 301 473 326
rect 549 325 729 326
rect 549 301 575 325
rect 692 324 729 325
rect 695 322 729 324
rect 697 320 729 322
rect 699 314 729 320
rect 218 270 311 286
rect 218 206 244 270
rect 699 284 826 314
rect 800 246 826 284
rect 888 292 918 356
rect 960 357 976 389
rect 1008 357 1026 389
rect 960 341 1026 357
rect 1062 457 1208 475
rect 1062 425 1162 457
rect 1194 425 1208 457
rect 1062 409 1208 425
rect 888 262 928 292
rect 902 246 928 262
rect 980 246 1006 341
rect 1062 292 1092 409
rect 1535 479 1561 515
rect 1497 465 1566 479
rect 1497 433 1511 465
rect 1543 433 1566 465
rect 1602 478 1628 515
rect 1602 444 1642 478
rect 1704 477 1730 515
rect 1497 417 1566 433
rect 1303 376 1329 391
rect 1300 367 1336 376
rect 1146 349 1336 367
rect 1146 317 1162 349
rect 1194 337 1336 349
rect 1405 369 1431 391
rect 1405 339 1530 369
rect 1194 317 1212 337
rect 1146 301 1212 317
rect 1052 262 1092 292
rect 1052 246 1078 262
rect 1176 245 1202 301
rect 1310 272 1462 291
rect 1310 261 1412 272
rect 1310 245 1336 261
rect 144 86 170 122
rect 218 73 244 122
rect 447 117 473 153
rect 549 117 575 153
rect 800 126 826 162
rect 902 126 928 162
rect 980 126 1006 162
rect 1052 73 1078 162
rect 1396 240 1412 261
rect 1444 240 1462 272
rect 1396 224 1462 240
rect 1504 201 1530 339
rect 1616 290 1642 444
rect 1689 459 1760 477
rect 1689 427 1703 459
rect 1735 427 1760 459
rect 1689 411 1760 427
rect 1582 272 1652 290
rect 1582 240 1602 272
rect 1634 240 1652 272
rect 1582 224 1652 240
rect 1582 201 1608 224
rect 1694 201 1720 411
rect 1806 363 1832 515
rect 1918 363 1944 412
rect 2213 363 2239 468
rect 2315 370 2341 412
rect 1766 345 2239 363
rect 1766 313 1782 345
rect 1814 313 2239 345
rect 1766 306 2239 313
rect 1765 297 2239 306
rect 2288 352 2354 370
rect 2288 320 2304 352
rect 2336 320 2354 352
rect 2288 304 2354 320
rect 1765 201 1791 297
rect 1973 266 1999 297
rect 2213 228 2239 297
rect 2321 266 2347 304
rect 1176 81 1202 117
rect 1310 81 1336 117
rect 1504 81 1530 117
rect 1582 81 1608 117
rect 1694 81 1720 117
rect 1765 81 1791 117
rect 1973 82 1999 118
rect 2213 82 2239 118
rect 2321 82 2347 118
rect 218 47 1078 73
<< polycont >>
rect 105 396 137 428
rect 105 328 137 360
rect 105 260 137 292
rect 261 422 293 454
rect 261 354 293 386
rect 446 349 478 381
rect 760 391 792 423
rect 976 425 1008 457
rect 579 339 611 371
rect 261 286 293 318
rect 976 357 1008 389
rect 1162 425 1194 457
rect 1511 433 1543 465
rect 1162 317 1194 349
rect 1412 240 1444 272
rect 1703 427 1735 459
rect 1602 240 1634 272
rect 1782 313 1814 345
rect 2304 320 2336 352
<< metal1 >>
rect 0 772 2496 800
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 608 772
rect 640 740 704 772
rect 736 740 800 772
rect 832 740 896 772
rect 928 740 992 772
rect 1024 740 1088 772
rect 1120 740 1184 772
rect 1216 740 1280 772
rect 1312 740 1376 772
rect 1408 740 1472 772
rect 1504 740 1568 772
rect 1600 740 1664 772
rect 1696 740 1760 772
rect 1792 740 1856 772
rect 1888 740 1952 772
rect 1984 740 2048 772
rect 2080 740 2144 772
rect 2176 740 2240 772
rect 2272 740 2336 772
rect 2368 740 2432 772
rect 2464 740 2496 772
rect 0 712 2496 740
rect 71 609 123 712
rect 275 622 327 712
rect 71 577 81 609
rect 113 577 123 609
rect 71 572 123 577
rect 173 609 225 619
rect 173 577 183 609
rect 215 577 225 609
rect 275 590 285 622
rect 317 590 327 622
rect 275 587 327 590
rect 479 620 531 712
rect 479 588 489 620
rect 521 588 531 620
rect 996 609 1048 712
rect 173 551 225 577
rect 711 564 764 582
rect 711 551 721 564
rect 173 532 721 551
rect 753 532 764 564
rect 809 577 936 583
rect 809 545 823 577
rect 855 545 936 577
rect 996 577 1006 609
rect 1038 577 1048 609
rect 996 575 1048 577
rect 1247 577 1283 712
rect 809 540 936 545
rect 173 525 764 532
rect 183 519 764 525
rect 88 428 147 483
rect 88 396 105 428
rect 137 396 147 428
rect 88 360 147 396
rect 88 328 105 360
rect 137 328 147 360
rect 88 292 147 328
rect 88 260 105 292
rect 137 260 147 292
rect 88 244 147 260
rect 183 190 215 519
rect 726 504 764 519
rect 904 539 936 540
rect 1105 562 1157 572
rect 1105 539 1119 562
rect 904 530 1119 539
rect 1151 530 1157 562
rect 904 507 1157 530
rect 1247 545 1249 577
rect 1281 545 1283 577
rect 1247 508 1283 545
rect 581 482 633 483
rect 251 454 305 472
rect 377 463 387 482
rect 251 442 261 454
rect 293 442 305 454
rect 251 402 260 442
rect 300 402 305 442
rect 251 386 305 402
rect 251 354 261 386
rect 293 354 305 386
rect 251 318 305 354
rect 251 286 261 318
rect 293 286 305 318
rect 251 270 305 286
rect 341 450 387 463
rect 419 450 429 482
rect 341 424 429 450
rect 581 450 591 482
rect 623 460 633 482
rect 726 472 868 504
rect 623 457 645 460
rect 623 456 649 457
rect 623 452 650 456
rect 623 450 655 452
rect 581 443 655 450
rect 581 434 703 443
rect 341 279 373 424
rect 581 423 800 434
rect 581 417 760 423
rect 628 409 760 417
rect 454 383 498 397
rect 409 381 498 383
rect 409 349 446 381
rect 478 349 498 381
rect 674 391 760 409
rect 792 391 800 423
rect 674 375 800 391
rect 409 315 498 349
rect 567 371 638 373
rect 567 339 579 371
rect 611 339 638 371
rect 567 329 638 339
rect 567 279 602 329
rect 674 294 706 375
rect 836 303 868 472
rect 341 247 602 279
rect 650 262 706 294
rect 753 271 868 303
rect 341 232 429 247
rect 341 204 393 232
rect 80 179 215 190
rect 355 200 393 204
rect 425 200 429 232
rect 650 211 683 262
rect 753 231 792 271
rect 904 235 936 507
rect 80 147 90 179
rect 122 152 215 179
rect 256 179 308 182
rect 122 147 132 152
rect 80 137 132 147
rect 256 147 266 179
rect 298 147 308 179
rect 355 163 429 200
rect 485 197 537 204
rect 485 165 495 197
rect 527 165 537 197
rect 256 44 308 147
rect 485 44 537 165
rect 584 199 683 211
rect 584 167 597 199
rect 629 167 683 199
rect 736 221 792 231
rect 736 189 746 221
rect 778 189 792 221
rect 736 179 792 189
rect 839 221 936 235
rect 972 457 1019 469
rect 972 425 976 457
rect 1008 425 1019 457
rect 972 389 1019 425
rect 972 357 976 389
rect 1008 357 1019 389
rect 972 262 1019 357
rect 1055 367 1087 507
rect 1247 476 1249 508
rect 1281 476 1283 508
rect 1123 465 1203 471
rect 1123 425 1132 465
rect 1172 457 1203 465
rect 1194 425 1203 457
rect 1123 409 1203 425
rect 1247 440 1283 476
rect 1247 408 1249 440
rect 1281 408 1283 440
rect 1247 398 1283 408
rect 1349 577 1385 587
rect 1349 545 1351 577
rect 1383 545 1385 577
rect 1349 506 1385 545
rect 1451 565 1613 575
rect 1451 533 1461 565
rect 1493 533 1613 565
rect 1451 523 1613 533
rect 1649 572 1683 712
rect 1850 609 1902 712
rect 1649 540 1650 572
rect 1682 540 1683 572
rect 1649 530 1683 540
rect 1742 572 1813 582
rect 1742 540 1752 572
rect 1784 540 1813 572
rect 1742 529 1813 540
rect 1349 474 1351 506
rect 1383 474 1385 506
rect 1349 437 1385 474
rect 1349 405 1351 437
rect 1383 405 1385 437
rect 1055 349 1206 367
rect 1349 358 1385 405
rect 1055 333 1162 349
rect 1148 317 1162 333
rect 1194 317 1206 349
rect 1148 301 1206 317
rect 1243 326 1385 358
rect 1428 465 1545 483
rect 1428 433 1511 465
rect 1543 433 1545 465
rect 1428 417 1545 433
rect 1243 262 1296 326
rect 1428 290 1460 417
rect 1581 363 1613 523
rect 1665 468 1745 477
rect 1665 428 1687 468
rect 1727 459 1745 468
rect 1665 427 1703 428
rect 1735 427 1745 459
rect 1665 411 1745 427
rect 1781 431 1813 529
rect 1850 577 1860 609
rect 1892 577 1902 609
rect 1850 513 1902 577
rect 1850 481 1860 513
rect 1892 481 1902 513
rect 1850 479 1902 481
rect 1958 622 2076 633
rect 1958 590 1966 622
rect 1998 590 2034 622
rect 2066 590 2076 622
rect 1958 539 2076 590
rect 1958 507 1966 539
rect 1998 507 2034 539
rect 2066 507 2076 539
rect 1958 458 2076 507
rect 1781 399 1920 431
rect 1958 426 1966 458
rect 1998 426 2034 458
rect 2066 426 2076 458
rect 1958 416 2076 426
rect 2149 621 2201 627
rect 2149 589 2159 621
rect 2191 589 2201 621
rect 2149 514 2201 589
rect 2149 482 2159 514
rect 2191 482 2201 514
rect 2251 622 2303 712
rect 2251 590 2261 622
rect 2293 590 2303 622
rect 2251 539 2303 590
rect 2251 507 2261 539
rect 2293 507 2303 539
rect 2251 504 2303 507
rect 2357 622 2429 632
rect 2357 590 2363 622
rect 2395 590 2429 622
rect 2357 539 2429 590
rect 2357 507 2363 539
rect 2395 507 2429 539
rect 972 230 1296 262
rect 839 189 848 221
rect 880 189 936 221
rect 1253 218 1296 230
rect 839 178 936 189
rect 584 153 683 167
rect 650 127 683 153
rect 1001 162 1216 194
rect 1253 186 1256 218
rect 1288 186 1296 218
rect 1253 176 1296 186
rect 1359 272 1460 290
rect 1359 240 1412 272
rect 1444 240 1460 272
rect 1359 224 1460 240
rect 1520 345 1824 363
rect 1520 329 1782 345
rect 1001 127 1038 162
rect 650 95 1038 127
rect 1184 139 1216 162
rect 1359 139 1393 224
rect 1520 177 1554 329
rect 1770 313 1782 329
rect 1814 313 1824 345
rect 1770 300 1824 313
rect 1592 272 1644 275
rect 1592 240 1602 272
rect 1634 258 1644 272
rect 1887 258 1920 399
rect 1634 240 1920 258
rect 1592 224 1920 240
rect 2018 252 2070 416
rect 1096 94 1106 126
rect 1138 94 1148 126
rect 1184 106 1393 139
rect 1432 172 1554 177
rect 1803 175 1855 224
rect 1432 140 1442 172
rect 1474 140 1554 172
rect 1432 134 1554 140
rect 1626 170 1678 175
rect 1626 138 1636 170
rect 1668 138 1678 170
rect 1096 44 1148 94
rect 1626 44 1678 138
rect 1803 143 1813 175
rect 1845 143 1855 175
rect 2018 220 2028 252
rect 2060 220 2070 252
rect 1803 133 1855 143
rect 1909 164 1961 172
rect 1909 132 1919 164
rect 1951 132 1961 164
rect 1909 44 1961 132
rect 2018 164 2070 220
rect 2018 132 2028 164
rect 2060 132 2070 164
rect 2149 370 2201 482
rect 2357 458 2429 507
rect 2357 426 2363 458
rect 2395 426 2429 458
rect 2357 416 2429 426
rect 2149 352 2354 370
rect 2149 320 2304 352
rect 2336 320 2354 352
rect 2149 304 2354 320
rect 2149 187 2202 304
rect 2395 256 2429 416
rect 2149 155 2159 187
rect 2191 155 2202 187
rect 2149 141 2202 155
rect 2257 252 2309 254
rect 2257 220 2267 252
rect 2299 220 2309 252
rect 2257 165 2309 220
rect 2018 121 2070 132
rect 2257 133 2267 165
rect 2299 133 2309 165
rect 2257 44 2309 133
rect 2355 252 2429 256
rect 2355 220 2369 252
rect 2401 220 2429 252
rect 2355 164 2429 220
rect 2355 132 2369 164
rect 2401 132 2429 164
rect 2355 129 2429 132
rect 0 16 2496 44
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 608 16
rect 640 -16 704 16
rect 736 -16 800 16
rect 832 -16 896 16
rect 928 -16 992 16
rect 1024 -16 1088 16
rect 1120 -16 1184 16
rect 1216 -16 1280 16
rect 1312 -16 1376 16
rect 1408 -16 1472 16
rect 1504 -16 1568 16
rect 1600 -16 1664 16
rect 1696 -16 1760 16
rect 1792 -16 1856 16
rect 1888 -16 1952 16
rect 1984 -16 2048 16
rect 2080 -16 2144 16
rect 2176 -16 2240 16
rect 2272 -16 2336 16
rect 2368 -16 2432 16
rect 2464 -16 2496 16
rect 0 -44 2496 -16
<< via1 >>
rect 260 422 261 442
rect 261 422 293 442
rect 293 422 300 442
rect 260 402 300 422
rect 1132 457 1172 465
rect 1132 425 1162 457
rect 1162 425 1172 457
rect 1687 459 1727 468
rect 1687 428 1703 459
rect 1703 428 1727 459
<< metal2 >>
rect 256 442 314 474
rect 256 402 260 442
rect 300 440 314 442
rect 1120 465 1178 474
rect 1120 440 1132 465
rect 300 425 1132 440
rect 1172 440 1178 465
rect 1655 468 1745 474
rect 1655 440 1687 468
rect 1172 428 1687 440
rect 1727 428 1745 468
rect 1172 425 1745 428
rect 300 402 1745 425
rect 256 400 1745 402
rect 256 393 314 400
<< labels >>
flabel metal2 s 256 393 314 474 0 FreeSans 400 0 0 0 RESET_B
port 1 nsew
flabel metal1 s 88 244 147 483 0 FreeSans 400 0 0 0 D
port 3 nsew
flabel metal1 s 1958 416 2076 633 0 FreeSans 400 0 0 0 Q_N
port 4 nsew
flabel metal1 s 409 315 498 383 0 FreeSans 400 0 0 0 CLK
port 5 nsew
flabel metal1 s 0 -44 2496 44 0 FreeSans 400 0 0 0 VSS
port 6 nsew
flabel metal1 s 0 712 2496 800 0 FreeSans 400 0 0 0 VDD
port 7 nsew
flabel metal1 s 2357 421 2429 627 0 FreeSans 400 0 0 0 Q
port 8 nsew
<< properties >>
string FIXED_BBOX 0 0 2496 756
string GDS_END 59514
string GDS_FILE ../gds/controller.gds
string GDS_START 43598
<< end >>
