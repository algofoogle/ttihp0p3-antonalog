magic
tech ihp-sg13g2
magscale 1 2
timestamp 1746816402
<< nwell >>
rect -48 350 624 834
<< pwell >>
rect 30 241 539 292
rect 30 56 550 241
rect -26 -56 602 56
<< nmos >>
rect 124 118 150 266
rect 226 118 252 266
rect 328 118 354 266
rect 430 118 456 266
<< pmos >>
rect 124 412 150 636
rect 208 412 234 636
rect 322 412 348 636
rect 436 412 462 636
<< ndiff >>
rect 56 241 124 266
rect 56 209 70 241
rect 102 209 124 241
rect 56 165 124 209
rect 56 133 70 165
rect 102 133 124 165
rect 56 118 124 133
rect 150 250 226 266
rect 150 218 172 250
rect 204 218 226 250
rect 150 165 226 218
rect 150 133 172 165
rect 204 133 226 165
rect 150 118 226 133
rect 252 195 328 266
rect 252 163 274 195
rect 306 163 328 195
rect 252 118 328 163
rect 354 251 430 266
rect 354 219 376 251
rect 408 219 430 251
rect 354 165 430 219
rect 354 133 376 165
rect 408 133 430 165
rect 354 118 430 133
rect 456 215 513 266
rect 456 186 524 215
rect 456 154 478 186
rect 510 154 524 186
rect 456 118 524 154
<< pdiff >>
rect 56 621 124 636
rect 56 589 70 621
rect 102 589 124 621
rect 56 540 124 589
rect 56 508 70 540
rect 102 508 124 540
rect 56 459 124 508
rect 56 427 70 459
rect 102 427 124 459
rect 56 412 124 427
rect 150 412 208 636
rect 234 412 322 636
rect 348 412 436 636
rect 462 621 534 636
rect 462 589 488 621
rect 520 589 534 621
rect 462 553 534 589
rect 462 521 488 553
rect 520 521 534 553
rect 462 483 534 521
rect 462 451 488 483
rect 520 451 534 483
rect 462 412 534 451
<< ndiffc >>
rect 70 209 102 241
rect 70 133 102 165
rect 172 218 204 250
rect 172 133 204 165
rect 274 163 306 195
rect 376 219 408 251
rect 376 133 408 165
rect 478 154 510 186
<< pdiffc >>
rect 70 589 102 621
rect 70 508 102 540
rect 70 427 102 459
rect 488 589 520 621
rect 488 521 520 553
rect 488 451 520 483
<< psubdiff >>
rect 0 16 576 30
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 576 16
rect 0 -30 576 -16
<< nsubdiff >>
rect 0 772 576 786
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 576 772
rect 0 726 576 740
<< psubdiffcont >>
rect 32 -16 64 16
rect 128 -16 160 16
rect 224 -16 256 16
rect 320 -16 352 16
rect 416 -16 448 16
rect 512 -16 544 16
<< nsubdiffcont >>
rect 32 740 64 772
rect 128 740 160 772
rect 224 740 256 772
rect 320 740 352 772
rect 416 740 448 772
rect 512 740 544 772
<< poly >>
rect 124 636 150 672
rect 208 636 234 672
rect 322 636 348 672
rect 436 636 462 672
rect 124 397 150 412
rect 208 397 234 412
rect 322 397 348 412
rect 436 397 462 412
rect 121 354 150 397
rect 52 337 150 354
rect 52 305 69 337
rect 101 305 150 337
rect 187 380 241 397
rect 187 363 252 380
rect 187 331 204 363
rect 236 331 252 363
rect 187 314 252 331
rect 288 363 354 397
rect 288 331 305 363
rect 337 331 354 363
rect 288 314 354 331
rect 390 363 469 397
rect 390 331 417 363
rect 449 331 469 363
rect 390 314 469 331
rect 52 288 150 305
rect 124 266 150 288
rect 226 266 252 314
rect 328 266 354 314
rect 430 266 456 314
rect 124 82 150 118
rect 226 82 252 118
rect 328 82 354 118
rect 430 82 456 118
<< polycont >>
rect 69 305 101 337
rect 204 331 236 363
rect 305 331 337 363
rect 417 331 449 363
<< metal1 >>
rect 0 772 576 800
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 576 772
rect 0 712 576 740
rect 60 621 112 712
rect 60 589 70 621
rect 102 589 112 621
rect 60 540 112 589
rect 60 508 70 540
rect 102 508 112 540
rect 60 459 112 508
rect 60 427 70 459
rect 102 427 112 459
rect 60 424 112 427
rect 39 337 126 366
rect 39 305 69 337
rect 101 305 126 337
rect 167 363 252 622
rect 445 621 540 640
rect 445 589 488 621
rect 520 589 540 621
rect 445 553 540 589
rect 445 521 488 553
rect 520 521 540 553
rect 445 483 540 521
rect 167 331 204 363
rect 236 331 252 363
rect 167 314 252 331
rect 288 363 348 474
rect 445 451 488 483
rect 520 451 540 483
rect 445 434 540 451
rect 288 331 305 363
rect 337 331 348 363
rect 288 314 348 331
rect 390 363 464 396
rect 390 331 417 363
rect 449 331 464 363
rect 390 314 464 331
rect 39 283 126 305
rect 501 278 540 434
rect 162 251 540 278
rect 162 250 376 251
rect 58 241 112 246
rect 58 209 70 241
rect 102 209 112 241
rect 58 165 112 209
rect 58 133 70 165
rect 102 133 112 165
rect 58 44 112 133
rect 162 218 172 250
rect 204 235 376 250
rect 204 218 214 235
rect 162 165 214 218
rect 366 219 376 235
rect 408 235 540 251
rect 408 219 418 235
rect 162 133 172 165
rect 204 133 214 165
rect 162 129 214 133
rect 264 195 316 199
rect 264 163 274 195
rect 306 163 316 195
rect 264 44 316 163
rect 366 165 418 219
rect 366 133 376 165
rect 408 133 418 165
rect 366 129 418 133
rect 468 186 520 193
rect 468 154 478 186
rect 510 154 520 186
rect 468 44 520 154
rect 0 16 576 44
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 576 16
rect 0 -44 576 -16
<< labels >>
flabel metal1 s 0 -44 576 44 0 FreeSans 400 0 0 0 VSS
port 2 nsew
flabel metal1 s 0 712 576 800 0 FreeSans 400 0 0 0 VDD
port 3 nsew
flabel metal1 s 167 314 252 622 0 FreeSans 400 0 0 0 B
port 4 nsew
flabel metal1 s 288 314 348 474 0 FreeSans 400 0 0 0 C
port 5 nsew
flabel metal1 s 445 434 540 640 0 FreeSans 400 0 0 0 Y
port 6 nsew
flabel metal1 s 39 283 126 366 0 FreeSans 400 0 0 0 A
port 7 nsew
flabel metal1 s 390 314 464 396 0 FreeSans 400 0 0 0 D
port 8 nsew
<< properties >>
string FIXED_BBOX 0 0 576 756
string GDS_END 190504
string GDS_FILE ../gds/controller.gds
string GDS_START 185062
<< end >>
