magic
tech ihp-sg13g2
timestamp 1747537721
<< nwell >>
rect -24 175 216 417
<< pwell >>
rect 2 28 193 144
rect -13 -28 205 28
<< nmos >>
rect 75 76 88 131
rect 133 57 146 131
<< pmos >>
rect 76 234 89 318
rect 129 206 142 318
<< ndiff >>
rect 15 123 75 131
rect 15 107 46 123
rect 62 107 75 123
rect 15 100 75 107
rect 48 76 75 100
rect 88 97 133 131
rect 88 81 102 97
rect 118 81 133 97
rect 88 76 133 81
rect 95 57 133 76
rect 146 122 180 131
rect 146 106 157 122
rect 173 106 180 122
rect 146 81 180 106
rect 146 65 157 81
rect 173 65 180 81
rect 146 57 180 65
<< pdiff >>
rect 40 310 76 318
rect 40 294 47 310
rect 63 294 76 310
rect 40 275 76 294
rect 40 259 47 275
rect 63 259 76 275
rect 40 234 76 259
rect 89 310 129 318
rect 89 294 101 310
rect 117 294 129 310
rect 89 234 129 294
rect 103 206 129 234
rect 142 310 178 318
rect 142 294 155 310
rect 171 294 178 310
rect 142 270 178 294
rect 142 254 155 270
rect 171 254 178 270
rect 142 232 178 254
rect 142 216 155 232
rect 171 216 178 232
rect 142 206 178 216
<< ndiffc >>
rect 46 107 62 123
rect 102 81 118 97
rect 157 106 173 122
rect 157 65 173 81
<< pdiffc >>
rect 47 294 63 310
rect 47 259 63 275
rect 101 294 117 310
rect 155 294 171 310
rect 155 254 171 270
rect 155 216 171 232
<< psubdiff >>
rect 0 8 192 15
rect 0 -8 16 8
rect 32 -8 64 8
rect 80 -8 112 8
rect 128 -8 160 8
rect 176 -8 192 8
rect 0 -15 192 -8
<< nsubdiff >>
rect 0 386 192 393
rect 0 370 16 386
rect 32 370 64 386
rect 80 370 112 386
rect 128 370 160 386
rect 176 370 192 386
rect 0 363 192 370
<< psubdiffcont >>
rect 16 -8 32 8
rect 64 -8 80 8
rect 112 -8 128 8
rect 160 -8 176 8
<< nsubdiffcont >>
rect 16 370 32 386
rect 64 370 80 386
rect 112 370 128 386
rect 160 370 176 386
<< poly >>
rect 76 318 89 336
rect 129 318 142 336
rect 76 224 89 234
rect 73 207 91 224
rect 73 198 88 207
rect 20 189 88 198
rect 129 196 142 206
rect 20 173 28 189
rect 44 173 62 189
rect 78 173 88 189
rect 128 183 146 196
rect 20 165 88 173
rect 75 131 88 165
rect 112 174 146 183
rect 112 158 120 174
rect 136 158 146 174
rect 112 150 146 158
rect 133 131 146 150
rect 75 58 88 76
rect 133 39 146 57
<< polycont >>
rect 28 173 44 189
rect 62 173 78 189
rect 120 158 136 174
<< metal1 >>
rect 0 386 192 400
rect 0 370 16 386
rect 32 370 64 386
rect 80 370 112 386
rect 128 370 160 386
rect 176 370 192 386
rect 0 356 192 370
rect 43 310 70 318
rect 43 294 47 310
rect 63 294 70 310
rect 43 275 70 294
rect 94 310 124 356
rect 94 294 101 310
rect 117 294 124 310
rect 94 284 124 294
rect 149 310 179 318
rect 149 294 155 310
rect 171 294 179 310
rect 43 259 47 275
rect 63 262 70 275
rect 149 270 179 294
rect 63 259 126 262
rect 43 244 126 259
rect 10 189 87 211
rect 10 173 28 189
rect 44 173 62 189
rect 78 173 87 189
rect 10 165 87 173
rect 109 183 126 244
rect 149 254 155 270
rect 171 254 179 270
rect 149 232 179 254
rect 149 216 155 232
rect 171 216 179 232
rect 149 202 179 216
rect 109 174 141 183
rect 109 158 120 174
rect 136 158 141 174
rect 109 150 141 158
rect 109 146 126 150
rect 31 129 126 146
rect 160 129 179 202
rect 31 123 70 129
rect 31 107 46 123
rect 62 107 70 123
rect 31 100 70 107
rect 150 122 179 129
rect 150 106 157 122
rect 173 106 179 122
rect 93 97 126 102
rect 93 81 102 97
rect 118 81 126 97
rect 93 22 126 81
rect 150 81 179 106
rect 150 65 157 81
rect 173 65 179 81
rect 150 55 179 65
rect 0 8 192 22
rect 0 -8 16 8
rect 32 -8 64 8
rect 80 -8 112 8
rect 128 -8 160 8
rect 176 -8 192 8
rect 0 -22 192 -8
<< labels >>
flabel metal1 s 0 -22 192 22 0 FreeSans 200 0 0 0 VSS
port 3 nsew
flabel metal1 s 0 356 192 400 0 FreeSans 200 0 0 0 VDD
port 2 nsew
<< properties >>
string FIXED_BBOX 0 0 192 378
string GDS_END 186940
string GDS_FILE ../gds/controller.gds
string GDS_START 183652
<< end >>
