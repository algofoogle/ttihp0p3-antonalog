magic
tech ihp-sg13g2
magscale 1 2
timestamp 1747537721
<< nwell >>
rect -48 350 912 834
<< pwell >>
rect 412 228 810 292
rect 30 56 810 228
rect -26 -56 890 56
<< nmos >>
rect 124 118 150 202
rect 226 118 326 202
rect 506 182 606 266
rect 690 118 716 266
<< pmos >>
rect 124 511 150 595
rect 226 436 326 636
rect 506 412 606 612
rect 688 412 714 636
<< ndiff >>
rect 438 234 506 266
rect 438 202 452 234
rect 484 202 506 234
rect 56 175 124 202
rect 56 143 70 175
rect 102 143 124 175
rect 56 118 124 143
rect 150 164 226 202
rect 150 132 172 164
rect 204 132 226 164
rect 150 118 226 132
rect 326 175 394 202
rect 438 182 506 202
rect 606 182 690 266
rect 326 143 348 175
rect 380 143 394 175
rect 622 165 690 182
rect 326 118 394 143
rect 622 133 636 165
rect 668 133 690 165
rect 622 118 690 133
rect 716 250 784 266
rect 716 218 738 250
rect 770 218 784 250
rect 716 164 784 218
rect 716 132 738 164
rect 770 132 784 164
rect 716 118 784 132
<< pdiff >>
rect 176 595 226 636
rect 56 571 124 595
rect 56 539 70 571
rect 102 539 124 571
rect 56 511 124 539
rect 150 568 226 595
rect 150 536 172 568
rect 204 536 226 568
rect 150 511 226 536
rect 176 436 226 511
rect 326 571 394 636
rect 620 621 688 636
rect 620 612 634 621
rect 326 539 348 571
rect 380 539 394 571
rect 326 436 394 539
rect 438 464 506 612
rect 438 432 452 464
rect 484 432 506 464
rect 438 412 506 432
rect 606 589 634 612
rect 666 589 688 621
rect 606 513 688 589
rect 606 481 630 513
rect 662 481 688 513
rect 606 412 688 481
rect 714 621 790 636
rect 714 589 744 621
rect 776 589 790 621
rect 714 545 790 589
rect 714 513 744 545
rect 776 513 790 545
rect 714 458 790 513
rect 714 426 744 458
rect 776 426 790 458
rect 714 412 790 426
<< ndiffc >>
rect 452 202 484 234
rect 70 143 102 175
rect 172 132 204 164
rect 348 143 380 175
rect 636 133 668 165
rect 738 218 770 250
rect 738 132 770 164
<< pdiffc >>
rect 70 539 102 571
rect 172 536 204 568
rect 348 539 380 571
rect 452 432 484 464
rect 634 589 666 621
rect 630 481 662 513
rect 744 589 776 621
rect 744 513 776 545
rect 744 426 776 458
<< psubdiff >>
rect 0 16 864 30
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 608 16
rect 640 -16 704 16
rect 736 -16 800 16
rect 832 -16 864 16
rect 0 -30 864 -16
<< nsubdiff >>
rect 0 772 864 786
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 608 772
rect 640 740 704 772
rect 736 740 800 772
rect 832 740 864 772
rect 0 726 864 740
<< psubdiffcont >>
rect 32 -16 64 16
rect 128 -16 160 16
rect 224 -16 256 16
rect 320 -16 352 16
rect 416 -16 448 16
rect 512 -16 544 16
rect 608 -16 640 16
rect 704 -16 736 16
rect 800 -16 832 16
<< nsubdiffcont >>
rect 32 740 64 772
rect 128 740 160 772
rect 224 740 256 772
rect 320 740 352 772
rect 416 740 448 772
rect 512 740 544 772
rect 608 740 640 772
rect 704 740 736 772
rect 800 740 832 772
<< poly >>
rect 226 636 326 672
rect 124 595 150 631
rect 124 348 150 511
rect 506 612 606 648
rect 688 636 714 672
rect 226 389 326 436
rect 226 357 248 389
rect 280 357 326 389
rect 506 370 606 412
rect 118 330 184 348
rect 118 298 134 330
rect 166 298 184 330
rect 118 282 184 298
rect 226 318 326 357
rect 226 286 248 318
rect 280 286 326 318
rect 463 352 607 370
rect 688 369 714 412
rect 463 320 479 352
rect 511 320 547 352
rect 579 320 607 352
rect 463 304 607 320
rect 649 351 722 369
rect 649 319 665 351
rect 697 319 722 351
rect 124 202 150 282
rect 226 202 326 286
rect 506 266 606 304
rect 649 303 722 319
rect 690 266 716 303
rect 506 146 606 182
rect 124 82 150 118
rect 226 82 326 118
rect 690 82 716 118
<< polycont >>
rect 248 357 280 389
rect 134 298 166 330
rect 248 286 280 318
rect 479 320 511 352
rect 547 320 579 352
rect 665 319 697 351
<< metal1 >>
rect 0 772 864 800
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 608 772
rect 640 740 704 772
rect 736 740 800 772
rect 832 740 864 772
rect 0 712 864 740
rect 60 571 112 576
rect 60 539 70 571
rect 102 539 112 571
rect 60 496 112 539
rect 162 568 214 712
rect 620 621 672 712
rect 620 589 634 621
rect 666 589 672 621
rect 162 536 172 568
rect 204 536 214 568
rect 162 533 214 536
rect 335 571 391 586
rect 335 539 348 571
rect 380 539 391 571
rect 335 523 391 539
rect 60 464 291 496
rect 57 330 183 416
rect 57 298 134 330
rect 166 298 183 330
rect 57 282 183 298
rect 235 389 291 464
rect 235 357 248 389
rect 280 357 291 389
rect 235 318 291 357
rect 235 286 248 318
rect 280 286 291 318
rect 235 241 291 286
rect 60 203 291 241
rect 344 362 391 523
rect 620 513 672 589
rect 620 481 630 513
rect 662 481 672 513
rect 620 479 672 481
rect 731 621 804 634
rect 731 589 744 621
rect 776 589 804 621
rect 731 545 804 589
rect 731 513 744 545
rect 776 513 804 545
rect 441 464 493 476
rect 441 432 452 464
rect 484 443 493 464
rect 731 458 804 513
rect 484 432 668 443
rect 441 409 668 432
rect 731 426 744 458
rect 776 426 804 458
rect 731 415 804 426
rect 630 369 668 409
rect 344 352 585 362
rect 344 320 479 352
rect 511 320 547 352
rect 579 320 585 352
rect 344 310 585 320
rect 630 351 707 369
rect 630 319 665 351
rect 697 319 707 351
rect 60 175 112 203
rect 60 143 70 175
rect 102 143 112 175
rect 344 175 391 310
rect 630 303 707 319
rect 630 247 668 303
rect 761 268 804 415
rect 441 234 668 247
rect 441 202 452 234
rect 484 209 668 234
rect 722 250 804 268
rect 722 218 738 250
rect 770 218 804 250
rect 484 202 494 209
rect 441 189 494 202
rect 60 138 112 143
rect 160 164 214 167
rect 160 132 172 164
rect 204 132 214 164
rect 344 143 348 175
rect 380 143 391 175
rect 344 133 391 143
rect 626 165 678 170
rect 626 133 636 165
rect 668 133 678 165
rect 160 44 214 132
rect 626 44 678 133
rect 722 164 804 218
rect 722 132 738 164
rect 770 132 804 164
rect 722 119 804 132
rect 0 16 864 44
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 608 16
rect 640 -16 704 16
rect 736 -16 800 16
rect 832 -16 864 16
rect 0 -44 864 -16
<< labels >>
flabel metal1 s 57 282 183 416 0 FreeSans 400 0 0 0 A
port 2 nsew
flabel metal1 s 0 712 864 800 0 FreeSans 400 0 0 0 VDD
port 3 nsew
flabel metal1 s 0 -44 864 44 0 FreeSans 400 0 0 0 VSS
port 4 nsew
flabel metal1 s 731 415 804 634 0 FreeSans 400 0 0 0 X
port 5 nsew
<< properties >>
string FIXED_BBOX 0 0 864 756
string GDS_END 57084
string GDS_FILE ../gds/controller.gds
string GDS_START 50868
<< end >>
