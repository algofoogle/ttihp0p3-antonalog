** sch_path: /home/anton/projects/antonalog--REPO/xschem/r2r_dac.sch
.subckt r2r_dac IN[7] IN[6] IN[5] IN[4] IN[3] IN[2] IN[1] IN[0] OUT GND
*.PININFO IN[7:0]:I GND:B OUT:O
XR0a wi0 IN[0] rhigh w=1.0e-6 l=6.0e-6 m=1 b=0
XR0b wJ0 wi0 rhigh w=1.0e-6 l=6.0e-6 m=1 b=0
XR1c wJ0 wJ1 rhigh w=1.0e-6 l=6.0e-6 m=1 b=0
XR0c wg0 wJ0 rhigh w=1.0e-6 l=6.0e-6 m=1 b=0
XR0d GND wg0 rhigh w=1.0e-6 l=6.0e-6 m=1 b=0
XR1a wi1 IN[1] rhigh w=1.0e-6 l=6.0e-6 m=1 b=0
XR1b wJ1 wi1 rhigh w=1.0e-6 l=6.0e-6 m=1 b=0
XR2c wJ1 wJ2 rhigh w=1.0e-6 l=6.0e-6 m=1 b=0
XR2a wi2 IN[2] rhigh w=1.0e-6 l=6.0e-6 m=1 b=0
XR2b wJ2 wi2 rhigh w=1.0e-6 l=6.0e-6 m=1 b=0
XR3c wJ2 wJ3 rhigh w=1.0e-6 l=6.0e-6 m=1 b=0
XR3a wi3 IN[3] rhigh w=1.0e-6 l=6.0e-6 m=1 b=0
XR3b wJ3 wi3 rhigh w=1.0e-6 l=6.0e-6 m=1 b=0
XR4c wJ3 wJ4 rhigh w=1.0e-6 l=6.0e-6 m=1 b=0
XR4a wi4 IN[4] rhigh w=1.0e-6 l=6.0e-6 m=1 b=0
XR4b wJ4 wi4 rhigh w=1.0e-6 l=6.0e-6 m=1 b=0
XR5c wJ4 wJ5 rhigh w=1.0e-6 l=6.0e-6 m=1 b=0
XR5a wi5 IN[5] rhigh w=1.0e-6 l=6.0e-6 m=1 b=0
XR5b wJ5 wi5 rhigh w=1.0e-6 l=6.0e-6 m=1 b=0
XR6c wJ5 wJ6 rhigh w=1.0e-6 l=6.0e-6 m=1 b=0
XR6a wi6 IN[6] rhigh w=1.0e-6 l=6.0e-6 m=1 b=0
XR6b wJ6 wi6 rhigh w=1.0e-6 l=6.0e-6 m=1 b=0
XR7c wJ6 OUT rhigh w=1.0e-6 l=6.0e-6 m=1 b=0
XR7a wi7 IN[7] rhigh w=1.0e-6 l=6.0e-6 m=1 b=0
XR7b OUT wi7 rhigh w=1.0e-6 l=6.0e-6 m=1 b=0
.ends
