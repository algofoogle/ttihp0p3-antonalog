magic
tech ihp-sg13g2
magscale 1 2
timestamp 1747056038
<< nwell >>
rect -48 350 816 834
<< pwell >>
rect 21 56 745 314
rect -26 -56 794 56
<< nmos >>
rect 115 140 141 288
rect 217 140 243 288
rect 319 140 345 288
rect 421 140 447 288
rect 523 140 549 288
rect 625 140 651 288
<< pmos >>
rect 115 412 141 636
rect 217 412 243 636
rect 319 412 345 636
rect 421 412 447 636
rect 523 412 549 636
rect 625 412 651 636
<< ndiff >>
rect 47 274 115 288
rect 47 242 61 274
rect 93 242 115 274
rect 47 186 115 242
rect 47 154 61 186
rect 93 154 115 186
rect 47 140 115 154
rect 141 186 217 288
rect 141 154 163 186
rect 195 154 217 186
rect 141 140 217 154
rect 243 274 319 288
rect 243 242 265 274
rect 297 242 319 274
rect 243 202 319 242
rect 243 170 265 202
rect 297 170 319 202
rect 243 140 319 170
rect 345 186 421 288
rect 345 154 367 186
rect 399 154 421 186
rect 345 140 421 154
rect 447 186 523 288
rect 447 154 469 186
rect 501 154 523 186
rect 447 140 523 154
rect 549 274 625 288
rect 549 242 571 274
rect 603 242 625 274
rect 549 186 625 242
rect 549 154 571 186
rect 603 154 625 186
rect 549 140 625 154
rect 651 274 719 288
rect 651 242 673 274
rect 705 242 719 274
rect 651 186 719 242
rect 651 154 673 186
rect 705 154 719 186
rect 651 140 719 154
<< pdiff >>
rect 47 622 115 636
rect 47 590 61 622
rect 93 590 115 622
rect 47 543 115 590
rect 47 511 61 543
rect 93 511 115 543
rect 47 412 115 511
rect 141 622 217 636
rect 141 590 163 622
rect 195 590 217 622
rect 141 412 217 590
rect 243 622 319 636
rect 243 590 265 622
rect 297 590 319 622
rect 243 543 319 590
rect 243 511 265 543
rect 297 511 319 543
rect 243 412 319 511
rect 345 622 421 636
rect 345 590 367 622
rect 399 590 421 622
rect 345 412 421 590
rect 447 622 523 636
rect 447 590 469 622
rect 501 590 523 622
rect 447 543 523 590
rect 447 511 469 543
rect 501 511 523 543
rect 447 412 523 511
rect 549 543 625 636
rect 549 511 571 543
rect 603 511 625 543
rect 549 458 625 511
rect 549 426 571 458
rect 603 426 625 458
rect 549 412 625 426
rect 651 622 719 636
rect 651 590 673 622
rect 705 590 719 622
rect 651 543 719 590
rect 651 511 673 543
rect 705 511 719 543
rect 651 412 719 511
<< ndiffc >>
rect 61 242 93 274
rect 61 154 93 186
rect 163 154 195 186
rect 265 242 297 274
rect 265 170 297 202
rect 367 154 399 186
rect 469 154 501 186
rect 571 242 603 274
rect 571 154 603 186
rect 673 242 705 274
rect 673 154 705 186
<< pdiffc >>
rect 61 590 93 622
rect 61 511 93 543
rect 163 590 195 622
rect 265 590 297 622
rect 265 511 297 543
rect 367 590 399 622
rect 469 590 501 622
rect 469 511 501 543
rect 571 511 603 543
rect 571 426 603 458
rect 673 590 705 622
rect 673 511 705 543
<< psubdiff >>
rect 0 16 768 30
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 608 16
rect 640 -16 704 16
rect 736 -16 768 16
rect 0 -30 768 -16
<< nsubdiff >>
rect 0 772 768 786
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 608 772
rect 640 740 704 772
rect 736 740 768 772
rect 0 726 768 740
<< psubdiffcont >>
rect 32 -16 64 16
rect 128 -16 160 16
rect 224 -16 256 16
rect 320 -16 352 16
rect 416 -16 448 16
rect 512 -16 544 16
rect 608 -16 640 16
rect 704 -16 736 16
<< nsubdiffcont >>
rect 32 740 64 772
rect 128 740 160 772
rect 224 740 256 772
rect 320 740 352 772
rect 416 740 448 772
rect 512 740 544 772
rect 608 740 640 772
rect 704 740 736 772
<< poly >>
rect 115 636 141 672
rect 217 636 243 672
rect 319 636 345 672
rect 421 636 447 672
rect 523 636 549 672
rect 625 636 651 672
rect 115 380 141 412
rect 217 380 243 412
rect 319 380 345 412
rect 421 380 447 412
rect 523 380 549 412
rect 625 380 651 412
rect 98 366 158 380
rect 98 334 112 366
rect 144 334 158 366
rect 98 320 158 334
rect 217 366 345 380
rect 217 334 231 366
rect 263 334 299 366
rect 331 334 345 366
rect 217 320 345 334
rect 404 366 464 380
rect 404 334 418 366
rect 450 334 464 366
rect 404 320 464 334
rect 523 366 717 380
rect 523 334 671 366
rect 703 334 717 366
rect 523 320 717 334
rect 115 288 141 320
rect 217 288 243 320
rect 319 288 345 320
rect 421 288 447 320
rect 523 288 549 320
rect 625 288 651 320
rect 115 104 141 140
rect 217 104 243 140
rect 319 104 345 140
rect 421 104 447 140
rect 523 104 549 140
rect 625 104 651 140
<< polycont >>
rect 112 334 144 366
rect 231 334 263 366
rect 299 334 331 366
rect 418 334 450 366
rect 671 334 703 366
<< metal1 >>
rect 0 772 768 800
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 608 772
rect 640 740 704 772
rect 736 740 768 772
rect 0 712 768 740
rect 51 622 103 632
rect 51 590 61 622
rect 93 590 103 622
rect 153 622 205 712
rect 153 590 163 622
rect 195 590 205 622
rect 255 622 307 632
rect 255 590 265 622
rect 297 590 307 622
rect 357 622 409 712
rect 357 590 367 622
rect 399 590 409 622
rect 459 622 715 632
rect 459 590 469 622
rect 501 590 673 622
rect 705 590 715 622
rect 51 553 103 590
rect 255 553 307 590
rect 459 580 715 590
rect 459 553 511 580
rect 51 543 511 553
rect 663 543 715 580
rect 51 511 61 543
rect 93 511 265 543
rect 297 511 469 543
rect 501 511 511 543
rect 51 501 511 511
rect 561 511 571 543
rect 603 511 613 543
rect 78 418 460 463
rect 78 366 154 418
rect 78 334 112 366
rect 144 334 154 366
rect 78 320 154 334
rect 217 366 345 380
rect 217 334 231 366
rect 263 334 299 366
rect 331 334 345 366
rect 217 314 345 334
rect 408 366 460 418
rect 408 334 418 366
rect 450 334 460 366
rect 408 320 460 334
rect 561 458 613 511
rect 663 511 673 543
rect 705 511 715 543
rect 663 501 715 511
rect 561 426 571 458
rect 603 426 613 458
rect 51 274 103 284
rect 561 278 613 426
rect 656 366 715 456
rect 656 334 671 366
rect 703 334 715 366
rect 656 325 715 334
rect 51 242 61 274
rect 93 242 103 274
rect 51 186 103 242
rect 255 274 613 278
rect 255 242 265 274
rect 297 242 571 274
rect 603 242 613 274
rect 255 232 613 242
rect 255 202 307 232
rect 51 154 61 186
rect 93 154 103 186
rect 51 44 103 154
rect 153 186 205 196
rect 153 154 163 186
rect 195 154 205 186
rect 255 170 265 202
rect 297 170 307 202
rect 357 186 409 196
rect 153 134 205 154
rect 357 154 367 186
rect 399 154 409 186
rect 357 134 409 154
rect 153 89 409 134
rect 459 186 511 196
rect 459 154 469 186
rect 501 154 511 186
rect 459 44 511 154
rect 561 186 613 232
rect 561 154 571 186
rect 603 154 613 186
rect 561 144 613 154
rect 663 274 715 284
rect 663 242 673 274
rect 705 242 715 274
rect 663 186 715 242
rect 663 154 673 186
rect 705 154 715 186
rect 663 44 715 154
rect 0 16 768 44
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 608 16
rect 640 -16 704 16
rect 736 -16 768 16
rect 0 -44 768 -16
<< labels >>
flabel metal1 s 561 144 613 543 0 FreeSans 400 0 0 0 Y
port 2 nsew
flabel metal1 s 78 320 154 463 0 FreeSans 400 0 0 0 A2
port 3 nsew
flabel metal1 s 0 712 768 800 0 FreeSans 400 0 0 0 VDD
port 4 nsew
flabel metal1 s 217 314 345 380 0 FreeSans 400 0 0 0 A1
port 5 nsew
flabel metal1 s 656 325 715 456 0 FreeSans 400 0 0 0 B1
port 6 nsew
flabel metal1 s 0 -44 768 44 0 FreeSans 400 0 0 0 VSS
port 7 nsew
<< properties >>
string FIXED_BBOX 0 0 768 756
string GDS_END 143476
string GDS_FILE ../gds/controller.gds
string GDS_START 137936
<< end >>
