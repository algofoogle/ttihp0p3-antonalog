magic
tech ihp-sg13g2
magscale 1 2
timestamp 1747537721
<< nwell >>
rect -48 350 528 834
<< pwell >>
rect 45 56 475 300
rect -26 -56 506 56
<< nmos >>
rect 139 120 165 274
rect 253 120 279 274
rect 355 120 381 274
<< pmos >>
rect 139 412 165 636
rect 228 412 254 636
rect 319 412 345 636
<< ndiff >>
rect 71 234 139 274
rect 71 202 85 234
rect 117 202 139 234
rect 71 166 139 202
rect 71 134 85 166
rect 117 134 139 166
rect 71 120 139 134
rect 165 252 253 274
rect 165 220 199 252
rect 231 220 253 252
rect 165 166 253 220
rect 165 134 199 166
rect 231 134 253 166
rect 165 120 253 134
rect 279 166 355 274
rect 279 134 301 166
rect 333 134 355 166
rect 279 120 355 134
rect 381 252 449 274
rect 381 220 403 252
rect 435 220 449 252
rect 381 166 449 220
rect 381 134 403 166
rect 435 134 449 166
rect 381 120 449 134
<< pdiff >>
rect 71 621 139 636
rect 71 589 85 621
rect 117 589 139 621
rect 71 551 139 589
rect 71 519 85 551
rect 117 519 139 551
rect 71 483 139 519
rect 71 451 85 483
rect 117 451 139 483
rect 71 412 139 451
rect 165 412 228 636
rect 254 412 319 636
rect 345 621 413 636
rect 345 589 367 621
rect 399 589 413 621
rect 345 553 413 589
rect 345 521 367 553
rect 399 521 413 553
rect 345 483 413 521
rect 345 451 367 483
rect 399 451 413 483
rect 345 412 413 451
<< ndiffc >>
rect 85 202 117 234
rect 85 134 117 166
rect 199 220 231 252
rect 199 134 231 166
rect 301 134 333 166
rect 403 220 435 252
rect 403 134 435 166
<< pdiffc >>
rect 85 589 117 621
rect 85 519 117 551
rect 85 451 117 483
rect 367 589 399 621
rect 367 521 399 553
rect 367 451 399 483
<< psubdiff >>
rect 0 16 480 30
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 480 16
rect 0 -30 480 -16
<< nsubdiff >>
rect 0 772 480 786
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 480 772
rect 0 726 480 740
<< psubdiffcont >>
rect 32 -16 64 16
rect 128 -16 160 16
rect 224 -16 256 16
rect 320 -16 352 16
rect 416 -16 448 16
<< nsubdiffcont >>
rect 32 740 64 772
rect 128 740 160 772
rect 224 740 256 772
rect 320 740 352 772
rect 416 740 448 772
<< poly >>
rect 139 636 165 672
rect 228 636 254 672
rect 319 636 345 672
rect 139 354 165 412
rect 228 370 254 412
rect 319 370 345 412
rect 65 337 165 354
rect 65 305 82 337
rect 114 305 165 337
rect 65 288 165 305
rect 215 353 281 370
rect 215 321 232 353
rect 264 321 281 353
rect 215 304 281 321
rect 319 353 419 370
rect 319 321 370 353
rect 402 321 419 353
rect 319 304 419 321
rect 139 274 165 288
rect 253 274 279 304
rect 355 274 381 304
rect 139 60 165 120
rect 253 60 279 120
rect 355 60 381 120
<< polycont >>
rect 82 305 114 337
rect 232 321 264 353
rect 370 321 402 353
<< metal1 >>
rect 0 772 480 800
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 480 772
rect 0 712 480 740
rect 72 621 122 712
rect 72 589 85 621
rect 117 589 122 621
rect 72 551 122 589
rect 72 519 85 551
rect 117 519 122 551
rect 357 621 409 626
rect 357 589 367 621
rect 399 589 409 621
rect 357 553 409 589
rect 357 533 367 553
rect 72 483 122 519
rect 72 451 85 483
rect 117 451 122 483
rect 72 441 122 451
rect 158 521 367 533
rect 399 521 409 553
rect 158 483 409 521
rect 158 451 367 483
rect 399 451 409 483
rect 158 434 409 451
rect 65 337 116 400
rect 65 305 82 337
rect 114 305 116 337
rect 65 292 116 305
rect 158 270 193 434
rect 230 353 307 389
rect 230 321 232 353
rect 264 321 307 353
rect 230 307 307 321
rect 353 353 419 389
rect 353 321 370 353
rect 402 321 419 353
rect 353 307 419 321
rect 158 252 445 270
rect 72 234 117 247
rect 72 202 85 234
rect 158 220 199 252
rect 231 220 403 252
rect 435 220 445 252
rect 72 166 117 202
rect 72 134 85 166
rect 72 44 117 134
rect 189 166 241 220
rect 189 134 199 166
rect 231 134 241 166
rect 189 131 241 134
rect 291 166 343 169
rect 291 134 301 166
rect 333 134 343 166
rect 291 44 343 134
rect 393 166 445 220
rect 393 134 403 166
rect 435 134 445 166
rect 393 131 445 134
rect 0 16 480 44
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 480 16
rect 0 -44 480 -16
<< labels >>
flabel metal1 s 65 292 116 400 0 FreeSans 400 0 0 0 A
port 2 nsew
flabel metal1 s 158 476 409 533 0 FreeSans 400 0 0 0 Y
port 3 nsew
flabel metal1 s 230 307 307 389 0 FreeSans 400 0 0 0 B
port 4 nsew
flabel metal1 s 353 307 419 389 0 FreeSans 400 0 0 0 C
port 5 nsew
flabel metal1 s 0 712 480 800 0 FreeSans 400 0 0 0 VDD
port 6 nsew
flabel metal1 s 0 -44 480 44 0 FreeSans 400 0 0 0 VSS
port 7 nsew
<< properties >>
string FIXED_BBOX 0 0 480 756
string GDS_END 103594
string GDS_FILE ../gds/controller.gds
string GDS_START 99078
<< end >>
