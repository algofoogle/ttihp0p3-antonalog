magic
tech ihp-sg13g2
timestamp 1747537721
<< nwell >>
rect -24 175 552 417
<< pwell >>
rect 16 28 528 146
rect -13 -28 541 28
<< nmos >>
rect 63 78 76 133
rect 129 59 142 133
rect 178 59 191 133
rect 235 59 248 133
rect 339 59 352 133
rect 392 59 405 133
rect 460 59 473 133
<< pmos >>
rect 63 206 76 290
rect 129 206 142 306
rect 209 206 222 306
rect 266 206 279 306
rect 339 206 352 306
rect 392 206 405 318
rect 460 206 473 318
<< ndiff >>
rect 29 113 63 133
rect 29 97 36 113
rect 52 97 63 113
rect 29 78 63 97
rect 76 126 129 133
rect 76 110 90 126
rect 106 110 129 126
rect 76 82 129 110
rect 76 78 90 82
rect 83 66 90 78
rect 106 66 129 82
rect 83 59 129 66
rect 142 59 178 133
rect 191 82 235 133
rect 191 66 206 82
rect 222 66 235 82
rect 191 59 235 66
rect 248 59 339 133
rect 352 82 392 133
rect 352 66 365 82
rect 381 66 392 82
rect 352 59 392 66
rect 405 124 460 133
rect 405 108 433 124
rect 449 108 460 124
rect 405 83 460 108
rect 405 67 433 83
rect 449 67 460 83
rect 405 59 460 67
rect 473 126 515 133
rect 473 110 492 126
rect 508 110 515 126
rect 473 82 515 110
rect 473 66 492 82
rect 508 66 515 82
rect 473 59 515 66
<< pdiff >>
rect 359 306 392 318
rect 91 290 129 306
rect 29 283 63 290
rect 29 267 36 283
rect 52 267 63 283
rect 29 235 63 267
rect 29 219 36 235
rect 52 219 63 235
rect 29 206 63 219
rect 76 280 129 290
rect 76 264 102 280
rect 118 264 129 280
rect 76 206 129 264
rect 142 206 209 306
rect 222 286 266 306
rect 222 270 235 286
rect 251 270 266 286
rect 222 229 266 270
rect 222 213 235 229
rect 251 213 266 229
rect 222 206 266 213
rect 279 206 339 306
rect 352 298 392 306
rect 352 282 365 298
rect 381 282 392 298
rect 352 263 392 282
rect 352 247 365 263
rect 381 247 392 263
rect 352 229 392 247
rect 352 213 365 229
rect 381 213 392 229
rect 352 206 392 213
rect 405 311 460 318
rect 405 295 433 311
rect 449 295 460 311
rect 405 269 460 295
rect 405 253 433 269
rect 449 253 460 269
rect 405 229 460 253
rect 405 213 433 229
rect 449 213 460 229
rect 405 206 460 213
rect 473 298 515 318
rect 473 282 492 298
rect 508 282 515 298
rect 473 263 515 282
rect 473 247 492 263
rect 508 247 515 263
rect 473 229 515 247
rect 473 213 492 229
rect 508 213 515 229
rect 473 206 515 213
<< ndiffc >>
rect 36 97 52 113
rect 90 110 106 126
rect 90 66 106 82
rect 206 66 222 82
rect 365 66 381 82
rect 433 108 449 124
rect 433 67 449 83
rect 492 110 508 126
rect 492 66 508 82
<< pdiffc >>
rect 36 267 52 283
rect 36 219 52 235
rect 102 264 118 280
rect 235 270 251 286
rect 235 213 251 229
rect 365 282 381 298
rect 365 247 381 263
rect 365 213 381 229
rect 433 295 449 311
rect 433 253 449 269
rect 433 213 449 229
rect 492 282 508 298
rect 492 247 508 263
rect 492 213 508 229
<< psubdiff >>
rect 0 8 528 15
rect 0 -8 16 8
rect 32 -8 64 8
rect 80 -8 112 8
rect 128 -8 160 8
rect 176 -8 208 8
rect 224 -8 256 8
rect 272 -8 304 8
rect 320 -8 352 8
rect 368 -8 400 8
rect 416 -8 448 8
rect 464 -8 496 8
rect 512 -8 528 8
rect 0 -15 528 -8
<< nsubdiff >>
rect 0 386 528 393
rect 0 370 16 386
rect 32 370 64 386
rect 80 370 112 386
rect 128 370 160 386
rect 176 370 208 386
rect 224 370 256 386
rect 272 370 304 386
rect 320 370 352 386
rect 368 370 400 386
rect 416 370 448 386
rect 464 370 496 386
rect 512 370 528 386
rect 0 363 528 370
<< psubdiffcont >>
rect 16 -8 32 8
rect 64 -8 80 8
rect 112 -8 128 8
rect 160 -8 176 8
rect 208 -8 224 8
rect 256 -8 272 8
rect 304 -8 320 8
rect 352 -8 368 8
rect 400 -8 416 8
rect 448 -8 464 8
rect 496 -8 512 8
<< nsubdiffcont >>
rect 16 370 32 386
rect 64 370 80 386
rect 112 370 128 386
rect 160 370 176 386
rect 208 370 224 386
rect 256 370 272 386
rect 304 370 320 386
rect 352 370 368 386
rect 400 370 416 386
rect 448 370 464 386
rect 496 370 512 386
<< poly >>
rect 63 290 76 308
rect 129 306 142 324
rect 209 306 222 324
rect 266 306 279 324
rect 339 306 352 324
rect 392 318 405 336
rect 460 318 473 336
rect 63 190 76 206
rect 129 190 142 206
rect 63 181 142 190
rect 63 165 70 181
rect 86 165 142 181
rect 209 177 222 206
rect 266 177 279 206
rect 339 187 352 206
rect 339 178 372 187
rect 63 157 142 165
rect 63 133 76 157
rect 129 133 142 157
rect 161 168 191 175
rect 161 152 168 168
rect 184 152 191 168
rect 161 145 191 152
rect 178 133 191 145
rect 209 168 248 177
rect 209 152 217 168
rect 233 152 248 168
rect 209 144 248 152
rect 266 168 299 177
rect 266 152 274 168
rect 290 152 299 168
rect 266 144 299 152
rect 339 162 347 178
rect 363 162 372 178
rect 339 154 372 162
rect 392 185 405 206
rect 460 185 473 206
rect 392 176 473 185
rect 392 160 401 176
rect 417 160 473 176
rect 235 133 248 144
rect 339 133 352 154
rect 392 152 473 160
rect 392 133 405 152
rect 460 133 473 152
rect 63 60 76 78
rect 129 41 142 59
rect 178 41 191 59
rect 235 41 248 59
rect 339 41 352 59
rect 392 41 405 59
rect 460 41 473 59
<< polycont >>
rect 70 165 86 181
rect 168 152 184 168
rect 217 152 233 168
rect 274 152 290 168
rect 347 162 363 178
rect 401 160 417 176
<< metal1 >>
rect 0 386 528 400
rect 0 370 16 386
rect 32 370 64 386
rect 80 370 112 386
rect 128 370 160 386
rect 176 370 208 386
rect 224 370 256 386
rect 272 370 304 386
rect 320 370 352 386
rect 368 370 400 386
rect 416 370 448 386
rect 464 370 496 386
rect 512 370 528 386
rect 0 356 528 370
rect 14 283 57 284
rect 14 267 36 283
rect 52 267 57 283
rect 14 246 57 267
rect 97 280 123 356
rect 97 264 102 280
rect 118 264 123 280
rect 148 312 342 329
rect 148 246 164 312
rect 14 235 164 246
rect 14 219 36 235
rect 52 230 164 235
rect 230 286 256 287
rect 230 270 235 286
rect 251 270 256 286
rect 52 219 57 230
rect 14 217 57 219
rect 230 229 256 270
rect 14 118 35 217
rect 230 213 235 229
rect 251 213 256 229
rect 182 212 256 213
rect 127 196 256 212
rect 127 195 191 196
rect 60 181 109 190
rect 60 165 70 181
rect 86 165 109 181
rect 60 150 109 165
rect 85 126 109 131
rect 14 113 57 118
rect 14 97 36 113
rect 52 97 57 113
rect 14 92 57 97
rect 85 110 90 126
rect 106 110 109 126
rect 85 82 109 110
rect 85 66 90 82
rect 106 66 109 82
rect 85 22 109 66
rect 127 83 143 195
rect 325 187 342 312
rect 363 298 383 356
rect 363 282 365 298
rect 381 282 383 298
rect 363 263 383 282
rect 363 247 365 263
rect 381 247 383 263
rect 363 229 383 247
rect 363 213 365 229
rect 381 213 383 229
rect 363 208 383 213
rect 413 311 468 320
rect 413 295 433 311
rect 449 295 468 311
rect 413 269 468 295
rect 413 253 433 269
rect 449 253 468 269
rect 413 229 468 253
rect 413 213 433 229
rect 449 213 468 229
rect 413 204 468 213
rect 490 298 510 356
rect 490 282 492 298
rect 508 282 510 298
rect 490 263 510 282
rect 490 247 492 263
rect 508 247 510 263
rect 490 229 510 247
rect 490 213 492 229
rect 508 213 510 229
rect 490 208 510 213
rect 325 178 372 187
rect 161 168 189 175
rect 161 152 168 168
rect 184 152 189 168
rect 161 144 189 152
rect 171 120 189 144
rect 209 168 248 178
rect 209 152 217 168
rect 233 152 248 168
rect 209 140 248 152
rect 269 168 299 178
rect 269 152 274 168
rect 290 152 299 168
rect 325 162 347 178
rect 363 162 372 178
rect 325 154 372 162
rect 394 176 424 185
rect 394 160 401 176
rect 417 160 424 176
rect 269 120 299 152
rect 394 152 424 160
rect 394 120 413 152
rect 451 131 468 204
rect 171 103 299 120
rect 319 103 413 120
rect 431 124 468 131
rect 431 108 433 124
rect 449 108 468 124
rect 319 83 336 103
rect 127 82 336 83
rect 127 66 206 82
rect 222 66 336 82
rect 127 61 336 66
rect 360 82 386 84
rect 360 66 365 82
rect 381 66 386 82
rect 360 22 386 66
rect 431 83 468 108
rect 431 67 433 83
rect 449 67 468 83
rect 431 57 468 67
rect 487 126 513 131
rect 487 110 492 126
rect 508 110 513 126
rect 487 82 513 110
rect 487 66 492 82
rect 508 66 513 82
rect 487 22 513 66
rect 0 8 528 22
rect 0 -8 16 8
rect 32 -8 64 8
rect 80 -8 112 8
rect 128 -8 160 8
rect 176 -8 208 8
rect 224 -8 256 8
rect 272 -8 304 8
rect 320 -8 352 8
rect 368 -8 400 8
rect 416 -8 448 8
rect 464 -8 496 8
rect 512 -8 528 8
rect 0 -22 528 -8
<< labels >>
flabel metal1 s 269 103 299 178 0 FreeSans 200 0 0 0 A1
port 2 nsew
flabel metal1 s 413 204 468 320 0 FreeSans 200 0 0 0 X
port 3 nsew
flabel metal1 s 60 150 109 190 0 FreeSans 200 0 0 0 S
port 4 nsew
flabel metal1 s 0 356 528 400 0 FreeSans 200 0 0 0 VDD
port 5 nsew
flabel metal1 s 0 -22 528 22 0 FreeSans 200 0 0 0 VSS
port 6 nsew
flabel metal1 s 209 140 248 178 0 FreeSans 200 0 0 0 A0
port 7 nsew
<< properties >>
string FIXED_BBOX 0 0 528 378
string GDS_END 199358
string GDS_FILE ../gds/controller.gds
string GDS_START 191706
<< end >>
