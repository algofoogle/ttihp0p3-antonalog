* NGSPICE file created from r2r_dac.ext - technology: ihp-sg13g2

.subckt rhigh a_0_1200# a_0_n86#
X0 a_0_1200# a_0_n86# rhigh l=6u w=1u
.ends

*.subckt resistors B rhigh_0[0]/a_0_1200# rhigh_0[23]/a_0_n86# rhigh_0[11]/a_0_1200#
.subckt resistors rhigh_0[0]/a_0_1200# rhigh_0[23]/a_0_n86# rhigh_0[11]/a_0_1200#
+ rhigh_0[6]/a_0_n86# rhigh_0[21]/a_0_1200# rhigh_0[1]/a_0_1200# rhigh_0[2]/a_0_n86#
+ rhigh_0[12]/a_0_1200# rhigh_0[18]/a_0_n86# rhigh_0[22]/a_0_1200# rhigh_0[2]/a_0_1200#
+ rhigh_0[14]/a_0_n86# rhigh_0[13]/a_0_1200# rhigh_0[10]/a_0_n86# rhigh_0[23]/a_0_1200#
+ rhigh_0[3]/a_0_1200# rhigh_0[24]/a_0_n86# rhigh_0[20]/a_0_n86# rhigh_0[7]/a_0_n86#
+ rhigh_0[14]/a_0_1200# rhigh_0[3]/a_0_n86# rhigh_0[24]/a_0_1200# rhigh_0[4]/a_0_1200#
+ rhigh_0[19]/a_0_n86# rhigh_0[15]/a_0_1200# rhigh_0[15]/a_0_n86# rhigh_0[5]/a_0_1200#
+ rhigh_0[11]/a_0_n86# rhigh_0[16]/a_0_1200# rhigh_0[8]/a_0_n86# rhigh_0[21]/a_0_n86#
+ rhigh_0[4]/a_0_n86# rhigh_0[6]/a_0_1200# rhigh_0[17]/a_0_1200# rhigh_0[0]/a_0_n86#
+ rhigh_0[18]/a_0_1200# rhigh_0[7]/a_0_1200# rhigh_0[16]/a_0_n86# rhigh_0[12]/a_0_n86#
+ rhigh_0[8]/a_0_1200# rhigh_0[19]/a_0_1200# rhigh_0[9]/a_0_n86# rhigh_0[22]/a_0_n86#
+ rhigh_0[9]/a_0_1200# rhigh_0[5]/a_0_n86# rhigh_0[1]/a_0_n86# rhigh_0[17]/a_0_n86#
+ rhigh_0[10]/a_0_1200# rhigh_0[13]/a_0_n86# rhigh_0[20]/a_0_1200#
Xrhigh_0[0] rhigh_0[0]/a_0_1200# rhigh_0[0]/a_0_n86# rhigh
Xrhigh_0[1] rhigh_0[1]/a_0_1200# rhigh_0[1]/a_0_n86# rhigh
Xrhigh_0[2] rhigh_0[2]/a_0_1200# rhigh_0[2]/a_0_n86# rhigh
Xrhigh_0[3] rhigh_0[3]/a_0_1200# rhigh_0[3]/a_0_n86# rhigh
Xrhigh_0[4] rhigh_0[4]/a_0_1200# rhigh_0[4]/a_0_n86# rhigh
Xrhigh_0[5] rhigh_0[5]/a_0_1200# rhigh_0[5]/a_0_n86# rhigh
Xrhigh_0[6] rhigh_0[6]/a_0_1200# rhigh_0[6]/a_0_n86# rhigh
Xrhigh_0[7] rhigh_0[7]/a_0_1200# rhigh_0[7]/a_0_n86# rhigh
Xrhigh_0[8] rhigh_0[8]/a_0_1200# rhigh_0[8]/a_0_n86# rhigh
Xrhigh_0[9] rhigh_0[9]/a_0_1200# rhigh_0[9]/a_0_n86# rhigh
Xrhigh_0[10] rhigh_0[10]/a_0_1200# rhigh_0[10]/a_0_n86# rhigh
Xrhigh_0[11] rhigh_0[11]/a_0_1200# rhigh_0[11]/a_0_n86# rhigh
Xrhigh_0[12] rhigh_0[12]/a_0_1200# rhigh_0[12]/a_0_n86# rhigh
Xrhigh_0[13] rhigh_0[13]/a_0_1200# rhigh_0[13]/a_0_n86# rhigh
Xrhigh_0[14] rhigh_0[14]/a_0_1200# rhigh_0[14]/a_0_n86# rhigh
Xrhigh_0[15] rhigh_0[15]/a_0_1200# rhigh_0[15]/a_0_n86# rhigh
Xrhigh_0[16] rhigh_0[16]/a_0_1200# rhigh_0[16]/a_0_n86# rhigh
Xrhigh_0[17] rhigh_0[17]/a_0_1200# rhigh_0[17]/a_0_n86# rhigh
Xrhigh_0[18] rhigh_0[18]/a_0_1200# rhigh_0[18]/a_0_n86# rhigh
Xrhigh_0[19] rhigh_0[19]/a_0_1200# rhigh_0[19]/a_0_n86# rhigh
Xrhigh_0[20] rhigh_0[20]/a_0_1200# rhigh_0[20]/a_0_n86# rhigh
Xrhigh_0[21] rhigh_0[21]/a_0_1200# rhigh_0[21]/a_0_n86# rhigh
Xrhigh_0[22] rhigh_0[22]/a_0_1200# rhigh_0[22]/a_0_n86# rhigh
Xrhigh_0[23] rhigh_0[23]/a_0_1200# rhigh_0[23]/a_0_n86# rhigh
Xrhigh_0[24] rhigh_0[24]/a_0_1200# rhigh_0[24]/a_0_n86# rhigh
.ends

.subckt r2r_dac IN[7] IN[6] IN[5] IN[4] IN[3] IN[2] IN[1] IN[0] OUT GND
Xresistors_0 wg0 wi7 wJ3 wi1 wi6 wg0 wJ0 IN[3] wi5 OUT wi0 wJ4 wJ3 wJ2 OUT wi0
+ wi7 wJ6 wJ2 wi4 IN[0] IN[7] wJ1 wJ6 wi4 IN[4] wJ1 wi3 wJ5 wJ2 IN[6] wJ0 IN[1] wJ5
+ GND IN[5] wJ1 wJ4 wi3 wi2 wJ5 IN[2] wJ6 wi2 wi1 wJ0 wi5 wJ3 wJ4 wi6 resistors
.ends

