magic
tech ihp-sg13g2
timestamp 1747537721
<< nwell >>
rect -24 175 312 417
<< pwell >>
rect 15 28 275 146
rect -13 -28 301 28
<< nmos >>
rect 62 59 75 133
rect 113 59 126 133
rect 164 59 177 133
rect 215 59 228 133
<< pmos >>
rect 62 206 75 318
rect 113 206 126 318
rect 164 206 177 318
rect 215 206 228 318
<< ndiff >>
rect 28 126 62 133
rect 28 110 35 126
rect 51 110 62 126
rect 28 82 62 110
rect 28 66 35 82
rect 51 66 62 82
rect 28 59 62 66
rect 75 126 113 133
rect 75 110 86 126
rect 102 110 113 126
rect 75 82 113 110
rect 75 66 86 82
rect 102 66 113 82
rect 75 59 113 66
rect 126 82 164 133
rect 126 66 137 82
rect 153 66 164 82
rect 126 59 164 66
rect 177 126 215 133
rect 177 110 188 126
rect 204 110 215 126
rect 177 82 215 110
rect 177 66 188 82
rect 204 66 215 82
rect 177 59 215 66
rect 228 82 262 133
rect 228 66 239 82
rect 255 66 262 82
rect 228 59 262 66
<< pdiff >>
rect 26 311 62 318
rect 26 295 35 311
rect 51 295 62 311
rect 26 275 62 295
rect 26 259 35 275
rect 51 259 62 275
rect 26 229 62 259
rect 26 213 35 229
rect 51 213 62 229
rect 26 206 62 213
rect 75 311 113 318
rect 75 295 86 311
rect 102 295 113 311
rect 75 275 113 295
rect 75 259 86 275
rect 102 259 113 275
rect 75 206 113 259
rect 126 311 164 318
rect 126 295 137 311
rect 153 295 164 311
rect 126 275 164 295
rect 126 259 137 275
rect 153 259 164 275
rect 126 229 164 259
rect 126 213 137 229
rect 153 213 164 229
rect 126 206 164 213
rect 177 229 215 318
rect 177 213 188 229
rect 204 213 215 229
rect 177 206 215 213
rect 228 311 262 318
rect 228 295 239 311
rect 255 295 262 311
rect 228 275 262 295
rect 228 259 239 275
rect 255 259 262 275
rect 228 206 262 259
<< ndiffc >>
rect 35 110 51 126
rect 35 66 51 82
rect 86 110 102 126
rect 86 66 102 82
rect 137 66 153 82
rect 188 110 204 126
rect 188 66 204 82
rect 239 66 255 82
<< pdiffc >>
rect 35 295 51 311
rect 35 259 51 275
rect 35 213 51 229
rect 86 295 102 311
rect 86 259 102 275
rect 137 295 153 311
rect 137 259 153 275
rect 137 213 153 229
rect 188 213 204 229
rect 239 295 255 311
rect 239 259 255 275
<< psubdiff >>
rect 0 8 288 15
rect 0 -8 16 8
rect 32 -8 64 8
rect 80 -8 112 8
rect 128 -8 160 8
rect 176 -8 208 8
rect 224 -8 256 8
rect 272 -8 288 8
rect 0 -15 288 -8
<< nsubdiff >>
rect 0 386 288 393
rect 0 370 16 386
rect 32 370 64 386
rect 80 370 112 386
rect 128 370 160 386
rect 176 370 208 386
rect 224 370 256 386
rect 272 370 288 386
rect 0 363 288 370
<< psubdiffcont >>
rect 16 -8 32 8
rect 64 -8 80 8
rect 112 -8 128 8
rect 160 -8 176 8
rect 208 -8 224 8
rect 256 -8 272 8
<< nsubdiffcont >>
rect 16 370 32 386
rect 64 370 80 386
rect 112 370 128 386
rect 160 370 176 386
rect 208 370 224 386
rect 256 370 272 386
<< poly >>
rect 62 318 75 336
rect 113 318 126 336
rect 164 318 177 336
rect 215 318 228 336
rect 62 184 75 206
rect 113 184 126 206
rect 62 176 126 184
rect 62 160 86 176
rect 102 160 126 176
rect 62 153 126 160
rect 62 133 75 153
rect 113 133 126 153
rect 164 184 177 206
rect 215 184 228 206
rect 164 176 228 184
rect 164 160 188 176
rect 204 160 228 176
rect 164 153 228 160
rect 164 133 177 153
rect 215 133 228 153
rect 62 41 75 59
rect 113 41 126 59
rect 164 41 177 59
rect 215 41 228 59
<< polycont >>
rect 86 160 102 176
rect 188 160 204 176
<< metal1 >>
rect 0 386 288 400
rect 0 370 16 386
rect 32 370 64 386
rect 80 370 112 386
rect 128 370 160 386
rect 176 370 208 386
rect 224 370 256 386
rect 272 370 288 386
rect 0 356 288 370
rect 30 311 56 317
rect 30 295 35 311
rect 51 295 56 311
rect 30 275 56 295
rect 30 259 35 275
rect 51 259 56 275
rect 30 236 56 259
rect 81 311 107 356
rect 81 295 86 311
rect 102 295 107 311
rect 81 275 107 295
rect 81 259 86 275
rect 102 259 107 275
rect 81 254 107 259
rect 132 311 260 320
rect 132 295 137 311
rect 153 295 239 311
rect 255 295 260 311
rect 132 286 260 295
rect 132 275 158 286
rect 132 259 137 275
rect 153 259 158 275
rect 234 275 260 286
rect 132 236 158 259
rect 30 229 158 236
rect 30 213 35 229
rect 51 213 137 229
rect 153 213 158 229
rect 30 205 158 213
rect 178 236 213 264
rect 234 259 239 275
rect 255 259 260 275
rect 234 254 260 259
rect 178 229 260 236
rect 178 213 188 229
rect 204 213 260 229
rect 178 205 260 213
rect 77 176 110 182
rect 77 160 86 176
rect 102 160 110 176
rect 77 152 110 160
rect 180 176 212 182
rect 180 160 188 176
rect 204 160 212 176
rect 180 152 212 160
rect 30 126 56 132
rect 234 131 260 205
rect 30 110 35 126
rect 51 110 56 126
rect 30 82 56 110
rect 30 66 35 82
rect 51 66 56 82
rect 30 22 56 66
rect 81 126 260 131
rect 81 110 86 126
rect 102 110 188 126
rect 204 110 260 126
rect 81 107 260 110
rect 81 82 106 107
rect 81 66 86 82
rect 102 66 106 82
rect 81 59 106 66
rect 132 82 158 86
rect 132 66 137 82
rect 153 66 158 82
rect 132 22 158 66
rect 183 82 208 107
rect 183 66 188 82
rect 204 66 208 82
rect 183 59 208 66
rect 234 82 260 86
rect 234 66 239 82
rect 255 66 260 82
rect 234 22 260 66
rect 0 8 288 22
rect 0 -8 16 8
rect 32 -8 64 8
rect 80 -8 112 8
rect 128 -8 160 8
rect 176 -8 208 8
rect 224 -8 256 8
rect 272 -8 288 8
rect 0 -22 288 -8
<< labels >>
flabel metal1 s 77 152 110 182 0 FreeSans 200 0 0 0 A
port 2 nsew
flabel metal1 s 0 356 288 400 0 FreeSans 200 0 0 0 VDD
port 3 nsew
flabel metal1 s 178 205 213 264 0 FreeSans 200 0 0 0 Y
port 4 nsew
flabel metal1 s 0 -22 288 22 0 FreeSans 200 0 0 0 VSS
port 5 nsew
flabel metal1 s 180 152 212 182 0 FreeSans 200 0 0 0 B
port 6 nsew
<< properties >>
string FIXED_BBOX 0 0 288 378
string GDS_END 153712
string GDS_FILE ../gds/controller.gds
string GDS_START 144890
<< end >>
