magic
tech ihp-sg13g2
magscale 1 2
timestamp 1747056038
<< nwell >>
rect -48 350 816 834
<< pwell >>
rect 22 56 746 314
rect -26 -56 794 56
<< nmos >>
rect 116 140 142 288
rect 218 140 244 288
rect 320 140 346 288
rect 524 140 550 288
rect 626 140 652 288
<< pmos >>
rect 116 412 142 636
rect 218 412 244 636
rect 320 412 346 636
rect 524 412 550 636
rect 626 412 652 636
<< ndiff >>
rect 48 274 116 288
rect 48 242 62 274
rect 94 242 116 274
rect 48 186 116 242
rect 48 154 62 186
rect 94 154 116 186
rect 48 140 116 154
rect 142 186 218 288
rect 142 154 164 186
rect 196 154 218 186
rect 142 140 218 154
rect 244 140 320 288
rect 346 186 414 288
rect 346 154 368 186
rect 400 154 414 186
rect 346 140 414 154
rect 456 186 524 288
rect 456 154 470 186
rect 502 154 524 186
rect 456 140 524 154
rect 550 140 626 288
rect 652 186 720 288
rect 652 154 674 186
rect 706 154 720 186
rect 652 140 720 154
<< pdiff >>
rect 48 622 116 636
rect 48 590 62 622
rect 94 590 116 622
rect 48 543 116 590
rect 48 511 62 543
rect 94 511 116 543
rect 48 458 116 511
rect 48 426 62 458
rect 94 426 116 458
rect 48 412 116 426
rect 142 622 218 636
rect 142 590 164 622
rect 196 590 218 622
rect 142 543 218 590
rect 142 511 164 543
rect 196 511 218 543
rect 142 412 218 511
rect 244 543 320 636
rect 244 511 266 543
rect 298 511 320 543
rect 244 412 320 511
rect 346 622 414 636
rect 346 590 368 622
rect 400 590 414 622
rect 346 412 414 590
rect 456 622 524 636
rect 456 590 470 622
rect 502 590 524 622
rect 456 412 524 590
rect 550 622 626 636
rect 550 590 572 622
rect 604 590 626 622
rect 550 543 626 590
rect 550 511 572 543
rect 604 511 626 543
rect 550 412 626 511
rect 652 622 720 636
rect 652 590 674 622
rect 706 590 720 622
rect 652 543 720 590
rect 652 511 674 543
rect 706 511 720 543
rect 652 412 720 511
<< ndiffc >>
rect 62 242 94 274
rect 62 154 94 186
rect 164 154 196 186
rect 368 154 400 186
rect 470 154 502 186
rect 674 154 706 186
<< pdiffc >>
rect 62 590 94 622
rect 62 511 94 543
rect 62 426 94 458
rect 164 590 196 622
rect 164 511 196 543
rect 266 511 298 543
rect 368 590 400 622
rect 470 590 502 622
rect 572 590 604 622
rect 572 511 604 543
rect 674 590 706 622
rect 674 511 706 543
<< psubdiff >>
rect 0 16 768 30
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 608 16
rect 640 -16 704 16
rect 736 -16 768 16
rect 0 -30 768 -16
<< nsubdiff >>
rect 0 772 768 786
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 608 772
rect 640 740 704 772
rect 736 740 768 772
rect 0 726 768 740
<< psubdiffcont >>
rect 32 -16 64 16
rect 128 -16 160 16
rect 224 -16 256 16
rect 320 -16 352 16
rect 416 -16 448 16
rect 512 -16 544 16
rect 608 -16 640 16
rect 704 -16 736 16
<< nsubdiffcont >>
rect 32 740 64 772
rect 128 740 160 772
rect 224 740 256 772
rect 320 740 352 772
rect 416 740 448 772
rect 512 740 544 772
rect 608 740 640 772
rect 704 740 736 772
<< poly >>
rect 116 636 142 672
rect 218 636 244 672
rect 320 636 346 672
rect 524 636 550 672
rect 626 636 652 672
rect 116 380 142 412
rect 218 380 244 412
rect 320 380 346 412
rect 524 380 550 412
rect 626 380 652 412
rect 52 366 142 380
rect 52 334 74 366
rect 106 334 142 366
rect 52 320 142 334
rect 201 366 261 380
rect 201 334 215 366
rect 247 334 261 366
rect 201 320 261 334
rect 320 366 410 380
rect 320 334 355 366
rect 387 334 410 366
rect 320 320 410 334
rect 460 366 550 380
rect 460 334 482 366
rect 514 334 550 366
rect 460 320 550 334
rect 609 366 669 380
rect 609 334 623 366
rect 655 334 669 366
rect 609 320 669 334
rect 116 288 142 320
rect 218 288 244 320
rect 320 288 346 320
rect 524 288 550 320
rect 626 288 652 320
rect 116 104 142 140
rect 218 104 244 140
rect 320 104 346 140
rect 524 104 550 140
rect 626 104 652 140
<< polycont >>
rect 74 334 106 366
rect 215 334 247 366
rect 355 334 387 366
rect 482 334 514 366
rect 623 334 655 366
<< metal1 >>
rect 0 772 768 800
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 608 772
rect 640 740 704 772
rect 736 740 768 772
rect 0 712 768 740
rect 52 622 104 632
rect 52 590 62 622
rect 94 590 104 622
rect 52 543 104 590
rect 52 511 62 543
rect 94 511 104 543
rect 52 458 104 511
rect 154 622 410 632
rect 154 590 164 622
rect 196 590 368 622
rect 400 590 410 622
rect 154 543 206 590
rect 358 580 410 590
rect 460 622 512 712
rect 460 590 470 622
rect 502 590 512 622
rect 460 580 512 590
rect 562 622 614 632
rect 562 590 572 622
rect 604 590 614 622
rect 154 511 164 543
rect 196 511 206 543
rect 154 501 206 511
rect 256 543 308 553
rect 562 543 614 590
rect 256 511 266 543
rect 298 511 572 543
rect 604 511 614 543
rect 256 501 614 511
rect 664 622 716 712
rect 664 590 674 622
rect 706 590 716 622
rect 664 543 716 590
rect 664 511 674 543
rect 706 511 716 543
rect 664 501 716 511
rect 52 426 62 458
rect 94 426 749 458
rect 52 416 749 426
rect 50 366 128 380
rect 50 334 74 366
rect 106 334 128 366
rect 50 314 128 334
rect 176 366 272 380
rect 176 334 215 366
rect 247 334 272 366
rect 176 314 272 334
rect 308 366 400 380
rect 308 334 355 366
rect 387 334 400 366
rect 308 314 400 334
rect 52 242 62 274
rect 94 242 308 274
rect 52 232 308 242
rect 344 232 400 314
rect 436 366 540 380
rect 436 334 482 366
rect 514 334 540 366
rect 436 314 540 334
rect 576 366 677 380
rect 576 334 623 366
rect 655 334 677 366
rect 576 314 677 334
rect 436 232 496 314
rect 713 274 749 416
rect 562 232 749 274
rect 52 186 104 232
rect 256 196 308 232
rect 562 196 614 232
rect 52 154 62 186
rect 94 154 104 186
rect 52 144 104 154
rect 154 186 206 196
rect 154 154 164 186
rect 196 154 206 186
rect 154 44 206 154
rect 256 186 614 196
rect 256 154 368 186
rect 400 154 470 186
rect 502 154 614 186
rect 256 144 614 154
rect 664 186 716 196
rect 664 154 674 186
rect 706 154 716 186
rect 664 44 716 154
rect 0 16 768 44
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 608 16
rect 640 -16 704 16
rect 736 -16 768 16
rect 0 -44 768 -16
<< labels >>
flabel metal1 s 0 -44 768 44 0 FreeSans 400 0 0 0 VSS
port 3 nsew
flabel metal1 s 0 712 768 800 0 FreeSans 400 0 0 0 VDD
port 5 nsew
flabel metal1 s 50 314 128 380 0 FreeSans 400 0 0 0 C1
port 6 nsew
flabel metal1 s 713 232 749 458 0 FreeSans 400 0 0 0 Y
port 7 nsew
flabel metal1 s 176 314 272 380 0 FreeSans 400 0 0 0 B2
port 8 nsew
flabel metal1 s 344 232 400 380 0 FreeSans 400 0 0 0 B1
port 9 nsew
flabel metal1 s 576 314 677 380 0 FreeSans 400 0 0 0 A2
port 10 nsew
flabel metal1 s 436 232 496 380 0 FreeSans 400 0 0 0 A1
port 11 nsew
<< properties >>
string FIXED_BBOX 0 0 768 756
string GDS_END 127946
string GDS_FILE ../gds/controller.gds
string GDS_START 122234
<< end >>
