magic
tech ihp-sg13g2
timestamp 1747537721
<< nwell >>
rect -24 175 360 417
<< pwell >>
rect 90 142 332 157
rect 79 28 332 142
rect -13 -28 349 28
<< nmos >>
rect 126 70 139 144
rect 183 80 196 144
rect 234 80 247 144
rect 272 80 285 144
<< pmos >>
rect 62 206 75 318
rect 166 218 179 318
rect 221 218 234 318
rect 272 218 285 318
<< ndiff >>
rect 103 129 126 144
rect 92 109 126 129
rect 92 93 99 109
rect 115 93 126 109
rect 92 70 126 93
rect 139 94 183 144
rect 139 78 150 94
rect 166 80 183 94
rect 196 104 234 144
rect 196 88 207 104
rect 223 88 234 104
rect 196 80 234 88
rect 247 80 272 144
rect 285 135 319 144
rect 285 119 296 135
rect 312 119 319 135
rect 285 80 319 119
rect 166 78 176 80
rect 139 70 176 78
<< pdiff >>
rect 28 309 62 318
rect 28 293 35 309
rect 51 293 62 309
rect 28 270 62 293
rect 28 254 35 270
rect 51 254 62 270
rect 28 231 62 254
rect 28 215 35 231
rect 51 215 62 231
rect 28 206 62 215
rect 75 309 109 318
rect 75 293 86 309
rect 102 293 109 309
rect 75 270 109 293
rect 75 254 86 270
rect 102 254 109 270
rect 75 231 109 254
rect 75 215 86 231
rect 102 215 109 231
rect 131 311 166 318
rect 131 295 138 311
rect 154 295 166 311
rect 131 276 166 295
rect 131 260 138 276
rect 154 260 166 276
rect 131 241 166 260
rect 131 225 138 241
rect 154 225 166 241
rect 131 218 166 225
rect 179 311 221 318
rect 179 295 190 311
rect 206 295 221 311
rect 179 276 221 295
rect 179 260 190 276
rect 206 260 221 276
rect 179 241 221 260
rect 179 225 190 241
rect 206 225 221 241
rect 179 218 221 225
rect 234 311 272 318
rect 234 295 245 311
rect 261 295 272 311
rect 234 275 272 295
rect 234 259 245 275
rect 261 259 272 275
rect 234 218 272 259
rect 285 311 319 318
rect 285 295 296 311
rect 312 295 319 311
rect 285 276 319 295
rect 285 260 296 276
rect 312 260 319 276
rect 285 241 319 260
rect 285 225 296 241
rect 312 225 319 241
rect 285 218 319 225
rect 75 206 109 215
<< ndiffc >>
rect 99 93 115 109
rect 150 78 166 94
rect 207 88 223 104
rect 296 119 312 135
<< pdiffc >>
rect 35 293 51 309
rect 35 254 51 270
rect 35 215 51 231
rect 86 293 102 309
rect 86 254 102 270
rect 86 215 102 231
rect 138 295 154 311
rect 138 260 154 276
rect 138 225 154 241
rect 190 295 206 311
rect 190 260 206 276
rect 190 225 206 241
rect 245 295 261 311
rect 245 259 261 275
rect 296 295 312 311
rect 296 260 312 276
rect 296 225 312 241
<< psubdiff >>
rect 0 8 336 15
rect 0 -8 16 8
rect 32 -8 64 8
rect 80 -8 112 8
rect 128 -8 160 8
rect 176 -8 208 8
rect 224 -8 256 8
rect 272 -8 304 8
rect 320 -8 336 8
rect 0 -15 336 -8
<< nsubdiff >>
rect 0 386 336 393
rect 0 370 16 386
rect 32 370 64 386
rect 80 370 112 386
rect 128 370 160 386
rect 176 370 208 386
rect 224 370 256 386
rect 272 370 304 386
rect 320 370 336 386
rect 0 363 336 370
<< psubdiffcont >>
rect 16 -8 32 8
rect 64 -8 80 8
rect 112 -8 128 8
rect 160 -8 176 8
rect 208 -8 224 8
rect 256 -8 272 8
rect 304 -8 320 8
<< nsubdiffcont >>
rect 16 370 32 386
rect 64 370 80 386
rect 112 370 128 386
rect 160 370 176 386
rect 208 370 224 386
rect 256 370 272 386
rect 304 370 320 386
<< poly >>
rect 62 318 75 336
rect 166 318 179 336
rect 221 318 234 336
rect 272 318 285 336
rect 166 210 179 218
rect 62 187 75 206
rect 166 191 200 210
rect 57 178 92 187
rect 57 162 68 178
rect 84 176 92 178
rect 84 162 139 176
rect 166 175 176 191
rect 192 175 200 191
rect 166 167 200 175
rect 221 200 234 218
rect 221 191 254 200
rect 221 175 230 191
rect 246 175 254 191
rect 221 167 254 175
rect 57 161 139 162
rect 57 154 92 161
rect 126 144 139 161
rect 183 144 196 167
rect 234 144 247 167
rect 272 144 285 218
rect 126 52 139 70
rect 183 62 196 80
rect 234 62 247 80
rect 272 70 285 80
rect 272 61 314 70
rect 272 45 290 61
rect 306 45 314 61
rect 272 37 314 45
<< polycont >>
rect 68 162 84 178
rect 176 175 192 191
rect 230 175 246 191
rect 290 45 306 61
<< metal1 >>
rect 0 386 336 400
rect 0 370 16 386
rect 32 370 64 386
rect 80 370 112 386
rect 128 370 160 386
rect 176 370 208 386
rect 224 370 256 386
rect 272 370 304 386
rect 320 370 336 386
rect 0 356 336 370
rect 20 309 56 310
rect 20 293 35 309
rect 51 293 56 309
rect 20 270 56 293
rect 20 254 35 270
rect 51 254 56 270
rect 20 231 56 254
rect 20 215 35 231
rect 51 215 56 231
rect 20 209 56 215
rect 81 309 107 356
rect 81 293 86 309
rect 102 293 107 309
rect 81 270 107 293
rect 81 254 86 270
rect 102 254 107 270
rect 81 231 107 254
rect 81 215 86 231
rect 102 215 107 231
rect 81 214 107 215
rect 133 311 159 312
rect 133 295 138 311
rect 154 295 159 311
rect 133 276 159 295
rect 133 260 138 276
rect 154 260 159 276
rect 133 241 159 260
rect 133 225 138 241
rect 154 225 159 241
rect 133 217 159 225
rect 185 311 211 312
rect 185 295 190 311
rect 206 295 211 311
rect 185 276 211 295
rect 185 260 190 276
rect 206 260 211 276
rect 185 241 211 260
rect 240 311 266 356
rect 240 295 245 311
rect 261 295 266 311
rect 240 275 266 295
rect 240 259 245 275
rect 261 259 266 275
rect 240 258 266 259
rect 291 311 317 312
rect 291 295 296 311
rect 312 295 317 311
rect 291 276 317 295
rect 291 260 296 276
rect 312 260 317 276
rect 185 225 190 241
rect 206 240 211 241
rect 291 241 317 260
rect 291 240 296 241
rect 206 225 296 240
rect 312 225 317 241
rect 185 221 317 225
rect 20 114 44 209
rect 133 187 157 217
rect 62 178 157 187
rect 62 162 68 178
rect 84 162 157 178
rect 62 154 157 162
rect 175 191 200 200
rect 175 175 176 191
rect 192 175 200 191
rect 175 157 200 175
rect 221 191 254 200
rect 221 175 230 191
rect 246 175 254 191
rect 221 156 254 175
rect 141 138 157 154
rect 141 122 227 138
rect 292 135 316 141
rect 292 131 296 135
rect 20 109 122 114
rect 20 93 99 109
rect 115 93 122 109
rect 202 104 227 122
rect 20 88 122 93
rect 145 94 171 96
rect 145 78 150 94
rect 166 78 171 94
rect 202 88 207 104
rect 223 88 227 104
rect 202 82 227 88
rect 245 119 296 131
rect 312 119 316 135
rect 245 114 316 119
rect 145 22 171 78
rect 245 22 261 114
rect 281 61 321 96
rect 281 45 290 61
rect 306 45 321 61
rect 281 40 321 45
rect 0 8 336 22
rect 0 -8 16 8
rect 32 -8 64 8
rect 80 -8 112 8
rect 128 -8 160 8
rect 176 -8 208 8
rect 224 -8 256 8
rect 272 -8 304 8
rect 320 -8 336 8
rect 0 -22 336 -8
<< labels >>
flabel metal1 s 175 157 200 200 0 FreeSans 200 0 0 0 B1
port 2 nsew
flabel metal1 s 28 209 56 310 0 FreeSans 200 0 0 0 X
port 3 nsew
flabel metal1 s 0 356 336 400 0 FreeSans 200 0 0 0 VDD
port 4 nsew
flabel metal1 s 0 -22 336 22 0 FreeSans 200 0 0 0 VSS
port 5 nsew
flabel metal1 s 221 156 254 200 0 FreeSans 200 0 0 0 A1
port 6 nsew
flabel metal1 s 281 40 321 96 0 FreeSans 200 0 0 0 A2
port 7 nsew
<< properties >>
string FIXED_BBOX 0 0 336 378
string GDS_END 89618
string GDS_FILE ../gds/controller.gds
string GDS_START 84462
<< end >>
