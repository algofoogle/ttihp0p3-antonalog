magic
tech ihp-sg13g2
magscale 1 2
timestamp 1747537721
<< nwell >>
rect -48 350 528 834
<< pwell >>
rect 16 56 465 296
rect -26 -56 506 56
<< nmos >>
rect 120 122 146 270
rect 239 122 265 270
rect 324 122 350 270
<< pmos >>
rect 120 426 146 650
rect 222 426 248 650
rect 324 426 350 650
<< ndiff >>
rect 42 182 120 270
rect 42 150 56 182
rect 88 150 120 182
rect 42 122 120 150
rect 146 122 239 270
rect 265 122 324 270
rect 350 252 439 270
rect 350 220 385 252
rect 417 220 439 252
rect 350 171 439 220
rect 350 139 372 171
rect 404 139 439 171
rect 350 122 439 139
<< pdiff >>
rect 52 635 120 650
rect 52 603 66 635
rect 98 603 120 635
rect 52 565 120 603
rect 52 533 66 565
rect 98 533 120 565
rect 52 481 120 533
rect 52 449 66 481
rect 98 449 120 481
rect 52 426 120 449
rect 146 635 222 650
rect 146 603 168 635
rect 200 603 222 635
rect 146 567 222 603
rect 146 535 168 567
rect 200 535 222 567
rect 146 497 222 535
rect 146 465 168 497
rect 200 465 222 497
rect 146 426 222 465
rect 248 635 324 650
rect 248 603 270 635
rect 302 603 324 635
rect 248 565 324 603
rect 248 533 270 565
rect 302 533 324 565
rect 248 426 324 533
rect 350 635 418 650
rect 350 603 372 635
rect 404 603 418 635
rect 350 554 418 603
rect 350 522 372 554
rect 404 522 418 554
rect 350 475 418 522
rect 350 443 372 475
rect 404 443 418 475
rect 350 426 418 443
<< ndiffc >>
rect 56 150 88 182
rect 385 220 417 252
rect 372 139 404 171
<< pdiffc >>
rect 66 603 98 635
rect 66 533 98 565
rect 66 449 98 481
rect 168 603 200 635
rect 168 535 200 567
rect 168 465 200 497
rect 270 603 302 635
rect 270 533 302 565
rect 372 603 404 635
rect 372 522 404 554
rect 372 443 404 475
<< psubdiff >>
rect 0 16 480 30
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 480 16
rect 0 -30 480 -16
<< nsubdiff >>
rect 0 772 480 786
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 480 772
rect 0 726 480 740
<< psubdiffcont >>
rect 32 -16 64 16
rect 128 -16 160 16
rect 224 -16 256 16
rect 320 -16 352 16
rect 416 -16 448 16
<< nsubdiffcont >>
rect 32 740 64 772
rect 128 740 160 772
rect 224 740 256 772
rect 320 740 352 772
rect 416 740 448 772
<< poly >>
rect 120 650 146 686
rect 222 650 248 686
rect 324 650 350 686
rect 120 374 146 426
rect 222 380 248 426
rect 72 360 146 374
rect 72 328 86 360
rect 118 328 146 360
rect 72 314 146 328
rect 205 363 265 380
rect 324 371 350 426
rect 205 331 219 363
rect 251 331 265 363
rect 205 317 265 331
rect 120 270 146 314
rect 239 270 265 317
rect 301 357 375 371
rect 301 325 320 357
rect 352 325 375 357
rect 301 311 375 325
rect 324 270 350 311
rect 120 86 146 122
rect 239 86 265 122
rect 324 86 350 122
<< polycont >>
rect 86 328 118 360
rect 219 331 251 363
rect 320 325 352 357
<< metal1 >>
rect 0 772 480 800
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 480 772
rect 0 712 480 740
rect 56 635 108 712
rect 56 603 66 635
rect 98 603 108 635
rect 56 565 108 603
rect 56 533 66 565
rect 98 533 108 565
rect 56 481 108 533
rect 56 449 66 481
rect 98 449 108 481
rect 56 434 108 449
rect 158 635 210 640
rect 158 603 168 635
rect 200 603 210 635
rect 158 567 210 603
rect 158 535 168 567
rect 200 535 210 567
rect 158 497 210 535
rect 260 635 312 712
rect 260 603 270 635
rect 302 603 312 635
rect 260 565 312 603
rect 260 533 270 565
rect 302 533 312 565
rect 260 515 312 533
rect 356 635 452 654
rect 356 603 372 635
rect 404 603 452 635
rect 356 554 452 603
rect 356 522 372 554
rect 404 522 452 554
rect 158 465 168 497
rect 200 479 210 497
rect 356 479 452 522
rect 200 475 452 479
rect 200 465 372 475
rect 158 443 372 465
rect 404 443 452 475
rect 158 436 452 443
rect 356 434 452 436
rect 72 360 138 397
rect 72 328 86 360
rect 118 328 138 360
rect 72 314 138 328
rect 190 363 265 400
rect 190 331 219 363
rect 251 331 265 363
rect 190 314 265 331
rect 307 357 374 398
rect 307 325 320 357
rect 352 325 374 357
rect 307 310 374 325
rect 410 272 452 434
rect 374 252 452 272
rect 374 220 385 252
rect 417 220 452 252
rect 374 202 452 220
rect 45 182 99 192
rect 45 150 56 182
rect 88 150 99 182
rect 45 44 99 150
rect 354 171 452 202
rect 354 139 372 171
rect 404 139 452 171
rect 354 124 452 139
rect 0 16 480 44
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 480 16
rect 0 -44 480 -16
<< labels >>
flabel metal1 s 0 712 480 800 0 FreeSans 400 0 0 0 VDD
port 2 nsew
flabel metal1 s 356 434 452 654 0 FreeSans 400 0 0 0 Y
port 3 nsew
flabel metal1 s 190 314 265 400 0 FreeSans 400 0 0 0 B
port 4 nsew
flabel metal1 s 72 314 138 397 0 FreeSans 400 0 0 0 C
port 5 nsew
flabel metal1 s 0 -44 480 44 0 FreeSans 400 0 0 0 VSS
port 6 nsew
flabel metal1 s 307 310 374 398 0 FreeSans 400 0 0 0 A
port 7 nsew
<< properties >>
string FIXED_BBOX 0 0 480 756
string GDS_END 122778
string GDS_FILE ../gds/controller.gds
string GDS_START 118150
<< end >>
