magic
tech ihp-sg13g2
magscale 1 2
timestamp 1746816402
<< nwell >>
rect -48 350 816 834
<< pwell >>
rect 21 56 772 304
rect -26 -56 794 56
<< nmos >>
rect 183 168 209 278
rect 336 168 362 278
rect 448 130 474 278
rect 522 130 548 278
rect 636 130 662 278
<< pmos >>
rect 151 436 177 636
rect 226 436 252 636
rect 448 412 474 636
rect 550 412 576 636
rect 652 412 678 636
<< ndiff >>
rect 47 224 183 278
rect 47 192 61 224
rect 93 192 129 224
rect 161 192 183 224
rect 47 168 183 192
rect 209 234 336 278
rect 209 202 231 234
rect 263 202 336 234
rect 209 168 336 202
rect 362 264 448 278
rect 362 232 390 264
rect 422 232 448 264
rect 362 177 448 232
rect 362 168 390 177
rect 376 145 390 168
rect 422 145 448 177
rect 376 130 448 145
rect 474 130 522 278
rect 548 256 636 278
rect 548 224 577 256
rect 609 224 636 256
rect 548 177 636 224
rect 548 145 577 177
rect 609 145 636 177
rect 548 130 636 145
rect 662 177 746 278
rect 662 145 684 177
rect 716 145 746 177
rect 662 130 746 145
<< pdiff >>
rect 79 621 151 636
rect 79 589 97 621
rect 129 589 151 621
rect 79 551 151 589
rect 79 519 97 551
rect 129 519 151 551
rect 79 482 151 519
rect 79 450 97 482
rect 129 450 151 482
rect 79 436 151 450
rect 177 436 226 636
rect 252 621 320 636
rect 252 589 274 621
rect 306 589 320 621
rect 252 552 320 589
rect 252 520 274 552
rect 306 520 320 552
rect 252 482 320 520
rect 252 450 274 482
rect 306 450 320 482
rect 252 436 320 450
rect 380 621 448 636
rect 380 589 394 621
rect 426 589 448 621
rect 380 550 448 589
rect 380 518 394 550
rect 426 518 448 550
rect 380 412 448 518
rect 474 621 550 636
rect 474 589 496 621
rect 528 589 550 621
rect 474 412 550 589
rect 576 621 652 636
rect 576 589 598 621
rect 630 589 652 621
rect 576 550 652 589
rect 576 518 598 550
rect 630 518 652 550
rect 576 412 652 518
rect 678 621 746 636
rect 678 589 700 621
rect 732 589 746 621
rect 678 551 746 589
rect 678 519 700 551
rect 732 519 746 551
rect 678 476 746 519
rect 678 444 700 476
rect 732 444 746 476
rect 678 412 746 444
<< ndiffc >>
rect 61 192 93 224
rect 129 192 161 224
rect 231 202 263 234
rect 390 232 422 264
rect 390 145 422 177
rect 577 224 609 256
rect 577 145 609 177
rect 684 145 716 177
<< pdiffc >>
rect 97 589 129 621
rect 97 519 129 551
rect 97 450 129 482
rect 274 589 306 621
rect 274 520 306 552
rect 274 450 306 482
rect 394 589 426 621
rect 394 518 426 550
rect 496 589 528 621
rect 598 589 630 621
rect 598 518 630 550
rect 700 589 732 621
rect 700 519 732 551
rect 700 444 732 476
<< psubdiff >>
rect 0 16 768 30
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 608 16
rect 640 -16 704 16
rect 736 -16 768 16
rect 0 -30 768 -16
<< nsubdiff >>
rect 0 772 768 786
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 608 772
rect 640 740 704 772
rect 736 740 768 772
rect 0 726 768 740
<< psubdiffcont >>
rect 32 -16 64 16
rect 128 -16 160 16
rect 224 -16 256 16
rect 320 -16 352 16
rect 416 -16 448 16
rect 512 -16 544 16
rect 608 -16 640 16
rect 704 -16 736 16
<< nsubdiffcont >>
rect 32 740 64 772
rect 128 740 160 772
rect 224 740 256 772
rect 320 740 352 772
rect 416 740 448 772
rect 512 740 544 772
rect 608 740 640 772
rect 704 740 736 772
<< poly >>
rect 151 636 177 673
rect 226 636 252 673
rect 448 636 474 673
rect 550 636 576 673
rect 652 636 678 673
rect 151 366 177 436
rect 226 412 252 436
rect 226 382 362 412
rect 448 396 474 412
rect 40 349 177 366
rect 40 317 54 349
rect 86 317 122 349
rect 154 330 177 349
rect 276 365 362 382
rect 276 333 310 365
rect 342 333 362 365
rect 154 317 209 330
rect 40 300 209 317
rect 276 316 362 333
rect 183 278 209 300
rect 336 278 362 316
rect 438 293 474 396
rect 550 396 576 412
rect 550 379 588 396
rect 448 278 474 293
rect 522 362 588 379
rect 652 373 678 412
rect 522 330 536 362
rect 568 330 588 362
rect 522 313 588 330
rect 624 356 690 373
rect 624 324 638 356
rect 670 324 690 356
rect 522 278 548 313
rect 624 307 690 324
rect 636 278 662 307
rect 183 94 209 168
rect 336 132 362 168
rect 448 94 474 130
rect 522 94 548 130
rect 636 94 662 130
rect 183 64 474 94
<< polycont >>
rect 54 317 86 349
rect 122 317 154 349
rect 310 333 342 365
rect 536 330 568 362
rect 638 324 670 356
<< metal1 >>
rect 0 772 768 800
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 608 772
rect 640 740 704 772
rect 736 740 768 772
rect 0 712 768 740
rect 87 621 139 712
rect 87 589 97 621
rect 129 589 139 621
rect 87 551 139 589
rect 87 519 97 551
rect 129 519 139 551
rect 87 482 139 519
rect 87 450 97 482
rect 129 450 139 482
rect 87 446 139 450
rect 206 621 310 631
rect 206 589 274 621
rect 306 589 310 621
rect 206 552 310 589
rect 206 520 274 552
rect 306 520 310 552
rect 206 482 310 520
rect 384 621 436 631
rect 384 589 394 621
rect 426 589 436 621
rect 384 550 436 589
rect 486 621 538 712
rect 486 589 496 621
rect 528 589 538 621
rect 486 579 538 589
rect 588 621 640 632
rect 588 589 598 621
rect 630 589 640 621
rect 384 518 394 550
rect 426 536 436 550
rect 588 550 640 589
rect 588 536 598 550
rect 426 518 598 536
rect 630 518 640 550
rect 384 504 640 518
rect 690 621 742 632
rect 690 589 700 621
rect 732 589 742 621
rect 690 551 742 589
rect 690 519 700 551
rect 732 519 742 551
rect 206 450 274 482
rect 306 468 310 482
rect 690 476 742 519
rect 306 450 654 468
rect 206 434 654 450
rect 29 349 164 383
rect 29 317 54 349
rect 86 317 122 349
rect 154 317 164 349
rect 29 290 164 317
rect 206 252 240 434
rect 622 374 654 434
rect 690 444 700 476
rect 732 444 742 476
rect 690 431 742 444
rect 295 365 586 374
rect 295 333 310 365
rect 342 362 586 365
rect 342 333 536 362
rect 295 330 536 333
rect 568 330 586 362
rect 295 307 586 330
rect 622 356 670 374
rect 622 324 638 356
rect 622 308 670 324
rect 380 264 432 268
rect 57 224 164 236
rect 57 192 61 224
rect 93 192 129 224
rect 161 192 164 224
rect 57 44 164 192
rect 206 234 280 252
rect 206 202 231 234
rect 263 202 280 234
rect 206 186 280 202
rect 380 232 390 264
rect 422 232 432 264
rect 706 263 742 431
rect 380 177 432 232
rect 380 145 390 177
rect 422 145 432 177
rect 380 44 432 145
rect 567 256 742 263
rect 567 224 577 256
rect 609 224 742 256
rect 567 221 742 224
rect 567 177 620 221
rect 567 145 577 177
rect 609 145 620 177
rect 567 134 620 145
rect 674 177 726 181
rect 674 145 684 177
rect 716 145 726 177
rect 674 44 726 145
rect 0 16 768 44
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 608 16
rect 640 -16 704 16
rect 736 -16 768 16
rect 0 -44 768 -16
<< labels >>
flabel metal1 s 690 431 742 632 0 FreeSans 400 0 0 0 X
port 2 nsew
flabel metal1 s 0 712 768 800 0 FreeSans 400 0 0 0 VDD
port 3 nsew
flabel metal1 s 295 307 586 374 0 FreeSans 400 0 0 0 B
port 4 nsew
flabel metal1 s 29 290 164 383 0 FreeSans 400 0 0 0 A
port 5 nsew
flabel metal1 s 0 -44 768 44 0 FreeSans 400 0 0 0 VSS
port 6 nsew
<< properties >>
string FIXED_BBOX 0 0 768 756
string GDS_END 92314
string GDS_FILE ../gds/controller.gds
string GDS_START 86964
<< end >>
