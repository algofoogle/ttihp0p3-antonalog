magic
tech ihp-sg13g2
magscale 1 2
timestamp 1747539407
<< metal1 >>
rect 576 27992 31392 28016
rect 576 27952 4352 27992
rect 4720 27952 12126 27992
rect 12494 27952 19900 27992
rect 20268 27952 27674 27992
rect 28042 27952 31392 27992
rect 576 27928 31392 27952
rect 11194 27740 11252 27741
rect 11194 27700 11203 27740
rect 11243 27700 11252 27740
rect 11194 27699 11252 27700
rect 22330 27740 22388 27741
rect 22330 27700 22339 27740
rect 22379 27700 22388 27740
rect 22330 27699 22388 27700
rect 25114 27740 25172 27741
rect 25114 27700 25123 27740
rect 25163 27700 25172 27740
rect 25114 27699 25172 27700
rect 25498 27740 25556 27741
rect 25498 27700 25507 27740
rect 25547 27700 25556 27740
rect 25498 27699 25556 27700
rect 3610 27656 3668 27657
rect 3610 27616 3619 27656
rect 3659 27616 3668 27656
rect 3610 27615 3668 27616
rect 6106 27656 6164 27657
rect 6106 27616 6115 27656
rect 6155 27616 6164 27656
rect 6106 27615 6164 27616
rect 8602 27656 8660 27657
rect 8602 27616 8611 27656
rect 8651 27616 8660 27656
rect 8602 27615 8660 27616
rect 11578 27656 11636 27657
rect 11578 27616 11587 27656
rect 11627 27616 11636 27656
rect 11578 27615 11636 27616
rect 14187 27656 14229 27665
rect 14187 27616 14188 27656
rect 14228 27616 14229 27656
rect 14187 27607 14229 27616
rect 16378 27656 16436 27657
rect 16378 27616 16387 27656
rect 16427 27616 16436 27656
rect 16378 27615 16436 27616
rect 17067 27656 17109 27665
rect 17067 27616 17068 27656
rect 17108 27616 17109 27656
rect 17067 27607 17109 27616
rect 18106 27656 18164 27657
rect 18106 27616 18115 27656
rect 18155 27616 18164 27656
rect 18106 27615 18164 27616
rect 22714 27656 22772 27657
rect 22714 27616 22723 27656
rect 22763 27616 22772 27656
rect 22714 27615 22772 27616
rect 25035 27656 25077 27665
rect 25035 27616 25036 27656
rect 25076 27616 25077 27656
rect 25035 27607 25077 27616
rect 25210 27656 25268 27657
rect 25210 27616 25219 27656
rect 25259 27616 25268 27656
rect 25210 27615 25268 27616
rect 25323 27656 25365 27665
rect 25323 27616 25324 27656
rect 25364 27616 25365 27656
rect 25323 27607 25365 27616
rect 25882 27656 25940 27657
rect 25882 27616 25891 27656
rect 25931 27616 25940 27656
rect 25882 27615 25940 27616
rect 28011 27656 28053 27665
rect 28011 27616 28012 27656
rect 28052 27616 28053 27656
rect 28011 27607 28053 27616
rect 28866 27647 28912 27656
rect 28866 27607 28867 27647
rect 28907 27607 28912 27647
rect 28866 27598 28912 27607
rect 29346 27647 29392 27656
rect 29346 27607 29347 27647
rect 29387 27607 29392 27647
rect 29346 27598 29392 27607
rect 29826 27647 29872 27656
rect 29826 27607 29827 27647
rect 29867 27607 29872 27647
rect 29826 27598 29872 27607
rect 3243 27572 3285 27581
rect 3243 27532 3244 27572
rect 3284 27532 3285 27572
rect 3243 27523 3285 27532
rect 5739 27572 5781 27581
rect 5739 27532 5740 27572
rect 5780 27532 5781 27572
rect 5739 27523 5781 27532
rect 8235 27572 8277 27581
rect 8235 27532 8236 27572
rect 8276 27532 8277 27572
rect 8235 27523 8277 27532
rect 16762 27572 16820 27573
rect 16762 27532 16771 27572
rect 16811 27532 16820 27572
rect 16762 27531 16820 27532
rect 17739 27572 17781 27581
rect 17739 27532 17740 27572
rect 17780 27532 17781 27572
rect 17739 27523 17781 27532
rect 29019 27572 29061 27581
rect 29019 27532 29020 27572
rect 29060 27532 29061 27572
rect 29019 27523 29061 27532
rect 29499 27572 29541 27581
rect 29499 27532 29500 27572
rect 29540 27532 29541 27572
rect 29499 27523 29541 27532
rect 29979 27572 30021 27581
rect 29979 27532 29980 27572
rect 30020 27532 30021 27572
rect 29979 27523 30021 27532
rect 30891 27572 30933 27581
rect 30891 27532 30892 27572
rect 30932 27532 30933 27572
rect 30891 27523 30933 27532
rect 3051 27488 3093 27497
rect 3051 27448 3052 27488
rect 3092 27448 3093 27488
rect 3051 27439 3093 27448
rect 13707 27488 13749 27497
rect 13707 27448 13708 27488
rect 13748 27448 13749 27488
rect 13707 27439 13749 27448
rect 20235 27488 20277 27497
rect 20235 27448 20236 27488
rect 20276 27448 20277 27488
rect 20235 27439 20277 27448
rect 20811 27488 20853 27497
rect 20811 27448 20812 27488
rect 20852 27448 20853 27488
rect 20811 27439 20853 27448
rect 30315 27488 30357 27497
rect 30315 27448 30316 27488
rect 30356 27448 30357 27488
rect 30315 27439 30357 27448
rect 31083 27488 31125 27497
rect 31083 27448 31084 27488
rect 31124 27448 31125 27488
rect 31083 27439 31125 27448
rect 5547 27404 5589 27413
rect 5547 27364 5548 27404
rect 5588 27364 5589 27404
rect 5547 27355 5589 27364
rect 8043 27404 8085 27413
rect 8043 27364 8044 27404
rect 8084 27364 8085 27404
rect 8043 27355 8085 27364
rect 10539 27404 10581 27413
rect 10539 27364 10540 27404
rect 10580 27364 10581 27404
rect 10539 27355 10581 27364
rect 13515 27404 13557 27413
rect 13515 27364 13516 27404
rect 13556 27364 13557 27404
rect 13515 27355 13557 27364
rect 14043 27404 14085 27413
rect 14043 27364 14044 27404
rect 14084 27364 14085 27404
rect 14043 27355 14085 27364
rect 14475 27404 14517 27413
rect 14475 27364 14476 27404
rect 14516 27364 14517 27404
rect 14475 27355 14517 27364
rect 16923 27404 16965 27413
rect 16923 27364 16924 27404
rect 16964 27364 16965 27404
rect 16923 27355 16965 27364
rect 20043 27404 20085 27413
rect 20043 27364 20044 27404
rect 20084 27364 20085 27404
rect 20043 27355 20085 27364
rect 24651 27404 24693 27413
rect 24651 27364 24652 27404
rect 24692 27364 24693 27404
rect 24651 27355 24693 27364
rect 27819 27404 27861 27413
rect 27819 27364 27820 27404
rect 27860 27364 27861 27404
rect 27819 27355 27861 27364
rect 28683 27404 28725 27413
rect 28683 27364 28684 27404
rect 28724 27364 28725 27404
rect 28683 27355 28725 27364
rect 30651 27404 30693 27413
rect 30651 27364 30652 27404
rect 30692 27364 30693 27404
rect 30651 27355 30693 27364
rect 576 27236 31392 27260
rect 576 27196 3112 27236
rect 3480 27196 10886 27236
rect 11254 27196 18660 27236
rect 19028 27196 26434 27236
rect 26802 27196 31392 27236
rect 576 27172 31392 27196
rect 11691 27068 11733 27077
rect 11691 27028 11692 27068
rect 11732 27028 11733 27068
rect 11691 27019 11733 27028
rect 14074 27068 14132 27069
rect 14074 27028 14083 27068
rect 14123 27028 14132 27068
rect 14074 27027 14132 27028
rect 16779 27068 16821 27077
rect 16779 27028 16780 27068
rect 16820 27028 16821 27068
rect 16779 27019 16821 27028
rect 17931 27068 17973 27077
rect 17931 27028 17932 27068
rect 17972 27028 17973 27068
rect 17931 27019 17973 27028
rect 26842 27068 26900 27069
rect 26842 27028 26851 27068
rect 26891 27028 26900 27068
rect 26842 27027 26900 27028
rect 2763 26984 2805 26993
rect 2763 26944 2764 26984
rect 2804 26944 2805 26984
rect 2763 26935 2805 26944
rect 3147 26984 3189 26993
rect 3147 26944 3148 26984
rect 3188 26944 3189 26984
rect 3147 26935 3189 26944
rect 3531 26984 3573 26993
rect 3531 26944 3532 26984
rect 3572 26944 3573 26984
rect 3531 26935 3573 26944
rect 3723 26984 3765 26993
rect 3723 26944 3724 26984
rect 3764 26944 3765 26984
rect 3723 26935 3765 26944
rect 5451 26984 5493 26993
rect 5451 26944 5452 26984
rect 5492 26944 5493 26984
rect 5451 26935 5493 26944
rect 6699 26984 6741 26993
rect 6699 26944 6700 26984
rect 6740 26944 6741 26984
rect 6699 26935 6741 26944
rect 9291 26984 9333 26993
rect 9291 26944 9292 26984
rect 9332 26944 9333 26984
rect 9291 26935 9333 26944
rect 11883 26984 11925 26993
rect 11883 26944 11884 26984
rect 11924 26944 11925 26984
rect 11883 26935 11925 26944
rect 13707 26984 13749 26993
rect 13707 26944 13708 26984
rect 13748 26944 13749 26984
rect 13707 26935 13749 26944
rect 15723 26984 15765 26993
rect 15723 26944 15724 26984
rect 15764 26944 15765 26984
rect 15723 26935 15765 26944
rect 17739 26984 17781 26993
rect 17739 26944 17740 26984
rect 17780 26944 17781 26984
rect 17739 26935 17781 26944
rect 24459 26984 24501 26993
rect 24459 26944 24460 26984
rect 24500 26944 24501 26984
rect 24459 26935 24501 26944
rect 27819 26984 27861 26993
rect 27819 26944 27820 26984
rect 27860 26944 27861 26984
rect 27819 26935 27861 26944
rect 8475 26900 8517 26909
rect 8475 26860 8476 26900
rect 8516 26860 8517 26900
rect 8475 26851 8517 26860
rect 15243 26900 15285 26909
rect 15243 26860 15244 26900
rect 15284 26860 15285 26900
rect 15243 26851 15285 26860
rect 23307 26900 23349 26909
rect 23307 26860 23308 26900
rect 23348 26860 23349 26900
rect 23307 26851 23349 26860
rect 24826 26900 24884 26901
rect 24826 26860 24835 26900
rect 24875 26860 24884 26900
rect 24826 26859 24884 26860
rect 28954 26900 29012 26901
rect 28954 26860 28963 26900
rect 29003 26860 29012 26900
rect 28954 26859 29012 26860
rect 3723 26816 3765 26825
rect 3723 26776 3724 26816
rect 3764 26776 3765 26816
rect 3723 26767 3765 26776
rect 3915 26816 3957 26825
rect 3915 26776 3916 26816
rect 3956 26776 3957 26816
rect 3915 26767 3957 26776
rect 6315 26816 6357 26825
rect 6315 26776 6316 26816
rect 6356 26776 6357 26816
rect 6315 26767 6357 26776
rect 7467 26816 7509 26825
rect 7467 26776 7468 26816
rect 7508 26776 7509 26816
rect 7467 26767 7509 26776
rect 8311 26816 8369 26817
rect 8311 26776 8320 26816
rect 8360 26776 8369 26816
rect 8311 26775 8369 26776
rect 10251 26816 10293 26825
rect 10251 26776 10252 26816
rect 10292 26776 10293 26816
rect 10251 26767 10293 26776
rect 10395 26816 10437 26825
rect 10395 26776 10396 26816
rect 10436 26776 10437 26816
rect 10395 26767 10437 26776
rect 10731 26816 10773 26825
rect 10731 26776 10732 26816
rect 10772 26776 10773 26816
rect 10731 26767 10773 26776
rect 10819 26816 10877 26817
rect 10819 26776 10828 26816
rect 10868 26776 10877 26816
rect 10819 26775 10877 26776
rect 11019 26816 11061 26825
rect 11019 26776 11020 26816
rect 11060 26776 11061 26816
rect 11019 26767 11061 26776
rect 12555 26816 12597 26825
rect 12555 26776 12556 26816
rect 12596 26776 12597 26816
rect 12555 26767 12597 26776
rect 12747 26816 12789 26825
rect 12747 26776 12748 26816
rect 12788 26776 12789 26816
rect 12747 26767 12789 26776
rect 14371 26816 14429 26817
rect 14371 26776 14380 26816
rect 14420 26776 14429 26816
rect 14371 26775 14429 26776
rect 14571 26816 14613 26825
rect 14571 26776 14572 26816
rect 14612 26776 14613 26816
rect 14571 26767 14613 26776
rect 16107 26816 16149 26825
rect 16107 26776 16108 26816
rect 16148 26776 16149 26816
rect 16107 26767 16149 26776
rect 17067 26816 17109 26825
rect 17067 26776 17068 26816
rect 17108 26776 17109 26816
rect 17067 26767 17109 26776
rect 17338 26816 17396 26817
rect 17338 26776 17347 26816
rect 17387 26776 17396 26816
rect 17338 26775 17396 26776
rect 18603 26816 18645 26825
rect 18603 26776 18604 26816
rect 18644 26776 18645 26816
rect 18603 26767 18645 26776
rect 19467 26816 19509 26825
rect 19467 26776 19468 26816
rect 19508 26776 19509 26816
rect 19467 26767 19509 26776
rect 20122 26816 20180 26817
rect 20122 26776 20131 26816
rect 20171 26776 20180 26816
rect 20122 26775 20180 26776
rect 23791 26816 23849 26817
rect 23791 26776 23800 26816
rect 23840 26776 23849 26816
rect 23791 26775 23849 26776
rect 23959 26816 24017 26817
rect 23959 26776 23968 26816
rect 24008 26776 24017 26816
rect 23959 26775 24017 26776
rect 25515 26816 25557 26825
rect 25515 26776 25516 26816
rect 25556 26776 25557 26816
rect 25515 26767 25557 26776
rect 25899 26816 25941 26825
rect 25899 26776 25900 26816
rect 25940 26776 25941 26816
rect 25899 26767 25941 26776
rect 26020 26816 26062 26825
rect 26020 26776 26021 26816
rect 26061 26776 26062 26816
rect 26020 26767 26062 26776
rect 26314 26816 26372 26817
rect 26314 26776 26323 26816
rect 26363 26776 26372 26816
rect 26314 26775 26372 26776
rect 27051 26816 27093 26825
rect 27051 26776 27052 26816
rect 27092 26776 27093 26816
rect 27051 26767 27093 26776
rect 27139 26816 27197 26817
rect 27139 26776 27148 26816
rect 27188 26776 27197 26816
rect 27139 26775 27197 26776
rect 27274 26816 27332 26817
rect 27274 26776 27283 26816
rect 27323 26776 27332 26816
rect 27274 26775 27332 26776
rect 28378 26816 28436 26817
rect 28378 26776 28387 26816
rect 28427 26776 28436 26816
rect 28378 26775 28436 26776
rect 28491 26816 28533 26825
rect 28491 26776 28492 26816
rect 28532 26776 28533 26816
rect 28491 26767 28533 26776
rect 30874 26816 30932 26817
rect 30874 26776 30883 26816
rect 30923 26776 30932 26816
rect 30874 26775 30932 26776
rect 8139 26732 8181 26741
rect 8139 26692 8140 26732
rect 8180 26692 8181 26732
rect 8139 26683 8181 26692
rect 10525 26732 10567 26741
rect 10525 26692 10526 26732
rect 10566 26692 10567 26732
rect 10525 26683 10567 26692
rect 14077 26732 14119 26741
rect 14077 26692 14078 26732
rect 14118 26692 14119 26732
rect 14077 26683 14119 26692
rect 17451 26732 17493 26741
rect 17451 26692 17452 26732
rect 17492 26692 17493 26732
rect 17451 26683 17493 26692
rect 18778 26732 18836 26733
rect 18778 26692 18787 26732
rect 18827 26692 18836 26732
rect 18778 26691 18836 26692
rect 19738 26732 19796 26733
rect 19738 26692 19747 26732
rect 19787 26692 19796 26732
rect 19738 26691 19796 26692
rect 25690 26732 25748 26733
rect 25690 26692 25699 26732
rect 25739 26692 25748 26732
rect 25690 26691 25748 26692
rect 26845 26732 26887 26741
rect 26845 26692 26846 26732
rect 26886 26692 26887 26732
rect 26845 26683 26887 26692
rect 31258 26732 31316 26733
rect 31258 26692 31267 26732
rect 31307 26692 31316 26732
rect 31258 26691 31316 26692
rect 4299 26648 4341 26657
rect 4299 26608 4300 26648
rect 4340 26608 4341 26648
rect 4299 26599 4341 26608
rect 4683 26648 4725 26657
rect 4683 26608 4684 26648
rect 4724 26608 4725 26648
rect 4683 26599 4725 26608
rect 5067 26648 5109 26657
rect 5067 26608 5068 26648
rect 5108 26608 5109 26648
rect 5067 26599 5109 26608
rect 5643 26648 5685 26657
rect 5643 26608 5644 26648
rect 5684 26608 5685 26648
rect 5643 26599 5685 26608
rect 7275 26648 7317 26657
rect 7275 26608 7276 26648
rect 7316 26608 7317 26648
rect 7275 26599 7317 26608
rect 8811 26648 8853 26657
rect 8811 26608 8812 26648
rect 8852 26608 8853 26648
rect 8811 26599 8853 26608
rect 10618 26648 10676 26649
rect 10618 26608 10627 26648
rect 10667 26608 10676 26648
rect 10618 26607 10676 26608
rect 13419 26648 13461 26657
rect 13419 26608 13420 26648
rect 13460 26608 13461 26648
rect 13419 26599 13461 26608
rect 14283 26648 14325 26657
rect 14283 26608 14284 26648
rect 14324 26608 14325 26648
rect 14283 26599 14325 26608
rect 22059 26648 22101 26657
rect 22059 26608 22060 26648
rect 22100 26608 22101 26648
rect 22059 26599 22101 26608
rect 23067 26648 23109 26657
rect 23067 26608 23068 26648
rect 23108 26608 23109 26648
rect 23067 26599 23109 26608
rect 23626 26648 23684 26649
rect 23626 26608 23635 26648
rect 23675 26608 23684 26648
rect 23626 26607 23684 26608
rect 24123 26648 24165 26657
rect 24123 26608 24124 26648
rect 24164 26608 24165 26648
rect 24123 26599 24165 26608
rect 26001 26648 26043 26657
rect 26001 26608 26002 26648
rect 26042 26608 26043 26648
rect 26001 26599 26043 26608
rect 26523 26648 26565 26657
rect 26523 26608 26524 26648
rect 26564 26608 26565 26648
rect 26523 26599 26565 26608
rect 27483 26648 27525 26657
rect 27483 26608 27484 26648
rect 27524 26608 27525 26648
rect 27483 26599 27525 26608
rect 28779 26648 28821 26657
rect 28779 26608 28780 26648
rect 28820 26608 28821 26648
rect 28779 26599 28821 26608
rect 576 26480 31392 26504
rect 576 26440 4352 26480
rect 4720 26440 12126 26480
rect 12494 26440 19900 26480
rect 20268 26440 27674 26480
rect 28042 26440 31392 26480
rect 576 26416 31392 26440
rect 4714 26312 4772 26313
rect 4714 26272 4723 26312
rect 4763 26272 4772 26312
rect 4714 26271 4772 26272
rect 7947 26312 7989 26321
rect 7947 26272 7948 26312
rect 7988 26272 7989 26312
rect 7947 26263 7989 26272
rect 8283 26312 8325 26321
rect 8283 26272 8284 26312
rect 8324 26272 8325 26312
rect 8283 26263 8325 26272
rect 8715 26312 8757 26321
rect 8715 26272 8716 26312
rect 8756 26272 8757 26312
rect 8715 26263 8757 26272
rect 9658 26312 9716 26313
rect 9658 26272 9667 26312
rect 9707 26272 9716 26312
rect 9658 26271 9716 26272
rect 9963 26312 10005 26321
rect 9963 26272 9964 26312
rect 10004 26272 10005 26312
rect 9963 26263 10005 26272
rect 11386 26312 11444 26313
rect 11386 26272 11395 26312
rect 11435 26272 11444 26312
rect 11386 26271 11444 26272
rect 11914 26312 11972 26313
rect 11914 26272 11923 26312
rect 11963 26272 11972 26312
rect 11914 26271 11972 26272
rect 15147 26312 15189 26321
rect 15147 26272 15148 26312
rect 15188 26272 15189 26312
rect 15147 26263 15189 26272
rect 17434 26312 17492 26313
rect 17434 26272 17443 26312
rect 17483 26272 17492 26312
rect 17434 26271 17492 26272
rect 18106 26312 18164 26313
rect 18106 26272 18115 26312
rect 18155 26272 18164 26312
rect 18106 26271 18164 26272
rect 18795 26312 18837 26321
rect 18795 26272 18796 26312
rect 18836 26272 18837 26312
rect 18795 26263 18837 26272
rect 19755 26312 19797 26321
rect 19755 26272 19756 26312
rect 19796 26272 19797 26312
rect 19755 26263 19797 26272
rect 23962 26312 24020 26313
rect 23962 26272 23971 26312
rect 24011 26272 24020 26312
rect 23962 26271 24020 26272
rect 26091 26312 26133 26321
rect 26091 26272 26092 26312
rect 26132 26272 26133 26312
rect 26091 26263 26133 26272
rect 30507 26312 30549 26321
rect 30507 26272 30508 26312
rect 30548 26272 30549 26312
rect 30507 26263 30549 26272
rect 5163 26228 5205 26237
rect 5163 26188 5164 26228
rect 5204 26188 5205 26228
rect 5163 26179 5205 26188
rect 5626 26228 5684 26229
rect 12826 26228 12884 26229
rect 5626 26188 5635 26228
rect 5675 26188 5684 26228
rect 5626 26187 5684 26188
rect 10434 26219 10480 26228
rect 10434 26179 10435 26219
rect 10475 26179 10480 26219
rect 12826 26188 12835 26228
rect 12875 26188 12884 26228
rect 12826 26187 12884 26188
rect 15531 26228 15573 26237
rect 15531 26188 15532 26228
rect 15572 26188 15573 26228
rect 15531 26179 15573 26188
rect 18589 26228 18631 26237
rect 18589 26188 18590 26228
rect 18630 26188 18631 26228
rect 18589 26179 18631 26188
rect 18682 26228 18740 26229
rect 18682 26188 18691 26228
rect 18731 26188 18740 26228
rect 18682 26187 18740 26188
rect 24075 26228 24117 26237
rect 24075 26188 24076 26228
rect 24116 26188 24117 26228
rect 24075 26179 24117 26188
rect 27850 26228 27908 26229
rect 27850 26188 27859 26228
rect 27899 26188 27908 26228
rect 27850 26187 27908 26188
rect 10434 26170 10480 26179
rect 3610 26144 3668 26145
rect 4570 26144 4628 26145
rect 3610 26104 3619 26144
rect 3659 26104 3668 26144
rect 3610 26103 3668 26104
rect 4479 26135 4521 26144
rect 4479 26095 4480 26135
rect 4520 26095 4521 26135
rect 4570 26104 4579 26144
rect 4619 26104 4628 26144
rect 4570 26103 4628 26104
rect 5067 26144 5109 26153
rect 5067 26104 5068 26144
rect 5108 26104 5109 26144
rect 5067 26095 5109 26104
rect 5259 26144 5301 26153
rect 5259 26104 5260 26144
rect 5300 26104 5301 26144
rect 5259 26095 5301 26104
rect 6010 26144 6068 26145
rect 6010 26104 6019 26144
rect 6059 26104 6068 26144
rect 6010 26103 6068 26104
rect 8139 26144 8181 26153
rect 8139 26104 8140 26144
rect 8180 26104 8181 26144
rect 8139 26095 8181 26104
rect 8424 26144 8466 26153
rect 8424 26104 8425 26144
rect 8465 26104 8466 26144
rect 8424 26095 8466 26104
rect 8542 26144 8600 26145
rect 8542 26104 8551 26144
rect 8591 26104 8600 26144
rect 8542 26103 8600 26104
rect 8668 26144 8726 26145
rect 8668 26104 8677 26144
rect 8717 26104 8726 26144
rect 8668 26103 8726 26104
rect 8899 26144 8957 26145
rect 8899 26104 8908 26144
rect 8948 26104 8957 26144
rect 8899 26103 8957 26104
rect 9039 26144 9097 26145
rect 9039 26104 9048 26144
rect 9088 26104 9097 26144
rect 9039 26103 9097 26104
rect 9148 26144 9206 26145
rect 9148 26104 9157 26144
rect 9197 26104 9206 26144
rect 9148 26103 9206 26104
rect 9771 26144 9813 26153
rect 9771 26104 9772 26144
rect 9812 26104 9813 26144
rect 9771 26095 9813 26104
rect 10138 26144 10196 26145
rect 10522 26144 10580 26145
rect 10138 26104 10147 26144
rect 10187 26104 10196 26144
rect 10138 26103 10196 26104
rect 10251 26135 10293 26144
rect 10251 26095 10252 26135
rect 10292 26095 10293 26135
rect 10522 26104 10531 26144
rect 10571 26104 10580 26144
rect 10522 26103 10580 26104
rect 10656 26144 10714 26145
rect 10656 26104 10665 26144
rect 10705 26104 10714 26144
rect 11307 26144 11349 26153
rect 10656 26103 10714 26104
rect 4479 26086 4521 26095
rect 10251 26086 10293 26095
rect 11067 26102 11109 26111
rect 11067 26062 11068 26102
rect 11108 26062 11109 26102
rect 11307 26104 11308 26144
rect 11348 26104 11349 26144
rect 11307 26095 11349 26104
rect 12079 26144 12137 26145
rect 12079 26104 12088 26144
rect 12128 26104 12137 26144
rect 12079 26103 12137 26104
rect 12228 26144 12286 26145
rect 12228 26104 12237 26144
rect 12277 26104 12286 26144
rect 12228 26103 12286 26104
rect 12398 26144 12440 26153
rect 12398 26104 12399 26144
rect 12439 26104 12440 26144
rect 12398 26095 12440 26104
rect 12682 26144 12740 26145
rect 12682 26104 12691 26144
rect 12731 26104 12740 26144
rect 12682 26103 12740 26104
rect 13210 26144 13268 26145
rect 13210 26104 13219 26144
rect 13259 26104 13268 26144
rect 13210 26103 13268 26104
rect 15435 26144 15477 26153
rect 15435 26104 15436 26144
rect 15476 26104 15477 26144
rect 15435 26095 15477 26104
rect 15627 26144 15669 26153
rect 15627 26104 15628 26144
rect 15668 26104 15669 26144
rect 15627 26095 15669 26104
rect 15994 26144 16052 26145
rect 15994 26104 16003 26144
rect 16043 26104 16052 26144
rect 15994 26103 16052 26104
rect 16107 26144 16149 26153
rect 16107 26104 16108 26144
rect 16148 26104 16149 26144
rect 16107 26095 16149 26104
rect 16546 26144 16604 26145
rect 16546 26104 16555 26144
rect 16595 26104 16604 26144
rect 16546 26103 16604 26104
rect 16779 26144 16821 26153
rect 16779 26104 16780 26144
rect 16820 26104 16821 26144
rect 16779 26095 16821 26104
rect 17547 26144 17589 26153
rect 17547 26104 17548 26144
rect 17588 26104 17589 26144
rect 17547 26095 17589 26104
rect 17931 26144 17973 26153
rect 17931 26104 17932 26144
rect 17972 26104 17973 26144
rect 17931 26095 17973 26104
rect 18219 26144 18261 26153
rect 19069 26144 19111 26153
rect 18219 26104 18220 26144
rect 18260 26104 18261 26144
rect 18219 26095 18261 26104
rect 18891 26135 18933 26144
rect 18891 26095 18892 26135
rect 18932 26095 18933 26135
rect 19069 26104 19070 26144
rect 19110 26104 19111 26144
rect 19069 26095 19111 26104
rect 19275 26144 19317 26153
rect 20427 26144 20469 26153
rect 19275 26104 19276 26144
rect 19316 26104 19317 26144
rect 19275 26095 19317 26104
rect 19371 26135 19413 26144
rect 19371 26095 19372 26135
rect 19412 26095 19413 26135
rect 20427 26104 20428 26144
rect 20468 26104 20469 26144
rect 20427 26095 20469 26104
rect 20715 26144 20757 26153
rect 20715 26104 20716 26144
rect 20756 26104 20757 26144
rect 20715 26095 20757 26104
rect 20944 26144 21002 26145
rect 20944 26104 20953 26144
rect 20993 26104 21002 26144
rect 20944 26103 21002 26104
rect 21771 26144 21813 26153
rect 21771 26104 21772 26144
rect 21812 26104 21813 26144
rect 21771 26095 21813 26104
rect 23872 26144 23914 26153
rect 25995 26144 26037 26153
rect 23872 26104 23873 26144
rect 23913 26104 23914 26144
rect 23872 26095 23914 26104
rect 24171 26135 24213 26144
rect 24171 26095 24172 26135
rect 24212 26095 24213 26135
rect 18891 26086 18933 26095
rect 19371 26086 19413 26095
rect 24171 26086 24213 26095
rect 24738 26135 24784 26144
rect 24738 26095 24739 26135
rect 24779 26095 24784 26135
rect 24738 26086 24784 26095
rect 25506 26135 25552 26144
rect 25506 26095 25507 26135
rect 25547 26095 25552 26135
rect 25995 26104 25996 26144
rect 26036 26104 26037 26144
rect 25995 26095 26037 26104
rect 26170 26144 26228 26145
rect 26170 26104 26179 26144
rect 26219 26104 26228 26144
rect 26170 26103 26228 26104
rect 26871 26144 26913 26153
rect 26871 26104 26872 26144
rect 26912 26104 26913 26144
rect 26871 26095 26913 26104
rect 27056 26144 27098 26153
rect 27056 26104 27057 26144
rect 27097 26104 27098 26144
rect 27056 26095 27098 26104
rect 27235 26144 27293 26145
rect 27235 26104 27244 26144
rect 27284 26104 27293 26144
rect 27235 26103 27293 26104
rect 27484 26144 27542 26145
rect 27484 26104 27493 26144
rect 27533 26104 27542 26144
rect 27484 26103 27542 26104
rect 28045 26144 28103 26145
rect 28045 26104 28054 26144
rect 28094 26104 28103 26144
rect 28045 26103 28103 26104
rect 28203 26144 28245 26153
rect 28203 26104 28204 26144
rect 28244 26104 28245 26144
rect 27357 26102 27415 26103
rect 25506 26086 25552 26095
rect 3994 26060 4052 26061
rect 3994 26020 4003 26060
rect 4043 26020 4052 26060
rect 11067 26053 11109 26062
rect 11194 26060 11252 26061
rect 3994 26019 4052 26020
rect 11194 26020 11203 26060
rect 11243 26020 11252 26060
rect 11194 26019 11252 26020
rect 12550 26060 12608 26061
rect 12550 26020 12559 26060
rect 12599 26020 12608 26060
rect 12550 26019 12608 26020
rect 16666 26060 16724 26061
rect 16666 26020 16675 26060
rect 16715 26020 16724 26060
rect 16666 26019 16724 26020
rect 16875 26060 16917 26069
rect 16875 26020 16876 26060
rect 16916 26020 16917 26060
rect 16875 26011 16917 26020
rect 20619 26060 20661 26069
rect 20619 26020 20620 26060
rect 20660 26020 20661 26060
rect 20619 26011 20661 26020
rect 20834 26060 20876 26069
rect 20834 26020 20835 26060
rect 20875 26020 20876 26060
rect 20834 26011 20876 26020
rect 24891 26060 24933 26069
rect 24891 26020 24892 26060
rect 24932 26020 24933 26060
rect 24891 26011 24933 26020
rect 25659 26060 25701 26069
rect 25659 26020 25660 26060
rect 25700 26020 25701 26060
rect 25659 26011 25701 26020
rect 26667 26060 26709 26069
rect 27357 26062 27366 26102
rect 27406 26062 27415 26102
rect 28203 26095 28245 26104
rect 28378 26144 28436 26145
rect 28378 26104 28387 26144
rect 28427 26104 28436 26144
rect 28378 26103 28436 26104
rect 28810 26144 28868 26145
rect 28810 26104 28819 26144
rect 28859 26104 28868 26144
rect 28810 26103 28868 26104
rect 29005 26144 29063 26145
rect 29005 26104 29014 26144
rect 29054 26104 29063 26144
rect 29005 26103 29063 26104
rect 29146 26144 29204 26145
rect 29146 26104 29155 26144
rect 29195 26104 29204 26144
rect 29146 26103 29204 26104
rect 29835 26144 29877 26153
rect 29835 26104 29836 26144
rect 29876 26104 29877 26144
rect 29835 26095 29877 26104
rect 30411 26144 30453 26153
rect 30411 26104 30412 26144
rect 30452 26104 30453 26144
rect 30411 26095 30453 26104
rect 30603 26144 30645 26153
rect 30603 26104 30604 26144
rect 30644 26104 30645 26144
rect 30603 26095 30645 26104
rect 27357 26061 27415 26062
rect 26667 26020 26668 26060
rect 26708 26020 26709 26060
rect 26667 26011 26709 26020
rect 30987 26060 31029 26069
rect 30987 26020 30988 26060
rect 31028 26020 31029 26060
rect 30987 26011 31029 26020
rect 1707 25976 1749 25985
rect 1707 25936 1708 25976
rect 1748 25936 1749 25976
rect 1707 25927 1749 25936
rect 4186 25976 4244 25977
rect 4186 25936 4195 25976
rect 4235 25936 4244 25976
rect 4186 25935 4244 25936
rect 9195 25976 9237 25985
rect 9195 25936 9196 25976
rect 9236 25936 9237 25976
rect 9195 25927 9237 25936
rect 12459 25976 12501 25985
rect 12459 25936 12460 25976
rect 12500 25936 12501 25976
rect 12459 25927 12501 25936
rect 16282 25976 16340 25977
rect 16282 25936 16291 25976
rect 16331 25936 16340 25976
rect 16282 25935 16340 25936
rect 18411 25976 18453 25985
rect 18411 25936 18412 25976
rect 18452 25936 18453 25976
rect 18411 25927 18453 25936
rect 22251 25976 22293 25985
rect 22251 25936 22252 25976
rect 22292 25936 22293 25976
rect 22251 25927 22293 25936
rect 26427 25976 26469 25985
rect 26427 25936 26428 25976
rect 26468 25936 26469 25976
rect 26427 25927 26469 25936
rect 27531 25976 27573 25985
rect 27531 25936 27532 25976
rect 27572 25936 27573 25976
rect 27531 25927 27573 25936
rect 30027 25976 30069 25985
rect 30027 25936 30028 25976
rect 30068 25936 30069 25976
rect 30027 25927 30069 25936
rect 30747 25976 30789 25985
rect 30747 25936 30748 25976
rect 30788 25936 30789 25976
rect 30747 25927 30789 25936
rect 10138 25892 10196 25893
rect 10138 25852 10147 25892
rect 10187 25852 10196 25892
rect 10138 25851 10196 25852
rect 19066 25892 19124 25893
rect 19066 25852 19075 25892
rect 19115 25852 19124 25892
rect 19066 25851 19124 25852
rect 21099 25892 21141 25901
rect 21099 25852 21100 25892
rect 21140 25852 21141 25892
rect 21099 25843 21141 25852
rect 26859 25892 26901 25901
rect 26859 25852 26860 25892
rect 26900 25852 26901 25892
rect 26859 25843 26901 25852
rect 28378 25892 28436 25893
rect 28378 25852 28387 25892
rect 28427 25852 28436 25892
rect 28378 25851 28436 25852
rect 576 25724 31392 25748
rect 576 25684 3112 25724
rect 3480 25684 10886 25724
rect 11254 25684 18660 25724
rect 19028 25684 26434 25724
rect 26802 25684 31392 25724
rect 576 25660 31392 25684
rect 5530 25556 5588 25557
rect 5530 25516 5539 25556
rect 5579 25516 5588 25556
rect 5530 25515 5588 25516
rect 9274 25556 9332 25557
rect 9274 25516 9283 25556
rect 9323 25516 9332 25556
rect 9274 25515 9332 25516
rect 10827 25556 10869 25565
rect 10827 25516 10828 25556
rect 10868 25516 10869 25556
rect 10827 25507 10869 25516
rect 12651 25556 12693 25565
rect 12651 25516 12652 25556
rect 12692 25516 12693 25556
rect 12651 25507 12693 25516
rect 16155 25556 16197 25565
rect 16155 25516 16156 25556
rect 16196 25516 16197 25556
rect 16155 25507 16197 25516
rect 19899 25556 19941 25565
rect 19899 25516 19900 25556
rect 19940 25516 19941 25556
rect 19899 25507 19941 25516
rect 25419 25556 25461 25565
rect 25419 25516 25420 25556
rect 25460 25516 25461 25556
rect 25419 25507 25461 25516
rect 5146 25472 5204 25473
rect 5146 25432 5155 25472
rect 5195 25432 5204 25472
rect 5146 25431 5204 25432
rect 6891 25472 6933 25481
rect 6891 25432 6892 25472
rect 6932 25432 6933 25472
rect 6891 25423 6933 25432
rect 13035 25472 13077 25481
rect 13035 25432 13036 25472
rect 13076 25432 13077 25472
rect 13035 25423 13077 25432
rect 14667 25472 14709 25481
rect 14667 25432 14668 25472
rect 14708 25432 14709 25472
rect 14667 25423 14709 25432
rect 24843 25472 24885 25481
rect 24843 25432 24844 25472
rect 24884 25432 24885 25472
rect 24843 25423 24885 25432
rect 26955 25472 26997 25481
rect 26955 25432 26956 25472
rect 26996 25432 26997 25472
rect 26955 25423 26997 25432
rect 28090 25472 28148 25473
rect 28090 25432 28099 25472
rect 28139 25432 28148 25472
rect 28090 25431 28148 25432
rect 11146 25388 11204 25389
rect 11146 25348 11155 25388
rect 11195 25348 11204 25388
rect 11146 25347 11204 25348
rect 23883 25388 23925 25397
rect 28570 25388 28628 25389
rect 23883 25348 23884 25388
rect 23924 25348 23925 25388
rect 25554 25379 25600 25388
rect 11338 25346 11396 25347
rect 4779 25329 4821 25338
rect 3130 25304 3188 25305
rect 3130 25264 3139 25304
rect 3179 25264 3188 25304
rect 3130 25263 3188 25264
rect 4480 25304 4522 25313
rect 4480 25264 4481 25304
rect 4521 25264 4522 25304
rect 4779 25289 4780 25329
rect 4820 25289 4821 25329
rect 4779 25280 4821 25289
rect 4971 25304 5013 25313
rect 4480 25255 4522 25264
rect 4971 25264 4972 25304
rect 5012 25264 5013 25304
rect 4971 25255 5013 25264
rect 5146 25304 5204 25305
rect 5146 25264 5155 25304
rect 5195 25264 5204 25304
rect 5146 25263 5204 25264
rect 5355 25304 5397 25313
rect 5355 25264 5356 25304
rect 5396 25264 5397 25304
rect 5355 25255 5397 25264
rect 5530 25304 5588 25305
rect 5530 25264 5539 25304
rect 5579 25264 5588 25304
rect 5530 25263 5588 25264
rect 6507 25304 6549 25313
rect 6507 25264 6508 25304
rect 6548 25264 6549 25304
rect 6507 25255 6549 25264
rect 8235 25304 8277 25313
rect 8235 25264 8236 25304
rect 8276 25264 8277 25304
rect 8235 25255 8277 25264
rect 9274 25304 9332 25305
rect 9274 25264 9283 25304
rect 9323 25264 9332 25304
rect 9274 25263 9332 25264
rect 9402 25304 9460 25305
rect 9402 25264 9411 25304
rect 9451 25264 9460 25304
rect 9402 25263 9460 25264
rect 9524 25304 9582 25305
rect 9524 25264 9533 25304
rect 9573 25264 9582 25304
rect 9524 25263 9582 25264
rect 9658 25304 9716 25305
rect 9658 25264 9667 25304
rect 9707 25264 9716 25304
rect 9658 25263 9716 25264
rect 9835 25304 9893 25305
rect 9835 25264 9844 25304
rect 9884 25264 9893 25304
rect 9835 25263 9893 25264
rect 10539 25304 10581 25313
rect 11338 25306 11347 25346
rect 11387 25306 11396 25346
rect 23883 25339 23925 25348
rect 24219 25346 24261 25355
rect 11338 25305 11396 25306
rect 10539 25264 10540 25304
rect 10580 25264 10581 25304
rect 10539 25255 10581 25264
rect 10653 25304 10711 25305
rect 10653 25264 10662 25304
rect 10702 25264 10711 25304
rect 10653 25263 10711 25264
rect 10780 25304 10838 25305
rect 10780 25264 10789 25304
rect 10829 25264 10838 25304
rect 10780 25263 10838 25264
rect 11479 25304 11537 25305
rect 11479 25264 11488 25304
rect 11528 25264 11537 25304
rect 11479 25263 11537 25264
rect 11979 25304 12021 25313
rect 11979 25264 11980 25304
rect 12020 25264 12021 25304
rect 11979 25255 12021 25264
rect 12346 25304 12404 25305
rect 12346 25264 12355 25304
rect 12395 25264 12404 25304
rect 12346 25263 12404 25264
rect 12662 25304 12704 25313
rect 12662 25264 12663 25304
rect 12703 25264 12704 25304
rect 12662 25255 12704 25264
rect 14283 25304 14325 25313
rect 14283 25264 14284 25304
rect 14324 25264 14325 25304
rect 14283 25255 14325 25264
rect 14475 25304 14517 25313
rect 14475 25264 14476 25304
rect 14516 25264 14517 25304
rect 14475 25255 14517 25264
rect 15339 25304 15381 25313
rect 15339 25264 15340 25304
rect 15380 25264 15381 25304
rect 15339 25255 15381 25264
rect 16491 25304 16533 25313
rect 16491 25264 16492 25304
rect 16532 25264 16533 25304
rect 16491 25255 16533 25264
rect 16779 25304 16821 25313
rect 16779 25264 16780 25304
rect 16820 25264 16821 25304
rect 16779 25255 16821 25264
rect 17338 25304 17396 25305
rect 17338 25264 17347 25304
rect 17387 25264 17396 25304
rect 17338 25263 17396 25264
rect 17461 25304 17503 25313
rect 17461 25264 17462 25304
rect 17502 25264 17503 25304
rect 17461 25255 17503 25264
rect 18108 25304 18150 25313
rect 18108 25264 18109 25304
rect 18149 25264 18150 25304
rect 18108 25255 18150 25264
rect 18219 25304 18261 25313
rect 18219 25264 18220 25304
rect 18260 25264 18261 25304
rect 18219 25255 18261 25264
rect 18699 25304 18741 25313
rect 18699 25264 18700 25304
rect 18740 25264 18741 25304
rect 18699 25255 18741 25264
rect 18891 25304 18933 25313
rect 18891 25264 18892 25304
rect 18932 25264 18933 25304
rect 18891 25255 18933 25264
rect 19371 25304 19413 25313
rect 19371 25264 19372 25304
rect 19412 25264 19413 25304
rect 19371 25255 19413 25264
rect 19659 25304 19701 25313
rect 19659 25264 19660 25304
rect 19700 25264 19701 25304
rect 19659 25255 19701 25264
rect 20043 25304 20085 25313
rect 20043 25264 20044 25304
rect 20084 25264 20085 25304
rect 20043 25255 20085 25264
rect 20331 25304 20373 25313
rect 20331 25264 20332 25304
rect 20372 25264 20373 25304
rect 20331 25255 20373 25264
rect 20602 25304 20660 25305
rect 20602 25264 20611 25304
rect 20651 25264 20660 25304
rect 20602 25263 20660 25264
rect 21562 25304 21620 25305
rect 21562 25264 21571 25304
rect 21611 25264 21620 25304
rect 21562 25263 21620 25264
rect 23979 25304 24021 25313
rect 23979 25264 23980 25304
rect 24020 25264 24021 25304
rect 23979 25255 24021 25264
rect 24098 25304 24140 25313
rect 24098 25264 24099 25304
rect 24139 25264 24140 25304
rect 24219 25306 24220 25346
rect 24260 25306 24261 25346
rect 24219 25297 24261 25306
rect 24394 25337 24436 25346
rect 24394 25297 24395 25337
rect 24435 25297 24436 25337
rect 25136 25339 25178 25348
rect 24651 25304 24693 25313
rect 24394 25288 24436 25297
rect 24546 25295 24592 25304
rect 24098 25255 24140 25264
rect 24546 25255 24547 25295
rect 24587 25255 24592 25295
rect 24651 25264 24652 25304
rect 24692 25264 24693 25304
rect 24651 25255 24693 25264
rect 24843 25304 24885 25313
rect 24843 25264 24844 25304
rect 24884 25264 24885 25304
rect 24843 25255 24885 25264
rect 24960 25304 25018 25305
rect 24960 25264 24969 25304
rect 25009 25264 25018 25304
rect 25136 25299 25137 25339
rect 25177 25299 25178 25339
rect 25554 25339 25555 25379
rect 25595 25339 25600 25379
rect 28570 25348 28579 25388
rect 28619 25348 28628 25388
rect 28570 25347 28628 25348
rect 25554 25330 25600 25339
rect 25136 25290 25178 25299
rect 25323 25304 25365 25313
rect 24960 25263 25018 25264
rect 25323 25264 25324 25304
rect 25364 25264 25365 25304
rect 25323 25255 25365 25264
rect 25654 25304 25712 25305
rect 25654 25264 25663 25304
rect 25703 25264 25712 25304
rect 25654 25263 25712 25264
rect 25899 25304 25941 25313
rect 25899 25264 25900 25304
rect 25940 25264 25941 25304
rect 25899 25255 25941 25264
rect 26362 25304 26420 25305
rect 26362 25264 26371 25304
rect 26411 25264 26420 25304
rect 26362 25263 26420 25264
rect 26475 25304 26517 25313
rect 26475 25264 26476 25304
rect 26516 25264 26517 25304
rect 26475 25255 26517 25264
rect 26859 25304 26901 25313
rect 26859 25264 26860 25304
rect 26900 25264 26901 25304
rect 26859 25255 26901 25264
rect 26973 25304 27031 25305
rect 26973 25264 26982 25304
rect 27022 25264 27031 25304
rect 26973 25263 27031 25264
rect 27100 25304 27158 25305
rect 27100 25264 27109 25304
rect 27149 25264 27158 25304
rect 27100 25263 27158 25264
rect 27802 25304 27860 25305
rect 27802 25264 27811 25304
rect 27851 25264 27860 25304
rect 27802 25263 27860 25264
rect 27909 25304 27967 25305
rect 27909 25264 27918 25304
rect 27958 25264 27967 25304
rect 27909 25263 27967 25264
rect 28438 25304 28480 25313
rect 28438 25264 28439 25304
rect 28479 25264 28480 25304
rect 28438 25255 28480 25264
rect 28683 25304 28725 25313
rect 28683 25264 28684 25304
rect 28724 25264 28725 25304
rect 28683 25255 28725 25264
rect 29338 25304 29396 25305
rect 29338 25264 29347 25304
rect 29387 25264 29396 25304
rect 29338 25263 29396 25264
rect 24546 25246 24592 25255
rect 3514 25220 3572 25221
rect 3514 25180 3523 25220
rect 3563 25180 3572 25220
rect 3514 25179 3572 25180
rect 11643 25220 11685 25229
rect 11643 25180 11644 25220
rect 11684 25180 11685 25220
rect 11643 25171 11685 25180
rect 14379 25220 14421 25229
rect 14379 25180 14380 25220
rect 14420 25180 14421 25220
rect 14379 25171 14421 25180
rect 20715 25220 20757 25229
rect 20715 25180 20716 25220
rect 20756 25180 20757 25220
rect 20715 25171 20757 25180
rect 21178 25220 21236 25221
rect 21178 25180 21187 25220
rect 21227 25180 21236 25220
rect 21178 25179 21236 25180
rect 26650 25220 26708 25221
rect 26650 25180 26659 25220
rect 26699 25180 26708 25220
rect 26650 25179 26708 25180
rect 28762 25220 28820 25221
rect 28762 25180 28771 25220
rect 28811 25180 28820 25220
rect 28762 25179 28820 25180
rect 28954 25220 29012 25221
rect 28954 25180 28963 25220
rect 29003 25180 29012 25220
rect 28954 25179 29012 25180
rect 1227 25136 1269 25145
rect 1227 25096 1228 25136
rect 1268 25096 1269 25136
rect 1227 25087 1269 25096
rect 4570 25136 4628 25137
rect 4570 25096 4579 25136
rect 4619 25096 4628 25136
rect 4570 25095 4628 25096
rect 4683 25136 4725 25145
rect 4683 25096 4684 25136
rect 4724 25096 4725 25136
rect 4683 25087 4725 25096
rect 5835 25136 5877 25145
rect 5835 25096 5836 25136
rect 5876 25096 5877 25136
rect 5835 25087 5877 25096
rect 7275 25136 7317 25145
rect 7275 25096 7276 25136
rect 7316 25096 7317 25136
rect 7275 25087 7317 25096
rect 8122 25136 8180 25137
rect 8122 25096 8131 25136
rect 8171 25096 8180 25136
rect 8122 25095 8180 25096
rect 8427 25136 8469 25145
rect 8427 25096 8428 25136
rect 8468 25096 8469 25136
rect 8427 25087 8469 25096
rect 12442 25136 12500 25137
rect 12442 25096 12451 25136
rect 12491 25096 12500 25136
rect 12442 25095 12500 25096
rect 16011 25136 16053 25145
rect 16011 25096 16012 25136
rect 16052 25096 16053 25136
rect 16011 25087 16053 25096
rect 17739 25136 17781 25145
rect 17739 25096 17740 25136
rect 17780 25096 17781 25136
rect 17739 25087 17781 25096
rect 17914 25136 17972 25137
rect 17914 25096 17923 25136
rect 17963 25096 17972 25136
rect 17914 25095 17972 25096
rect 18874 25136 18932 25137
rect 18874 25096 18883 25136
rect 18923 25096 18932 25136
rect 18874 25095 18932 25096
rect 19162 25136 19220 25137
rect 19162 25096 19171 25136
rect 19211 25096 19220 25136
rect 19162 25095 19220 25096
rect 21051 25136 21093 25145
rect 21051 25096 21052 25136
rect 21092 25096 21093 25136
rect 21051 25087 21093 25096
rect 23499 25136 23541 25145
rect 23499 25096 23500 25136
rect 23540 25096 23541 25136
rect 23499 25087 23541 25096
rect 24363 25136 24405 25145
rect 24363 25096 24364 25136
rect 24404 25096 24405 25136
rect 24363 25087 24405 25096
rect 25419 25136 25461 25145
rect 25419 25096 25420 25136
rect 25460 25096 25461 25136
rect 25419 25087 25461 25096
rect 26379 25136 26421 25145
rect 26379 25096 26380 25136
rect 26420 25096 26421 25136
rect 26379 25087 26421 25096
rect 31275 25136 31317 25145
rect 31275 25096 31276 25136
rect 31316 25096 31317 25136
rect 31275 25087 31317 25096
rect 576 24968 31392 24992
rect 576 24928 4352 24968
rect 4720 24928 12126 24968
rect 12494 24928 19900 24968
rect 20268 24928 27674 24968
rect 28042 24928 31392 24968
rect 576 24904 31392 24928
rect 4090 24800 4148 24801
rect 4090 24760 4099 24800
rect 4139 24760 4148 24800
rect 4090 24759 4148 24760
rect 4971 24800 5013 24809
rect 4971 24760 4972 24800
rect 5012 24760 5013 24800
rect 4971 24751 5013 24760
rect 5547 24800 5589 24809
rect 5547 24760 5548 24800
rect 5588 24760 5589 24800
rect 5547 24751 5589 24760
rect 8139 24800 8181 24809
rect 8139 24760 8140 24800
rect 8180 24760 8181 24800
rect 8139 24751 8181 24760
rect 8890 24800 8948 24801
rect 8890 24760 8899 24800
rect 8939 24760 8948 24800
rect 8890 24759 8948 24760
rect 9195 24800 9237 24809
rect 9195 24760 9196 24800
rect 9236 24760 9237 24800
rect 9195 24751 9237 24760
rect 10618 24800 10676 24801
rect 10618 24760 10627 24800
rect 10667 24760 10676 24800
rect 10618 24759 10676 24760
rect 14746 24800 14804 24801
rect 14746 24760 14755 24800
rect 14795 24760 14804 24800
rect 14746 24759 14804 24760
rect 16810 24800 16868 24801
rect 16810 24760 16819 24800
rect 16859 24760 16868 24800
rect 16810 24759 16868 24760
rect 17818 24800 17876 24801
rect 17818 24760 17827 24800
rect 17867 24760 17876 24800
rect 17818 24759 17876 24760
rect 17931 24800 17973 24809
rect 17931 24760 17932 24800
rect 17972 24760 17973 24800
rect 17931 24751 17973 24760
rect 21195 24800 21237 24809
rect 21195 24760 21196 24800
rect 21236 24760 21237 24800
rect 21195 24751 21237 24760
rect 23499 24800 23541 24809
rect 23499 24760 23500 24800
rect 23540 24760 23541 24800
rect 23499 24751 23541 24760
rect 25323 24800 25365 24809
rect 25323 24760 25324 24800
rect 25364 24760 25365 24800
rect 25323 24751 25365 24760
rect 26379 24800 26421 24809
rect 26379 24760 26380 24800
rect 26420 24760 26421 24800
rect 26379 24751 26421 24760
rect 27051 24800 27093 24809
rect 27051 24760 27052 24800
rect 27092 24760 27093 24800
rect 27051 24751 27093 24760
rect 28090 24800 28148 24801
rect 28090 24760 28099 24800
rect 28139 24760 28148 24800
rect 28090 24759 28148 24760
rect 28875 24800 28917 24809
rect 28875 24760 28876 24800
rect 28916 24760 28917 24800
rect 28875 24751 28917 24760
rect 18038 24716 18080 24725
rect 25210 24716 25268 24717
rect 10050 24707 10096 24716
rect 10050 24667 10051 24707
rect 10091 24667 10096 24707
rect 18038 24676 18039 24716
rect 18079 24676 18080 24716
rect 18038 24667 18080 24676
rect 19554 24707 19600 24716
rect 19554 24667 19555 24707
rect 19595 24667 19600 24707
rect 25210 24676 25219 24716
rect 25259 24676 25268 24716
rect 25210 24675 25268 24676
rect 10050 24658 10096 24667
rect 19554 24658 19600 24667
rect 28289 24659 28347 24660
rect 2187 24632 2229 24641
rect 2187 24592 2188 24632
rect 2228 24592 2229 24632
rect 2187 24583 2229 24592
rect 4203 24632 4245 24641
rect 4203 24592 4204 24632
rect 4244 24592 4245 24632
rect 4203 24583 4245 24592
rect 4587 24632 4629 24641
rect 4587 24592 4588 24632
rect 4628 24592 4629 24632
rect 4587 24583 4629 24592
rect 4779 24632 4821 24641
rect 4779 24592 4780 24632
rect 4820 24592 4821 24632
rect 4779 24583 4821 24592
rect 5146 24632 5204 24633
rect 5146 24592 5155 24632
rect 5195 24592 5204 24632
rect 5146 24591 5204 24592
rect 5451 24632 5493 24641
rect 5451 24592 5452 24632
rect 5492 24592 5493 24632
rect 5451 24583 5493 24592
rect 5626 24632 5684 24633
rect 5626 24592 5635 24632
rect 5675 24592 5684 24632
rect 5626 24591 5684 24592
rect 6202 24632 6260 24633
rect 6202 24592 6211 24632
rect 6251 24592 6260 24632
rect 6202 24591 6260 24592
rect 8292 24632 8350 24633
rect 8292 24592 8301 24632
rect 8341 24592 8350 24632
rect 8292 24591 8350 24592
rect 8448 24632 8490 24641
rect 8448 24592 8449 24632
rect 8489 24592 8490 24632
rect 8448 24583 8490 24592
rect 8740 24632 8782 24641
rect 8740 24592 8741 24632
rect 8781 24592 8782 24632
rect 8740 24583 8782 24592
rect 9003 24632 9045 24641
rect 9003 24592 9004 24632
rect 9044 24592 9045 24632
rect 9003 24583 9045 24592
rect 9754 24632 9812 24633
rect 10146 24632 10204 24633
rect 9754 24592 9763 24632
rect 9803 24592 9812 24632
rect 9754 24591 9812 24592
rect 9867 24623 9909 24632
rect 9867 24583 9868 24623
rect 9908 24583 9909 24623
rect 10146 24592 10155 24632
rect 10195 24592 10204 24632
rect 10146 24591 10204 24592
rect 10315 24632 10373 24633
rect 10315 24592 10324 24632
rect 10364 24592 10373 24632
rect 10315 24591 10373 24592
rect 10906 24632 10964 24633
rect 10906 24592 10915 24632
rect 10955 24592 10964 24632
rect 10906 24591 10964 24592
rect 11446 24632 11488 24641
rect 11446 24592 11447 24632
rect 11487 24592 11488 24632
rect 11446 24583 11488 24592
rect 11691 24632 11733 24641
rect 11691 24592 11692 24632
rect 11732 24592 11733 24632
rect 11691 24583 11733 24592
rect 12346 24632 12404 24633
rect 12346 24592 12355 24632
rect 12395 24592 12404 24632
rect 12346 24591 12404 24592
rect 14422 24632 14464 24641
rect 14422 24592 14423 24632
rect 14463 24592 14464 24632
rect 14422 24583 14464 24592
rect 14554 24632 14612 24633
rect 14554 24592 14563 24632
rect 14603 24592 14612 24632
rect 14554 24591 14612 24592
rect 14667 24632 14709 24641
rect 16107 24632 16149 24641
rect 14667 24592 14668 24632
rect 14708 24592 14709 24632
rect 14667 24583 14709 24592
rect 14946 24623 14992 24632
rect 14946 24583 14947 24623
rect 14987 24583 14992 24623
rect 16107 24592 16108 24632
rect 16148 24592 16149 24632
rect 16107 24583 16149 24592
rect 16975 24632 17033 24633
rect 16975 24592 16984 24632
rect 17024 24592 17033 24632
rect 16975 24591 17033 24592
rect 17722 24632 17780 24633
rect 17722 24592 17731 24632
rect 17771 24592 17780 24632
rect 17722 24591 17780 24592
rect 18214 24627 18256 24636
rect 18214 24587 18215 24627
rect 18255 24587 18256 24627
rect 9867 24574 9909 24583
rect 14946 24574 14992 24583
rect 18214 24578 18256 24587
rect 18411 24632 18453 24641
rect 18411 24592 18412 24632
rect 18452 24592 18453 24632
rect 18411 24583 18453 24592
rect 18699 24632 18741 24641
rect 18699 24592 18700 24632
rect 18740 24592 18741 24632
rect 18699 24583 18741 24592
rect 18987 24632 19029 24641
rect 18987 24592 18988 24632
rect 19028 24592 19029 24632
rect 18987 24583 19029 24592
rect 19131 24632 19173 24641
rect 19131 24592 19132 24632
rect 19172 24592 19173 24632
rect 19131 24583 19173 24592
rect 19258 24632 19316 24633
rect 19642 24632 19700 24633
rect 19258 24592 19267 24632
rect 19307 24592 19316 24632
rect 19258 24591 19316 24592
rect 19371 24623 19413 24632
rect 19371 24583 19372 24623
rect 19412 24583 19413 24623
rect 19642 24592 19651 24632
rect 19691 24592 19700 24632
rect 19642 24591 19700 24592
rect 19776 24632 19834 24633
rect 19776 24592 19785 24632
rect 19825 24592 19834 24632
rect 19776 24591 19834 24592
rect 19995 24632 20037 24641
rect 19995 24592 19996 24632
rect 20036 24592 20037 24632
rect 19995 24583 20037 24592
rect 20296 24632 20338 24641
rect 20296 24592 20297 24632
rect 20337 24592 20338 24632
rect 20296 24583 20338 24592
rect 20458 24632 20516 24633
rect 20458 24592 20467 24632
rect 20507 24592 20516 24632
rect 20458 24591 20516 24592
rect 21867 24632 21909 24641
rect 21867 24592 21868 24632
rect 21908 24592 21909 24632
rect 21867 24583 21909 24592
rect 22827 24632 22869 24641
rect 22827 24592 22828 24632
rect 22868 24592 22869 24632
rect 22827 24583 22869 24592
rect 23595 24632 23637 24641
rect 23595 24592 23596 24632
rect 23636 24592 23637 24632
rect 23595 24583 23637 24592
rect 24324 24632 24382 24633
rect 24324 24592 24333 24632
rect 24373 24592 24382 24632
rect 24324 24591 24382 24592
rect 24494 24632 24536 24641
rect 24494 24592 24495 24632
rect 24535 24592 24536 24632
rect 24494 24583 24536 24592
rect 24772 24632 24814 24641
rect 24772 24592 24773 24632
rect 24813 24592 24814 24632
rect 24772 24583 24814 24592
rect 25117 24632 25159 24641
rect 25950 24632 25992 24641
rect 26187 24632 26229 24641
rect 25117 24592 25118 24632
rect 25158 24592 25159 24632
rect 25117 24583 25159 24592
rect 25417 24629 25475 24630
rect 25417 24589 25426 24629
rect 25466 24589 25475 24629
rect 25417 24588 25475 24589
rect 25848 24623 25890 24632
rect 25848 24583 25849 24623
rect 25889 24583 25890 24623
rect 25950 24592 25951 24632
rect 25991 24592 25992 24632
rect 25950 24583 25992 24592
rect 26082 24623 26128 24632
rect 26082 24583 26083 24623
rect 26123 24583 26128 24623
rect 26187 24592 26188 24632
rect 26228 24592 26229 24632
rect 26187 24583 26229 24592
rect 26368 24632 26410 24641
rect 26368 24592 26369 24632
rect 26409 24592 26410 24632
rect 26368 24583 26410 24592
rect 26576 24632 26618 24641
rect 26576 24592 26577 24632
rect 26617 24592 26618 24632
rect 26576 24583 26618 24592
rect 26955 24632 26997 24641
rect 26955 24592 26956 24632
rect 26996 24592 26997 24632
rect 26955 24583 26997 24592
rect 27130 24632 27188 24633
rect 27130 24592 27139 24632
rect 27179 24592 27188 24632
rect 27130 24591 27188 24592
rect 27435 24632 27477 24641
rect 27435 24592 27436 24632
rect 27476 24592 27477 24632
rect 27435 24583 27477 24592
rect 27627 24632 27669 24641
rect 27627 24592 27628 24632
rect 27668 24592 27669 24632
rect 27627 24583 27669 24592
rect 27915 24632 27957 24641
rect 27915 24592 27916 24632
rect 27956 24592 27957 24632
rect 27915 24583 27957 24592
rect 28107 24632 28149 24641
rect 28107 24592 28108 24632
rect 28148 24592 28149 24632
rect 28289 24619 28298 24659
rect 28338 24619 28347 24659
rect 28289 24618 28347 24619
rect 28491 24632 28533 24641
rect 28107 24583 28149 24592
rect 28491 24592 28492 24632
rect 28532 24592 28533 24632
rect 28491 24583 28533 24592
rect 29547 24632 29589 24641
rect 29547 24592 29548 24632
rect 29588 24592 29589 24632
rect 29547 24583 29589 24592
rect 30795 24632 30837 24641
rect 30795 24592 30796 24632
rect 30836 24592 30837 24632
rect 30795 24583 30837 24592
rect 19371 24574 19413 24583
rect 25848 24574 25890 24583
rect 26082 24574 26128 24583
rect 5835 24548 5877 24557
rect 5835 24508 5836 24548
rect 5876 24508 5877 24548
rect 5835 24499 5877 24508
rect 8619 24548 8661 24557
rect 8619 24508 8620 24548
rect 8660 24508 8661 24548
rect 8619 24499 8661 24508
rect 10522 24548 10580 24549
rect 10522 24508 10531 24548
rect 10571 24508 10580 24548
rect 10522 24507 10580 24508
rect 11098 24548 11156 24549
rect 11098 24508 11107 24548
rect 11147 24508 11156 24548
rect 11098 24507 11156 24508
rect 11578 24548 11636 24549
rect 11578 24508 11587 24548
rect 11627 24508 11636 24548
rect 11578 24507 11636 24508
rect 11787 24548 11829 24557
rect 11787 24508 11788 24548
rect 11828 24508 11829 24548
rect 11787 24499 11829 24508
rect 11979 24548 12021 24557
rect 11979 24508 11980 24548
rect 12020 24508 12021 24548
rect 11979 24499 12021 24508
rect 15099 24548 15141 24557
rect 15099 24508 15100 24548
rect 15140 24508 15141 24548
rect 15099 24499 15141 24508
rect 18315 24548 18357 24557
rect 18315 24508 18316 24548
rect 18356 24508 18357 24548
rect 18315 24499 18357 24508
rect 20139 24548 20181 24557
rect 20139 24508 20140 24548
rect 20180 24508 20181 24548
rect 20139 24499 20181 24508
rect 22138 24548 22196 24549
rect 22138 24508 22147 24548
rect 22187 24508 22196 24548
rect 22138 24507 22196 24508
rect 23499 24548 23541 24557
rect 23499 24508 23500 24548
rect 23540 24508 23541 24548
rect 23499 24499 23541 24508
rect 24651 24548 24693 24557
rect 24651 24508 24652 24548
rect 24692 24508 24693 24548
rect 24651 24499 24693 24508
rect 27723 24548 27765 24557
rect 27723 24508 27724 24548
rect 27764 24508 27765 24548
rect 27723 24499 27765 24508
rect 28395 24548 28437 24557
rect 28395 24508 28396 24548
rect 28436 24508 28437 24548
rect 28395 24499 28437 24508
rect 1899 24464 1941 24473
rect 1899 24424 1900 24464
rect 1940 24424 1941 24464
rect 1899 24415 1941 24424
rect 3051 24464 3093 24473
rect 3051 24424 3052 24464
rect 3092 24424 3093 24464
rect 3051 24415 3093 24424
rect 4395 24464 4437 24473
rect 4395 24424 4396 24464
rect 4436 24424 4437 24464
rect 4395 24415 4437 24424
rect 5199 24464 5241 24473
rect 5199 24424 5200 24464
rect 5240 24424 5241 24464
rect 5199 24415 5241 24424
rect 8523 24464 8565 24473
rect 8523 24424 8524 24464
rect 8564 24424 8565 24464
rect 8523 24415 8565 24424
rect 14283 24464 14325 24473
rect 14283 24424 14284 24464
rect 14324 24424 14325 24464
rect 14283 24415 14325 24424
rect 17163 24464 17205 24473
rect 17163 24424 17164 24464
rect 17204 24424 17205 24464
rect 17163 24415 17205 24424
rect 20235 24464 20277 24473
rect 20235 24424 20236 24464
rect 20276 24424 20277 24464
rect 20235 24415 20277 24424
rect 23019 24464 23061 24473
rect 23019 24424 23020 24464
rect 23060 24424 23061 24464
rect 23019 24415 23061 24424
rect 24555 24464 24597 24473
rect 24555 24424 24556 24464
rect 24596 24424 24597 24464
rect 24555 24415 24597 24424
rect 29931 24464 29973 24473
rect 29931 24424 29932 24464
rect 29972 24424 29973 24464
rect 29931 24415 29973 24424
rect 30987 24464 31029 24473
rect 30987 24424 30988 24464
rect 31028 24424 31029 24464
rect 30987 24415 31029 24424
rect 2859 24380 2901 24389
rect 2859 24340 2860 24380
rect 2900 24340 2901 24380
rect 2859 24331 2901 24340
rect 4587 24380 4629 24389
rect 4587 24340 4588 24380
rect 4628 24340 4629 24380
rect 4587 24331 4629 24340
rect 9754 24380 9812 24381
rect 9754 24340 9763 24380
rect 9803 24340 9812 24380
rect 9754 24339 9812 24340
rect 13899 24380 13941 24389
rect 13899 24340 13900 24380
rect 13940 24340 13941 24380
rect 13899 24331 13941 24340
rect 15435 24380 15477 24389
rect 15435 24340 15436 24380
rect 15476 24340 15477 24380
rect 15435 24331 15477 24340
rect 19258 24380 19316 24381
rect 19258 24340 19267 24380
rect 19307 24340 19316 24380
rect 19258 24339 19316 24340
rect 25899 24380 25941 24389
rect 25899 24340 25900 24380
rect 25940 24340 25941 24380
rect 25899 24331 25941 24340
rect 27130 24380 27188 24381
rect 27130 24340 27139 24380
rect 27179 24340 27188 24380
rect 27130 24339 27188 24340
rect 30123 24380 30165 24389
rect 30123 24340 30124 24380
rect 30164 24340 30165 24380
rect 30123 24331 30165 24340
rect 576 24212 31392 24236
rect 576 24172 3112 24212
rect 3480 24172 10886 24212
rect 11254 24172 18660 24212
rect 19028 24172 26434 24212
rect 26802 24172 31392 24212
rect 576 24148 31392 24172
rect 5242 24044 5300 24045
rect 5242 24004 5251 24044
rect 5291 24004 5300 24044
rect 5242 24003 5300 24004
rect 7930 24044 7988 24045
rect 7930 24004 7939 24044
rect 7979 24004 7988 24044
rect 7930 24003 7988 24004
rect 9291 24044 9333 24053
rect 9291 24004 9292 24044
rect 9332 24004 9333 24044
rect 9291 23995 9333 24004
rect 9675 24044 9717 24053
rect 9675 24004 9676 24044
rect 9716 24004 9717 24044
rect 9675 23995 9717 24004
rect 12267 24044 12309 24053
rect 12267 24004 12268 24044
rect 12308 24004 12309 24044
rect 12267 23995 12309 24004
rect 18603 24044 18645 24053
rect 18603 24004 18604 24044
rect 18644 24004 18645 24044
rect 18603 23995 18645 24004
rect 19450 24044 19508 24045
rect 19450 24004 19459 24044
rect 19499 24004 19508 24044
rect 19450 24003 19508 24004
rect 28203 24044 28245 24053
rect 28203 24004 28204 24044
rect 28244 24004 28245 24044
rect 28203 23995 28245 24004
rect 31275 24044 31317 24053
rect 31275 24004 31276 24044
rect 31316 24004 31317 24044
rect 31275 23995 31317 24004
rect 3147 23960 3189 23969
rect 3147 23920 3148 23960
rect 3188 23920 3189 23960
rect 3147 23911 3189 23920
rect 6219 23960 6261 23969
rect 6219 23920 6220 23960
rect 6260 23920 6261 23960
rect 6219 23911 6261 23920
rect 7083 23960 7125 23969
rect 7083 23920 7084 23960
rect 7124 23920 7125 23960
rect 7083 23911 7125 23920
rect 9099 23960 9141 23969
rect 9099 23920 9100 23960
rect 9140 23920 9141 23960
rect 9099 23911 9141 23920
rect 11962 23960 12020 23961
rect 27531 23960 27573 23969
rect 11962 23920 11971 23960
rect 12011 23920 12020 23960
rect 11962 23919 12020 23920
rect 18859 23951 18901 23960
rect 18859 23911 18860 23951
rect 18900 23911 18901 23951
rect 27531 23920 27532 23960
rect 27572 23920 27573 23960
rect 27531 23911 27573 23920
rect 18859 23902 18901 23911
rect 2938 23876 2996 23877
rect 2938 23836 2947 23876
rect 2987 23836 2996 23876
rect 2938 23835 2996 23836
rect 4234 23876 4292 23877
rect 12538 23876 12596 23877
rect 4234 23836 4243 23876
rect 4283 23836 4292 23876
rect 4234 23835 4292 23836
rect 5010 23867 5056 23876
rect 5010 23827 5011 23867
rect 5051 23827 5056 23867
rect 12538 23836 12547 23876
rect 12587 23836 12596 23876
rect 12538 23835 12596 23836
rect 14506 23876 14564 23877
rect 14506 23836 14515 23876
rect 14555 23836 14564 23876
rect 14506 23835 14564 23836
rect 15435 23876 15477 23885
rect 15435 23836 15436 23876
rect 15476 23836 15477 23876
rect 15435 23827 15477 23836
rect 19803 23876 19845 23885
rect 19803 23836 19804 23876
rect 19844 23836 19845 23876
rect 19803 23827 19845 23836
rect 23098 23876 23156 23877
rect 23098 23836 23107 23876
rect 23147 23836 23156 23876
rect 23098 23835 23156 23836
rect 24699 23876 24741 23885
rect 24699 23836 24700 23876
rect 24740 23836 24741 23876
rect 24699 23827 24741 23836
rect 28971 23876 29013 23885
rect 28971 23836 28972 23876
rect 29012 23836 29013 23876
rect 28971 23827 29013 23836
rect 5010 23818 5056 23827
rect 2554 23792 2612 23793
rect 3819 23792 3861 23801
rect 2554 23752 2563 23792
rect 2603 23752 2612 23792
rect 2554 23751 2612 23752
rect 3531 23783 3573 23792
rect 3531 23743 3532 23783
rect 3572 23743 3573 23783
rect 3819 23752 3820 23792
rect 3860 23752 3861 23792
rect 3819 23743 3861 23752
rect 4429 23792 4487 23793
rect 4429 23752 4438 23792
rect 4478 23752 4487 23792
rect 4429 23751 4487 23752
rect 4874 23792 4916 23801
rect 4874 23752 4875 23792
rect 4915 23752 4916 23792
rect 4874 23743 4916 23752
rect 5104 23792 5162 23793
rect 5104 23752 5113 23792
rect 5153 23752 5162 23792
rect 5104 23751 5162 23752
rect 5539 23792 5597 23793
rect 5539 23752 5548 23792
rect 5588 23752 5597 23792
rect 5539 23751 5597 23752
rect 6891 23792 6933 23801
rect 6891 23752 6892 23792
rect 6932 23752 6933 23792
rect 6891 23743 6933 23752
rect 7936 23792 7978 23801
rect 7936 23752 7937 23792
rect 7977 23752 7978 23792
rect 7936 23743 7978 23752
rect 8227 23792 8285 23793
rect 8227 23752 8236 23792
rect 8276 23752 8285 23792
rect 8227 23751 8285 23752
rect 8523 23792 8565 23801
rect 8523 23752 8524 23792
rect 8564 23752 8565 23792
rect 8523 23743 8565 23752
rect 8715 23792 8757 23801
rect 8715 23752 8716 23792
rect 8756 23752 8757 23792
rect 8715 23743 8757 23752
rect 9291 23792 9333 23801
rect 9291 23752 9292 23792
rect 9332 23752 9333 23792
rect 9291 23743 9333 23752
rect 9483 23792 9525 23801
rect 9483 23752 9484 23792
rect 9524 23752 9525 23792
rect 9483 23743 9525 23752
rect 9675 23792 9717 23801
rect 9675 23752 9676 23792
rect 9716 23752 9717 23792
rect 9675 23743 9717 23752
rect 9867 23792 9909 23801
rect 9867 23752 9868 23792
rect 9908 23752 9909 23792
rect 9867 23743 9909 23752
rect 10683 23792 10725 23801
rect 10683 23752 10684 23792
rect 10724 23752 10725 23792
rect 10683 23743 10725 23752
rect 10923 23792 10965 23801
rect 10923 23752 10924 23792
rect 10964 23752 10965 23792
rect 10923 23743 10965 23752
rect 11787 23792 11829 23801
rect 11787 23752 11788 23792
rect 11828 23752 11829 23792
rect 11787 23743 11829 23752
rect 11962 23792 12020 23793
rect 11962 23752 11971 23792
rect 12011 23752 12020 23792
rect 11962 23751 12020 23752
rect 12154 23792 12196 23801
rect 12154 23752 12155 23792
rect 12195 23752 12196 23792
rect 12154 23743 12196 23752
rect 12363 23792 12405 23801
rect 12363 23752 12364 23792
rect 12404 23752 12405 23792
rect 12363 23743 12405 23752
rect 13227 23792 13269 23801
rect 13227 23752 13228 23792
rect 13268 23752 13269 23792
rect 13227 23743 13269 23752
rect 14187 23792 14229 23801
rect 14187 23752 14188 23792
rect 14228 23752 14229 23792
rect 14187 23743 14229 23752
rect 14671 23792 14729 23793
rect 14671 23752 14680 23792
rect 14720 23752 14729 23792
rect 14671 23751 14729 23752
rect 15046 23792 15088 23801
rect 15046 23752 15047 23792
rect 15087 23752 15088 23792
rect 15046 23743 15088 23752
rect 15243 23792 15285 23801
rect 15243 23752 15244 23792
rect 15284 23752 15285 23792
rect 15243 23743 15285 23752
rect 15802 23792 15860 23793
rect 15802 23752 15811 23792
rect 15851 23752 15860 23792
rect 15802 23751 15860 23752
rect 17931 23792 17973 23801
rect 17931 23752 17932 23792
rect 17972 23752 17973 23792
rect 17931 23743 17973 23752
rect 18874 23792 18932 23793
rect 18874 23752 18883 23792
rect 18923 23752 18932 23792
rect 18874 23751 18932 23752
rect 19275 23792 19317 23801
rect 19275 23752 19276 23792
rect 19316 23752 19317 23792
rect 19275 23743 19317 23752
rect 19450 23792 19508 23793
rect 19450 23752 19459 23792
rect 19499 23752 19508 23792
rect 19450 23751 19508 23752
rect 19639 23792 19697 23793
rect 19639 23752 19648 23792
rect 19688 23752 19697 23792
rect 19639 23751 19697 23752
rect 22714 23792 22772 23793
rect 22714 23752 22723 23792
rect 22763 23752 22772 23792
rect 22714 23751 22772 23752
rect 23451 23792 23493 23801
rect 23451 23752 23452 23792
rect 23492 23752 23493 23792
rect 23451 23743 23493 23752
rect 23595 23792 23637 23801
rect 23595 23752 23596 23792
rect 23636 23752 23637 23792
rect 23595 23743 23637 23752
rect 24267 23792 24309 23801
rect 24267 23752 24268 23792
rect 24308 23752 24309 23792
rect 24267 23743 24309 23752
rect 24355 23792 24413 23793
rect 24355 23752 24364 23792
rect 24404 23752 24413 23792
rect 24355 23751 24413 23752
rect 24490 23792 24548 23793
rect 24490 23752 24499 23792
rect 24539 23752 24548 23792
rect 24490 23751 24548 23752
rect 24982 23792 25024 23801
rect 24982 23752 24983 23792
rect 25023 23752 25024 23792
rect 24982 23743 25024 23752
rect 25114 23792 25172 23793
rect 25114 23752 25123 23792
rect 25163 23752 25172 23792
rect 25114 23751 25172 23752
rect 25225 23792 25267 23801
rect 25225 23752 25226 23792
rect 25266 23752 25267 23792
rect 25225 23743 25267 23752
rect 25515 23792 25557 23801
rect 25515 23752 25516 23792
rect 25556 23752 25557 23792
rect 25515 23743 25557 23752
rect 25649 23792 25707 23793
rect 25649 23752 25658 23792
rect 25698 23752 25707 23792
rect 25649 23751 25707 23752
rect 26187 23792 26229 23801
rect 26187 23752 26188 23792
rect 26228 23752 26229 23792
rect 26187 23743 26229 23752
rect 26379 23792 26421 23801
rect 26379 23752 26380 23792
rect 26420 23752 26421 23792
rect 26379 23743 26421 23752
rect 26667 23792 26709 23801
rect 26667 23752 26668 23792
rect 26708 23752 26709 23792
rect 26667 23743 26709 23752
rect 27243 23792 27285 23801
rect 27243 23752 27244 23792
rect 27284 23752 27285 23792
rect 27243 23743 27285 23752
rect 27418 23792 27476 23793
rect 27418 23752 27427 23792
rect 27467 23752 27476 23792
rect 27418 23751 27476 23752
rect 27531 23792 27573 23801
rect 27531 23752 27532 23792
rect 27572 23752 27573 23792
rect 27531 23743 27573 23752
rect 27867 23792 27909 23801
rect 27867 23752 27868 23792
rect 27908 23752 27909 23792
rect 27867 23743 27909 23752
rect 28002 23792 28060 23793
rect 28002 23752 28011 23792
rect 28051 23752 28060 23792
rect 28002 23751 28060 23752
rect 28378 23792 28436 23793
rect 28378 23752 28387 23792
rect 28427 23752 28436 23792
rect 28378 23751 28436 23752
rect 28697 23792 28739 23801
rect 28697 23752 28698 23792
rect 28738 23752 28739 23792
rect 28697 23743 28739 23752
rect 29338 23792 29396 23793
rect 29338 23752 29347 23792
rect 29387 23752 29396 23792
rect 29338 23751 29396 23752
rect 3531 23734 3573 23743
rect 634 23708 692 23709
rect 634 23668 643 23708
rect 683 23668 692 23708
rect 634 23667 692 23668
rect 3435 23708 3477 23717
rect 3435 23668 3436 23708
rect 3476 23668 3477 23708
rect 3435 23659 3477 23668
rect 4779 23708 4821 23717
rect 4779 23668 4780 23708
rect 4820 23668 4821 23708
rect 4779 23659 4821 23668
rect 5248 23708 5290 23717
rect 5248 23668 5249 23708
rect 5289 23668 5290 23708
rect 5248 23659 5290 23668
rect 10042 23708 10100 23709
rect 10042 23668 10051 23708
rect 10091 23668 10100 23708
rect 10042 23667 10100 23668
rect 13498 23708 13556 23709
rect 13498 23668 13507 23708
rect 13547 23668 13556 23708
rect 13498 23667 13556 23668
rect 24061 23708 24103 23717
rect 24061 23668 24062 23708
rect 24102 23668 24103 23708
rect 24061 23659 24103 23668
rect 24154 23708 24212 23709
rect 24154 23668 24163 23708
rect 24203 23668 24212 23708
rect 24154 23667 24212 23668
rect 28587 23708 28629 23717
rect 28587 23668 28588 23708
rect 28628 23668 28629 23708
rect 28587 23659 28629 23668
rect 5451 23624 5493 23633
rect 5451 23584 5452 23624
rect 5492 23584 5493 23624
rect 5451 23575 5493 23584
rect 8139 23624 8181 23633
rect 8139 23584 8140 23624
rect 8180 23584 8181 23624
rect 8139 23575 8181 23584
rect 8698 23624 8756 23625
rect 8698 23584 8707 23624
rect 8747 23584 8756 23624
rect 8698 23583 8756 23584
rect 11595 23624 11637 23633
rect 11595 23584 11596 23624
rect 11636 23584 11637 23624
rect 11595 23575 11637 23584
rect 15226 23624 15284 23625
rect 15226 23584 15235 23624
rect 15275 23584 15284 23624
rect 15226 23583 15284 23584
rect 17739 23624 17781 23633
rect 17739 23584 17740 23624
rect 17780 23584 17781 23624
rect 17739 23575 17781 23584
rect 19066 23624 19124 23625
rect 19066 23584 19075 23624
rect 19115 23584 19124 23624
rect 19066 23583 19124 23584
rect 20811 23624 20853 23633
rect 20811 23584 20812 23624
rect 20852 23584 20853 23624
rect 20811 23575 20853 23584
rect 23290 23624 23348 23625
rect 23290 23584 23299 23624
rect 23339 23584 23348 23624
rect 23290 23583 23348 23584
rect 24267 23624 24309 23633
rect 24267 23584 24268 23624
rect 24308 23584 24309 23624
rect 24267 23575 24309 23584
rect 25306 23624 25364 23625
rect 25306 23584 25315 23624
rect 25355 23584 25364 23624
rect 25306 23583 25364 23584
rect 25803 23624 25845 23633
rect 25803 23584 25804 23624
rect 25844 23584 25845 23624
rect 25803 23575 25845 23584
rect 26187 23624 26229 23633
rect 26187 23584 26188 23624
rect 26228 23584 26229 23624
rect 26187 23575 26229 23584
rect 26554 23624 26612 23625
rect 26554 23584 26563 23624
rect 26603 23584 26612 23624
rect 26554 23583 26612 23584
rect 26859 23624 26901 23633
rect 26859 23584 26860 23624
rect 26900 23584 26901 23624
rect 26859 23575 26901 23584
rect 27915 23624 27957 23633
rect 27915 23584 27916 23624
rect 27956 23584 27957 23624
rect 27915 23575 27957 23584
rect 28474 23624 28532 23625
rect 28474 23584 28483 23624
rect 28523 23584 28532 23624
rect 28474 23583 28532 23584
rect 576 23456 31392 23480
rect 576 23416 4352 23456
rect 4720 23416 12126 23456
rect 12494 23416 19900 23456
rect 20268 23416 27674 23456
rect 28042 23416 31392 23456
rect 576 23392 31392 23416
rect 4858 23288 4916 23289
rect 4858 23248 4867 23288
rect 4907 23248 4916 23288
rect 4858 23247 4916 23248
rect 5067 23288 5109 23297
rect 5067 23248 5068 23288
rect 5108 23248 5109 23288
rect 5067 23239 5109 23248
rect 11355 23288 11397 23297
rect 11355 23248 11356 23288
rect 11396 23248 11397 23288
rect 11355 23239 11397 23248
rect 12555 23288 12597 23297
rect 12555 23248 12556 23288
rect 12596 23248 12597 23288
rect 12555 23239 12597 23248
rect 15531 23288 15573 23297
rect 15531 23248 15532 23288
rect 15572 23248 15573 23288
rect 15531 23239 15573 23248
rect 16522 23288 16580 23289
rect 16522 23248 16531 23288
rect 16571 23248 16580 23288
rect 16522 23247 16580 23248
rect 20410 23288 20468 23289
rect 20410 23248 20419 23288
rect 20459 23248 20468 23288
rect 20410 23247 20468 23248
rect 23595 23288 23637 23297
rect 23595 23248 23596 23288
rect 23636 23248 23637 23288
rect 23595 23239 23637 23248
rect 27754 23288 27812 23289
rect 27754 23248 27763 23288
rect 27803 23248 27812 23288
rect 27754 23247 27812 23248
rect 31275 23288 31317 23297
rect 31275 23248 31276 23288
rect 31316 23248 31317 23288
rect 31275 23239 31317 23248
rect 5530 23204 5588 23205
rect 5530 23164 5539 23204
rect 5579 23164 5588 23204
rect 5530 23163 5588 23164
rect 8410 23204 8468 23205
rect 8410 23164 8419 23204
rect 8459 23164 8468 23204
rect 8410 23163 8468 23164
rect 11050 23204 11108 23205
rect 11050 23164 11059 23204
rect 11099 23164 11108 23204
rect 11050 23163 11108 23164
rect 26562 23195 26608 23204
rect 26562 23155 26563 23195
rect 26603 23155 26608 23195
rect 26562 23146 26608 23155
rect 2283 23120 2325 23129
rect 2283 23080 2284 23120
rect 2324 23080 2325 23120
rect 2283 23071 2325 23080
rect 3147 23120 3189 23129
rect 3147 23080 3148 23120
rect 3188 23080 3189 23120
rect 3147 23071 3189 23080
rect 3531 23120 3573 23129
rect 3531 23080 3532 23120
rect 3572 23080 3573 23120
rect 3531 23071 3573 23080
rect 4683 23120 4725 23129
rect 4683 23080 4684 23120
rect 4724 23080 4725 23120
rect 4683 23071 4725 23080
rect 4875 23120 4917 23129
rect 4875 23080 4876 23120
rect 4916 23080 4917 23120
rect 4875 23071 4917 23080
rect 5163 23120 5205 23129
rect 5163 23080 5164 23120
rect 5204 23080 5205 23120
rect 5163 23071 5205 23080
rect 5392 23120 5450 23121
rect 5392 23080 5401 23120
rect 5441 23080 5450 23120
rect 5392 23079 5450 23080
rect 5914 23120 5972 23121
rect 5914 23080 5923 23120
rect 5963 23080 5972 23120
rect 5914 23079 5972 23080
rect 8043 23120 8085 23129
rect 8043 23080 8044 23120
rect 8084 23080 8085 23120
rect 8043 23071 8085 23080
rect 8794 23120 8852 23121
rect 8794 23080 8803 23120
rect 8843 23080 8852 23120
rect 8794 23079 8852 23080
rect 11215 23120 11273 23121
rect 11215 23080 11224 23120
rect 11264 23080 11273 23120
rect 11215 23079 11273 23080
rect 11773 23120 11815 23129
rect 11773 23080 11774 23120
rect 11814 23080 11815 23120
rect 11773 23071 11815 23080
rect 11885 23120 11927 23129
rect 11885 23080 11886 23120
rect 11926 23080 11927 23120
rect 11885 23071 11927 23080
rect 12075 23120 12117 23129
rect 12075 23080 12076 23120
rect 12116 23080 12117 23120
rect 12075 23071 12117 23080
rect 12267 23120 12309 23129
rect 12267 23080 12268 23120
rect 12308 23080 12309 23120
rect 12508 23120 12566 23121
rect 12267 23071 12309 23080
rect 12411 23099 12453 23108
rect 12411 23059 12412 23099
rect 12452 23059 12453 23099
rect 12508 23080 12517 23120
rect 12557 23080 12566 23120
rect 12508 23079 12566 23080
rect 12747 23120 12789 23129
rect 12747 23080 12748 23120
rect 12788 23080 12789 23120
rect 12747 23071 12789 23080
rect 12862 23120 12920 23121
rect 12862 23080 12871 23120
rect 12911 23080 12920 23120
rect 12862 23079 12920 23080
rect 12987 23120 13029 23129
rect 12987 23080 12988 23120
rect 13028 23080 13029 23120
rect 12987 23071 13029 23080
rect 13594 23120 13652 23121
rect 13594 23080 13603 23120
rect 13643 23080 13652 23120
rect 13594 23079 13652 23080
rect 16717 23120 16775 23121
rect 16717 23080 16726 23120
rect 16766 23080 16775 23120
rect 16717 23079 16775 23080
rect 17355 23120 17397 23129
rect 17787 23120 17829 23129
rect 17355 23080 17356 23120
rect 17396 23080 17397 23120
rect 17355 23071 17397 23080
rect 17634 23111 17680 23120
rect 17634 23071 17635 23111
rect 17675 23071 17680 23111
rect 17787 23080 17788 23120
rect 17828 23080 17829 23120
rect 17787 23071 17829 23080
rect 18298 23120 18356 23121
rect 18298 23080 18307 23120
rect 18347 23080 18356 23120
rect 18298 23079 18356 23080
rect 18411 23120 18453 23129
rect 18411 23080 18412 23120
rect 18452 23080 18453 23120
rect 18411 23071 18453 23080
rect 19035 23120 19077 23129
rect 19035 23080 19036 23120
rect 19076 23080 19077 23120
rect 19035 23071 19077 23080
rect 19179 23120 19221 23129
rect 19179 23080 19180 23120
rect 19220 23080 19221 23120
rect 19179 23071 19221 23080
rect 19834 23120 19892 23121
rect 19834 23080 19843 23120
rect 19883 23080 19892 23120
rect 19834 23079 19892 23080
rect 19947 23120 19989 23129
rect 19947 23080 19948 23120
rect 19988 23080 19989 23120
rect 19947 23071 19989 23080
rect 20571 23120 20613 23129
rect 20571 23080 20572 23120
rect 20612 23080 20613 23120
rect 20571 23071 20613 23080
rect 20715 23120 20757 23129
rect 20715 23080 20716 23120
rect 20756 23080 20757 23120
rect 20715 23071 20757 23080
rect 21291 23120 21333 23129
rect 21291 23080 21292 23120
rect 21332 23080 21333 23120
rect 21291 23071 21333 23080
rect 21520 23120 21578 23121
rect 21520 23080 21529 23120
rect 21569 23080 21578 23120
rect 21520 23079 21578 23080
rect 21670 23120 21712 23129
rect 21670 23080 21671 23120
rect 21711 23080 21712 23120
rect 21670 23071 21712 23080
rect 21867 23120 21909 23129
rect 21867 23080 21868 23120
rect 21908 23080 21909 23120
rect 21867 23071 21909 23080
rect 22251 23120 22293 23129
rect 22251 23080 22252 23120
rect 22292 23080 22293 23120
rect 22251 23071 22293 23080
rect 22923 23120 22965 23129
rect 22923 23080 22924 23120
rect 22964 23080 22965 23120
rect 22923 23071 22965 23080
rect 23499 23120 23541 23129
rect 23499 23080 23500 23120
rect 23540 23080 23541 23120
rect 23499 23071 23541 23080
rect 23674 23120 23732 23121
rect 23674 23080 23683 23120
rect 23723 23080 23732 23120
rect 23674 23079 23732 23080
rect 24171 23120 24213 23129
rect 24171 23080 24172 23120
rect 24212 23080 24213 23120
rect 24171 23071 24213 23080
rect 24459 23120 24501 23129
rect 24459 23080 24460 23120
rect 24500 23080 24501 23120
rect 24459 23071 24501 23080
rect 24634 23120 24692 23121
rect 24634 23080 24643 23120
rect 24683 23080 24692 23120
rect 24634 23079 24692 23080
rect 25210 23120 25268 23121
rect 25210 23080 25219 23120
rect 25259 23080 25268 23120
rect 25210 23079 25268 23080
rect 25498 23120 25556 23121
rect 25498 23080 25507 23120
rect 25547 23080 25556 23120
rect 25498 23079 25556 23080
rect 25803 23120 25845 23129
rect 25803 23080 25804 23120
rect 25844 23080 25845 23120
rect 25803 23071 25845 23080
rect 25995 23120 26037 23129
rect 25995 23080 25996 23120
rect 26036 23080 26037 23120
rect 25995 23071 26037 23080
rect 26277 23120 26335 23121
rect 26650 23120 26708 23121
rect 26277 23080 26286 23120
rect 26326 23080 26335 23120
rect 26277 23079 26335 23080
rect 26379 23111 26421 23120
rect 26379 23071 26380 23111
rect 26420 23071 26421 23111
rect 26650 23080 26659 23120
rect 26699 23080 26708 23120
rect 26650 23079 26708 23080
rect 26827 23120 26885 23121
rect 26827 23080 26836 23120
rect 26876 23080 26885 23120
rect 26827 23079 26885 23080
rect 27147 23120 27189 23129
rect 27147 23080 27148 23120
rect 27188 23080 27189 23120
rect 27147 23071 27189 23080
rect 27339 23120 27381 23129
rect 27339 23080 27340 23120
rect 27380 23080 27381 23120
rect 27339 23071 27381 23080
rect 27919 23120 27977 23121
rect 27919 23080 27928 23120
rect 27968 23080 27977 23120
rect 27919 23079 27977 23080
rect 28107 23120 28149 23129
rect 28107 23080 28108 23120
rect 28148 23080 28149 23120
rect 28107 23071 28149 23080
rect 28779 23120 28821 23129
rect 28779 23080 28780 23120
rect 28820 23080 28821 23120
rect 28779 23071 28821 23080
rect 28971 23120 29013 23129
rect 28971 23080 28972 23120
rect 29012 23080 29013 23120
rect 28971 23071 29013 23080
rect 29338 23120 29396 23121
rect 29338 23080 29347 23120
rect 29387 23080 29396 23120
rect 29338 23079 29396 23080
rect 17634 23062 17680 23071
rect 26379 23062 26421 23071
rect 12411 23050 12453 23059
rect 5282 23036 5324 23045
rect 5282 22996 5283 23036
rect 5323 22996 5324 23036
rect 5282 22987 5324 22996
rect 7467 23036 7509 23045
rect 7467 22996 7468 23036
rect 7508 22996 7509 23036
rect 7467 22987 7509 22996
rect 10347 23036 10389 23045
rect 10347 22996 10348 23036
rect 10388 22996 10389 23036
rect 10347 22987 10389 22996
rect 11595 23036 11637 23045
rect 11595 22996 11596 23036
rect 11636 22996 11637 23036
rect 11595 22987 11637 22996
rect 13227 23036 13269 23045
rect 13227 22996 13228 23036
rect 13268 22996 13269 23036
rect 13227 22987 13269 22996
rect 21195 23036 21237 23045
rect 21195 22996 21196 23036
rect 21236 22996 21237 23036
rect 21195 22987 21237 22996
rect 21410 23036 21452 23045
rect 21410 22996 21411 23036
rect 21451 22996 21452 23036
rect 21410 22987 21452 22996
rect 24315 23036 24357 23045
rect 24315 22996 24316 23036
rect 24356 22996 24357 23036
rect 24315 22987 24357 22996
rect 25035 23036 25077 23045
rect 25035 22996 25036 23036
rect 25076 22996 25077 23036
rect 25035 22987 25077 22996
rect 25611 23036 25653 23045
rect 25611 22996 25612 23036
rect 25652 22996 25653 23036
rect 25611 22987 25653 22996
rect 2091 22952 2133 22961
rect 2091 22912 2092 22952
rect 2132 22912 2133 22952
rect 2091 22903 2133 22912
rect 7851 22952 7893 22961
rect 7851 22912 7852 22952
rect 7892 22912 7893 22952
rect 7851 22903 7893 22912
rect 10731 22952 10773 22961
rect 10731 22912 10732 22952
rect 10772 22912 10773 22952
rect 10731 22903 10773 22912
rect 11979 22952 12021 22961
rect 11979 22912 11980 22952
rect 12020 22912 12021 22952
rect 11979 22903 12021 22912
rect 13035 22952 13077 22961
rect 13035 22912 13036 22952
rect 13076 22912 13077 22952
rect 13035 22903 13077 22912
rect 18586 22952 18644 22953
rect 18586 22912 18595 22952
rect 18635 22912 18644 22952
rect 18586 22911 18644 22912
rect 24634 22952 24692 22953
rect 24634 22912 24643 22952
rect 24683 22912 24692 22952
rect 24634 22911 24692 22912
rect 2955 22868 2997 22877
rect 2955 22828 2956 22868
rect 2996 22828 2997 22868
rect 2955 22819 2997 22828
rect 3771 22868 3813 22877
rect 3771 22828 3772 22868
rect 3812 22828 3813 22868
rect 3771 22819 3813 22828
rect 8187 22868 8229 22877
rect 8187 22828 8188 22868
rect 8228 22828 8229 22868
rect 8187 22819 8229 22828
rect 16954 22868 17012 22869
rect 16954 22828 16963 22868
rect 17003 22828 17012 22868
rect 16954 22827 17012 22828
rect 19066 22868 19124 22869
rect 19066 22828 19075 22868
rect 19115 22828 19124 22868
rect 19066 22827 19124 22828
rect 20122 22868 20180 22869
rect 20122 22828 20131 22868
rect 20171 22828 20180 22868
rect 20122 22827 20180 22828
rect 21771 22868 21813 22877
rect 21771 22828 21772 22868
rect 21812 22828 21813 22868
rect 21771 22819 21813 22828
rect 25803 22868 25845 22877
rect 25803 22828 25804 22868
rect 25844 22828 25845 22868
rect 25803 22819 25845 22828
rect 26266 22868 26324 22869
rect 26266 22828 26275 22868
rect 26315 22828 26324 22868
rect 26266 22827 26324 22828
rect 27243 22868 27285 22877
rect 27243 22828 27244 22868
rect 27284 22828 27285 22868
rect 27243 22819 27285 22828
rect 30891 22868 30933 22877
rect 30891 22828 30892 22868
rect 30932 22828 30933 22868
rect 30891 22819 30933 22828
rect 576 22700 31392 22724
rect 576 22660 3112 22700
rect 3480 22660 10886 22700
rect 11254 22660 18660 22700
rect 19028 22660 26434 22700
rect 26802 22660 31392 22700
rect 576 22636 31392 22660
rect 843 22532 885 22541
rect 843 22492 844 22532
rect 884 22492 885 22532
rect 843 22483 885 22492
rect 14842 22532 14900 22533
rect 14842 22492 14851 22532
rect 14891 22492 14900 22532
rect 14842 22491 14900 22492
rect 19371 22532 19413 22541
rect 19371 22492 19372 22532
rect 19412 22492 19413 22532
rect 19371 22483 19413 22492
rect 24651 22532 24693 22541
rect 24651 22492 24652 22532
rect 24692 22492 24693 22532
rect 24651 22483 24693 22492
rect 25594 22532 25652 22533
rect 25594 22492 25603 22532
rect 25643 22492 25652 22532
rect 25594 22491 25652 22492
rect 4011 22448 4053 22457
rect 4011 22408 4012 22448
rect 4052 22408 4053 22448
rect 4011 22399 4053 22408
rect 6507 22448 6549 22457
rect 6507 22408 6508 22448
rect 6548 22408 6549 22448
rect 6507 22399 6549 22408
rect 11355 22448 11397 22457
rect 11355 22408 11356 22448
rect 11396 22408 11397 22448
rect 11355 22399 11397 22408
rect 12939 22448 12981 22457
rect 25210 22448 25268 22449
rect 12939 22408 12940 22448
rect 12980 22408 12981 22448
rect 12939 22399 12981 22408
rect 24987 22439 25029 22448
rect 24987 22399 24988 22439
rect 25028 22399 25029 22439
rect 25210 22408 25219 22448
rect 25259 22408 25268 22448
rect 25210 22407 25268 22408
rect 27051 22448 27093 22457
rect 27051 22408 27052 22448
rect 27092 22408 27093 22448
rect 27051 22399 27093 22408
rect 28474 22448 28532 22449
rect 28474 22408 28483 22448
rect 28523 22408 28532 22448
rect 28474 22407 28532 22408
rect 24987 22390 25029 22399
rect 7515 22364 7557 22373
rect 7515 22324 7516 22364
rect 7556 22324 7557 22364
rect 7515 22315 7557 22324
rect 8506 22364 8564 22365
rect 8506 22324 8515 22364
rect 8555 22324 8564 22364
rect 8506 22323 8564 22324
rect 22929 22364 22971 22373
rect 22929 22324 22930 22364
rect 22970 22324 22971 22364
rect 22929 22315 22971 22324
rect 30682 22364 30740 22365
rect 30682 22324 30691 22364
rect 30731 22324 30740 22364
rect 30682 22323 30740 22324
rect 30891 22364 30933 22373
rect 30891 22324 30892 22364
rect 30932 22324 30933 22364
rect 25890 22313 25936 22322
rect 30891 22315 30933 22324
rect 2746 22280 2804 22281
rect 2746 22240 2755 22280
rect 2795 22240 2804 22280
rect 2746 22239 2804 22240
rect 3610 22280 3668 22281
rect 3610 22240 3619 22280
rect 3659 22240 3668 22280
rect 3610 22239 3668 22240
rect 4282 22280 4340 22281
rect 4282 22240 4291 22280
rect 4331 22240 4340 22280
rect 4282 22239 4340 22240
rect 4395 22280 4437 22289
rect 4395 22240 4396 22280
rect 4436 22240 4437 22280
rect 4395 22231 4437 22240
rect 4971 22280 5013 22289
rect 4971 22240 4972 22280
rect 5012 22240 5013 22280
rect 4971 22231 5013 22240
rect 5835 22280 5877 22289
rect 5835 22240 5836 22280
rect 5876 22240 5877 22280
rect 5835 22231 5877 22240
rect 6027 22280 6069 22289
rect 6027 22240 6028 22280
rect 6068 22240 6069 22280
rect 6027 22231 6069 22240
rect 7659 22280 7701 22289
rect 7659 22240 7660 22280
rect 7700 22240 7701 22280
rect 7659 22231 7701 22240
rect 8374 22280 8416 22289
rect 8374 22240 8375 22280
rect 8415 22240 8416 22280
rect 8374 22231 8416 22240
rect 8619 22280 8661 22289
rect 8619 22240 8620 22280
rect 8660 22240 8661 22280
rect 8619 22231 8661 22240
rect 10155 22280 10197 22289
rect 10155 22240 10156 22280
rect 10196 22240 10197 22280
rect 10155 22231 10197 22240
rect 10443 22280 10485 22289
rect 10443 22240 10444 22280
rect 10484 22240 10485 22280
rect 10443 22231 10485 22240
rect 10812 22280 10854 22289
rect 10812 22240 10813 22280
rect 10853 22240 10854 22280
rect 10812 22231 10854 22240
rect 10923 22280 10965 22289
rect 10923 22240 10924 22280
rect 10964 22240 10965 22280
rect 10923 22231 10965 22240
rect 11499 22280 11541 22289
rect 11499 22240 11500 22280
rect 11540 22240 11541 22280
rect 11499 22231 11541 22240
rect 12171 22280 12213 22289
rect 12171 22240 12172 22280
rect 12212 22240 12213 22280
rect 12171 22231 12213 22240
rect 12315 22280 12357 22289
rect 12315 22240 12316 22280
rect 12356 22240 12357 22280
rect 12315 22231 12357 22240
rect 12751 22280 12809 22281
rect 12751 22240 12760 22280
rect 12800 22240 12809 22280
rect 12751 22239 12809 22240
rect 12925 22280 12967 22289
rect 12925 22240 12926 22280
rect 12966 22240 12967 22280
rect 12925 22231 12967 22240
rect 13035 22280 13077 22289
rect 13035 22240 13036 22280
rect 13076 22240 13077 22280
rect 13035 22231 13077 22240
rect 13237 22280 13279 22289
rect 13237 22240 13238 22280
rect 13278 22240 13279 22280
rect 13237 22231 13279 22240
rect 15243 22280 15285 22289
rect 15243 22240 15244 22280
rect 15284 22240 15285 22280
rect 15243 22231 15285 22240
rect 16090 22280 16148 22281
rect 16090 22240 16099 22280
rect 16139 22240 16148 22280
rect 16090 22239 16148 22240
rect 18699 22280 18741 22289
rect 18699 22240 18700 22280
rect 18740 22240 18741 22280
rect 18699 22231 18741 22240
rect 19066 22280 19124 22281
rect 19066 22240 19075 22280
rect 19115 22240 19124 22280
rect 19066 22239 19124 22240
rect 19179 22280 19221 22289
rect 19179 22240 19180 22280
rect 19220 22240 19221 22280
rect 19179 22231 19221 22240
rect 21099 22280 21141 22289
rect 21099 22240 21100 22280
rect 21140 22240 21141 22280
rect 21099 22231 21141 22240
rect 21291 22280 21333 22289
rect 21291 22240 21292 22280
rect 21332 22240 21333 22280
rect 21291 22231 21333 22240
rect 21430 22280 21472 22289
rect 21430 22240 21431 22280
rect 21471 22240 21472 22280
rect 21430 22231 21472 22240
rect 21562 22280 21620 22281
rect 21562 22240 21571 22280
rect 21611 22240 21620 22280
rect 21562 22239 21620 22240
rect 21675 22280 21717 22289
rect 21675 22240 21676 22280
rect 21716 22240 21717 22280
rect 21675 22231 21717 22240
rect 22138 22280 22196 22281
rect 22138 22240 22147 22280
rect 22187 22240 22196 22280
rect 22138 22239 22196 22240
rect 22251 22280 22293 22289
rect 22251 22240 22252 22280
rect 22292 22240 22293 22280
rect 22251 22231 22293 22240
rect 23019 22280 23061 22289
rect 23019 22240 23020 22280
rect 23060 22240 23061 22280
rect 23019 22231 23061 22240
rect 23499 22280 23541 22289
rect 23499 22240 23500 22280
rect 23540 22240 23541 22280
rect 23499 22231 23541 22240
rect 23691 22280 23733 22289
rect 23691 22240 23692 22280
rect 23732 22240 23733 22280
rect 23691 22231 23733 22240
rect 24459 22280 24501 22289
rect 24459 22240 24460 22280
rect 24500 22240 24501 22280
rect 24459 22231 24501 22240
rect 24762 22280 24804 22289
rect 24762 22240 24763 22280
rect 24803 22240 24804 22280
rect 24762 22231 24804 22240
rect 25018 22280 25076 22281
rect 25018 22240 25027 22280
rect 25067 22240 25076 22280
rect 25890 22273 25891 22313
rect 25931 22273 25936 22313
rect 25890 22264 25936 22273
rect 25987 22280 26045 22281
rect 25018 22239 25076 22240
rect 25987 22240 25996 22280
rect 26036 22240 26045 22280
rect 25987 22239 26045 22240
rect 26554 22280 26612 22281
rect 26554 22240 26563 22280
rect 26603 22240 26612 22280
rect 26554 22239 26612 22240
rect 26746 22280 26804 22281
rect 26746 22240 26755 22280
rect 26795 22240 26804 22280
rect 26746 22239 26804 22240
rect 27178 22280 27236 22281
rect 27178 22240 27187 22280
rect 27227 22240 27236 22280
rect 27178 22239 27236 22240
rect 27382 22280 27424 22289
rect 27382 22240 27383 22280
rect 27423 22240 27424 22280
rect 27382 22231 27424 22240
rect 27496 22280 27554 22281
rect 27496 22240 27505 22280
rect 27545 22240 27554 22280
rect 27496 22239 27554 22240
rect 27627 22280 27669 22289
rect 27627 22240 27628 22280
rect 27668 22240 27669 22280
rect 27627 22231 27669 22240
rect 28186 22280 28244 22281
rect 28186 22240 28195 22280
rect 28235 22240 28244 22280
rect 28186 22239 28244 22240
rect 28299 22280 28341 22289
rect 28299 22240 28300 22280
rect 28340 22240 28341 22280
rect 28299 22231 28341 22240
rect 29451 22280 29493 22289
rect 29451 22240 29452 22280
rect 29492 22240 29493 22280
rect 29451 22231 29493 22240
rect 30411 22280 30453 22289
rect 30411 22240 30412 22280
rect 30452 22240 30453 22280
rect 30411 22231 30453 22240
rect 30550 22280 30592 22289
rect 30550 22240 30551 22280
rect 30591 22240 30592 22280
rect 30550 22231 30592 22240
rect 30795 22280 30837 22289
rect 30795 22240 30796 22280
rect 30836 22240 30837 22280
rect 30795 22231 30837 22240
rect 31083 22280 31125 22289
rect 31083 22240 31084 22280
rect 31124 22240 31125 22280
rect 31083 22231 31125 22240
rect 31275 22280 31317 22289
rect 31275 22240 31276 22280
rect 31316 22240 31317 22280
rect 31275 22231 31317 22240
rect 3130 22196 3188 22197
rect 3130 22156 3139 22196
rect 3179 22156 3188 22196
rect 3130 22155 3188 22156
rect 4491 22196 4533 22205
rect 4491 22156 4492 22196
rect 4532 22156 4533 22196
rect 4491 22147 4533 22156
rect 4601 22196 4643 22205
rect 4601 22156 4602 22196
rect 4642 22156 4643 22196
rect 4601 22147 4643 22156
rect 5931 22196 5973 22205
rect 5931 22156 5932 22196
rect 5972 22156 5973 22196
rect 5931 22147 5973 22156
rect 8698 22196 8756 22197
rect 8698 22156 8707 22196
rect 8747 22156 8756 22196
rect 8698 22155 8756 22156
rect 12586 22196 12644 22197
rect 12586 22156 12595 22196
rect 12635 22156 12644 22196
rect 12586 22155 12644 22156
rect 16491 22196 16533 22205
rect 16491 22156 16492 22196
rect 16532 22156 16533 22196
rect 16491 22147 16533 22156
rect 19385 22196 19427 22205
rect 19385 22156 19386 22196
rect 19426 22156 19427 22196
rect 19385 22147 19427 22156
rect 29722 22196 29780 22197
rect 29722 22156 29731 22196
rect 29771 22156 29780 22196
rect 29722 22155 29780 22156
rect 31179 22196 31221 22205
rect 31179 22156 31180 22196
rect 31220 22156 31221 22196
rect 31179 22147 31221 22156
rect 5643 22112 5685 22121
rect 5643 22072 5644 22112
rect 5684 22072 5685 22112
rect 5643 22063 5685 22072
rect 9946 22112 10004 22113
rect 9946 22072 9955 22112
rect 9995 22072 10004 22112
rect 9946 22071 10004 22072
rect 10618 22112 10676 22113
rect 10618 22072 10627 22112
rect 10667 22072 10676 22112
rect 10618 22071 10676 22072
rect 18586 22112 18644 22113
rect 18586 22072 18595 22112
rect 18635 22072 18644 22112
rect 18586 22071 18644 22072
rect 18891 22112 18933 22121
rect 18891 22072 18892 22112
rect 18932 22072 18933 22112
rect 18891 22063 18933 22072
rect 21274 22112 21332 22113
rect 21274 22072 21283 22112
rect 21323 22072 21332 22112
rect 21274 22071 21332 22072
rect 21754 22112 21812 22113
rect 21754 22072 21763 22112
rect 21803 22072 21812 22112
rect 21754 22071 21812 22072
rect 22539 22112 22581 22121
rect 22539 22072 22540 22112
rect 22580 22072 22581 22112
rect 22539 22063 22581 22072
rect 22714 22112 22772 22113
rect 22714 22072 22723 22112
rect 22763 22072 22772 22112
rect 22714 22071 22772 22072
rect 23674 22112 23732 22113
rect 23674 22072 23683 22112
rect 23723 22072 23732 22112
rect 23674 22071 23732 22072
rect 26098 22112 26156 22113
rect 26098 22072 26107 22112
rect 26147 22072 26156 22112
rect 26098 22071 26156 22072
rect 27339 22112 27381 22121
rect 27339 22072 27340 22112
rect 27380 22072 27381 22112
rect 27339 22063 27381 22072
rect 28779 22112 28821 22121
rect 28779 22072 28780 22112
rect 28820 22072 28821 22112
rect 28779 22063 28821 22072
rect 576 21944 31392 21968
rect 576 21904 4352 21944
rect 4720 21904 12126 21944
rect 12494 21904 19900 21944
rect 20268 21904 27674 21944
rect 28042 21904 31392 21944
rect 576 21880 31392 21904
rect 7755 21776 7797 21785
rect 7755 21736 7756 21776
rect 7796 21736 7797 21776
rect 7755 21727 7797 21736
rect 16570 21776 16628 21777
rect 16570 21736 16579 21776
rect 16619 21736 16628 21776
rect 16570 21735 16628 21736
rect 17338 21776 17396 21777
rect 17338 21736 17347 21776
rect 17387 21736 17396 21776
rect 17338 21735 17396 21736
rect 18171 21776 18213 21785
rect 18171 21736 18172 21776
rect 18212 21736 18213 21776
rect 18171 21727 18213 21736
rect 20026 21776 20084 21777
rect 20026 21736 20035 21776
rect 20075 21736 20084 21776
rect 20026 21735 20084 21736
rect 20266 21776 20324 21777
rect 20266 21736 20275 21776
rect 20315 21736 20324 21776
rect 20266 21735 20324 21736
rect 21963 21776 22005 21785
rect 21963 21736 21964 21776
rect 22004 21736 22005 21776
rect 21963 21727 22005 21736
rect 22779 21776 22821 21785
rect 22779 21736 22780 21776
rect 22820 21736 22821 21776
rect 22779 21727 22821 21736
rect 24939 21776 24981 21785
rect 24939 21736 24940 21776
rect 24980 21736 24981 21776
rect 24939 21727 24981 21736
rect 25498 21776 25556 21777
rect 25498 21736 25507 21776
rect 25547 21736 25556 21776
rect 25498 21735 25556 21736
rect 28971 21776 29013 21785
rect 28971 21736 28972 21776
rect 29012 21736 29013 21776
rect 28971 21727 29013 21736
rect 29914 21776 29972 21777
rect 29914 21736 29923 21776
rect 29963 21736 29972 21776
rect 29914 21735 29972 21736
rect 30459 21776 30501 21785
rect 30459 21736 30460 21776
rect 30500 21736 30501 21776
rect 30459 21727 30501 21736
rect 4186 21692 4244 21693
rect 4186 21652 4195 21692
rect 4235 21652 4244 21692
rect 4186 21651 4244 21652
rect 5434 21692 5492 21693
rect 5434 21652 5443 21692
rect 5483 21652 5492 21692
rect 5434 21651 5492 21652
rect 21387 21692 21429 21701
rect 21387 21652 21388 21692
rect 21428 21652 21429 21692
rect 21387 21643 21429 21652
rect 29821 21692 29863 21701
rect 29821 21652 29822 21692
rect 29862 21652 29863 21692
rect 29821 21643 29863 21652
rect 30027 21692 30069 21701
rect 30027 21652 30028 21692
rect 30068 21652 30069 21692
rect 30027 21643 30069 21652
rect 30922 21692 30980 21693
rect 30922 21652 30931 21692
rect 30971 21652 30980 21692
rect 30922 21651 30980 21652
rect 1707 21608 1749 21617
rect 1707 21568 1708 21608
rect 1748 21568 1749 21608
rect 1707 21559 1749 21568
rect 4107 21608 4149 21617
rect 4107 21568 4108 21608
rect 4148 21568 4149 21608
rect 4107 21559 4149 21568
rect 4282 21608 4340 21609
rect 4282 21568 4291 21608
rect 4331 21568 4340 21608
rect 4570 21608 4628 21609
rect 4282 21567 4340 21568
rect 4393 21576 4451 21577
rect 4393 21536 4402 21576
rect 4442 21536 4451 21576
rect 4570 21568 4579 21608
rect 4619 21568 4628 21608
rect 4570 21567 4628 21568
rect 4860 21608 4918 21609
rect 4860 21568 4869 21608
rect 4909 21568 4918 21608
rect 4860 21567 4918 21568
rect 5067 21608 5109 21617
rect 5067 21568 5068 21608
rect 5108 21568 5109 21608
rect 5067 21559 5109 21568
rect 5259 21608 5301 21617
rect 5259 21568 5260 21608
rect 5300 21568 5301 21608
rect 5259 21559 5301 21568
rect 5818 21608 5876 21609
rect 5818 21568 5827 21608
rect 5867 21568 5876 21608
rect 5818 21567 5876 21568
rect 9195 21608 9237 21617
rect 9195 21568 9196 21608
rect 9236 21568 9237 21608
rect 9195 21559 9237 21568
rect 9771 21608 9813 21617
rect 11883 21608 11925 21617
rect 9771 21568 9772 21608
rect 9812 21568 9813 21608
rect 9771 21559 9813 21568
rect 11586 21599 11632 21608
rect 11586 21559 11587 21599
rect 11627 21559 11632 21599
rect 11883 21568 11884 21608
rect 11924 21568 11925 21608
rect 11883 21559 11925 21568
rect 13323 21608 13365 21617
rect 13323 21568 13324 21608
rect 13364 21568 13365 21608
rect 13323 21559 13365 21568
rect 13611 21608 13653 21617
rect 13611 21568 13612 21608
rect 13652 21568 13653 21608
rect 13611 21559 13653 21568
rect 16858 21608 16916 21609
rect 16858 21568 16867 21608
rect 16907 21568 16916 21608
rect 16858 21567 16916 21568
rect 17626 21608 17684 21609
rect 19371 21608 19413 21617
rect 17626 21568 17635 21608
rect 17675 21568 17684 21608
rect 17626 21567 17684 21568
rect 18018 21599 18064 21608
rect 18018 21559 18019 21599
rect 18059 21559 18064 21599
rect 19371 21568 19372 21608
rect 19412 21568 19413 21608
rect 19371 21559 19413 21568
rect 19947 21608 19989 21617
rect 19947 21568 19948 21608
rect 19988 21568 19989 21608
rect 19947 21559 19989 21568
rect 20331 21608 20373 21617
rect 20331 21568 20332 21608
rect 20372 21568 20373 21608
rect 20331 21559 20373 21568
rect 20986 21608 21044 21609
rect 20986 21568 20995 21608
rect 21035 21568 21044 21608
rect 20986 21567 21044 21568
rect 21867 21608 21909 21617
rect 21867 21568 21868 21608
rect 21908 21568 21909 21608
rect 21867 21559 21909 21568
rect 22042 21608 22100 21609
rect 22042 21568 22051 21608
rect 22091 21568 22100 21608
rect 22042 21567 22100 21568
rect 22923 21608 22965 21617
rect 22923 21568 22924 21608
rect 22964 21568 22965 21608
rect 22923 21559 22965 21568
rect 24651 21608 24693 21617
rect 24651 21568 24652 21608
rect 24692 21568 24693 21608
rect 24651 21559 24693 21568
rect 24779 21605 24821 21614
rect 24779 21565 24780 21605
rect 24820 21565 24821 21605
rect 11586 21550 11632 21559
rect 18018 21550 18064 21559
rect 24779 21556 24821 21565
rect 25611 21608 25653 21617
rect 25611 21568 25612 21608
rect 25652 21568 25653 21608
rect 25611 21559 25653 21568
rect 25995 21608 26037 21617
rect 25995 21568 25996 21608
rect 26036 21568 26037 21608
rect 25995 21559 26037 21568
rect 26187 21608 26229 21617
rect 26187 21568 26188 21608
rect 26228 21568 26229 21608
rect 26187 21559 26229 21568
rect 26376 21608 26434 21609
rect 26376 21568 26385 21608
rect 26425 21568 26434 21608
rect 26376 21567 26434 21568
rect 26506 21608 26564 21609
rect 26506 21568 26515 21608
rect 26555 21568 26564 21608
rect 26506 21567 26564 21568
rect 26619 21608 26661 21617
rect 27147 21608 27189 21617
rect 26619 21568 26620 21608
rect 26660 21568 26661 21608
rect 26619 21559 26661 21568
rect 26718 21599 26760 21608
rect 26718 21559 26719 21599
rect 26759 21559 26760 21599
rect 27147 21568 27148 21608
rect 27188 21568 27189 21608
rect 27147 21559 27189 21568
rect 27322 21608 27380 21609
rect 27322 21568 27331 21608
rect 27371 21568 27380 21608
rect 27322 21567 27380 21568
rect 27514 21608 27572 21609
rect 27514 21568 27523 21608
rect 27563 21568 27572 21608
rect 27514 21567 27572 21568
rect 27819 21608 27861 21617
rect 27819 21568 27820 21608
rect 27860 21568 27861 21608
rect 27819 21559 27861 21568
rect 28107 21608 28149 21617
rect 28107 21568 28108 21608
rect 28148 21568 28149 21608
rect 28107 21559 28149 21568
rect 28298 21608 28340 21617
rect 28298 21568 28299 21608
rect 28339 21568 28340 21608
rect 28298 21559 28340 21568
rect 28474 21608 28532 21609
rect 28474 21568 28483 21608
rect 28523 21568 28532 21608
rect 28474 21567 28532 21568
rect 28587 21608 28629 21617
rect 28587 21568 28588 21608
rect 28628 21568 28629 21608
rect 28587 21559 28629 21568
rect 29643 21608 29685 21617
rect 31087 21608 31145 21609
rect 29643 21568 29644 21608
rect 29684 21568 29685 21608
rect 29643 21559 29685 21568
rect 30123 21599 30165 21608
rect 30123 21559 30124 21599
rect 30164 21559 30165 21599
rect 26718 21550 26760 21559
rect 30123 21550 30165 21559
rect 30306 21599 30352 21608
rect 30306 21559 30307 21599
rect 30347 21559 30352 21599
rect 31087 21568 31096 21608
rect 31136 21568 31145 21608
rect 31087 21567 31145 21568
rect 30306 21550 30352 21559
rect 4393 21535 4451 21536
rect 9681 21524 9723 21533
rect 9681 21484 9682 21524
rect 9722 21484 9723 21524
rect 9681 21475 9723 21484
rect 11770 21524 11828 21525
rect 11770 21484 11779 21524
rect 11819 21484 11828 21524
rect 11770 21483 11828 21484
rect 12363 21524 12405 21533
rect 12363 21484 12364 21524
rect 12404 21484 12405 21524
rect 12363 21475 12405 21484
rect 16059 21524 16101 21533
rect 16059 21484 16060 21524
rect 16100 21484 16101 21524
rect 16059 21475 16101 21484
rect 16299 21524 16341 21533
rect 16299 21484 16300 21524
rect 16340 21484 16341 21524
rect 16299 21475 16341 21484
rect 16474 21524 16532 21525
rect 16474 21484 16483 21524
rect 16523 21484 16532 21524
rect 16474 21483 16532 21484
rect 17050 21524 17108 21525
rect 17050 21484 17059 21524
rect 17099 21484 17108 21524
rect 17050 21483 17108 21484
rect 17242 21524 17300 21525
rect 17242 21484 17251 21524
rect 17291 21484 17300 21524
rect 17242 21483 17300 21484
rect 17818 21524 17876 21525
rect 17818 21484 17827 21524
rect 17867 21484 17876 21524
rect 17818 21483 17876 21484
rect 25131 21524 25173 21533
rect 25131 21484 25132 21524
rect 25172 21484 25173 21524
rect 25131 21475 25173 21484
rect 2571 21440 2613 21449
rect 2571 21400 2572 21440
rect 2612 21400 2613 21440
rect 2571 21391 2613 21400
rect 4875 21440 4917 21449
rect 4875 21400 4876 21440
rect 4916 21400 4917 21440
rect 4875 21391 4917 21400
rect 14475 21440 14517 21449
rect 14475 21400 14476 21440
rect 14516 21400 14517 21440
rect 14475 21391 14517 21400
rect 16570 21440 16628 21441
rect 16570 21400 16579 21440
rect 16619 21400 16628 21440
rect 16570 21399 16628 21400
rect 19755 21440 19797 21449
rect 19755 21400 19756 21440
rect 19796 21400 19797 21440
rect 19755 21391 19797 21400
rect 20523 21440 20565 21449
rect 20523 21400 20524 21440
rect 20564 21400 20565 21440
rect 20523 21391 20565 21400
rect 22443 21440 22485 21449
rect 22443 21400 22444 21440
rect 22484 21400 22485 21440
rect 22443 21391 22485 21400
rect 25371 21440 25413 21449
rect 25371 21400 25372 21440
rect 25412 21400 25413 21440
rect 25371 21391 25413 21400
rect 27819 21440 27861 21449
rect 27819 21400 27820 21440
rect 27860 21400 27861 21440
rect 27819 21391 27861 21400
rect 2379 21356 2421 21365
rect 2379 21316 2380 21356
rect 2420 21316 2421 21356
rect 2379 21307 2421 21316
rect 5067 21356 5109 21365
rect 5067 21316 5068 21356
rect 5108 21316 5109 21356
rect 5067 21307 5109 21316
rect 7371 21356 7413 21365
rect 7371 21316 7372 21356
rect 7412 21316 7413 21356
rect 7371 21307 7413 21316
rect 7755 21356 7797 21365
rect 7755 21316 7756 21356
rect 7796 21316 7797 21356
rect 7755 21307 7797 21316
rect 8794 21356 8852 21357
rect 8794 21316 8803 21356
rect 8843 21316 8852 21356
rect 8794 21315 8852 21316
rect 9658 21356 9716 21357
rect 9658 21316 9667 21356
rect 9707 21316 9716 21356
rect 9658 21315 9716 21316
rect 12123 21356 12165 21365
rect 12123 21316 12124 21356
rect 12164 21316 12165 21356
rect 12123 21307 12165 21316
rect 12987 21356 13029 21365
rect 12987 21316 12988 21356
rect 13028 21316 13029 21356
rect 12987 21307 13029 21316
rect 19179 21356 19221 21365
rect 19179 21316 19180 21356
rect 19220 21316 19221 21356
rect 19179 21307 19221 21316
rect 21195 21356 21237 21365
rect 21195 21316 21196 21356
rect 21236 21316 21237 21356
rect 21195 21307 21237 21316
rect 25803 21356 25845 21365
rect 25803 21316 25804 21356
rect 25844 21316 25845 21356
rect 25803 21307 25845 21316
rect 25995 21356 26037 21365
rect 25995 21316 25996 21356
rect 26036 21316 26037 21356
rect 25995 21307 26037 21316
rect 26667 21356 26709 21365
rect 26667 21316 26668 21356
rect 26708 21316 26709 21356
rect 26667 21307 26709 21316
rect 27322 21356 27380 21357
rect 27322 21316 27331 21356
rect 27371 21316 27380 21356
rect 27322 21315 27380 21316
rect 28587 21356 28629 21365
rect 28587 21316 28588 21356
rect 28628 21316 28629 21356
rect 28587 21307 28629 21316
rect 576 21188 31392 21212
rect 576 21148 3112 21188
rect 3480 21148 10886 21188
rect 11254 21148 18660 21188
rect 19028 21148 26434 21188
rect 26802 21148 31392 21188
rect 576 21124 31392 21148
rect 651 21020 693 21029
rect 651 20980 652 21020
rect 692 20980 693 21020
rect 651 20971 693 20980
rect 6219 21020 6261 21029
rect 6219 20980 6220 21020
rect 6260 20980 6261 21020
rect 6219 20971 6261 20980
rect 15723 21020 15765 21029
rect 15723 20980 15724 21020
rect 15764 20980 15765 21020
rect 15723 20971 15765 20980
rect 23691 21020 23733 21029
rect 23691 20980 23692 21020
rect 23732 20980 23733 21020
rect 23691 20971 23733 20980
rect 25899 21020 25941 21029
rect 25899 20980 25900 21020
rect 25940 20980 25941 21020
rect 25899 20971 25941 20980
rect 26859 21020 26901 21029
rect 26859 20980 26860 21020
rect 26900 20980 26901 21020
rect 26859 20971 26901 20980
rect 28203 21020 28245 21029
rect 28203 20980 28204 21020
rect 28244 20980 28245 21020
rect 28203 20971 28245 20980
rect 31275 21020 31317 21029
rect 31275 20980 31276 21020
rect 31316 20980 31317 21020
rect 31275 20971 31317 20980
rect 3771 20936 3813 20945
rect 3771 20896 3772 20936
rect 3812 20896 3813 20936
rect 3771 20887 3813 20896
rect 9243 20936 9285 20945
rect 9243 20896 9244 20936
rect 9284 20896 9285 20936
rect 9243 20887 9285 20896
rect 11674 20936 11732 20937
rect 11674 20896 11683 20936
rect 11723 20896 11732 20936
rect 11674 20895 11732 20896
rect 13227 20936 13269 20945
rect 13227 20896 13228 20936
rect 13268 20896 13269 20936
rect 13227 20887 13269 20896
rect 25035 20936 25077 20945
rect 25035 20896 25036 20936
rect 25076 20896 25077 20936
rect 25035 20887 25077 20896
rect 26667 20936 26709 20945
rect 26667 20896 26668 20936
rect 26708 20896 26709 20936
rect 26667 20887 26709 20896
rect 4474 20852 4532 20853
rect 4474 20812 4483 20852
rect 4523 20812 4532 20852
rect 4474 20811 4532 20812
rect 5434 20852 5492 20853
rect 5434 20812 5443 20852
rect 5483 20812 5492 20852
rect 5434 20811 5492 20812
rect 8122 20852 8180 20853
rect 8122 20812 8131 20852
rect 8171 20812 8180 20852
rect 8122 20811 8180 20812
rect 9003 20852 9045 20861
rect 9003 20812 9004 20852
rect 9044 20812 9045 20852
rect 9003 20803 9045 20812
rect 10347 20852 10389 20861
rect 10347 20812 10348 20852
rect 10388 20812 10389 20852
rect 10347 20803 10389 20812
rect 10810 20852 10868 20853
rect 10810 20812 10819 20852
rect 10859 20812 10868 20852
rect 10810 20811 10868 20812
rect 11386 20852 11444 20853
rect 11386 20812 11395 20852
rect 11435 20812 11444 20852
rect 11386 20811 11444 20812
rect 11578 20852 11636 20853
rect 11578 20812 11587 20852
rect 11627 20812 11636 20852
rect 11578 20811 11636 20812
rect 12154 20852 12212 20853
rect 12154 20812 12163 20852
rect 12203 20812 12212 20852
rect 12154 20811 12212 20812
rect 13419 20852 13461 20861
rect 13419 20812 13420 20852
rect 13460 20812 13461 20852
rect 13419 20803 13461 20812
rect 15339 20852 15381 20861
rect 15339 20812 15340 20852
rect 15380 20812 15381 20852
rect 15339 20803 15381 20812
rect 16299 20852 16341 20861
rect 16299 20812 16300 20852
rect 16340 20812 16341 20852
rect 16299 20803 16341 20812
rect 17259 20852 17301 20861
rect 17259 20812 17260 20852
rect 17300 20812 17301 20852
rect 17259 20803 17301 20812
rect 17835 20852 17877 20861
rect 17835 20812 17836 20852
rect 17876 20812 17877 20852
rect 17835 20803 17877 20812
rect 19306 20852 19364 20853
rect 19306 20812 19315 20852
rect 19355 20812 19364 20852
rect 19306 20811 19364 20812
rect 20642 20852 20684 20861
rect 20642 20812 20643 20852
rect 20683 20812 20684 20852
rect 20642 20803 20684 20812
rect 20986 20852 21044 20853
rect 20986 20812 20995 20852
rect 21035 20812 21044 20852
rect 20986 20811 21044 20812
rect 25611 20852 25653 20861
rect 27418 20852 27476 20853
rect 25611 20812 25612 20852
rect 25652 20812 25653 20852
rect 25611 20803 25653 20812
rect 25746 20843 25792 20852
rect 25746 20803 25747 20843
rect 25787 20803 25792 20843
rect 27418 20812 27427 20852
rect 27467 20812 27476 20852
rect 27418 20811 27476 20812
rect 28971 20852 29013 20861
rect 28971 20812 28972 20852
rect 29012 20812 29013 20852
rect 25746 20794 25792 20803
rect 26371 20801 26413 20810
rect 28971 20803 29013 20812
rect 2554 20768 2612 20769
rect 2554 20728 2563 20768
rect 2603 20728 2612 20768
rect 2554 20727 2612 20728
rect 3147 20768 3189 20777
rect 3147 20728 3148 20768
rect 3188 20728 3189 20768
rect 3147 20719 3189 20728
rect 3531 20768 3573 20777
rect 3531 20728 3532 20768
rect 3572 20728 3573 20768
rect 3531 20719 3573 20728
rect 4683 20768 4725 20777
rect 4683 20728 4684 20768
rect 4724 20728 4725 20768
rect 4683 20719 4725 20728
rect 5302 20768 5344 20777
rect 5302 20728 5303 20768
rect 5343 20728 5344 20768
rect 5302 20719 5344 20728
rect 5547 20768 5589 20777
rect 5547 20728 5548 20768
rect 5588 20728 5589 20768
rect 5547 20719 5589 20728
rect 6891 20768 6933 20777
rect 6891 20728 6892 20768
rect 6932 20728 6933 20768
rect 6891 20719 6933 20728
rect 8002 20768 8060 20769
rect 8002 20728 8011 20768
rect 8051 20728 8060 20768
rect 8002 20727 8060 20728
rect 8235 20768 8277 20777
rect 8235 20728 8236 20768
rect 8276 20728 8277 20768
rect 8235 20719 8277 20728
rect 10443 20768 10485 20777
rect 10443 20728 10444 20768
rect 10484 20728 10485 20768
rect 10443 20719 10485 20728
rect 10562 20768 10604 20777
rect 10562 20728 10563 20768
rect 10603 20728 10604 20768
rect 10562 20719 10604 20728
rect 10672 20768 10730 20769
rect 10672 20728 10681 20768
rect 10721 20728 10730 20768
rect 10672 20727 10730 20728
rect 11194 20768 11252 20769
rect 11194 20728 11203 20768
rect 11243 20728 11252 20768
rect 11194 20727 11252 20728
rect 11962 20768 12020 20769
rect 11962 20728 11971 20768
rect 12011 20728 12020 20768
rect 11962 20727 12020 20728
rect 12555 20768 12597 20777
rect 12555 20728 12556 20768
rect 12596 20728 12597 20768
rect 12555 20719 12597 20728
rect 12826 20768 12884 20769
rect 12826 20728 12835 20768
rect 12875 20728 12884 20768
rect 12826 20727 12884 20728
rect 13786 20768 13844 20769
rect 13786 20728 13795 20768
rect 13835 20728 13844 20768
rect 13786 20727 13844 20728
rect 15958 20768 16000 20777
rect 15958 20728 15959 20768
rect 15999 20728 16000 20768
rect 15958 20719 16000 20728
rect 16090 20768 16148 20769
rect 16090 20728 16099 20768
rect 16139 20728 16148 20768
rect 16090 20727 16148 20728
rect 16203 20768 16245 20777
rect 16203 20728 16204 20768
rect 16244 20728 16245 20768
rect 16203 20719 16245 20728
rect 17434 20768 17492 20769
rect 17434 20728 17443 20768
rect 17483 20728 17492 20768
rect 17434 20727 17492 20728
rect 17722 20768 17780 20769
rect 17722 20728 17731 20768
rect 17771 20728 17780 20768
rect 17722 20727 17780 20728
rect 17962 20768 18020 20769
rect 17962 20728 17971 20768
rect 18011 20728 18020 20768
rect 17962 20727 18020 20728
rect 19501 20768 19559 20769
rect 19501 20728 19510 20768
rect 19550 20728 19559 20768
rect 19501 20727 19559 20728
rect 19659 20768 19701 20777
rect 19659 20728 19660 20768
rect 19700 20728 19701 20768
rect 19659 20719 19701 20728
rect 19851 20768 19893 20777
rect 19851 20728 19852 20768
rect 19892 20728 19893 20768
rect 19851 20719 19893 20728
rect 20523 20768 20565 20777
rect 20523 20728 20524 20768
rect 20564 20728 20565 20768
rect 20523 20719 20565 20728
rect 20740 20768 20782 20777
rect 20740 20728 20741 20768
rect 20781 20728 20782 20768
rect 20740 20719 20782 20728
rect 20866 20768 20924 20769
rect 20866 20728 20875 20768
rect 20915 20728 20924 20768
rect 20866 20727 20924 20728
rect 21099 20768 21141 20777
rect 21099 20728 21100 20768
rect 21140 20728 21141 20768
rect 21099 20719 21141 20728
rect 21754 20768 21812 20769
rect 21754 20728 21763 20768
rect 21803 20728 21812 20768
rect 21754 20727 21812 20728
rect 23883 20768 23925 20777
rect 23883 20728 23884 20768
rect 23924 20728 23925 20768
rect 23883 20719 23925 20728
rect 24555 20768 24597 20777
rect 24555 20728 24556 20768
rect 24596 20728 24597 20768
rect 24555 20719 24597 20728
rect 24826 20768 24884 20769
rect 24826 20728 24835 20768
rect 24875 20728 24884 20768
rect 24826 20727 24884 20728
rect 25515 20768 25557 20777
rect 25515 20728 25516 20768
rect 25556 20728 25557 20768
rect 25515 20719 25557 20728
rect 25846 20768 25904 20769
rect 25846 20728 25855 20768
rect 25895 20728 25904 20768
rect 25846 20727 25904 20728
rect 26091 20768 26133 20777
rect 26091 20728 26092 20768
rect 26132 20728 26133 20768
rect 26091 20719 26133 20728
rect 26245 20768 26303 20769
rect 26245 20728 26254 20768
rect 26294 20728 26303 20768
rect 26371 20761 26372 20801
rect 26412 20761 26413 20801
rect 26371 20752 26413 20761
rect 26465 20768 26523 20769
rect 26245 20727 26303 20728
rect 26465 20728 26474 20768
rect 26514 20728 26523 20768
rect 26465 20727 26523 20728
rect 26902 20768 26944 20777
rect 27147 20768 27189 20777
rect 26902 20728 26903 20768
rect 26943 20728 26944 20768
rect 26902 20719 26944 20728
rect 27042 20759 27088 20768
rect 27042 20719 27043 20759
rect 27083 20719 27088 20759
rect 27147 20728 27148 20768
rect 27188 20728 27189 20768
rect 27147 20719 27189 20728
rect 27286 20768 27328 20777
rect 27286 20728 27287 20768
rect 27327 20728 27328 20768
rect 27286 20719 27328 20728
rect 27531 20768 27573 20777
rect 27531 20728 27532 20768
rect 27572 20728 27573 20768
rect 27531 20719 27573 20728
rect 27819 20768 27861 20777
rect 27819 20728 27820 20768
rect 27860 20728 27861 20768
rect 27819 20719 27861 20728
rect 28012 20768 28070 20769
rect 28012 20728 28021 20768
rect 28061 20728 28070 20768
rect 28012 20727 28070 20728
rect 28203 20768 28245 20777
rect 28203 20728 28204 20768
rect 28244 20728 28245 20768
rect 28203 20719 28245 20728
rect 28491 20768 28533 20777
rect 28491 20728 28492 20768
rect 28532 20728 28533 20768
rect 28491 20719 28533 20728
rect 29338 20768 29396 20769
rect 29338 20728 29347 20768
rect 29387 20728 29396 20768
rect 29338 20727 29396 20728
rect 27042 20710 27088 20719
rect 2938 20684 2996 20685
rect 2938 20644 2947 20684
rect 2987 20644 2996 20684
rect 2938 20643 2996 20644
rect 4282 20684 4340 20685
rect 4282 20644 4291 20684
rect 4331 20644 4340 20684
rect 4282 20643 4340 20644
rect 9243 20684 9285 20693
rect 9243 20644 9244 20684
rect 9284 20644 9285 20684
rect 9243 20635 9285 20644
rect 12939 20684 12981 20693
rect 12939 20644 12940 20684
rect 12980 20644 12981 20684
rect 12939 20635 12981 20644
rect 19755 20684 19797 20693
rect 19755 20644 19756 20684
rect 19796 20644 19797 20684
rect 19755 20635 19797 20644
rect 20427 20684 20469 20693
rect 20427 20644 20428 20684
rect 20468 20644 20469 20684
rect 20427 20635 20469 20644
rect 21178 20684 21236 20685
rect 21178 20644 21187 20684
rect 21227 20644 21236 20684
rect 21178 20643 21236 20644
rect 21370 20684 21428 20685
rect 21370 20644 21379 20684
rect 21419 20644 21428 20684
rect 21370 20643 21428 20644
rect 5626 20600 5684 20601
rect 5626 20560 5635 20600
rect 5675 20560 5684 20600
rect 5626 20559 5684 20560
rect 8314 20600 8372 20601
rect 8314 20560 8323 20600
rect 8363 20560 8372 20600
rect 8314 20559 8372 20560
rect 10906 20600 10964 20601
rect 10906 20560 10915 20600
rect 10955 20560 10964 20600
rect 10906 20559 10964 20560
rect 18171 20600 18213 20609
rect 18171 20560 18172 20600
rect 18212 20560 18213 20600
rect 18171 20551 18213 20560
rect 27610 20600 27668 20601
rect 27610 20560 27619 20600
rect 27659 20560 27668 20600
rect 27610 20559 27668 20560
rect 27819 20600 27861 20609
rect 27819 20560 27820 20600
rect 27860 20560 27861 20600
rect 27819 20551 27861 20560
rect 576 20432 31392 20456
rect 576 20392 4352 20432
rect 4720 20392 12126 20432
rect 12494 20392 19900 20432
rect 20268 20392 27674 20432
rect 28042 20392 31392 20432
rect 576 20368 31392 20392
rect 12730 20264 12788 20265
rect 12730 20224 12739 20264
rect 12779 20224 12788 20264
rect 12730 20223 12788 20224
rect 13402 20264 13460 20265
rect 13402 20224 13411 20264
rect 13451 20224 13460 20264
rect 13402 20223 13460 20224
rect 15706 20264 15764 20265
rect 15706 20224 15715 20264
rect 15755 20224 15764 20264
rect 15706 20223 15764 20224
rect 16779 20264 16821 20273
rect 16779 20224 16780 20264
rect 16820 20224 16821 20264
rect 16779 20215 16821 20224
rect 17530 20264 17588 20265
rect 17530 20224 17539 20264
rect 17579 20224 17588 20264
rect 17530 20223 17588 20224
rect 17739 20264 17781 20273
rect 17739 20224 17740 20264
rect 17780 20224 17781 20264
rect 17739 20215 17781 20224
rect 20379 20264 20421 20273
rect 20379 20224 20380 20264
rect 20420 20224 20421 20264
rect 20379 20215 20421 20224
rect 25018 20264 25076 20265
rect 25018 20224 25027 20264
rect 25067 20224 25076 20264
rect 25018 20223 25076 20224
rect 26859 20264 26901 20273
rect 26859 20224 26860 20264
rect 26900 20224 26901 20264
rect 26859 20215 26901 20224
rect 27130 20264 27188 20265
rect 27130 20224 27139 20264
rect 27179 20224 27188 20264
rect 27130 20223 27188 20224
rect 2667 20180 2709 20189
rect 2667 20140 2668 20180
rect 2708 20140 2709 20180
rect 2667 20131 2709 20140
rect 6699 20180 6741 20189
rect 6699 20140 6700 20180
rect 6740 20140 6741 20180
rect 6699 20131 6741 20140
rect 8698 20180 8756 20181
rect 8698 20140 8707 20180
rect 8747 20140 8756 20180
rect 8698 20139 8756 20140
rect 14362 20180 14420 20181
rect 14362 20140 14371 20180
rect 14411 20140 14420 20180
rect 14362 20139 14420 20140
rect 16491 20180 16533 20189
rect 16491 20140 16492 20180
rect 16532 20140 16533 20180
rect 16491 20131 16533 20140
rect 29626 20180 29684 20181
rect 29626 20140 29635 20180
rect 29675 20140 29684 20180
rect 29626 20139 29684 20140
rect 1803 20096 1845 20105
rect 1803 20056 1804 20096
rect 1844 20056 1845 20096
rect 1803 20047 1845 20056
rect 2032 20096 2090 20097
rect 2032 20056 2041 20096
rect 2081 20056 2090 20096
rect 2032 20055 2090 20056
rect 2283 20096 2325 20105
rect 2283 20056 2284 20096
rect 2324 20056 2325 20096
rect 2283 20047 2325 20056
rect 2554 20096 2612 20097
rect 2554 20056 2563 20096
rect 2603 20056 2612 20096
rect 2554 20055 2612 20056
rect 3370 20096 3428 20097
rect 3370 20056 3379 20096
rect 3419 20056 3428 20096
rect 3370 20055 3428 20056
rect 3565 20096 3623 20097
rect 3565 20056 3574 20096
rect 3614 20056 3623 20096
rect 3565 20055 3623 20056
rect 3819 20096 3861 20105
rect 3819 20056 3820 20096
rect 3860 20056 3861 20096
rect 3819 20047 3861 20056
rect 4048 20096 4106 20097
rect 4048 20056 4057 20096
rect 4097 20056 4106 20096
rect 4048 20055 4106 20056
rect 4299 20096 4341 20105
rect 4299 20056 4300 20096
rect 4340 20056 4341 20096
rect 4299 20047 4341 20056
rect 4491 20096 4533 20105
rect 4491 20056 4492 20096
rect 4532 20056 4533 20096
rect 4491 20047 4533 20056
rect 5146 20096 5204 20097
rect 5146 20056 5155 20096
rect 5195 20056 5204 20096
rect 5146 20055 5204 20056
rect 5914 20096 5972 20097
rect 5914 20056 5923 20096
rect 5963 20056 5972 20096
rect 5914 20055 5972 20056
rect 6493 20096 6535 20105
rect 7083 20096 7125 20105
rect 6493 20056 6494 20096
rect 6534 20056 6535 20096
rect 6493 20047 6535 20056
rect 6795 20087 6837 20096
rect 6795 20047 6796 20087
rect 6836 20047 6837 20087
rect 7083 20056 7084 20096
rect 7124 20056 7125 20096
rect 7083 20047 7125 20056
rect 7275 20096 7317 20105
rect 7275 20056 7276 20096
rect 7316 20056 7317 20096
rect 7275 20047 7317 20056
rect 7738 20096 7796 20097
rect 7738 20056 7747 20096
rect 7787 20056 7796 20096
rect 7738 20055 7796 20056
rect 8986 20096 9044 20097
rect 10443 20096 10485 20105
rect 8986 20056 8995 20096
rect 9035 20056 9044 20096
rect 8986 20055 9044 20056
rect 9378 20087 9424 20096
rect 9378 20047 9379 20087
rect 9419 20047 9424 20087
rect 10443 20056 10444 20096
rect 10484 20056 10485 20096
rect 10443 20047 10485 20056
rect 10635 20096 10677 20105
rect 10635 20056 10636 20096
rect 10676 20056 10677 20096
rect 10635 20047 10677 20056
rect 11002 20096 11060 20097
rect 11002 20056 11011 20096
rect 11051 20056 11060 20096
rect 11002 20055 11060 20056
rect 11290 20096 11348 20097
rect 11290 20056 11299 20096
rect 11339 20056 11348 20096
rect 11290 20055 11348 20056
rect 13210 20096 13268 20097
rect 13210 20056 13219 20096
rect 13259 20056 13268 20096
rect 13210 20055 13268 20056
rect 13786 20096 13844 20097
rect 13786 20056 13795 20096
rect 13835 20056 13844 20096
rect 13786 20055 13844 20056
rect 15051 20096 15093 20105
rect 15051 20056 15052 20096
rect 15092 20056 15093 20096
rect 15051 20047 15093 20056
rect 15819 20096 15861 20105
rect 15819 20056 15820 20096
rect 15860 20056 15861 20096
rect 15562 20054 15620 20055
rect 6795 20038 6837 20047
rect 9378 20038 9424 20047
rect 1707 20012 1749 20021
rect 3723 20012 3765 20021
rect 4587 20012 4629 20021
rect 1707 19972 1708 20012
rect 1748 19972 1749 20012
rect 1707 19963 1749 19972
rect 1938 20003 1984 20012
rect 1938 19963 1939 20003
rect 1979 19963 1984 20003
rect 3723 19972 3724 20012
rect 3764 19972 3765 20012
rect 3723 19963 3765 19972
rect 3954 20003 4000 20012
rect 3954 19963 3955 20003
rect 3995 19963 4000 20003
rect 4587 19972 4588 20012
rect 4628 19972 4629 20012
rect 4587 19963 4629 19972
rect 4971 20012 5013 20021
rect 4971 19972 4972 20012
rect 5012 19972 5013 20012
rect 4971 19963 5013 19972
rect 5547 20012 5589 20021
rect 5547 19972 5548 20012
rect 5588 19972 5589 20012
rect 5547 19963 5589 19972
rect 5739 20012 5781 20021
rect 5739 19972 5740 20012
rect 5780 19972 5781 20012
rect 5739 19963 5781 19972
rect 6315 20012 6357 20021
rect 6315 19972 6316 20012
rect 6356 19972 6357 20012
rect 6315 19963 6357 19972
rect 7563 20012 7605 20021
rect 7563 19972 7564 20012
rect 7604 19972 7605 20012
rect 7563 19963 7605 19972
rect 8139 20012 8181 20021
rect 8139 19972 8140 20012
rect 8180 19972 8181 20012
rect 8139 19963 8181 19972
rect 8602 20012 8660 20013
rect 8602 19972 8611 20012
rect 8651 19972 8660 20012
rect 8602 19971 8660 19972
rect 9178 20012 9236 20013
rect 9178 19972 9187 20012
rect 9227 19972 9236 20012
rect 9178 19971 9236 19972
rect 9531 20012 9573 20021
rect 9531 19972 9532 20012
rect 9572 19972 9573 20012
rect 9531 19963 9573 19972
rect 10827 20012 10869 20021
rect 10827 19972 10828 20012
rect 10868 19972 10869 20012
rect 10827 19963 10869 19972
rect 11403 20012 11445 20021
rect 11403 19972 11404 20012
rect 11444 19972 11445 20012
rect 11403 19963 11445 19972
rect 13035 20012 13077 20021
rect 13035 19972 13036 20012
rect 13076 19972 13077 20012
rect 13035 19963 13077 19972
rect 13707 20012 13749 20021
rect 15562 20014 15571 20054
rect 15611 20014 15620 20054
rect 15819 20047 15861 20056
rect 16395 20096 16437 20105
rect 16395 20056 16396 20096
rect 16436 20056 16437 20096
rect 16395 20047 16437 20056
rect 16570 20096 16628 20097
rect 16570 20056 16579 20096
rect 16619 20056 16628 20096
rect 16570 20055 16628 20056
rect 16874 20096 16916 20105
rect 16874 20056 16875 20096
rect 16915 20056 16916 20096
rect 16874 20047 16916 20056
rect 17106 20096 17148 20105
rect 17106 20056 17107 20096
rect 17147 20056 17148 20096
rect 17106 20047 17148 20056
rect 17211 20096 17253 20105
rect 17211 20056 17212 20096
rect 17252 20056 17253 20096
rect 17211 20047 17253 20056
rect 17451 20096 17493 20105
rect 17451 20056 17452 20096
rect 17492 20056 17493 20096
rect 17451 20047 17493 20056
rect 17835 20096 17877 20105
rect 17835 20056 17836 20096
rect 17876 20056 17877 20096
rect 17835 20047 17877 20056
rect 17954 20096 17996 20105
rect 17954 20056 17955 20096
rect 17995 20056 17996 20096
rect 17954 20047 17996 20056
rect 18064 20096 18122 20097
rect 19275 20096 19317 20105
rect 18064 20056 18073 20096
rect 18113 20056 18122 20096
rect 18064 20055 18122 20056
rect 18498 20087 18544 20096
rect 18498 20047 18499 20087
rect 18539 20047 18544 20087
rect 19275 20056 19276 20096
rect 19316 20056 19317 20096
rect 19275 20047 19317 20056
rect 19467 20096 19509 20105
rect 19467 20056 19468 20096
rect 19508 20056 19509 20096
rect 19467 20047 19509 20056
rect 19702 20096 19744 20105
rect 19702 20056 19703 20096
rect 19743 20056 19744 20096
rect 19702 20047 19744 20056
rect 19947 20096 19989 20105
rect 19947 20056 19948 20096
rect 19988 20056 19989 20096
rect 19947 20047 19989 20056
rect 20235 20096 20277 20105
rect 20235 20056 20236 20096
rect 20276 20056 20277 20096
rect 20235 20047 20277 20056
rect 20698 20096 20756 20097
rect 20698 20056 20707 20096
rect 20747 20056 20756 20096
rect 20698 20055 20756 20056
rect 20986 20096 21044 20097
rect 24459 20096 24501 20105
rect 20986 20056 20995 20096
rect 21035 20056 21044 20096
rect 20986 20055 21044 20056
rect 21282 20087 21328 20096
rect 21282 20047 21283 20087
rect 21323 20047 21328 20087
rect 24459 20056 24460 20096
rect 24500 20056 24501 20096
rect 24459 20047 24501 20056
rect 24634 20096 24692 20097
rect 24634 20056 24643 20096
rect 24683 20056 24692 20096
rect 24634 20055 24692 20056
rect 24747 20096 24789 20105
rect 24747 20056 24748 20096
rect 24788 20056 24789 20096
rect 24747 20047 24789 20056
rect 25018 20096 25076 20097
rect 25018 20056 25027 20096
rect 25067 20056 25076 20096
rect 25018 20055 25076 20056
rect 25306 20096 25364 20097
rect 25306 20056 25315 20096
rect 25355 20056 25364 20096
rect 25306 20055 25364 20056
rect 25498 20096 25556 20097
rect 25498 20056 25507 20096
rect 25547 20056 25556 20096
rect 25498 20055 25556 20056
rect 25690 20096 25748 20097
rect 25690 20056 25699 20096
rect 25739 20056 25748 20096
rect 25690 20055 25748 20056
rect 26571 20096 26613 20105
rect 26571 20056 26572 20096
rect 26612 20056 26613 20096
rect 26571 20047 26613 20056
rect 27051 20096 27093 20105
rect 27051 20056 27052 20096
rect 27092 20056 27093 20096
rect 27051 20047 27093 20056
rect 27298 20096 27356 20097
rect 27298 20056 27307 20096
rect 27347 20056 27356 20096
rect 27298 20055 27356 20056
rect 27531 20096 27573 20105
rect 27531 20056 27532 20096
rect 27572 20056 27573 20096
rect 27531 20047 27573 20056
rect 28186 20096 28244 20097
rect 28186 20056 28195 20096
rect 28235 20056 28244 20096
rect 28186 20055 28244 20056
rect 28299 20096 28341 20105
rect 28299 20056 28300 20096
rect 28340 20056 28341 20096
rect 28299 20047 28341 20056
rect 29451 20096 29493 20105
rect 29451 20056 29452 20096
rect 29492 20056 29493 20096
rect 29451 20047 29493 20056
rect 30315 20096 30357 20105
rect 30987 20096 31029 20105
rect 30315 20056 30316 20096
rect 30356 20056 30357 20096
rect 30315 20047 30357 20056
rect 30498 20087 30544 20096
rect 30498 20047 30499 20087
rect 30539 20047 30544 20087
rect 30987 20056 30988 20096
rect 31028 20056 31029 20096
rect 30987 20047 31029 20056
rect 31179 20096 31221 20105
rect 31179 20056 31180 20096
rect 31220 20056 31221 20096
rect 31179 20047 31221 20056
rect 18498 20038 18544 20047
rect 21282 20038 21328 20047
rect 30498 20038 30544 20047
rect 15562 20013 15620 20014
rect 13707 19972 13708 20012
rect 13748 19972 13749 20012
rect 13707 19963 13749 19972
rect 15370 20012 15428 20013
rect 15370 19972 15379 20012
rect 15419 19972 15428 20012
rect 15370 19971 15428 19972
rect 16994 20012 17036 20021
rect 16994 19972 16995 20012
rect 17035 19972 17036 20012
rect 16994 19963 17036 19972
rect 17338 20012 17396 20013
rect 17338 19972 17347 20012
rect 17387 19972 17396 20012
rect 17338 19971 17396 19972
rect 18651 20012 18693 20021
rect 18651 19972 18652 20012
rect 18692 19972 18693 20012
rect 18651 19963 18693 19972
rect 19834 20012 19892 20013
rect 19834 19972 19843 20012
rect 19883 19972 19892 20012
rect 19834 19971 19892 19972
rect 20043 20012 20085 20021
rect 20043 19972 20044 20012
rect 20084 19972 20085 20012
rect 20043 19963 20085 19972
rect 20523 20012 20565 20021
rect 20523 19972 20524 20012
rect 20564 19972 20565 20012
rect 20523 19963 20565 19972
rect 21099 20012 21141 20021
rect 21099 19972 21100 20012
rect 21140 19972 21141 20012
rect 21099 19963 21141 19972
rect 21435 20012 21477 20021
rect 21435 19972 21436 20012
rect 21476 19972 21477 20012
rect 21435 19963 21477 19972
rect 26427 20012 26469 20021
rect 26427 19972 26428 20012
rect 26468 19972 26469 20012
rect 26427 19963 26469 19972
rect 27418 20012 27476 20013
rect 27418 19972 27427 20012
rect 27467 19972 27476 20012
rect 27418 19971 27476 19972
rect 27627 20012 27669 20021
rect 27627 19972 27628 20012
rect 27668 19972 27669 20012
rect 27627 19963 27669 19972
rect 30651 20012 30693 20021
rect 30651 19972 30652 20012
rect 30692 19972 30693 20012
rect 30651 19963 30693 19972
rect 1938 19954 1984 19963
rect 3954 19954 4000 19963
rect 2955 19928 2997 19937
rect 2955 19888 2956 19928
rect 2996 19888 2997 19928
rect 2955 19879 2997 19888
rect 5451 19928 5493 19937
rect 5451 19888 5452 19928
rect 5492 19888 5493 19928
rect 5451 19879 5493 19888
rect 6219 19928 6261 19937
rect 6219 19888 6220 19928
rect 6260 19888 6261 19928
rect 6219 19879 6261 19888
rect 7066 19928 7124 19929
rect 7066 19888 7075 19928
rect 7115 19888 7124 19928
rect 7066 19887 7124 19888
rect 8043 19928 8085 19937
rect 8043 19888 8044 19928
rect 8084 19888 8085 19928
rect 8043 19879 8085 19888
rect 16011 19928 16053 19937
rect 16011 19888 16012 19928
rect 16052 19888 16053 19928
rect 16011 19879 16053 19888
rect 21003 19928 21045 19937
rect 21003 19888 21004 19928
rect 21044 19888 21045 19928
rect 21003 19879 21045 19888
rect 26283 19928 26325 19937
rect 26283 19888 26284 19928
rect 26324 19888 26325 19928
rect 26283 19879 26325 19888
rect 28474 19928 28532 19929
rect 28474 19888 28483 19928
rect 28523 19888 28532 19928
rect 28474 19887 28532 19888
rect 6490 19844 6548 19845
rect 6490 19804 6499 19844
rect 6539 19804 6548 19844
rect 6490 19803 6548 19804
rect 10443 19844 10485 19853
rect 10443 19804 10444 19844
rect 10484 19804 10485 19844
rect 10443 19795 10485 19804
rect 19275 19844 19317 19853
rect 19275 19804 19276 19844
rect 19316 19804 19317 19844
rect 19275 19795 19317 19804
rect 24747 19844 24789 19853
rect 24747 19804 24748 19844
rect 24788 19804 24789 19844
rect 24747 19795 24789 19804
rect 28779 19844 28821 19853
rect 28779 19804 28780 19844
rect 28820 19804 28821 19844
rect 28779 19795 28821 19804
rect 30987 19844 31029 19853
rect 30987 19804 30988 19844
rect 31028 19804 31029 19844
rect 30987 19795 31029 19804
rect 576 19676 31392 19700
rect 576 19636 3112 19676
rect 3480 19636 10886 19676
rect 11254 19636 18660 19676
rect 19028 19636 26434 19676
rect 26802 19636 31392 19676
rect 576 19612 31392 19636
rect 4155 19508 4197 19517
rect 4155 19468 4156 19508
rect 4196 19468 4197 19508
rect 4155 19459 4197 19468
rect 16186 19508 16244 19509
rect 16186 19468 16195 19508
rect 16235 19468 16244 19508
rect 16186 19467 16244 19468
rect 16666 19508 16724 19509
rect 16666 19468 16675 19508
rect 16715 19468 16724 19508
rect 16666 19467 16724 19468
rect 17626 19508 17684 19509
rect 17626 19468 17635 19508
rect 17675 19468 17684 19508
rect 17626 19467 17684 19468
rect 19467 19508 19509 19517
rect 19467 19468 19468 19508
rect 19508 19468 19509 19508
rect 19467 19459 19509 19468
rect 26170 19508 26228 19509
rect 26170 19468 26179 19508
rect 26219 19468 26228 19508
rect 26170 19467 26228 19468
rect 28971 19508 29013 19517
rect 28971 19468 28972 19508
rect 29012 19468 29013 19508
rect 28971 19459 29013 19468
rect 8139 19424 8181 19433
rect 8139 19384 8140 19424
rect 8180 19384 8181 19424
rect 8139 19375 8181 19384
rect 11979 19424 12021 19433
rect 11979 19384 11980 19424
rect 12020 19384 12021 19424
rect 11979 19375 12021 19384
rect 15051 19424 15093 19433
rect 15051 19384 15052 19424
rect 15092 19384 15093 19424
rect 15051 19375 15093 19384
rect 21291 19424 21333 19433
rect 21291 19384 21292 19424
rect 21332 19384 21333 19424
rect 21291 19375 21333 19384
rect 23002 19424 23060 19425
rect 23002 19384 23011 19424
rect 23051 19384 23060 19424
rect 23002 19383 23060 19384
rect 23386 19424 23444 19425
rect 23386 19384 23395 19424
rect 23435 19384 23444 19424
rect 23386 19383 23444 19384
rect 24555 19424 24597 19433
rect 24555 19384 24556 19424
rect 24596 19384 24597 19424
rect 24555 19375 24597 19384
rect 1131 19340 1173 19349
rect 1131 19300 1132 19340
rect 1172 19300 1173 19340
rect 1131 19291 1173 19300
rect 1707 19340 1749 19349
rect 1707 19300 1708 19340
rect 1748 19300 1749 19340
rect 1707 19291 1749 19300
rect 3170 19340 3212 19349
rect 3170 19300 3171 19340
rect 3211 19300 3212 19340
rect 3170 19291 3212 19300
rect 4395 19340 4437 19349
rect 4395 19300 4396 19340
rect 4436 19300 4437 19340
rect 4395 19291 4437 19300
rect 5835 19340 5877 19349
rect 5835 19300 5836 19340
rect 5876 19300 5877 19340
rect 7252 19340 7294 19349
rect 5835 19291 5877 19300
rect 7131 19298 7173 19307
rect 1885 19289 1943 19290
rect 1306 19256 1364 19257
rect 1306 19216 1315 19256
rect 1355 19216 1364 19256
rect 1885 19249 1894 19289
rect 1934 19249 1943 19289
rect 1885 19248 1943 19249
rect 2198 19256 2240 19265
rect 1306 19215 1364 19216
rect 2198 19216 2199 19256
rect 2239 19216 2240 19256
rect 2198 19207 2240 19216
rect 2461 19256 2503 19265
rect 2461 19216 2462 19256
rect 2502 19216 2503 19256
rect 2461 19207 2503 19216
rect 2755 19256 2813 19257
rect 2755 19216 2764 19256
rect 2804 19216 2813 19256
rect 2755 19215 2813 19216
rect 3051 19256 3093 19265
rect 3051 19216 3052 19256
rect 3092 19216 3093 19256
rect 3051 19207 3093 19216
rect 3268 19256 3310 19265
rect 3268 19216 3269 19256
rect 3309 19216 3310 19256
rect 3268 19207 3310 19216
rect 3435 19256 3477 19265
rect 3435 19216 3436 19256
rect 3476 19216 3477 19256
rect 3435 19207 3477 19216
rect 3610 19256 3668 19257
rect 3610 19216 3619 19256
rect 3659 19216 3668 19256
rect 3610 19215 3668 19216
rect 5506 19256 5564 19257
rect 5506 19216 5515 19256
rect 5555 19216 5564 19256
rect 5506 19215 5564 19216
rect 5626 19256 5684 19257
rect 5626 19216 5635 19256
rect 5675 19216 5684 19256
rect 5626 19215 5684 19216
rect 5739 19256 5781 19265
rect 5739 19216 5740 19256
rect 5780 19216 5781 19256
rect 5739 19207 5781 19216
rect 6123 19256 6165 19265
rect 6123 19216 6124 19256
rect 6164 19216 6165 19256
rect 6123 19207 6165 19216
rect 6307 19256 6349 19265
rect 6307 19216 6308 19256
rect 6348 19216 6349 19256
rect 6307 19207 6349 19216
rect 6658 19256 6716 19257
rect 6658 19216 6667 19256
rect 6707 19216 6716 19256
rect 6658 19215 6716 19216
rect 6778 19256 6836 19257
rect 6778 19216 6787 19256
rect 6827 19216 6836 19256
rect 6778 19215 6836 19216
rect 6891 19256 6933 19265
rect 6891 19216 6892 19256
rect 6932 19216 6933 19256
rect 7131 19258 7132 19298
rect 7172 19258 7173 19298
rect 7252 19300 7253 19340
rect 7293 19300 7294 19340
rect 7252 19291 7294 19300
rect 7467 19340 7509 19349
rect 7467 19300 7468 19340
rect 7508 19300 7509 19340
rect 7467 19291 7509 19300
rect 7659 19340 7701 19349
rect 7659 19300 7660 19340
rect 7700 19300 7701 19340
rect 7659 19291 7701 19300
rect 8235 19340 8277 19349
rect 8235 19300 8236 19340
rect 8276 19300 8277 19340
rect 8235 19291 8277 19300
rect 8930 19340 8972 19349
rect 8930 19300 8931 19340
rect 8971 19300 8972 19340
rect 8930 19291 8972 19300
rect 9850 19340 9908 19341
rect 9850 19300 9859 19340
rect 9899 19300 9908 19340
rect 9850 19299 9908 19300
rect 10522 19340 10580 19341
rect 10522 19300 10531 19340
rect 10571 19300 10580 19340
rect 10522 19299 10580 19300
rect 10923 19340 10965 19349
rect 13419 19340 13461 19349
rect 10923 19300 10924 19340
rect 10964 19300 10965 19340
rect 10923 19291 10965 19300
rect 11154 19331 11200 19340
rect 11154 19291 11155 19331
rect 11195 19291 11200 19331
rect 13419 19300 13420 19340
rect 13460 19300 13461 19340
rect 13419 19291 13461 19300
rect 19930 19340 19988 19341
rect 19930 19300 19939 19340
rect 19979 19300 19988 19340
rect 19930 19299 19988 19300
rect 20410 19340 20468 19341
rect 20410 19300 20419 19340
rect 20459 19300 20468 19340
rect 20410 19299 20468 19300
rect 20619 19340 20661 19349
rect 20619 19300 20620 19340
rect 20660 19300 20661 19340
rect 20619 19291 20661 19300
rect 20811 19340 20853 19349
rect 20811 19300 20812 19340
rect 20852 19300 20853 19340
rect 20811 19291 20853 19300
rect 21387 19340 21429 19349
rect 21387 19300 21388 19340
rect 21428 19300 21429 19340
rect 21387 19291 21429 19300
rect 23290 19340 23348 19341
rect 23290 19300 23299 19340
rect 23339 19300 23348 19340
rect 23290 19299 23348 19300
rect 23547 19340 23589 19349
rect 23547 19300 23548 19340
rect 23588 19300 23589 19340
rect 23547 19291 23589 19300
rect 25035 19340 25077 19349
rect 25035 19300 25036 19340
rect 25076 19300 25077 19340
rect 11154 19282 11200 19291
rect 24271 19289 24313 19298
rect 25035 19291 25077 19300
rect 31258 19340 31316 19341
rect 31258 19300 31267 19340
rect 31307 19300 31316 19340
rect 31258 19299 31316 19300
rect 7131 19249 7173 19258
rect 7371 19256 7413 19265
rect 6891 19207 6933 19216
rect 7371 19216 7372 19256
rect 7412 19216 7413 19256
rect 7371 19207 7413 19216
rect 7834 19256 7892 19257
rect 7834 19216 7843 19256
rect 7883 19216 7892 19256
rect 7834 19215 7892 19216
rect 8811 19256 8853 19265
rect 8811 19216 8812 19256
rect 8852 19216 8853 19256
rect 8811 19207 8853 19216
rect 9040 19256 9098 19257
rect 9040 19216 9049 19256
rect 9089 19216 9098 19256
rect 9040 19215 9098 19216
rect 9271 19256 9329 19257
rect 9271 19216 9280 19256
rect 9320 19216 9329 19256
rect 9271 19215 9329 19216
rect 9718 19256 9760 19265
rect 9718 19216 9719 19256
rect 9759 19216 9760 19256
rect 9718 19207 9760 19216
rect 9963 19256 10005 19265
rect 9963 19216 9964 19256
rect 10004 19216 10005 19256
rect 9963 19207 10005 19216
rect 10390 19256 10432 19265
rect 10390 19216 10391 19256
rect 10431 19216 10432 19256
rect 10390 19207 10432 19216
rect 10635 19256 10677 19265
rect 10635 19216 10636 19256
rect 10676 19216 10677 19256
rect 10635 19207 10677 19216
rect 11019 19256 11061 19265
rect 11019 19216 11020 19256
rect 11060 19216 11061 19256
rect 11019 19207 11061 19216
rect 11248 19256 11306 19257
rect 11248 19216 11257 19256
rect 11297 19216 11306 19256
rect 11248 19215 11306 19216
rect 11499 19256 11541 19265
rect 11499 19216 11500 19256
rect 11540 19216 11541 19256
rect 11499 19207 11541 19216
rect 11618 19256 11660 19265
rect 11618 19216 11619 19256
rect 11659 19216 11660 19256
rect 11618 19207 11660 19216
rect 11728 19256 11786 19257
rect 11728 19216 11737 19256
rect 11777 19216 11786 19256
rect 11728 19215 11786 19216
rect 11883 19256 11925 19265
rect 11883 19216 11884 19256
rect 11924 19216 11925 19256
rect 11883 19207 11925 19216
rect 12075 19256 12117 19265
rect 12075 19216 12076 19256
rect 12116 19216 12117 19256
rect 12075 19207 12117 19216
rect 12267 19256 12309 19265
rect 12267 19216 12268 19256
rect 12308 19216 12309 19256
rect 12267 19207 12309 19216
rect 12459 19256 12501 19265
rect 12459 19216 12460 19256
rect 12500 19216 12501 19256
rect 12459 19207 12501 19216
rect 13131 19256 13173 19265
rect 13131 19216 13132 19256
rect 13172 19216 13173 19256
rect 13131 19207 13173 19216
rect 13323 19256 13365 19265
rect 13323 19216 13324 19256
rect 13364 19216 13365 19256
rect 13323 19207 13365 19216
rect 13803 19256 13845 19265
rect 13803 19216 13804 19256
rect 13844 19216 13845 19256
rect 13803 19207 13845 19216
rect 14410 19256 14468 19257
rect 14410 19216 14419 19256
rect 14459 19216 14468 19256
rect 14410 19215 14468 19216
rect 14605 19256 14663 19257
rect 15051 19256 15093 19265
rect 14605 19216 14614 19256
rect 14654 19216 14663 19256
rect 14605 19215 14663 19216
rect 14754 19247 14800 19256
rect 14754 19207 14755 19247
rect 14795 19207 14800 19247
rect 15051 19216 15052 19256
rect 15092 19216 15093 19256
rect 15051 19207 15093 19216
rect 15435 19256 15477 19265
rect 15435 19216 15436 19256
rect 15476 19216 15477 19256
rect 15435 19207 15477 19216
rect 16011 19256 16053 19265
rect 16011 19216 16012 19256
rect 16052 19216 16053 19256
rect 16011 19207 16053 19216
rect 16186 19256 16244 19257
rect 16186 19216 16195 19256
rect 16235 19216 16244 19256
rect 16186 19215 16244 19216
rect 16963 19256 17021 19257
rect 16963 19216 16972 19256
rect 17012 19216 17021 19256
rect 16963 19215 17021 19216
rect 17259 19256 17301 19265
rect 17259 19216 17260 19256
rect 17300 19216 17301 19256
rect 17259 19207 17301 19216
rect 17378 19256 17420 19265
rect 17378 19216 17379 19256
rect 17419 19216 17420 19256
rect 17378 19207 17420 19216
rect 17488 19256 17546 19257
rect 17488 19216 17497 19256
rect 17537 19216 17546 19256
rect 17488 19215 17546 19216
rect 17929 19256 17987 19257
rect 17929 19216 17938 19256
rect 17978 19216 17987 19256
rect 17929 19215 17987 19216
rect 19162 19256 19220 19257
rect 19162 19216 19171 19256
rect 19211 19216 19220 19256
rect 19162 19215 19220 19216
rect 19478 19256 19520 19265
rect 19478 19216 19479 19256
rect 19519 19216 19520 19256
rect 19478 19207 19520 19216
rect 19798 19256 19840 19265
rect 19798 19216 19799 19256
rect 19839 19216 19840 19256
rect 19798 19207 19840 19216
rect 20043 19256 20085 19265
rect 20043 19216 20044 19256
rect 20084 19216 20085 19256
rect 20043 19207 20085 19216
rect 20278 19256 20320 19265
rect 20278 19216 20279 19256
rect 20319 19216 20320 19256
rect 20278 19207 20320 19216
rect 20523 19256 20565 19265
rect 20523 19216 20524 19256
rect 20564 19216 20565 19256
rect 20523 19207 20565 19216
rect 20986 19256 21044 19257
rect 20986 19216 20995 19256
rect 21035 19216 21044 19256
rect 20986 19215 21044 19216
rect 21514 19256 21572 19257
rect 21514 19216 21523 19256
rect 21563 19216 21572 19256
rect 21514 19215 21572 19216
rect 22714 19256 22772 19257
rect 22714 19216 22723 19256
rect 22763 19216 22772 19256
rect 22714 19215 22772 19216
rect 22827 19256 22869 19265
rect 22827 19216 22828 19256
rect 22868 19216 22869 19256
rect 22827 19207 22869 19216
rect 23681 19256 23739 19257
rect 23681 19216 23690 19256
rect 23730 19216 23739 19256
rect 23681 19215 23739 19216
rect 24154 19256 24212 19257
rect 24154 19216 24163 19256
rect 24203 19216 24212 19256
rect 24271 19249 24272 19289
rect 24312 19249 24313 19289
rect 24271 19240 24313 19249
rect 25210 19256 25268 19257
rect 24154 19215 24212 19216
rect 25210 19216 25219 19256
rect 25259 19216 25268 19256
rect 25210 19215 25268 19216
rect 25882 19256 25940 19257
rect 25882 19216 25891 19256
rect 25931 19216 25940 19256
rect 25882 19215 25940 19216
rect 25995 19256 26037 19265
rect 25995 19216 25996 19256
rect 26036 19216 26037 19256
rect 25995 19207 26037 19216
rect 26475 19256 26517 19265
rect 26475 19216 26476 19256
rect 26516 19216 26517 19256
rect 26475 19207 26517 19216
rect 28107 19256 28149 19265
rect 28107 19216 28108 19256
rect 28148 19216 28149 19256
rect 28107 19207 28149 19216
rect 28282 19256 28340 19257
rect 28282 19216 28291 19256
rect 28331 19216 28340 19256
rect 28282 19215 28340 19216
rect 30874 19256 30932 19257
rect 30874 19216 30883 19256
rect 30923 19216 30932 19256
rect 30874 19215 30932 19216
rect 14754 19198 14800 19207
rect 1611 19172 1653 19181
rect 1611 19132 1612 19172
rect 1652 19132 1653 19172
rect 1611 19123 1653 19132
rect 2554 19172 2612 19173
rect 2554 19132 2563 19172
rect 2603 19132 2612 19172
rect 2554 19131 2612 19132
rect 6010 19172 6068 19173
rect 6010 19132 6019 19172
rect 6059 19132 6068 19172
rect 6010 19131 6068 19132
rect 8715 19172 8757 19181
rect 8715 19132 8716 19172
rect 8756 19132 8757 19172
rect 8715 19123 8757 19132
rect 11403 19172 11445 19181
rect 11403 19132 11404 19172
rect 11444 19132 11445 19172
rect 11403 19123 11445 19132
rect 13594 19172 13652 19173
rect 13594 19132 13603 19172
rect 13643 19132 13652 19172
rect 13594 19131 13652 19132
rect 16107 19172 16149 19181
rect 16107 19132 16108 19172
rect 16148 19132 16149 19172
rect 16107 19123 16149 19132
rect 16669 19172 16711 19181
rect 16669 19132 16670 19172
rect 16710 19132 16711 19172
rect 16669 19123 16711 19132
rect 17629 19172 17671 19181
rect 17629 19132 17630 19172
rect 17670 19132 17671 19172
rect 17629 19123 17671 19132
rect 27147 19172 27189 19181
rect 27147 19132 27148 19172
rect 27188 19132 27189 19172
rect 27147 19123 27189 19132
rect 28598 19172 28640 19181
rect 28598 19132 28599 19172
rect 28639 19132 28640 19172
rect 28598 19123 28640 19132
rect 1978 19088 2036 19089
rect 1978 19048 1987 19088
rect 2027 19048 2036 19088
rect 1978 19047 2036 19048
rect 2091 19088 2133 19097
rect 2091 19048 2092 19088
rect 2132 19048 2133 19088
rect 2091 19039 2133 19048
rect 2667 19088 2709 19097
rect 2667 19048 2668 19088
rect 2708 19048 2709 19088
rect 2667 19039 2709 19048
rect 2955 19088 2997 19097
rect 2955 19048 2956 19088
rect 2996 19048 2997 19088
rect 2955 19039 2997 19048
rect 3531 19088 3573 19097
rect 3531 19048 3532 19088
rect 3572 19048 3573 19088
rect 3531 19039 3573 19048
rect 6970 19088 7028 19089
rect 6970 19048 6979 19088
rect 7019 19048 7028 19088
rect 6970 19047 7028 19048
rect 9435 19088 9477 19097
rect 9435 19048 9436 19088
rect 9476 19048 9477 19088
rect 9435 19039 9477 19048
rect 10042 19088 10100 19089
rect 10042 19048 10051 19088
rect 10091 19048 10100 19088
rect 10042 19047 10100 19048
rect 10714 19088 10772 19089
rect 10714 19048 10723 19088
rect 10763 19048 10772 19088
rect 10714 19047 10772 19048
rect 12363 19088 12405 19097
rect 12363 19048 12364 19088
rect 12404 19048 12405 19088
rect 12363 19039 12405 19048
rect 13882 19088 13940 19089
rect 13882 19048 13891 19088
rect 13931 19048 13940 19088
rect 13882 19047 13940 19048
rect 15322 19088 15380 19089
rect 15322 19048 15331 19088
rect 15371 19048 15380 19088
rect 15322 19047 15380 19048
rect 15610 19088 15668 19089
rect 15610 19048 15619 19088
rect 15659 19048 15668 19088
rect 15610 19047 15668 19048
rect 16875 19088 16917 19097
rect 16875 19048 16876 19088
rect 16916 19048 16917 19088
rect 16875 19039 16917 19048
rect 17163 19088 17205 19097
rect 17163 19048 17164 19088
rect 17204 19048 17205 19088
rect 17163 19039 17205 19048
rect 17835 19088 17877 19097
rect 17835 19048 17836 19088
rect 17876 19048 17877 19088
rect 17835 19039 17877 19048
rect 19258 19088 19316 19089
rect 19258 19048 19267 19088
rect 19307 19048 19316 19088
rect 19258 19047 19316 19048
rect 20122 19088 20180 19089
rect 20122 19048 20131 19088
rect 20171 19048 20180 19088
rect 20122 19047 20180 19048
rect 21723 19088 21765 19097
rect 21723 19048 21724 19088
rect 21764 19048 21765 19088
rect 21723 19039 21765 19048
rect 23115 19088 23157 19097
rect 23115 19048 23116 19088
rect 23156 19048 23157 19088
rect 23115 19039 23157 19048
rect 23386 19088 23444 19089
rect 24730 19088 24788 19089
rect 23386 19048 23395 19088
rect 23435 19048 23444 19088
rect 23386 19047 23444 19048
rect 24066 19079 24112 19088
rect 24066 19039 24067 19079
rect 24107 19039 24112 19079
rect 24730 19048 24739 19088
rect 24779 19048 24788 19088
rect 24730 19047 24788 19048
rect 27435 19088 27477 19097
rect 27435 19048 27436 19088
rect 27476 19048 27477 19088
rect 27435 19039 27477 19048
rect 28378 19088 28436 19089
rect 28378 19048 28387 19088
rect 28427 19048 28436 19088
rect 28378 19047 28436 19048
rect 28491 19088 28533 19097
rect 28491 19048 28492 19088
rect 28532 19048 28533 19088
rect 28491 19039 28533 19048
rect 28971 19088 29013 19097
rect 28971 19048 28972 19088
rect 29012 19048 29013 19088
rect 28971 19039 29013 19048
rect 24066 19030 24112 19039
rect 576 18920 31392 18944
rect 576 18880 4352 18920
rect 4720 18880 12126 18920
rect 12494 18880 19900 18920
rect 20268 18880 27674 18920
rect 28042 18880 31392 18920
rect 576 18856 31392 18880
rect 1402 18752 1460 18753
rect 1402 18712 1411 18752
rect 1451 18712 1460 18752
rect 1402 18711 1460 18712
rect 1882 18752 1940 18753
rect 1882 18712 1891 18752
rect 1931 18712 1940 18752
rect 1882 18711 1940 18712
rect 3051 18752 3093 18761
rect 3051 18712 3052 18752
rect 3092 18712 3093 18752
rect 3051 18703 3093 18712
rect 4203 18752 4245 18761
rect 4203 18712 4204 18752
rect 4244 18712 4245 18752
rect 4203 18703 4245 18712
rect 5242 18752 5300 18753
rect 5242 18712 5251 18752
rect 5291 18712 5300 18752
rect 5242 18711 5300 18712
rect 6411 18752 6453 18761
rect 6411 18712 6412 18752
rect 6452 18712 6453 18752
rect 6411 18703 6453 18712
rect 7275 18752 7317 18761
rect 7275 18712 7276 18752
rect 7316 18712 7317 18752
rect 7275 18703 7317 18712
rect 8890 18752 8948 18753
rect 8890 18712 8899 18752
rect 8939 18712 8948 18752
rect 8890 18711 8948 18712
rect 9243 18752 9285 18761
rect 9243 18712 9244 18752
rect 9284 18712 9285 18752
rect 9243 18703 9285 18712
rect 11019 18752 11061 18761
rect 11019 18712 11020 18752
rect 11060 18712 11061 18752
rect 11019 18703 11061 18712
rect 11307 18752 11349 18761
rect 11307 18712 11308 18752
rect 11348 18712 11349 18752
rect 11307 18703 11349 18712
rect 13882 18752 13940 18753
rect 13882 18712 13891 18752
rect 13931 18712 13940 18752
rect 13882 18711 13940 18712
rect 16683 18752 16725 18761
rect 16683 18712 16684 18752
rect 16724 18712 16725 18752
rect 16683 18703 16725 18712
rect 17914 18752 17972 18753
rect 17914 18712 17923 18752
rect 17963 18712 17972 18752
rect 17914 18711 17972 18712
rect 18394 18752 18452 18753
rect 18394 18712 18403 18752
rect 18443 18712 18452 18752
rect 18394 18711 18452 18712
rect 19354 18752 19412 18753
rect 19354 18712 19363 18752
rect 19403 18712 19412 18752
rect 19354 18711 19412 18712
rect 22923 18752 22965 18761
rect 22923 18712 22924 18752
rect 22964 18712 22965 18752
rect 22923 18703 22965 18712
rect 27754 18752 27812 18753
rect 27754 18712 27763 18752
rect 27803 18712 27812 18752
rect 27754 18711 27812 18712
rect 28971 18752 29013 18761
rect 28971 18712 28972 18752
rect 29012 18712 29013 18752
rect 28971 18703 29013 18712
rect 2091 18668 2133 18677
rect 2091 18628 2092 18668
rect 2132 18628 2133 18668
rect 2091 18619 2133 18628
rect 2557 18668 2599 18677
rect 2557 18628 2558 18668
rect 2598 18628 2599 18668
rect 2557 18619 2599 18628
rect 2650 18668 2708 18669
rect 2650 18628 2659 18668
rect 2699 18628 2708 18668
rect 2650 18627 2708 18628
rect 3997 18668 4039 18677
rect 3997 18628 3998 18668
rect 4038 18628 4039 18668
rect 3997 18619 4039 18628
rect 7659 18668 7701 18677
rect 7659 18628 7660 18668
rect 7700 18628 7701 18668
rect 7659 18619 7701 18628
rect 8170 18668 8228 18669
rect 8170 18628 8179 18668
rect 8219 18628 8228 18668
rect 8170 18627 8228 18628
rect 8797 18668 8839 18677
rect 8797 18628 8798 18668
rect 8838 18628 8839 18668
rect 8797 18619 8839 18628
rect 9003 18668 9045 18677
rect 9003 18628 9004 18668
rect 9044 18628 9045 18668
rect 9003 18619 9045 18628
rect 13594 18668 13652 18669
rect 13594 18628 13603 18668
rect 13643 18628 13652 18668
rect 13594 18627 13652 18628
rect 16971 18668 17013 18677
rect 16971 18628 16972 18668
rect 17012 18628 17013 18668
rect 16971 18619 17013 18628
rect 18507 18668 18549 18677
rect 18507 18628 18508 18668
rect 18548 18628 18549 18668
rect 18507 18619 18549 18628
rect 19755 18668 19797 18677
rect 19755 18628 19756 18668
rect 19796 18628 19797 18668
rect 19755 18619 19797 18628
rect 20314 18668 20372 18669
rect 20314 18628 20323 18668
rect 20363 18628 20372 18668
rect 20314 18627 20372 18628
rect 21387 18668 21429 18677
rect 21387 18628 21388 18668
rect 21428 18628 21429 18668
rect 21387 18619 21429 18628
rect 24442 18668 24500 18669
rect 24442 18628 24451 18668
rect 24491 18628 24500 18668
rect 24442 18627 24500 18628
rect 27322 18668 27380 18669
rect 27322 18628 27331 18668
rect 27371 18628 27380 18668
rect 27322 18627 27380 18628
rect 1078 18584 1120 18593
rect 1078 18544 1079 18584
rect 1119 18544 1120 18584
rect 1078 18535 1120 18544
rect 1323 18584 1365 18593
rect 1323 18544 1324 18584
rect 1364 18544 1365 18584
rect 1803 18584 1845 18593
rect 1323 18535 1365 18544
rect 1563 18542 1605 18551
rect 1563 18502 1564 18542
rect 1604 18502 1605 18542
rect 1803 18544 1804 18584
rect 1844 18544 1845 18584
rect 1803 18535 1845 18544
rect 2187 18584 2229 18593
rect 2187 18544 2188 18584
rect 2228 18544 2229 18584
rect 2187 18535 2229 18544
rect 2416 18584 2474 18585
rect 2416 18544 2425 18584
rect 2465 18544 2474 18584
rect 2416 18543 2474 18544
rect 2763 18584 2805 18593
rect 3147 18584 3189 18593
rect 2763 18544 2764 18584
rect 2804 18544 2805 18584
rect 2763 18535 2805 18544
rect 2859 18575 2901 18584
rect 2859 18535 2860 18575
rect 2900 18535 2901 18575
rect 3147 18544 3148 18584
rect 3188 18544 3189 18584
rect 3147 18535 3189 18544
rect 3266 18584 3308 18593
rect 4930 18584 4988 18585
rect 3266 18544 3267 18584
rect 3307 18544 3308 18584
rect 4299 18575 4341 18584
rect 3266 18535 3308 18544
rect 3387 18542 3429 18551
rect 2859 18526 2901 18535
rect 1210 18500 1268 18501
rect 1210 18460 1219 18500
rect 1259 18460 1268 18500
rect 1563 18493 1605 18502
rect 1690 18500 1748 18501
rect 1210 18459 1268 18460
rect 1690 18460 1699 18500
rect 1739 18460 1748 18500
rect 1690 18459 1748 18460
rect 2091 18500 2133 18509
rect 2091 18460 2092 18500
rect 2132 18460 2133 18500
rect 2091 18451 2133 18460
rect 2306 18500 2348 18509
rect 2306 18460 2307 18500
rect 2347 18460 2348 18500
rect 3387 18502 3388 18542
rect 3428 18502 3429 18542
rect 4299 18535 4300 18575
rect 4340 18535 4341 18575
rect 4930 18544 4939 18584
rect 4979 18544 4988 18584
rect 4930 18543 4988 18544
rect 5163 18584 5205 18593
rect 5163 18544 5164 18584
rect 5204 18544 5205 18584
rect 4299 18526 4341 18535
rect 4810 18542 4868 18543
rect 3387 18493 3429 18502
rect 3819 18500 3861 18509
rect 4810 18502 4819 18542
rect 4859 18502 4868 18542
rect 5163 18535 5205 18544
rect 5547 18584 5589 18593
rect 5547 18544 5548 18584
rect 5588 18544 5589 18584
rect 5547 18535 5589 18544
rect 5764 18584 5806 18593
rect 5764 18544 5765 18584
rect 5805 18544 5806 18584
rect 5764 18535 5806 18544
rect 5920 18584 5962 18593
rect 5920 18544 5921 18584
rect 5961 18544 5962 18584
rect 5920 18535 5962 18544
rect 6123 18584 6165 18593
rect 6507 18584 6549 18593
rect 6123 18544 6124 18584
rect 6164 18544 6165 18584
rect 6123 18535 6165 18544
rect 6219 18575 6261 18584
rect 6219 18535 6220 18575
rect 6260 18535 6261 18575
rect 6507 18544 6508 18584
rect 6548 18544 6549 18584
rect 6507 18535 6549 18544
rect 6736 18584 6794 18585
rect 6736 18544 6745 18584
rect 6785 18544 6794 18584
rect 6736 18543 6794 18544
rect 7179 18584 7221 18593
rect 7179 18544 7180 18584
rect 7220 18544 7221 18584
rect 7179 18535 7221 18544
rect 7370 18584 7412 18593
rect 7370 18544 7371 18584
rect 7411 18544 7412 18584
rect 7370 18535 7412 18544
rect 7546 18584 7604 18585
rect 7546 18544 7555 18584
rect 7595 18544 7604 18584
rect 7546 18543 7604 18544
rect 7862 18584 7904 18593
rect 7862 18544 7863 18584
rect 7903 18544 7904 18584
rect 7862 18535 7904 18544
rect 8365 18584 8423 18585
rect 8365 18544 8374 18584
rect 8414 18544 8423 18584
rect 8365 18543 8423 18544
rect 8523 18584 8565 18593
rect 10731 18584 10773 18593
rect 8523 18544 8524 18584
rect 8564 18544 8565 18584
rect 8523 18535 8565 18544
rect 9099 18575 9141 18584
rect 9099 18535 9100 18575
rect 9140 18535 9141 18575
rect 10731 18544 10732 18584
rect 10772 18544 10773 18584
rect 10731 18535 10773 18544
rect 10865 18584 10923 18585
rect 10865 18544 10874 18584
rect 10914 18544 10923 18584
rect 10865 18543 10923 18544
rect 11211 18584 11253 18593
rect 11211 18544 11212 18584
rect 11252 18544 11253 18584
rect 11211 18535 11253 18544
rect 11386 18584 11444 18585
rect 11386 18544 11395 18584
rect 11435 18544 11444 18584
rect 11386 18543 11444 18544
rect 12685 18584 12743 18585
rect 12685 18544 12694 18584
rect 12734 18544 12743 18584
rect 12685 18543 12743 18544
rect 13323 18584 13365 18593
rect 13323 18544 13324 18584
rect 13364 18544 13365 18584
rect 13323 18535 13365 18544
rect 13803 18584 13845 18593
rect 13803 18544 13804 18584
rect 13844 18544 13845 18584
rect 13803 18535 13845 18544
rect 14667 18584 14709 18593
rect 14667 18544 14668 18584
rect 14708 18544 14709 18584
rect 14667 18535 14709 18544
rect 14859 18584 14901 18593
rect 14859 18544 14860 18584
rect 14900 18544 14901 18584
rect 14859 18535 14901 18544
rect 16203 18584 16245 18593
rect 16203 18544 16204 18584
rect 16244 18544 16245 18584
rect 16203 18535 16245 18544
rect 16372 18584 16414 18593
rect 16372 18544 16373 18584
rect 16413 18544 16414 18584
rect 16372 18535 16414 18544
rect 16491 18584 16533 18593
rect 16491 18544 16492 18584
rect 16532 18544 16533 18584
rect 16491 18535 16533 18544
rect 16858 18584 16916 18585
rect 16858 18544 16867 18584
rect 16907 18544 16916 18584
rect 16858 18543 16916 18544
rect 17174 18584 17216 18593
rect 17174 18544 17175 18584
rect 17215 18544 17216 18584
rect 17174 18535 17216 18544
rect 17290 18584 17348 18585
rect 17290 18544 17299 18584
rect 17339 18544 17348 18584
rect 17290 18543 17348 18544
rect 17818 18584 17876 18585
rect 17818 18544 17827 18584
rect 17867 18544 17876 18584
rect 17818 18543 17876 18544
rect 18134 18584 18176 18593
rect 18134 18544 18135 18584
rect 18175 18544 18176 18584
rect 18134 18535 18176 18544
rect 18301 18584 18343 18593
rect 19030 18584 19072 18593
rect 18301 18544 18302 18584
rect 18342 18544 18343 18584
rect 18301 18535 18343 18544
rect 18603 18575 18645 18584
rect 18603 18535 18604 18575
rect 18644 18535 18645 18575
rect 19030 18544 19031 18584
rect 19071 18544 19072 18584
rect 19030 18535 19072 18544
rect 19273 18584 19315 18593
rect 19273 18544 19274 18584
rect 19314 18544 19315 18584
rect 19273 18535 19315 18544
rect 19546 18584 19604 18585
rect 19546 18544 19555 18584
rect 19595 18544 19604 18584
rect 19546 18543 19604 18544
rect 19659 18584 19701 18593
rect 19659 18544 19660 18584
rect 19700 18544 19701 18584
rect 19659 18535 19701 18544
rect 19862 18584 19904 18593
rect 19862 18544 19863 18584
rect 19903 18544 19904 18584
rect 19862 18535 19904 18544
rect 19995 18584 20037 18593
rect 19995 18544 19996 18584
rect 20036 18544 20037 18584
rect 19995 18535 20037 18544
rect 20122 18584 20180 18585
rect 20122 18544 20131 18584
rect 20171 18544 20180 18584
rect 20122 18543 20180 18544
rect 20235 18584 20277 18593
rect 20235 18544 20236 18584
rect 20276 18544 20277 18584
rect 20235 18535 20277 18544
rect 21082 18584 21140 18585
rect 21082 18544 21091 18584
rect 21131 18544 21140 18584
rect 21082 18543 21140 18544
rect 22906 18584 22964 18585
rect 22906 18544 22915 18584
rect 22955 18544 22964 18584
rect 22906 18543 22964 18544
rect 23019 18584 23061 18593
rect 23019 18544 23020 18584
rect 23060 18544 23061 18584
rect 23019 18535 23061 18544
rect 24363 18584 24405 18593
rect 24363 18544 24364 18584
rect 24404 18544 24405 18584
rect 24363 18535 24405 18544
rect 24555 18584 24597 18593
rect 24555 18544 24556 18584
rect 24596 18544 24597 18584
rect 24555 18535 24597 18544
rect 26938 18584 26996 18585
rect 26938 18544 26947 18584
rect 26987 18544 26996 18584
rect 26938 18543 26996 18544
rect 27946 18584 28004 18585
rect 27946 18544 27955 18584
rect 27995 18544 28004 18584
rect 27946 18543 28004 18544
rect 28066 18584 28124 18585
rect 28066 18544 28075 18584
rect 28115 18544 28124 18584
rect 28522 18584 28580 18585
rect 28066 18543 28124 18544
rect 28367 18542 28409 18551
rect 28522 18544 28531 18584
rect 28571 18544 28580 18584
rect 28522 18543 28580 18544
rect 28779 18584 28821 18593
rect 28779 18544 28780 18584
rect 28820 18544 28821 18584
rect 6219 18526 6261 18535
rect 9099 18526 9141 18535
rect 18603 18526 18645 18535
rect 4810 18501 4868 18502
rect 2306 18451 2348 18460
rect 3819 18460 3820 18500
rect 3860 18460 3861 18500
rect 3819 18451 3861 18460
rect 4618 18500 4676 18501
rect 4618 18460 4627 18500
rect 4667 18460 4676 18500
rect 4618 18459 4676 18460
rect 5050 18500 5108 18501
rect 5050 18460 5059 18500
rect 5099 18460 5108 18500
rect 5050 18459 5108 18460
rect 5451 18500 5493 18509
rect 6626 18500 6668 18509
rect 5451 18460 5452 18500
rect 5492 18460 5493 18500
rect 5451 18451 5493 18460
rect 5682 18491 5728 18500
rect 5682 18451 5683 18491
rect 5723 18451 5728 18491
rect 6626 18460 6627 18500
rect 6667 18460 6668 18500
rect 6626 18451 6668 18460
rect 9483 18500 9525 18509
rect 9483 18460 9484 18500
rect 9524 18460 9525 18500
rect 9483 18451 9525 18460
rect 12490 18500 12548 18501
rect 12490 18460 12499 18500
rect 12539 18460 12548 18500
rect 12490 18459 12548 18460
rect 17499 18500 17541 18509
rect 17499 18460 17500 18500
rect 17540 18460 17541 18500
rect 17499 18451 17541 18460
rect 19162 18500 19220 18501
rect 19162 18460 19171 18500
rect 19211 18460 19220 18500
rect 19162 18459 19220 18460
rect 20907 18500 20949 18509
rect 20907 18460 20908 18500
rect 20948 18460 20949 18500
rect 20907 18451 20949 18460
rect 21483 18500 21525 18509
rect 21483 18460 21484 18500
rect 21524 18460 21525 18500
rect 21483 18451 21525 18460
rect 21867 18500 21909 18509
rect 21867 18460 21868 18500
rect 21908 18460 21909 18500
rect 21867 18451 21909 18460
rect 28203 18500 28245 18509
rect 28203 18460 28204 18500
rect 28244 18460 28245 18500
rect 28367 18502 28368 18542
rect 28408 18502 28409 18542
rect 28779 18535 28821 18544
rect 30874 18584 30932 18585
rect 30874 18544 30883 18584
rect 30923 18544 30932 18584
rect 30874 18543 30932 18544
rect 28367 18493 28409 18502
rect 28635 18500 28677 18509
rect 28203 18451 28245 18460
rect 28635 18460 28636 18500
rect 28676 18460 28677 18500
rect 28635 18451 28677 18460
rect 31258 18500 31316 18501
rect 31258 18460 31267 18500
rect 31307 18460 31316 18500
rect 31258 18459 31316 18460
rect 5682 18442 5728 18451
rect 23211 18416 23253 18425
rect 23211 18376 23212 18416
rect 23252 18376 23253 18416
rect 23211 18367 23253 18376
rect 25419 18416 25461 18425
rect 25419 18376 25420 18416
rect 25460 18376 25461 18416
rect 25419 18367 25461 18376
rect 28299 18416 28341 18425
rect 28299 18376 28300 18416
rect 28340 18376 28341 18416
rect 28299 18367 28341 18376
rect 3579 18332 3621 18341
rect 3579 18292 3580 18332
rect 3620 18292 3621 18332
rect 3579 18283 3621 18292
rect 3994 18332 4052 18333
rect 3994 18292 4003 18332
rect 4043 18292 4052 18332
rect 3994 18291 4052 18292
rect 5914 18332 5972 18333
rect 5914 18292 5923 18332
rect 5963 18292 5972 18332
rect 5914 18291 5972 18292
rect 7851 18332 7893 18341
rect 7851 18292 7852 18332
rect 7892 18292 7893 18332
rect 7851 18283 7893 18292
rect 13131 18332 13173 18341
rect 13131 18292 13132 18332
rect 13172 18292 13173 18332
rect 13131 18283 13173 18292
rect 14763 18332 14805 18341
rect 14763 18292 14764 18332
rect 14804 18292 14805 18332
rect 14763 18283 14805 18292
rect 17163 18332 17205 18341
rect 17163 18292 17164 18332
rect 17204 18292 17205 18332
rect 17163 18283 17205 18292
rect 18123 18332 18165 18341
rect 18123 18292 18124 18332
rect 18164 18292 18165 18332
rect 18123 18283 18165 18292
rect 21627 18332 21669 18341
rect 21627 18292 21628 18332
rect 21668 18292 21669 18332
rect 21627 18283 21669 18292
rect 25035 18332 25077 18341
rect 25035 18292 25036 18332
rect 25076 18292 25077 18332
rect 25035 18283 25077 18292
rect 576 18164 31392 18188
rect 576 18124 3112 18164
rect 3480 18124 10886 18164
rect 11254 18124 18660 18164
rect 19028 18124 26434 18164
rect 26802 18124 31392 18164
rect 576 18100 31392 18124
rect 1402 17996 1460 17997
rect 1402 17956 1411 17996
rect 1451 17956 1460 17996
rect 1402 17955 1460 17956
rect 2170 17996 2228 17997
rect 2170 17956 2179 17996
rect 2219 17956 2228 17996
rect 2170 17955 2228 17956
rect 5739 17996 5781 18005
rect 5739 17956 5740 17996
rect 5780 17956 5781 17996
rect 5739 17947 5781 17956
rect 7546 17996 7604 17997
rect 7546 17956 7555 17996
rect 7595 17956 7604 17996
rect 7546 17955 7604 17956
rect 8859 17996 8901 18005
rect 8859 17956 8860 17996
rect 8900 17956 8901 17996
rect 8859 17947 8901 17956
rect 16299 17996 16341 18005
rect 16299 17956 16300 17996
rect 16340 17956 16341 17996
rect 16299 17947 16341 17956
rect 18219 17996 18261 18005
rect 18219 17956 18220 17996
rect 18260 17956 18261 17996
rect 18219 17947 18261 17956
rect 19755 17996 19797 18005
rect 19755 17956 19756 17996
rect 19796 17956 19797 17996
rect 19755 17947 19797 17956
rect 22635 17996 22677 18005
rect 22635 17956 22636 17996
rect 22676 17956 22677 17996
rect 22635 17947 22677 17956
rect 27723 17996 27765 18005
rect 27723 17956 27724 17996
rect 27764 17956 27765 17996
rect 27723 17947 27765 17956
rect 30699 17996 30741 18005
rect 30699 17956 30700 17996
rect 30740 17956 30741 17996
rect 30699 17947 30741 17956
rect 29835 17912 29877 17921
rect 29835 17872 29836 17912
rect 29876 17872 29877 17912
rect 29835 17863 29877 17872
rect 30891 17912 30933 17921
rect 30891 17872 30892 17912
rect 30932 17872 30933 17912
rect 30891 17863 30933 17872
rect 2986 17828 3044 17829
rect 2986 17788 2995 17828
rect 3035 17788 3044 17828
rect 2986 17787 3044 17788
rect 4107 17828 4149 17837
rect 9771 17828 9813 17837
rect 4107 17788 4108 17828
rect 4148 17788 4149 17828
rect 4107 17779 4149 17788
rect 4530 17819 4576 17828
rect 4530 17779 4531 17819
rect 4571 17779 4576 17819
rect 9771 17788 9772 17828
rect 9812 17788 9813 17828
rect 9771 17779 9813 17788
rect 10827 17828 10869 17837
rect 10827 17788 10828 17828
rect 10868 17788 10869 17828
rect 10827 17779 10869 17788
rect 11722 17828 11780 17829
rect 11722 17788 11731 17828
rect 11771 17788 11780 17828
rect 11722 17787 11780 17788
rect 4530 17770 4576 17779
rect 1699 17744 1757 17745
rect 1699 17704 1708 17744
rect 1748 17704 1757 17744
rect 1699 17703 1757 17704
rect 2176 17744 2218 17753
rect 2176 17704 2177 17744
rect 2217 17704 2218 17744
rect 2176 17695 2218 17704
rect 2467 17744 2525 17745
rect 2467 17704 2476 17744
rect 2516 17704 2525 17744
rect 2467 17703 2525 17704
rect 3181 17744 3239 17745
rect 3181 17704 3190 17744
rect 3230 17704 3239 17744
rect 3181 17703 3239 17704
rect 3619 17744 3677 17745
rect 3619 17704 3628 17744
rect 3668 17704 3677 17744
rect 3619 17703 3677 17704
rect 3771 17744 3813 17753
rect 3771 17704 3772 17744
rect 3812 17704 3813 17744
rect 3771 17695 3813 17704
rect 3898 17744 3956 17745
rect 3898 17704 3907 17744
rect 3947 17704 3956 17744
rect 3898 17703 3956 17704
rect 4011 17744 4053 17753
rect 4011 17704 4012 17744
rect 4052 17704 4053 17744
rect 4011 17695 4053 17704
rect 4395 17744 4437 17753
rect 4395 17704 4396 17744
rect 4436 17704 4437 17744
rect 4395 17695 4437 17704
rect 4624 17744 4682 17745
rect 4624 17704 4633 17744
rect 4673 17704 4682 17744
rect 4624 17703 4682 17704
rect 4875 17744 4917 17753
rect 4875 17704 4876 17744
rect 4916 17704 4917 17744
rect 4875 17695 4917 17704
rect 4994 17744 5036 17753
rect 4994 17704 4995 17744
rect 5035 17704 5036 17744
rect 4994 17695 5036 17704
rect 5104 17744 5162 17745
rect 5104 17704 5113 17744
rect 5153 17704 5162 17744
rect 5104 17703 5162 17704
rect 5739 17744 5781 17753
rect 5739 17704 5740 17744
rect 5780 17704 5781 17744
rect 5739 17695 5781 17704
rect 5931 17744 5973 17753
rect 5931 17704 5932 17744
rect 5972 17704 5973 17744
rect 5931 17695 5973 17704
rect 6603 17744 6645 17753
rect 6603 17704 6604 17744
rect 6644 17704 6645 17744
rect 6603 17695 6645 17704
rect 6794 17744 6836 17753
rect 6794 17704 6795 17744
rect 6835 17704 6836 17744
rect 6794 17695 6836 17704
rect 6987 17744 7029 17753
rect 6987 17704 6988 17744
rect 7028 17704 7029 17744
rect 6987 17695 7029 17704
rect 7162 17744 7220 17745
rect 7162 17704 7171 17744
rect 7211 17704 7220 17744
rect 7162 17703 7220 17704
rect 7371 17744 7413 17753
rect 7371 17704 7372 17744
rect 7412 17704 7413 17744
rect 7371 17695 7413 17704
rect 7546 17744 7604 17745
rect 7546 17704 7555 17744
rect 7595 17704 7604 17744
rect 7546 17703 7604 17704
rect 8074 17744 8132 17745
rect 8074 17704 8083 17744
rect 8123 17704 8132 17744
rect 8074 17703 8132 17704
rect 8269 17744 8327 17745
rect 8269 17704 8278 17744
rect 8318 17704 8327 17744
rect 8269 17703 8327 17704
rect 9003 17744 9045 17753
rect 9003 17704 9004 17744
rect 9044 17704 9045 17744
rect 9003 17695 9045 17704
rect 9291 17744 9333 17753
rect 9291 17704 9292 17744
rect 9332 17704 9333 17744
rect 9291 17695 9333 17704
rect 9410 17744 9452 17753
rect 9410 17704 9411 17744
rect 9451 17704 9452 17744
rect 9410 17695 9452 17704
rect 9520 17744 9578 17745
rect 9520 17704 9529 17744
rect 9569 17704 9578 17744
rect 9520 17703 9578 17704
rect 9675 17744 9717 17753
rect 9675 17704 9676 17744
rect 9716 17704 9717 17744
rect 9675 17695 9717 17704
rect 9867 17744 9909 17753
rect 9867 17704 9868 17744
rect 9908 17704 9909 17744
rect 9867 17695 9909 17704
rect 10347 17744 10389 17753
rect 10347 17704 10348 17744
rect 10388 17704 10389 17744
rect 10347 17695 10389 17704
rect 10539 17744 10581 17753
rect 10539 17704 10540 17744
rect 10580 17704 10581 17744
rect 10539 17695 10581 17704
rect 10731 17744 10773 17753
rect 10731 17704 10732 17744
rect 10772 17704 10773 17744
rect 10731 17695 10773 17704
rect 10923 17744 10965 17753
rect 10923 17704 10924 17744
rect 10964 17704 10965 17744
rect 10923 17695 10965 17704
rect 11062 17744 11104 17753
rect 11062 17704 11063 17744
rect 11103 17704 11104 17744
rect 11062 17695 11104 17704
rect 11194 17744 11252 17745
rect 11194 17704 11203 17744
rect 11243 17704 11252 17744
rect 11194 17703 11252 17704
rect 11307 17744 11349 17753
rect 11307 17704 11308 17744
rect 11348 17704 11349 17744
rect 11307 17695 11349 17704
rect 11917 17744 11975 17745
rect 11917 17704 11926 17744
rect 11966 17704 11975 17744
rect 11917 17703 11975 17704
rect 13114 17744 13172 17745
rect 13114 17704 13123 17744
rect 13163 17704 13172 17744
rect 13114 17703 13172 17704
rect 13419 17744 13461 17753
rect 13419 17704 13420 17744
rect 13460 17704 13461 17744
rect 13419 17695 13461 17704
rect 14797 17744 14855 17745
rect 14797 17704 14806 17744
rect 14846 17704 14855 17744
rect 14797 17703 14855 17704
rect 15147 17744 15189 17753
rect 15147 17704 15148 17744
rect 15188 17704 15189 17744
rect 15147 17695 15189 17704
rect 15435 17744 15477 17753
rect 15435 17704 15436 17744
rect 15476 17704 15477 17744
rect 15435 17695 15477 17704
rect 15627 17744 15669 17753
rect 15627 17704 15628 17744
rect 15668 17704 15669 17744
rect 15627 17695 15669 17704
rect 15994 17744 16052 17745
rect 15994 17704 16003 17744
rect 16043 17704 16052 17744
rect 15994 17703 16052 17704
rect 16491 17744 16533 17753
rect 16491 17704 16492 17744
rect 16532 17704 16533 17744
rect 16491 17695 16533 17704
rect 16683 17744 16725 17753
rect 16683 17704 16684 17744
rect 16724 17704 16725 17744
rect 16683 17695 16725 17704
rect 17547 17744 17589 17753
rect 17547 17704 17548 17744
rect 17588 17704 17589 17744
rect 17547 17695 17589 17704
rect 17716 17744 17758 17753
rect 17716 17704 17717 17744
rect 17757 17704 17758 17744
rect 17716 17695 17758 17704
rect 17914 17744 17972 17745
rect 17914 17704 17923 17744
rect 17963 17704 17972 17744
rect 17914 17703 17972 17704
rect 18230 17744 18272 17753
rect 18230 17704 18231 17744
rect 18271 17704 18272 17744
rect 18230 17695 18272 17704
rect 19450 17744 19508 17745
rect 19450 17704 19459 17744
rect 19499 17704 19508 17744
rect 19450 17703 19508 17704
rect 19769 17744 19811 17753
rect 19769 17704 19770 17744
rect 19810 17704 19811 17744
rect 19769 17695 19811 17704
rect 22635 17744 22677 17753
rect 22635 17704 22636 17744
rect 22676 17704 22677 17744
rect 22635 17695 22677 17704
rect 22938 17744 22980 17753
rect 23403 17744 23445 17753
rect 22938 17704 22939 17744
rect 22979 17704 22980 17744
rect 22938 17695 22980 17704
rect 23106 17735 23152 17744
rect 23106 17695 23107 17735
rect 23147 17695 23152 17735
rect 23403 17704 23404 17744
rect 23444 17704 23445 17744
rect 23403 17695 23445 17704
rect 24171 17744 24213 17753
rect 24171 17704 24172 17744
rect 24212 17704 24213 17744
rect 24171 17695 24213 17704
rect 24459 17744 24501 17753
rect 24459 17704 24460 17744
rect 24500 17704 24501 17744
rect 24459 17695 24501 17704
rect 24843 17744 24885 17753
rect 24843 17704 24844 17744
rect 24884 17704 24885 17744
rect 24843 17695 24885 17704
rect 24987 17744 25029 17753
rect 24987 17704 24988 17744
rect 25028 17704 25029 17744
rect 24987 17695 25029 17704
rect 25899 17744 25941 17753
rect 25899 17704 25900 17744
rect 25940 17704 25941 17744
rect 25899 17695 25941 17704
rect 26091 17744 26133 17753
rect 26091 17704 26092 17744
rect 26132 17704 26133 17744
rect 26091 17695 26133 17704
rect 27627 17744 27669 17753
rect 27627 17704 27628 17744
rect 27668 17704 27669 17744
rect 27627 17695 27669 17704
rect 27819 17744 27861 17753
rect 27819 17704 27820 17744
rect 27860 17704 27861 17744
rect 27819 17695 27861 17704
rect 28395 17744 28437 17753
rect 28395 17704 28396 17744
rect 28436 17704 28437 17744
rect 28395 17695 28437 17704
rect 28570 17744 28628 17745
rect 28570 17704 28579 17744
rect 28619 17704 28628 17744
rect 28570 17703 28628 17704
rect 29259 17744 29301 17753
rect 29259 17704 29260 17744
rect 29300 17704 29301 17744
rect 29259 17695 29301 17704
rect 30027 17744 30069 17753
rect 30027 17704 30028 17744
rect 30068 17704 30069 17744
rect 30027 17695 30069 17704
rect 23106 17686 23152 17695
rect 1408 17660 1450 17669
rect 1408 17620 1409 17660
rect 1449 17620 1450 17660
rect 1408 17611 1450 17620
rect 3328 17660 3370 17669
rect 3328 17620 3329 17660
rect 3369 17620 3370 17660
rect 3328 17611 3370 17620
rect 4299 17660 4341 17669
rect 4299 17620 4300 17660
rect 4340 17620 4341 17660
rect 4299 17611 4341 17620
rect 6699 17660 6741 17669
rect 6699 17620 6700 17660
rect 6740 17620 6741 17660
rect 6699 17611 6741 17620
rect 9195 17660 9237 17669
rect 9195 17620 9196 17660
rect 9236 17620 9237 17660
rect 9195 17611 9237 17620
rect 11386 17660 11444 17661
rect 11386 17620 11395 17660
rect 11435 17620 11444 17660
rect 11386 17619 11444 17620
rect 12939 17660 12981 17669
rect 12939 17620 12940 17660
rect 12980 17620 12981 17660
rect 12939 17611 12981 17620
rect 15531 17660 15573 17669
rect 15531 17620 15532 17660
rect 15572 17620 15573 17660
rect 15531 17611 15573 17620
rect 16313 17660 16355 17669
rect 16313 17620 16314 17660
rect 16354 17620 16355 17660
rect 16313 17611 16355 17620
rect 16587 17660 16629 17669
rect 16587 17620 16588 17660
rect 16628 17620 16629 17660
rect 16587 17611 16629 17620
rect 23211 17660 23253 17669
rect 23211 17620 23212 17660
rect 23252 17620 23253 17660
rect 23211 17611 23253 17620
rect 24634 17660 24692 17661
rect 24634 17620 24643 17660
rect 24683 17620 24692 17660
rect 24634 17619 24692 17620
rect 28491 17660 28533 17669
rect 28491 17620 28492 17660
rect 28532 17620 28533 17660
rect 28491 17611 28533 17620
rect 1611 17576 1653 17585
rect 1611 17536 1612 17576
rect 1652 17536 1653 17576
rect 1611 17527 1653 17536
rect 2379 17576 2421 17585
rect 2379 17536 2380 17576
rect 2420 17536 2421 17576
rect 2379 17527 2421 17536
rect 3418 17576 3476 17577
rect 3418 17536 3427 17576
rect 3467 17536 3476 17576
rect 3418 17535 3476 17536
rect 3531 17576 3573 17585
rect 3531 17536 3532 17576
rect 3572 17536 3573 17576
rect 3531 17527 3573 17536
rect 4779 17576 4821 17585
rect 4779 17536 4780 17576
rect 4820 17536 4821 17576
rect 4779 17527 4821 17536
rect 7083 17576 7125 17585
rect 7083 17536 7084 17576
rect 7124 17536 7125 17576
rect 7083 17527 7125 17536
rect 10443 17576 10485 17585
rect 10443 17536 10444 17576
rect 10484 17536 10485 17576
rect 10443 17527 10485 17536
rect 14602 17576 14660 17577
rect 14602 17536 14611 17576
rect 14651 17536 14660 17576
rect 14602 17535 14660 17536
rect 14955 17576 14997 17585
rect 14955 17536 14956 17576
rect 14996 17536 14997 17576
rect 14955 17527 14997 17536
rect 15226 17576 15284 17577
rect 15226 17536 15235 17576
rect 15275 17536 15284 17576
rect 15226 17535 15284 17536
rect 16090 17576 16148 17577
rect 16090 17536 16099 17576
rect 16139 17536 16148 17576
rect 16090 17535 16148 17536
rect 17643 17576 17685 17585
rect 17643 17536 17644 17576
rect 17684 17536 17685 17576
rect 17643 17527 17685 17536
rect 18010 17576 18068 17577
rect 18010 17536 18019 17576
rect 18059 17536 18068 17576
rect 18010 17535 18068 17536
rect 19546 17576 19604 17577
rect 19546 17536 19555 17576
rect 19595 17536 19604 17576
rect 19546 17535 19604 17536
rect 23962 17576 24020 17577
rect 23962 17536 23971 17576
rect 24011 17536 24020 17576
rect 23962 17535 24020 17536
rect 24939 17576 24981 17585
rect 24939 17536 24940 17576
rect 24980 17536 24981 17576
rect 24939 17527 24981 17536
rect 25995 17576 26037 17585
rect 25995 17536 25996 17576
rect 26036 17536 26037 17576
rect 25995 17527 26037 17536
rect 29146 17576 29204 17577
rect 29146 17536 29155 17576
rect 29195 17536 29204 17576
rect 29146 17535 29204 17536
rect 29451 17576 29493 17585
rect 29451 17536 29452 17576
rect 29492 17536 29493 17576
rect 29451 17527 29493 17536
rect 576 17408 31392 17432
rect 576 17368 4352 17408
rect 4720 17368 12126 17408
rect 12494 17368 19900 17408
rect 20268 17368 27674 17408
rect 28042 17368 31392 17408
rect 576 17344 31392 17368
rect 5163 17240 5205 17249
rect 5163 17200 5164 17240
rect 5204 17200 5205 17240
rect 5163 17191 5205 17200
rect 6171 17240 6213 17249
rect 6171 17200 6172 17240
rect 6212 17200 6213 17240
rect 6171 17191 6213 17200
rect 9099 17240 9141 17249
rect 9099 17200 9100 17240
rect 9140 17200 9141 17240
rect 9099 17191 9141 17200
rect 11098 17240 11156 17241
rect 11098 17200 11107 17240
rect 11147 17200 11156 17240
rect 11098 17199 11156 17200
rect 11578 17240 11636 17241
rect 11578 17200 11587 17240
rect 11627 17200 11636 17240
rect 11578 17199 11636 17200
rect 13411 17240 13469 17241
rect 13411 17200 13420 17240
rect 13460 17200 13469 17240
rect 13411 17199 13469 17200
rect 16858 17240 16916 17241
rect 16858 17200 16867 17240
rect 16907 17200 16916 17240
rect 16858 17199 16916 17200
rect 18970 17240 19028 17241
rect 18970 17200 18979 17240
rect 19019 17200 19028 17240
rect 18970 17199 19028 17200
rect 25738 17240 25796 17241
rect 25738 17200 25747 17240
rect 25787 17200 25796 17240
rect 25738 17199 25796 17200
rect 29355 17240 29397 17249
rect 29355 17200 29356 17240
rect 29396 17200 29397 17240
rect 29355 17191 29397 17200
rect 640 17156 682 17165
rect 640 17116 641 17156
rect 681 17116 682 17156
rect 640 17107 682 17116
rect 1899 17156 1941 17165
rect 1899 17116 1900 17156
rect 1940 17116 1941 17156
rect 1899 17107 1941 17116
rect 4858 17156 4916 17157
rect 4858 17116 4867 17156
rect 4907 17116 4916 17156
rect 4858 17115 4916 17116
rect 6586 17156 6644 17157
rect 6586 17116 6595 17156
rect 6635 17116 6644 17156
rect 6586 17115 6644 17116
rect 8331 17156 8373 17165
rect 10810 17156 10868 17157
rect 8331 17116 8332 17156
rect 8372 17116 8373 17156
rect 8331 17107 8373 17116
rect 9186 17147 9232 17156
rect 9186 17107 9187 17147
rect 9227 17107 9232 17147
rect 10810 17116 10819 17156
rect 10859 17116 10868 17156
rect 10810 17115 10868 17116
rect 11005 17156 11047 17165
rect 11005 17116 11006 17156
rect 11046 17116 11047 17156
rect 11005 17107 11047 17116
rect 11211 17156 11253 17165
rect 11211 17116 11212 17156
rect 11252 17116 11253 17156
rect 11211 17107 11253 17116
rect 11691 17156 11733 17165
rect 20410 17156 20468 17157
rect 11691 17116 11692 17156
rect 11732 17116 11733 17156
rect 11691 17107 11733 17116
rect 18114 17147 18160 17156
rect 18114 17107 18115 17147
rect 18155 17107 18160 17147
rect 20410 17116 20419 17156
rect 20459 17116 20468 17156
rect 20410 17115 20468 17116
rect 24267 17156 24309 17165
rect 24267 17116 24268 17156
rect 24308 17116 24309 17156
rect 24267 17107 24309 17116
rect 24473 17156 24515 17165
rect 24473 17116 24474 17156
rect 24514 17116 24515 17156
rect 24473 17107 24515 17116
rect 9186 17098 9232 17107
rect 18114 17098 18160 17107
rect 843 17072 885 17081
rect 1306 17072 1364 17073
rect 843 17032 844 17072
rect 884 17032 885 17072
rect 843 17023 885 17032
rect 939 17063 981 17072
rect 939 17023 940 17063
rect 980 17023 981 17063
rect 1306 17032 1315 17072
rect 1355 17032 1364 17072
rect 1306 17031 1364 17032
rect 1995 17072 2037 17081
rect 1995 17032 1996 17072
rect 2036 17032 2037 17072
rect 1995 17023 2037 17032
rect 2224 17072 2282 17073
rect 2224 17032 2233 17072
rect 2273 17032 2282 17072
rect 2224 17031 2282 17032
rect 2379 17072 2421 17081
rect 2379 17032 2380 17072
rect 2420 17032 2421 17072
rect 2379 17023 2421 17032
rect 2552 17072 2594 17081
rect 2552 17032 2553 17072
rect 2593 17032 2594 17072
rect 2552 17023 2594 17032
rect 2763 17072 2805 17081
rect 2763 17032 2764 17072
rect 2804 17032 2805 17072
rect 2763 17023 2805 17032
rect 2938 17072 2996 17073
rect 2938 17032 2947 17072
rect 2987 17032 2996 17072
rect 2938 17031 2996 17032
rect 4186 17072 4244 17073
rect 4186 17032 4195 17072
rect 4235 17032 4244 17072
rect 4186 17031 4244 17032
rect 4534 17072 4576 17081
rect 4534 17032 4535 17072
rect 4575 17032 4576 17072
rect 4534 17023 4576 17032
rect 4779 17072 4821 17081
rect 4779 17032 4780 17072
rect 4820 17032 4821 17072
rect 4779 17023 4821 17032
rect 5062 17072 5104 17081
rect 5062 17032 5063 17072
rect 5103 17032 5104 17072
rect 5062 17023 5104 17032
rect 5242 17072 5300 17073
rect 5242 17032 5251 17072
rect 5291 17032 5300 17072
rect 5242 17031 5300 17032
rect 6027 17072 6069 17081
rect 6027 17032 6028 17072
rect 6068 17032 6069 17072
rect 6027 17023 6069 17032
rect 6987 17072 7029 17081
rect 6987 17032 6988 17072
rect 7028 17032 7029 17072
rect 6987 17023 7029 17032
rect 8139 17072 8181 17081
rect 8139 17032 8140 17072
rect 8180 17032 8181 17072
rect 8139 17023 8181 17032
rect 8442 17072 8484 17081
rect 8442 17032 8443 17072
rect 8483 17032 8484 17072
rect 8442 17023 8484 17032
rect 8890 17072 8948 17073
rect 9270 17072 9328 17073
rect 8890 17032 8899 17072
rect 8939 17032 8948 17072
rect 8890 17031 8948 17032
rect 9003 17063 9045 17072
rect 9003 17023 9004 17063
rect 9044 17023 9045 17063
rect 9270 17032 9279 17072
rect 9319 17032 9328 17072
rect 9270 17031 9328 17032
rect 9451 17072 9509 17073
rect 9451 17032 9460 17072
rect 9500 17032 9509 17072
rect 9451 17031 9509 17032
rect 10498 17072 10556 17073
rect 10498 17032 10507 17072
rect 10547 17032 10556 17072
rect 10498 17031 10556 17032
rect 10731 17072 10773 17081
rect 10731 17032 10732 17072
rect 10772 17032 10773 17072
rect 11482 17072 11540 17073
rect 10731 17023 10773 17032
rect 11297 17047 11339 17056
rect 939 17014 981 17023
rect 9003 17014 9045 17023
rect 11297 17007 11298 17047
rect 11338 17007 11339 17047
rect 11482 17032 11491 17072
rect 11531 17032 11540 17072
rect 11482 17031 11540 17032
rect 11798 17072 11840 17081
rect 11798 17032 11799 17072
rect 11839 17032 11840 17072
rect 11798 17023 11840 17032
rect 12459 17072 12501 17081
rect 12459 17032 12460 17072
rect 12500 17032 12501 17072
rect 12459 17023 12501 17032
rect 12778 17072 12836 17073
rect 12778 17032 12787 17072
rect 12827 17032 12836 17072
rect 12778 17031 12836 17032
rect 13018 17072 13076 17073
rect 13018 17032 13027 17072
rect 13067 17032 13076 17072
rect 13018 17031 13076 17032
rect 13563 17072 13605 17081
rect 13563 17032 13564 17072
rect 13604 17032 13605 17072
rect 13563 17023 13605 17032
rect 13899 17072 13941 17081
rect 13899 17032 13900 17072
rect 13940 17032 13941 17072
rect 13899 17023 13941 17032
rect 14863 17072 14921 17073
rect 15994 17072 16052 17073
rect 14863 17032 14872 17072
rect 14912 17032 14921 17072
rect 14863 17031 14921 17032
rect 15234 17063 15280 17072
rect 15234 17023 15235 17063
rect 15275 17023 15280 17063
rect 15994 17032 16003 17072
rect 16043 17032 16052 17072
rect 15994 17031 16052 17032
rect 16299 17072 16341 17081
rect 16299 17032 16300 17072
rect 16340 17032 16341 17072
rect 16299 17023 16341 17032
rect 16779 17072 16821 17081
rect 16779 17032 16780 17072
rect 16820 17032 16821 17072
rect 16779 17023 16821 17032
rect 17355 17072 17397 17081
rect 17355 17032 17356 17072
rect 17396 17032 17397 17072
rect 17355 17023 17397 17032
rect 17658 17072 17700 17081
rect 17658 17032 17659 17072
rect 17699 17032 17700 17072
rect 17658 17023 17700 17032
rect 17818 17072 17876 17073
rect 18205 17072 18247 17081
rect 17818 17032 17827 17072
rect 17867 17032 17876 17072
rect 17818 17031 17876 17032
rect 17931 17063 17973 17072
rect 17931 17023 17932 17063
rect 17972 17023 17973 17063
rect 18205 17032 18206 17072
rect 18246 17032 18247 17072
rect 18205 17023 18247 17032
rect 18378 17072 18436 17073
rect 18378 17032 18387 17072
rect 18427 17032 18436 17072
rect 18378 17031 18436 17032
rect 18619 17072 18677 17073
rect 18619 17032 18628 17072
rect 18668 17032 18677 17072
rect 18619 17031 18677 17032
rect 18778 17072 18836 17073
rect 18778 17032 18787 17072
rect 18827 17032 18836 17072
rect 18778 17031 18836 17032
rect 18903 17072 18945 17081
rect 18903 17032 18904 17072
rect 18944 17032 18945 17072
rect 18903 17023 18945 17032
rect 19066 17072 19124 17073
rect 19066 17032 19075 17072
rect 19115 17032 19124 17072
rect 19066 17031 19124 17032
rect 19188 17072 19246 17073
rect 19188 17032 19197 17072
rect 19237 17032 19246 17072
rect 19188 17031 19246 17032
rect 19851 17072 19893 17081
rect 19851 17032 19852 17072
rect 19892 17032 19893 17072
rect 19851 17023 19893 17032
rect 20086 17072 20128 17081
rect 20086 17032 20087 17072
rect 20127 17032 20128 17072
rect 20086 17023 20128 17032
rect 20331 17072 20373 17081
rect 20331 17032 20332 17072
rect 20372 17032 20373 17072
rect 20331 17023 20373 17032
rect 20619 17072 20661 17081
rect 20619 17032 20620 17072
rect 20660 17032 20661 17072
rect 20619 17023 20661 17032
rect 20794 17072 20852 17073
rect 20794 17032 20803 17072
rect 20843 17032 20852 17072
rect 20794 17031 20852 17032
rect 21387 17072 21429 17081
rect 21387 17032 21388 17072
rect 21428 17032 21429 17072
rect 21387 17023 21429 17032
rect 21508 17072 21566 17073
rect 21508 17032 21517 17072
rect 21557 17032 21566 17072
rect 21508 17031 21566 17032
rect 21771 17072 21813 17081
rect 21771 17032 21772 17072
rect 21812 17032 21813 17072
rect 21771 17023 21813 17032
rect 22539 17072 22581 17081
rect 23691 17072 23733 17081
rect 22539 17032 22540 17072
rect 22580 17032 22581 17072
rect 22539 17023 22581 17032
rect 22818 17063 22864 17072
rect 22818 17023 22819 17063
rect 22859 17023 22864 17063
rect 23691 17032 23692 17072
rect 23732 17032 23733 17072
rect 23691 17023 23733 17032
rect 23866 17072 23924 17073
rect 23866 17032 23875 17072
rect 23915 17032 23924 17072
rect 23866 17031 23924 17032
rect 23979 17072 24021 17081
rect 23979 17032 23980 17072
rect 24020 17032 24021 17072
rect 23979 17023 24021 17032
rect 24165 17072 24223 17073
rect 24165 17032 24174 17072
rect 24214 17032 24223 17072
rect 24165 17031 24223 17032
rect 25323 17072 25365 17081
rect 25323 17032 25324 17072
rect 25364 17032 25365 17072
rect 25323 17023 25365 17032
rect 25933 17072 25991 17073
rect 25933 17032 25942 17072
rect 25982 17032 25991 17072
rect 25933 17031 25991 17032
rect 28570 17072 28628 17073
rect 28570 17032 28579 17072
rect 28619 17032 28628 17072
rect 28570 17031 28628 17032
rect 30027 17072 30069 17081
rect 30027 17032 30028 17072
rect 30068 17032 30069 17072
rect 30027 17023 30069 17032
rect 15234 17014 15280 17023
rect 17931 17014 17973 17023
rect 22818 17014 22864 17023
rect 11297 16998 11339 17007
rect 1131 16988 1173 16997
rect 1131 16948 1132 16988
rect 1172 16948 1173 16988
rect 1131 16939 1173 16948
rect 1707 16988 1749 16997
rect 3802 16988 3860 16989
rect 1707 16948 1708 16988
rect 1748 16948 1749 16988
rect 1707 16939 1749 16948
rect 2130 16979 2176 16988
rect 2130 16939 2131 16979
rect 2171 16939 2176 16979
rect 3802 16948 3811 16988
rect 3851 16948 3860 16988
rect 3802 16947 3860 16948
rect 4378 16988 4436 16989
rect 4378 16948 4387 16988
rect 4427 16948 4436 16988
rect 4378 16947 4436 16948
rect 4666 16988 4724 16989
rect 4666 16948 4675 16988
rect 4715 16948 4724 16988
rect 4666 16947 4724 16948
rect 10618 16988 10676 16989
rect 10618 16948 10627 16988
rect 10667 16948 10676 16988
rect 10618 16947 10676 16948
rect 14698 16988 14756 16989
rect 14698 16948 14707 16988
rect 14747 16948 14756 16988
rect 14698 16947 14756 16948
rect 15387 16988 15429 16997
rect 15387 16948 15388 16988
rect 15428 16948 15429 16988
rect 15387 16939 15429 16948
rect 20218 16988 20276 16989
rect 20218 16948 20227 16988
rect 20267 16948 20276 16988
rect 20218 16947 20276 16948
rect 22971 16988 23013 16997
rect 22971 16948 22972 16988
rect 23012 16948 23013 16988
rect 22971 16939 23013 16948
rect 27034 16988 27092 16989
rect 27034 16948 27043 16988
rect 27083 16948 27092 16988
rect 27034 16947 27092 16948
rect 28954 16988 29012 16989
rect 28954 16948 28963 16988
rect 29003 16948 29012 16988
rect 28954 16947 29012 16948
rect 2130 16930 2176 16939
rect 1611 16904 1653 16913
rect 1611 16864 1612 16904
rect 1652 16864 1653 16904
rect 1611 16855 1653 16864
rect 3898 16904 3956 16905
rect 3898 16864 3907 16904
rect 3947 16864 3956 16904
rect 3898 16863 3956 16864
rect 13114 16904 13172 16905
rect 13114 16864 13123 16904
rect 13163 16864 13172 16904
rect 13114 16863 13172 16864
rect 16587 16904 16629 16913
rect 16587 16864 16588 16904
rect 16628 16864 16629 16904
rect 16587 16855 16629 16864
rect 19450 16904 19508 16905
rect 19450 16864 19459 16904
rect 19499 16864 19508 16904
rect 19450 16863 19508 16864
rect 20794 16904 20852 16905
rect 20794 16864 20803 16904
rect 20843 16864 20852 16904
rect 20794 16863 20852 16864
rect 21099 16904 21141 16913
rect 21099 16864 21100 16904
rect 21140 16864 21141 16904
rect 21099 16855 21141 16864
rect 30411 16904 30453 16913
rect 30411 16864 30412 16904
rect 30452 16864 30453 16904
rect 30411 16855 30453 16864
rect 30603 16904 30645 16913
rect 30603 16864 30604 16904
rect 30644 16864 30645 16904
rect 30603 16855 30645 16864
rect 634 16820 692 16821
rect 634 16780 643 16820
rect 683 16780 692 16820
rect 634 16779 692 16780
rect 2379 16820 2421 16829
rect 2379 16780 2380 16820
rect 2420 16780 2421 16820
rect 2379 16771 2421 16780
rect 2938 16820 2996 16821
rect 2938 16780 2947 16820
rect 2987 16780 2996 16820
rect 2938 16779 2996 16780
rect 12651 16820 12693 16829
rect 12651 16780 12652 16820
rect 12692 16780 12693 16820
rect 12651 16771 12693 16780
rect 13690 16820 13748 16821
rect 13690 16780 13699 16820
rect 13739 16780 13748 16820
rect 13690 16779 13748 16780
rect 15819 16820 15861 16829
rect 15819 16780 15820 16820
rect 15860 16780 15861 16820
rect 15819 16771 15861 16780
rect 17547 16820 17589 16829
rect 17547 16780 17548 16820
rect 17588 16780 17589 16820
rect 17547 16771 17589 16780
rect 17818 16820 17876 16821
rect 17818 16780 17827 16820
rect 17867 16780 17876 16820
rect 17818 16779 17876 16780
rect 22138 16820 22196 16821
rect 22138 16780 22147 16820
rect 22187 16780 22196 16820
rect 22138 16779 22196 16780
rect 23979 16820 24021 16829
rect 23979 16780 23980 16820
rect 24020 16780 24021 16820
rect 23979 16771 24021 16780
rect 24459 16820 24501 16829
rect 24459 16780 24460 16820
rect 24500 16780 24501 16820
rect 24459 16771 24501 16780
rect 24922 16820 24980 16821
rect 24922 16780 24931 16820
rect 24971 16780 24980 16820
rect 24922 16779 24980 16780
rect 26667 16820 26709 16829
rect 26667 16780 26668 16820
rect 26708 16780 26709 16820
rect 26667 16771 26709 16780
rect 576 16652 31392 16676
rect 576 16612 3112 16652
rect 3480 16612 10886 16652
rect 11254 16612 18660 16652
rect 19028 16612 26434 16652
rect 26802 16612 31392 16652
rect 576 16588 31392 16612
rect 2650 16484 2708 16485
rect 2650 16444 2659 16484
rect 2699 16444 2708 16484
rect 2650 16443 2708 16444
rect 4299 16484 4341 16493
rect 4299 16444 4300 16484
rect 4340 16444 4341 16484
rect 4299 16435 4341 16444
rect 6682 16484 6740 16485
rect 6682 16444 6691 16484
rect 6731 16444 6740 16484
rect 6682 16443 6740 16444
rect 7354 16484 7412 16485
rect 7354 16444 7363 16484
rect 7403 16444 7412 16484
rect 7354 16443 7412 16444
rect 9963 16484 10005 16493
rect 9963 16444 9964 16484
rect 10004 16444 10005 16484
rect 9963 16435 10005 16444
rect 12058 16484 12116 16485
rect 12058 16444 12067 16484
rect 12107 16444 12116 16484
rect 12058 16443 12116 16444
rect 16090 16484 16148 16485
rect 16090 16444 16099 16484
rect 16139 16444 16148 16484
rect 16090 16443 16148 16444
rect 16587 16484 16629 16493
rect 16587 16444 16588 16484
rect 16628 16444 16629 16484
rect 16587 16435 16629 16444
rect 17818 16484 17876 16485
rect 17818 16444 17827 16484
rect 17867 16444 17876 16484
rect 17818 16443 17876 16444
rect 24555 16484 24597 16493
rect 24555 16444 24556 16484
rect 24596 16444 24597 16484
rect 24555 16435 24597 16444
rect 26091 16484 26133 16493
rect 26091 16444 26092 16484
rect 26132 16444 26133 16484
rect 26091 16435 26133 16444
rect 28971 16484 29013 16493
rect 28971 16444 28972 16484
rect 29012 16444 29013 16484
rect 28971 16435 29013 16444
rect 29355 16484 29397 16493
rect 29355 16444 29356 16484
rect 29396 16444 29397 16484
rect 29355 16435 29397 16444
rect 9003 16400 9045 16409
rect 9003 16360 9004 16400
rect 9044 16360 9045 16400
rect 9003 16351 9045 16360
rect 22827 16400 22869 16409
rect 22827 16360 22828 16400
rect 22868 16360 22869 16400
rect 22827 16351 22869 16360
rect 28395 16400 28437 16409
rect 28395 16360 28396 16400
rect 28436 16360 28437 16400
rect 28395 16351 28437 16360
rect 1419 16316 1461 16325
rect 1419 16276 1420 16316
rect 1460 16276 1461 16316
rect 1419 16267 1461 16276
rect 1611 16316 1653 16325
rect 6970 16316 7028 16317
rect 1611 16276 1612 16316
rect 1652 16276 1653 16316
rect 1611 16267 1653 16276
rect 1842 16307 1888 16316
rect 1842 16267 1843 16307
rect 1883 16267 1888 16307
rect 6970 16276 6979 16316
rect 7019 16276 7028 16316
rect 6970 16275 7028 16276
rect 7179 16316 7221 16325
rect 7179 16276 7180 16316
rect 7220 16276 7221 16316
rect 1842 16258 1888 16267
rect 5578 16274 5636 16275
rect 1078 16232 1120 16241
rect 1078 16192 1079 16232
rect 1119 16192 1120 16232
rect 1078 16183 1120 16192
rect 1210 16232 1268 16233
rect 1210 16192 1219 16232
rect 1259 16192 1268 16232
rect 1210 16191 1268 16192
rect 1323 16232 1365 16241
rect 1323 16192 1324 16232
rect 1364 16192 1365 16232
rect 1323 16183 1365 16192
rect 1707 16232 1749 16241
rect 1707 16192 1708 16232
rect 1748 16192 1749 16232
rect 1707 16183 1749 16192
rect 1936 16232 1994 16233
rect 1936 16192 1945 16232
rect 1985 16192 1994 16232
rect 1936 16191 1994 16192
rect 2187 16232 2229 16241
rect 2187 16192 2188 16232
rect 2228 16192 2229 16232
rect 2187 16183 2229 16192
rect 2306 16232 2348 16241
rect 2306 16192 2307 16232
rect 2347 16192 2348 16232
rect 2306 16183 2348 16192
rect 2416 16232 2474 16233
rect 2416 16192 2425 16232
rect 2465 16192 2474 16232
rect 2416 16191 2474 16192
rect 2947 16232 3005 16233
rect 2947 16192 2956 16232
rect 2996 16192 3005 16232
rect 2947 16191 3005 16192
rect 3994 16232 4052 16233
rect 3994 16192 4003 16232
rect 4043 16192 4052 16232
rect 3994 16191 4052 16192
rect 4313 16232 4355 16241
rect 4313 16192 4314 16232
rect 4354 16192 4355 16232
rect 4313 16183 4355 16192
rect 4480 16232 4522 16241
rect 5578 16234 5587 16274
rect 5627 16234 5636 16274
rect 7179 16267 7221 16276
rect 10731 16316 10773 16325
rect 10731 16276 10732 16316
rect 10772 16276 10773 16316
rect 10731 16267 10773 16276
rect 19306 16316 19364 16317
rect 19306 16276 19315 16316
rect 19355 16276 19364 16316
rect 19306 16275 19364 16276
rect 21483 16316 21525 16325
rect 21483 16276 21484 16316
rect 21524 16276 21525 16316
rect 19498 16274 19556 16275
rect 5578 16233 5636 16234
rect 4480 16192 4481 16232
rect 4521 16192 4522 16232
rect 4480 16183 4522 16192
rect 4777 16232 4835 16233
rect 4777 16192 4786 16232
rect 4826 16192 4835 16232
rect 4777 16191 4835 16192
rect 5386 16232 5444 16233
rect 5386 16192 5395 16232
rect 5435 16192 5444 16232
rect 5386 16191 5444 16192
rect 5755 16232 5813 16233
rect 5755 16192 5764 16232
rect 5804 16192 5813 16232
rect 5755 16191 5813 16192
rect 5936 16232 5978 16241
rect 5936 16192 5937 16232
rect 5977 16192 5978 16232
rect 5936 16183 5978 16192
rect 6058 16232 6116 16233
rect 6058 16192 6067 16232
rect 6107 16192 6116 16232
rect 6058 16191 6116 16192
rect 6170 16232 6228 16233
rect 6170 16192 6179 16232
rect 6219 16192 6228 16232
rect 6170 16191 6228 16192
rect 6298 16232 6356 16233
rect 6298 16192 6307 16232
rect 6347 16192 6356 16232
rect 6298 16191 6356 16192
rect 6507 16232 6549 16241
rect 6507 16192 6508 16232
rect 6548 16192 6549 16232
rect 6507 16183 6549 16192
rect 6682 16232 6740 16233
rect 6682 16192 6691 16232
rect 6731 16192 6740 16232
rect 6682 16191 6740 16192
rect 6838 16232 6880 16241
rect 6838 16192 6839 16232
rect 6879 16192 6880 16232
rect 6838 16183 6880 16192
rect 7083 16232 7125 16241
rect 7083 16192 7084 16232
rect 7124 16192 7125 16232
rect 7083 16183 7125 16192
rect 7346 16232 7404 16233
rect 7346 16192 7355 16232
rect 7395 16192 7404 16232
rect 7346 16191 7404 16192
rect 7510 16232 7568 16233
rect 7510 16192 7519 16232
rect 7559 16192 7568 16232
rect 7510 16191 7568 16192
rect 7638 16232 7696 16233
rect 7638 16192 7647 16232
rect 7687 16192 7696 16232
rect 7638 16191 7696 16192
rect 7738 16232 7796 16233
rect 7738 16192 7747 16232
rect 7787 16192 7796 16232
rect 7738 16191 7796 16192
rect 7915 16232 7973 16233
rect 7915 16192 7924 16232
rect 7964 16192 7973 16232
rect 7915 16191 7973 16192
rect 8749 16232 8807 16233
rect 8749 16192 8758 16232
rect 8798 16192 8807 16232
rect 8749 16191 8807 16192
rect 9178 16232 9236 16233
rect 9178 16192 9187 16232
rect 9227 16192 9236 16232
rect 9178 16191 9236 16192
rect 9483 16232 9525 16241
rect 9483 16192 9484 16232
rect 9524 16192 9525 16232
rect 9483 16183 9525 16192
rect 9658 16232 9716 16233
rect 9658 16192 9667 16232
rect 9707 16192 9716 16232
rect 9658 16191 9716 16192
rect 10390 16232 10432 16241
rect 10390 16192 10391 16232
rect 10431 16192 10432 16232
rect 10390 16183 10432 16192
rect 10522 16232 10580 16233
rect 10522 16192 10531 16232
rect 10571 16192 10580 16232
rect 10522 16191 10580 16192
rect 10635 16232 10677 16241
rect 10635 16192 10636 16232
rect 10676 16192 10677 16232
rect 10635 16183 10677 16192
rect 11917 16232 11975 16233
rect 11917 16192 11926 16232
rect 11966 16192 11975 16232
rect 11917 16191 11975 16192
rect 12267 16232 12309 16241
rect 12267 16192 12268 16232
rect 12308 16192 12309 16232
rect 12267 16183 12309 16192
rect 12355 16232 12413 16233
rect 12355 16192 12364 16232
rect 12404 16192 12413 16232
rect 12355 16191 12413 16192
rect 13035 16232 13077 16241
rect 13035 16192 13036 16232
rect 13076 16192 13077 16232
rect 13035 16183 13077 16192
rect 13154 16232 13196 16241
rect 13154 16192 13155 16232
rect 13195 16192 13196 16232
rect 13154 16183 13196 16192
rect 13264 16232 13322 16233
rect 13264 16192 13273 16232
rect 13313 16192 13322 16232
rect 13264 16191 13322 16192
rect 13741 16232 13799 16233
rect 13741 16192 13750 16232
rect 13790 16192 13799 16232
rect 13741 16191 13799 16192
rect 14859 16232 14901 16241
rect 14859 16192 14860 16232
rect 14900 16192 14901 16232
rect 14859 16183 14901 16192
rect 15243 16232 15285 16241
rect 15243 16192 15244 16232
rect 15284 16192 15285 16232
rect 15243 16183 15285 16192
rect 15562 16232 15620 16233
rect 15562 16192 15571 16232
rect 15611 16192 15620 16232
rect 15562 16191 15620 16192
rect 16096 16232 16138 16241
rect 16096 16192 16097 16232
rect 16137 16192 16138 16232
rect 16096 16183 16138 16192
rect 16387 16232 16445 16233
rect 16387 16192 16396 16232
rect 16436 16192 16445 16232
rect 16387 16191 16445 16192
rect 16587 16232 16629 16241
rect 16587 16192 16588 16232
rect 16628 16192 16629 16232
rect 16587 16183 16629 16192
rect 16779 16232 16821 16241
rect 16779 16192 16780 16232
rect 16820 16192 16821 16232
rect 16779 16183 16821 16192
rect 17643 16232 17685 16241
rect 19498 16234 19507 16274
rect 19547 16234 19556 16274
rect 21483 16267 21525 16276
rect 23578 16316 23636 16317
rect 23578 16276 23587 16316
rect 23627 16276 23636 16316
rect 27819 16316 27861 16325
rect 23578 16275 23636 16276
rect 26763 16274 26805 16283
rect 19498 16233 19556 16234
rect 17643 16192 17644 16232
rect 17684 16192 17685 16232
rect 17643 16183 17685 16192
rect 17818 16232 17876 16233
rect 17818 16192 17827 16232
rect 17867 16192 17876 16232
rect 17818 16191 17876 16192
rect 19659 16232 19701 16241
rect 19659 16192 19660 16232
rect 19700 16192 19701 16232
rect 19659 16183 19701 16192
rect 19851 16232 19893 16241
rect 19851 16192 19852 16232
rect 19892 16192 19893 16232
rect 19851 16183 19893 16192
rect 20506 16232 20564 16233
rect 20506 16192 20515 16232
rect 20555 16192 20564 16232
rect 20506 16191 20564 16192
rect 20995 16232 21053 16233
rect 20995 16192 21004 16232
rect 21044 16192 21053 16232
rect 20995 16191 21053 16192
rect 21579 16232 21621 16241
rect 21579 16192 21580 16232
rect 21620 16192 21621 16232
rect 21579 16183 21621 16192
rect 21963 16232 22005 16241
rect 21963 16192 21964 16232
rect 22004 16192 22005 16232
rect 21963 16183 22005 16192
rect 22073 16232 22131 16233
rect 22073 16192 22082 16232
rect 22122 16192 22131 16232
rect 22073 16191 22131 16192
rect 22870 16232 22912 16241
rect 23115 16232 23157 16241
rect 22870 16192 22871 16232
rect 22911 16192 22912 16232
rect 22870 16183 22912 16192
rect 23010 16223 23056 16232
rect 23010 16183 23011 16223
rect 23051 16183 23056 16223
rect 23115 16192 23116 16232
rect 23156 16192 23157 16232
rect 23115 16183 23157 16192
rect 23446 16232 23488 16241
rect 23446 16192 23447 16232
rect 23487 16192 23488 16232
rect 23446 16183 23488 16192
rect 23691 16232 23733 16241
rect 23691 16192 23692 16232
rect 23732 16192 23733 16232
rect 23691 16183 23733 16192
rect 23931 16232 23973 16241
rect 23931 16192 23932 16232
rect 23972 16192 23973 16232
rect 23931 16183 23973 16192
rect 24058 16232 24116 16233
rect 24058 16192 24067 16232
rect 24107 16192 24116 16232
rect 24058 16191 24116 16192
rect 24171 16232 24213 16241
rect 24171 16192 24172 16232
rect 24212 16192 24213 16232
rect 24171 16183 24213 16192
rect 24459 16232 24501 16241
rect 24459 16192 24460 16232
rect 24500 16192 24501 16232
rect 24459 16183 24501 16192
rect 25786 16232 25844 16233
rect 25786 16192 25795 16232
rect 25835 16192 25844 16232
rect 25786 16191 25844 16192
rect 26427 16232 26469 16241
rect 26427 16192 26428 16232
rect 26468 16192 26469 16232
rect 26427 16183 26469 16192
rect 26619 16232 26661 16241
rect 26619 16192 26620 16232
rect 26660 16192 26661 16232
rect 26763 16234 26764 16274
rect 26804 16234 26805 16274
rect 27819 16276 27820 16316
rect 27860 16276 27861 16316
rect 27819 16267 27861 16276
rect 31258 16316 31316 16317
rect 31258 16276 31267 16316
rect 31307 16276 31316 16316
rect 31258 16275 31316 16276
rect 26763 16225 26805 16234
rect 26955 16232 26997 16241
rect 26619 16183 26661 16192
rect 26955 16192 26956 16232
rect 26996 16192 26997 16232
rect 26955 16183 26997 16192
rect 27147 16232 27189 16241
rect 27147 16192 27148 16232
rect 27188 16192 27189 16232
rect 27147 16183 27189 16192
rect 28011 16232 28053 16241
rect 28011 16192 28012 16232
rect 28052 16192 28053 16232
rect 28011 16183 28053 16192
rect 28203 16232 28245 16241
rect 28203 16192 28204 16232
rect 28244 16192 28245 16232
rect 28203 16183 28245 16192
rect 30874 16232 30932 16233
rect 30874 16192 30883 16232
rect 30923 16192 30932 16232
rect 30874 16191 30932 16192
rect 23010 16174 23056 16183
rect 2653 16148 2695 16157
rect 2653 16108 2654 16148
rect 2694 16108 2695 16148
rect 2653 16099 2695 16108
rect 4570 16148 4628 16149
rect 4570 16108 4579 16148
rect 4619 16108 4628 16148
rect 4570 16107 4628 16108
rect 9771 16148 9813 16157
rect 9771 16108 9772 16148
rect 9812 16108 9813 16148
rect 9771 16099 9813 16108
rect 9974 16148 10016 16157
rect 9974 16108 9975 16148
rect 10015 16108 10016 16148
rect 9974 16099 10016 16108
rect 12061 16148 12103 16157
rect 12061 16108 12062 16148
rect 12102 16108 12103 16148
rect 12061 16099 12103 16108
rect 15435 16148 15477 16157
rect 15435 16108 15436 16148
rect 15476 16108 15477 16148
rect 15435 16099 15477 16108
rect 19755 16148 19797 16157
rect 19755 16108 19756 16148
rect 19796 16108 19797 16148
rect 19755 16099 19797 16108
rect 23770 16148 23828 16149
rect 23770 16108 23779 16148
rect 23819 16108 23828 16148
rect 23770 16107 23828 16108
rect 26102 16148 26144 16157
rect 26102 16108 26103 16148
rect 26143 16108 26144 16148
rect 26102 16099 26144 16108
rect 2091 16064 2133 16073
rect 2091 16024 2092 16064
rect 2132 16024 2133 16064
rect 2091 16015 2133 16024
rect 2859 16064 2901 16073
rect 2859 16024 2860 16064
rect 2900 16024 2901 16064
rect 2859 16015 2901 16024
rect 4090 16064 4148 16065
rect 4090 16024 4099 16064
rect 4139 16024 4148 16064
rect 4090 16023 4148 16024
rect 4683 16064 4725 16073
rect 4683 16024 4684 16064
rect 4724 16024 4725 16064
rect 4683 16015 4725 16024
rect 5818 16064 5876 16065
rect 5818 16024 5827 16064
rect 5867 16024 5876 16064
rect 5818 16023 5876 16024
rect 8554 16064 8612 16065
rect 8554 16024 8563 16064
rect 8603 16024 8612 16064
rect 8554 16023 8612 16024
rect 11722 16064 11780 16065
rect 11722 16024 11731 16064
rect 11771 16024 11780 16064
rect 11722 16023 11780 16024
rect 12267 16064 12309 16073
rect 12267 16024 12268 16064
rect 12308 16024 12309 16064
rect 12267 16015 12309 16024
rect 12939 16064 12981 16073
rect 12939 16024 12940 16064
rect 12980 16024 12981 16064
rect 12939 16015 12981 16024
rect 13546 16064 13604 16065
rect 13546 16024 13555 16064
rect 13595 16024 13604 16064
rect 13546 16023 13604 16024
rect 14667 16064 14709 16073
rect 14667 16024 14668 16064
rect 14708 16024 14709 16064
rect 14667 16015 14709 16024
rect 16299 16064 16341 16073
rect 16299 16024 16300 16064
rect 16340 16024 16341 16064
rect 16299 16015 16341 16024
rect 20331 16064 20373 16073
rect 20331 16024 20332 16064
rect 20372 16024 20373 16064
rect 20331 16015 20373 16024
rect 24250 16064 24308 16065
rect 24250 16024 24259 16064
rect 24299 16024 24308 16064
rect 24250 16023 24308 16024
rect 25882 16064 25940 16065
rect 25882 16024 25891 16064
rect 25931 16024 25940 16064
rect 25882 16023 25940 16024
rect 26266 16064 26324 16065
rect 26266 16024 26275 16064
rect 26315 16024 26324 16064
rect 26266 16023 26324 16024
rect 26859 16064 26901 16073
rect 26859 16024 26860 16064
rect 26900 16024 26901 16064
rect 26859 16015 26901 16024
rect 28107 16064 28149 16073
rect 28107 16024 28108 16064
rect 28148 16024 28149 16064
rect 28107 16015 28149 16024
rect 576 15896 31392 15920
rect 576 15856 4352 15896
rect 4720 15856 12126 15896
rect 12494 15856 19900 15896
rect 20268 15856 27674 15896
rect 28042 15856 31392 15896
rect 576 15832 31392 15856
rect 2955 15728 2997 15737
rect 2955 15688 2956 15728
rect 2996 15688 2997 15728
rect 2955 15679 2997 15688
rect 4587 15728 4629 15737
rect 4587 15688 4588 15728
rect 4628 15688 4629 15728
rect 4587 15679 4629 15688
rect 6315 15728 6357 15737
rect 6315 15688 6316 15728
rect 6356 15688 6357 15728
rect 6315 15679 6357 15688
rect 8427 15728 8469 15737
rect 8427 15688 8428 15728
rect 8468 15688 8469 15728
rect 8427 15679 8469 15688
rect 9274 15728 9332 15729
rect 9274 15688 9283 15728
rect 9323 15688 9332 15728
rect 9274 15687 9332 15688
rect 11674 15728 11732 15729
rect 11674 15688 11683 15728
rect 11723 15688 11732 15728
rect 11674 15687 11732 15688
rect 13419 15728 13461 15737
rect 13419 15688 13420 15728
rect 13460 15688 13461 15728
rect 13419 15679 13461 15688
rect 15051 15728 15093 15737
rect 15051 15688 15052 15728
rect 15092 15688 15093 15728
rect 15051 15679 15093 15688
rect 15610 15728 15668 15729
rect 15610 15688 15619 15728
rect 15659 15688 15668 15728
rect 15610 15687 15668 15688
rect 16090 15728 16148 15729
rect 16090 15688 16099 15728
rect 16139 15688 16148 15728
rect 16090 15687 16148 15688
rect 16762 15728 16820 15729
rect 16762 15688 16771 15728
rect 16811 15688 16820 15728
rect 16762 15687 16820 15688
rect 17355 15728 17397 15737
rect 17355 15688 17356 15728
rect 17396 15688 17397 15728
rect 17355 15679 17397 15688
rect 18130 15728 18188 15729
rect 18130 15688 18139 15728
rect 18179 15688 18188 15728
rect 18130 15687 18188 15688
rect 18586 15728 18644 15729
rect 18586 15688 18595 15728
rect 18635 15688 18644 15728
rect 18586 15687 18644 15688
rect 21099 15728 21141 15737
rect 21099 15688 21100 15728
rect 21140 15688 21141 15728
rect 21099 15679 21141 15688
rect 23691 15728 23733 15737
rect 23691 15688 23692 15728
rect 23732 15688 23733 15728
rect 23691 15679 23733 15688
rect 24699 15728 24741 15737
rect 24699 15688 24700 15728
rect 24740 15688 24741 15728
rect 24699 15679 24741 15688
rect 24939 15728 24981 15737
rect 24939 15688 24940 15728
rect 24980 15688 24981 15728
rect 24939 15679 24981 15688
rect 26859 15728 26901 15737
rect 26859 15688 26860 15728
rect 26900 15688 26901 15728
rect 26859 15679 26901 15688
rect 27226 15728 27284 15729
rect 27226 15688 27235 15728
rect 27275 15688 27284 15728
rect 27226 15687 27284 15688
rect 3370 15644 3428 15645
rect 3370 15604 3379 15644
rect 3419 15604 3428 15644
rect 3370 15603 3428 15604
rect 8907 15644 8949 15653
rect 8907 15604 8908 15644
rect 8948 15604 8949 15644
rect 8907 15595 8949 15604
rect 12747 15644 12789 15653
rect 12747 15604 12748 15644
rect 12788 15604 12789 15644
rect 12747 15595 12789 15604
rect 14650 15644 14708 15645
rect 14650 15604 14659 15644
rect 14699 15604 14708 15644
rect 14650 15603 14708 15604
rect 14845 15644 14887 15653
rect 17152 15644 17194 15653
rect 14845 15604 14846 15644
rect 14886 15604 14887 15644
rect 14845 15595 14887 15604
rect 16578 15635 16624 15644
rect 16578 15595 16579 15635
rect 16619 15595 16624 15635
rect 17152 15604 17153 15644
rect 17193 15604 17194 15644
rect 17152 15595 17194 15604
rect 27339 15644 27381 15653
rect 27339 15604 27340 15644
rect 27380 15604 27381 15644
rect 27339 15595 27381 15604
rect 31258 15644 31316 15645
rect 31258 15604 31267 15644
rect 31307 15604 31316 15644
rect 31258 15603 31316 15604
rect 16578 15586 16624 15595
rect 1803 15560 1845 15569
rect 1803 15520 1804 15560
rect 1844 15520 1845 15560
rect 1803 15511 1845 15520
rect 2091 15560 2133 15569
rect 2091 15520 2092 15560
rect 2132 15520 2133 15560
rect 2091 15511 2133 15520
rect 2749 15560 2791 15569
rect 3535 15560 3593 15561
rect 2749 15520 2750 15560
rect 2790 15520 2791 15560
rect 2749 15511 2791 15520
rect 3051 15551 3093 15560
rect 3051 15511 3052 15551
rect 3092 15511 3093 15551
rect 3535 15520 3544 15560
rect 3584 15520 3593 15560
rect 3535 15519 3593 15520
rect 3819 15560 3861 15569
rect 3819 15520 3820 15560
rect 3860 15520 3861 15560
rect 3819 15511 3861 15520
rect 4186 15560 4244 15561
rect 4186 15520 4195 15560
rect 4235 15520 4244 15560
rect 5451 15560 5493 15569
rect 4186 15519 4244 15520
rect 4293 15533 4351 15534
rect 3051 15502 3093 15511
rect 4293 15493 4302 15533
rect 4342 15493 4351 15533
rect 5451 15520 5452 15560
rect 5492 15520 5493 15560
rect 5451 15511 5493 15520
rect 5700 15560 5758 15561
rect 5700 15520 5709 15560
rect 5749 15520 5758 15560
rect 6154 15560 6212 15561
rect 5700 15519 5758 15520
rect 5863 15518 5905 15527
rect 6154 15520 6163 15560
rect 6203 15520 6212 15560
rect 6154 15519 6212 15520
rect 6411 15560 6453 15569
rect 6411 15520 6412 15560
rect 6452 15520 6453 15560
rect 4293 15492 4351 15493
rect 3675 15476 3717 15485
rect 3675 15436 3676 15476
rect 3716 15436 3717 15476
rect 3675 15427 3717 15436
rect 5595 15476 5637 15485
rect 5595 15436 5596 15476
rect 5636 15436 5637 15476
rect 5863 15478 5864 15518
rect 5904 15478 5905 15518
rect 6411 15511 6453 15520
rect 6530 15560 6572 15569
rect 6530 15520 6531 15560
rect 6571 15520 6572 15560
rect 6530 15511 6572 15520
rect 6640 15560 6698 15561
rect 6640 15520 6649 15560
rect 6689 15520 6698 15560
rect 6640 15519 6698 15520
rect 7323 15560 7365 15569
rect 7323 15520 7324 15560
rect 7364 15520 7365 15560
rect 7786 15560 7844 15561
rect 7323 15511 7365 15520
rect 7467 15518 7509 15527
rect 7786 15520 7795 15560
rect 7835 15520 7844 15560
rect 7786 15519 7844 15520
rect 8139 15560 8181 15569
rect 8139 15520 8140 15560
rect 8180 15520 8181 15560
rect 8811 15560 8853 15569
rect 5863 15469 5905 15478
rect 6027 15476 6069 15485
rect 5595 15427 5637 15436
rect 6027 15436 6028 15476
rect 6068 15436 6069 15476
rect 7467 15478 7468 15518
rect 7508 15478 7509 15518
rect 8139 15511 8181 15520
rect 8273 15528 8331 15529
rect 8273 15488 8282 15528
rect 8322 15488 8331 15528
rect 8811 15520 8812 15560
rect 8852 15520 8853 15560
rect 8811 15511 8853 15520
rect 9003 15560 9045 15569
rect 9003 15520 9004 15560
rect 9044 15520 9045 15560
rect 9003 15511 9045 15520
rect 9254 15560 9312 15561
rect 9254 15520 9263 15560
rect 9303 15520 9312 15560
rect 9254 15519 9312 15520
rect 9370 15560 9428 15561
rect 9370 15520 9379 15560
rect 9419 15520 9428 15560
rect 9370 15519 9428 15520
rect 9514 15560 9572 15561
rect 9514 15520 9523 15560
rect 9563 15520 9572 15560
rect 9514 15519 9572 15520
rect 9658 15560 9716 15561
rect 9658 15520 9667 15560
rect 9707 15520 9716 15560
rect 10059 15560 10101 15569
rect 9658 15519 9716 15520
rect 9771 15549 9813 15558
rect 9771 15509 9772 15549
rect 9812 15509 9813 15549
rect 10059 15520 10060 15560
rect 10100 15520 10101 15560
rect 10059 15511 10101 15520
rect 10251 15560 10293 15569
rect 10251 15520 10252 15560
rect 10292 15520 10293 15560
rect 10251 15511 10293 15520
rect 11350 15560 11392 15569
rect 11350 15520 11351 15560
rect 11391 15520 11392 15560
rect 11350 15511 11392 15520
rect 11595 15560 11637 15569
rect 11595 15520 11596 15560
rect 11636 15520 11637 15560
rect 11595 15511 11637 15520
rect 12132 15560 12190 15561
rect 12132 15520 12141 15560
rect 12181 15520 12190 15560
rect 12132 15519 12190 15520
rect 12302 15560 12344 15569
rect 12302 15520 12303 15560
rect 12343 15520 12344 15560
rect 12302 15511 12344 15520
rect 12843 15560 12885 15569
rect 12843 15520 12844 15560
rect 12884 15520 12885 15560
rect 12586 15518 12644 15519
rect 9771 15500 9813 15509
rect 8273 15487 8331 15488
rect 7467 15469 7509 15478
rect 7659 15476 7701 15485
rect 6027 15427 6069 15436
rect 7659 15436 7660 15476
rect 7700 15436 7701 15476
rect 7659 15427 7701 15436
rect 11482 15476 11540 15477
rect 11482 15436 11491 15476
rect 11531 15436 11540 15476
rect 11482 15435 11540 15436
rect 12459 15476 12501 15485
rect 12586 15478 12595 15518
rect 12635 15478 12644 15518
rect 12843 15511 12885 15520
rect 13072 15560 13130 15561
rect 13072 15520 13081 15560
rect 13121 15520 13130 15560
rect 13072 15519 13130 15520
rect 13210 15560 13268 15561
rect 13210 15520 13219 15560
rect 13259 15520 13268 15560
rect 13210 15519 13268 15520
rect 13323 15560 13365 15569
rect 13323 15520 13324 15560
rect 13364 15520 13365 15560
rect 13323 15511 13365 15520
rect 13526 15560 13568 15569
rect 13526 15520 13527 15560
rect 13567 15520 13568 15560
rect 13526 15511 13568 15520
rect 14326 15560 14368 15569
rect 14326 15520 14327 15560
rect 14367 15520 14368 15560
rect 14326 15511 14368 15520
rect 14571 15560 14613 15569
rect 15286 15560 15328 15569
rect 14571 15520 14572 15560
rect 14612 15520 14613 15560
rect 14571 15511 14613 15520
rect 15147 15551 15189 15560
rect 15147 15511 15148 15551
rect 15188 15511 15189 15551
rect 15286 15520 15287 15560
rect 15327 15520 15328 15560
rect 15286 15511 15328 15520
rect 15531 15560 15573 15569
rect 15531 15520 15532 15560
rect 15572 15520 15573 15560
rect 15531 15511 15573 15520
rect 15766 15560 15808 15569
rect 15766 15520 15767 15560
rect 15807 15520 15808 15560
rect 15766 15511 15808 15520
rect 16011 15560 16053 15569
rect 16011 15520 16012 15560
rect 16052 15520 16053 15560
rect 16011 15511 16053 15520
rect 16282 15560 16340 15561
rect 16669 15560 16711 15569
rect 16282 15520 16291 15560
rect 16331 15520 16340 15560
rect 16282 15519 16340 15520
rect 16395 15551 16437 15560
rect 16395 15511 16396 15551
rect 16436 15511 16437 15551
rect 16669 15520 16670 15560
rect 16710 15520 16711 15560
rect 16669 15511 16711 15520
rect 16843 15560 16901 15561
rect 18010 15560 18068 15561
rect 16843 15520 16852 15560
rect 16892 15520 16901 15560
rect 16843 15519 16901 15520
rect 17451 15551 17493 15560
rect 17451 15511 17452 15551
rect 17492 15511 17493 15551
rect 15147 15502 15189 15511
rect 16395 15502 16437 15511
rect 17451 15502 17493 15511
rect 17919 15551 17961 15560
rect 17919 15511 17920 15551
rect 17960 15511 17961 15551
rect 18010 15520 18019 15560
rect 18059 15520 18068 15560
rect 18010 15519 18068 15520
rect 18274 15560 18332 15561
rect 18274 15520 18283 15560
rect 18323 15520 18332 15560
rect 18274 15519 18332 15520
rect 18507 15560 18549 15569
rect 18507 15520 18508 15560
rect 18548 15520 18549 15560
rect 18507 15511 18549 15520
rect 19642 15560 19700 15561
rect 19642 15520 19651 15560
rect 19691 15520 19700 15560
rect 19642 15519 19700 15520
rect 20890 15560 20948 15561
rect 20890 15520 20899 15560
rect 20939 15520 20948 15560
rect 20890 15519 20948 15520
rect 23595 15560 23637 15569
rect 23595 15520 23596 15560
rect 23636 15520 23637 15560
rect 23595 15511 23637 15520
rect 23787 15560 23829 15569
rect 23787 15520 23788 15560
rect 23828 15520 23829 15560
rect 23787 15511 23829 15520
rect 24034 15560 24092 15561
rect 24034 15520 24043 15560
rect 24083 15520 24092 15560
rect 24034 15519 24092 15520
rect 24267 15560 24309 15569
rect 24267 15520 24268 15560
rect 24308 15520 24309 15560
rect 24267 15511 24309 15520
rect 24843 15560 24885 15569
rect 24843 15520 24844 15560
rect 24884 15520 24885 15560
rect 24843 15511 24885 15520
rect 24987 15560 25029 15569
rect 24987 15520 24988 15560
rect 25028 15520 25029 15560
rect 24987 15511 25029 15520
rect 25366 15560 25408 15569
rect 25611 15560 25653 15569
rect 25366 15520 25367 15560
rect 25407 15520 25408 15560
rect 25366 15511 25408 15520
rect 25506 15551 25552 15560
rect 25506 15511 25507 15551
rect 25547 15511 25552 15551
rect 25611 15520 25612 15560
rect 25652 15520 25653 15560
rect 25611 15511 25653 15520
rect 26043 15560 26085 15569
rect 26043 15520 26044 15560
rect 26084 15520 26085 15560
rect 26043 15511 26085 15520
rect 26222 15560 26264 15569
rect 26222 15520 26223 15560
rect 26263 15520 26264 15560
rect 26222 15511 26264 15520
rect 26500 15560 26542 15569
rect 26500 15520 26501 15560
rect 26541 15520 26542 15560
rect 26500 15511 26542 15520
rect 26656 15560 26698 15569
rect 27130 15560 27188 15561
rect 26656 15520 26657 15560
rect 26697 15520 26698 15560
rect 26656 15511 26698 15520
rect 26955 15551 26997 15560
rect 26955 15511 26956 15551
rect 26996 15511 26997 15551
rect 27130 15520 27139 15560
rect 27179 15520 27188 15560
rect 27130 15519 27188 15520
rect 27446 15560 27488 15569
rect 27446 15520 27447 15560
rect 27487 15520 27488 15560
rect 27446 15511 27488 15520
rect 28779 15560 28821 15569
rect 28779 15520 28780 15560
rect 28820 15520 28821 15560
rect 28779 15511 28821 15520
rect 30874 15560 30932 15561
rect 30874 15520 30883 15560
rect 30923 15520 30932 15560
rect 30874 15519 30932 15520
rect 17919 15502 17961 15511
rect 25506 15502 25552 15511
rect 26955 15502 26997 15511
rect 12586 15477 12644 15478
rect 14458 15476 14516 15477
rect 12459 15436 12460 15476
rect 12500 15436 12501 15476
rect 12459 15427 12501 15436
rect 12978 15467 13024 15476
rect 12978 15427 12979 15467
rect 13019 15427 13024 15467
rect 14458 15436 14467 15476
rect 14507 15436 14516 15476
rect 14458 15435 14516 15436
rect 15418 15476 15476 15477
rect 15418 15436 15427 15476
rect 15467 15436 15476 15476
rect 15418 15435 15476 15436
rect 15898 15476 15956 15477
rect 15898 15436 15907 15476
rect 15947 15436 15956 15476
rect 15898 15435 15956 15436
rect 18394 15476 18452 15477
rect 18394 15436 18403 15476
rect 18443 15436 18452 15476
rect 18394 15435 18452 15436
rect 24154 15476 24212 15477
rect 24154 15436 24163 15476
rect 24203 15436 24212 15476
rect 24154 15435 24212 15436
rect 24363 15476 24405 15485
rect 24363 15436 24364 15476
rect 24404 15436 24405 15476
rect 24363 15427 24405 15436
rect 26379 15476 26421 15485
rect 26379 15436 26380 15476
rect 26420 15436 26421 15476
rect 26379 15427 26421 15436
rect 12978 15418 13024 15427
rect 1803 15392 1845 15401
rect 1803 15352 1804 15392
rect 1844 15352 1845 15392
rect 1803 15343 1845 15352
rect 5931 15392 5973 15401
rect 5931 15352 5932 15392
rect 5972 15352 5973 15392
rect 5931 15343 5973 15352
rect 7563 15392 7605 15401
rect 7563 15352 7564 15392
rect 7604 15352 7605 15392
rect 7563 15343 7605 15352
rect 10042 15392 10100 15393
rect 10042 15352 10051 15392
rect 10091 15352 10100 15392
rect 10042 15351 10100 15352
rect 12363 15392 12405 15401
rect 12363 15352 12364 15392
rect 12404 15352 12405 15392
rect 12363 15343 12405 15352
rect 26283 15392 26325 15401
rect 26283 15352 26284 15392
rect 26324 15352 26325 15392
rect 26283 15343 26325 15352
rect 2746 15308 2804 15309
rect 2746 15268 2755 15308
rect 2795 15268 2804 15308
rect 2746 15267 2804 15268
rect 14842 15308 14900 15309
rect 14842 15268 14851 15308
rect 14891 15268 14900 15308
rect 14842 15267 14900 15268
rect 17146 15308 17204 15309
rect 17146 15268 17155 15308
rect 17195 15268 17204 15308
rect 17146 15267 17204 15268
rect 17626 15308 17684 15309
rect 17626 15268 17635 15308
rect 17675 15268 17684 15308
rect 17626 15267 17684 15268
rect 20043 15308 20085 15317
rect 20043 15268 20044 15308
rect 20084 15268 20085 15308
rect 20043 15259 20085 15268
rect 21291 15308 21333 15317
rect 21291 15268 21292 15308
rect 21332 15268 21333 15308
rect 21291 15259 21333 15268
rect 25323 15308 25365 15317
rect 25323 15268 25324 15308
rect 25364 15268 25365 15308
rect 25323 15259 25365 15268
rect 26650 15308 26708 15309
rect 26650 15268 26659 15308
rect 26699 15268 26708 15308
rect 26650 15267 26708 15268
rect 28107 15308 28149 15317
rect 28107 15268 28108 15308
rect 28148 15268 28149 15308
rect 28107 15259 28149 15268
rect 28971 15308 29013 15317
rect 28971 15268 28972 15308
rect 29012 15268 29013 15308
rect 28971 15259 29013 15268
rect 29355 15308 29397 15317
rect 29355 15268 29356 15308
rect 29396 15268 29397 15308
rect 29355 15259 29397 15268
rect 576 15140 31392 15164
rect 576 15100 3112 15140
rect 3480 15100 10886 15140
rect 11254 15100 18660 15140
rect 19028 15100 26434 15140
rect 26802 15100 31392 15140
rect 576 15076 31392 15100
rect 3994 14972 4052 14973
rect 3994 14932 4003 14972
rect 4043 14932 4052 14972
rect 3994 14931 4052 14932
rect 7162 14972 7220 14973
rect 7162 14932 7171 14972
rect 7211 14932 7220 14972
rect 7162 14931 7220 14932
rect 7947 14972 7989 14981
rect 7947 14932 7948 14972
rect 7988 14932 7989 14972
rect 7947 14923 7989 14932
rect 9850 14972 9908 14973
rect 9850 14932 9859 14972
rect 9899 14932 9908 14972
rect 9850 14931 9908 14932
rect 11499 14972 11541 14981
rect 11499 14932 11500 14972
rect 11540 14932 11541 14972
rect 11499 14923 11541 14932
rect 12987 14972 13029 14981
rect 12987 14932 12988 14972
rect 13028 14932 13029 14972
rect 12987 14923 13029 14932
rect 18010 14972 18068 14973
rect 18010 14932 18019 14972
rect 18059 14932 18068 14972
rect 18010 14931 18068 14932
rect 18490 14972 18548 14973
rect 18490 14932 18499 14972
rect 18539 14932 18548 14972
rect 18490 14931 18548 14932
rect 24267 14972 24309 14981
rect 24267 14932 24268 14972
rect 24308 14932 24309 14972
rect 24267 14923 24309 14932
rect 24939 14972 24981 14981
rect 24939 14932 24940 14972
rect 24980 14932 24981 14972
rect 24939 14923 24981 14932
rect 27994 14972 28052 14973
rect 27994 14932 28003 14972
rect 28043 14932 28052 14972
rect 27994 14931 28052 14932
rect 28378 14972 28436 14973
rect 28378 14932 28387 14972
rect 28427 14932 28436 14972
rect 28378 14931 28436 14932
rect 4875 14888 4917 14897
rect 4875 14848 4876 14888
rect 4916 14848 4917 14888
rect 4875 14839 4917 14848
rect 6682 14888 6740 14889
rect 10347 14888 10389 14897
rect 6682 14848 6691 14888
rect 6731 14848 6740 14888
rect 6682 14847 6740 14848
rect 6939 14879 6981 14888
rect 6939 14839 6940 14879
rect 6980 14839 6981 14879
rect 10347 14848 10348 14888
rect 10388 14848 10389 14888
rect 10347 14839 10389 14848
rect 20043 14888 20085 14897
rect 20043 14848 20044 14888
rect 20084 14848 20085 14888
rect 20043 14839 20085 14848
rect 26667 14888 26709 14897
rect 26667 14848 26668 14888
rect 26708 14848 26709 14888
rect 26667 14839 26709 14848
rect 27226 14888 27284 14889
rect 27226 14848 27235 14888
rect 27275 14848 27284 14888
rect 27226 14847 27284 14848
rect 30699 14888 30741 14897
rect 30699 14848 30700 14888
rect 30740 14848 30741 14888
rect 30699 14839 30741 14848
rect 31083 14888 31125 14897
rect 31083 14848 31084 14888
rect 31124 14848 31125 14888
rect 31083 14839 31125 14848
rect 6939 14830 6981 14839
rect 4514 14804 4556 14813
rect 4514 14764 4515 14804
rect 4555 14764 4556 14804
rect 4514 14755 4556 14764
rect 10251 14804 10293 14813
rect 10251 14764 10252 14804
rect 10292 14764 10293 14804
rect 10251 14755 10293 14764
rect 11050 14804 11108 14805
rect 11050 14764 11059 14804
rect 11099 14764 11108 14804
rect 11050 14763 11108 14764
rect 14114 14804 14156 14813
rect 14114 14764 14115 14804
rect 14155 14764 14156 14804
rect 14114 14755 14156 14764
rect 14786 14804 14828 14813
rect 14786 14764 14787 14804
rect 14827 14764 14828 14804
rect 14786 14755 14828 14764
rect 16610 14804 16652 14813
rect 16610 14764 16611 14804
rect 16651 14764 16652 14804
rect 16610 14755 16652 14764
rect 21483 14804 21525 14813
rect 21483 14764 21484 14804
rect 21524 14764 21525 14804
rect 21483 14755 21525 14764
rect 24651 14804 24693 14813
rect 24651 14764 24652 14804
rect 24692 14764 24693 14804
rect 24211 14753 24253 14762
rect 24651 14755 24693 14764
rect 25323 14804 25365 14813
rect 28401 14804 28443 14813
rect 25323 14764 25324 14804
rect 25364 14764 25365 14804
rect 25323 14755 25365 14764
rect 25554 14795 25600 14804
rect 25554 14755 25555 14795
rect 25595 14755 25600 14795
rect 28401 14764 28402 14804
rect 28442 14764 28443 14804
rect 28401 14755 28443 14764
rect 6187 14731 6229 14740
rect 1227 14720 1269 14729
rect 1227 14680 1228 14720
rect 1268 14680 1269 14720
rect 1227 14671 1269 14680
rect 1371 14720 1413 14729
rect 1371 14680 1372 14720
rect 1412 14680 1413 14720
rect 1371 14671 1413 14680
rect 2379 14720 2421 14729
rect 3051 14720 3093 14729
rect 2379 14680 2380 14720
rect 2420 14680 2421 14720
rect 2379 14671 2421 14680
rect 2754 14711 2800 14720
rect 2754 14671 2755 14711
rect 2795 14671 2800 14711
rect 3051 14680 3052 14720
rect 3092 14680 3093 14720
rect 3051 14671 3093 14680
rect 3706 14720 3764 14721
rect 3706 14680 3715 14720
rect 3755 14680 3764 14720
rect 3706 14679 3764 14680
rect 3819 14720 3861 14729
rect 3819 14680 3820 14720
rect 3860 14680 3861 14720
rect 3819 14671 3861 14680
rect 4404 14720 4446 14729
rect 4404 14680 4405 14720
rect 4445 14680 4446 14720
rect 4404 14671 4446 14680
rect 4635 14720 4677 14729
rect 4635 14680 4636 14720
rect 4676 14680 4677 14720
rect 4971 14720 5013 14729
rect 4635 14671 4677 14680
rect 4774 14701 4816 14710
rect 2754 14662 2800 14671
rect 4774 14661 4775 14701
rect 4815 14661 4816 14701
rect 4971 14680 4972 14720
rect 5012 14680 5013 14720
rect 4971 14671 5013 14680
rect 5755 14720 5813 14721
rect 5755 14680 5764 14720
rect 5804 14680 5813 14720
rect 5755 14679 5813 14680
rect 5936 14720 5978 14729
rect 5936 14680 5937 14720
rect 5977 14680 5978 14720
rect 5936 14671 5978 14680
rect 6058 14720 6116 14721
rect 6058 14680 6067 14720
rect 6107 14680 6116 14720
rect 6187 14691 6188 14731
rect 6228 14691 6229 14731
rect 7387 14731 7429 14740
rect 6187 14682 6229 14691
rect 6298 14720 6356 14721
rect 6058 14679 6116 14680
rect 6298 14680 6307 14720
rect 6347 14680 6356 14720
rect 6298 14679 6356 14680
rect 6507 14720 6549 14729
rect 6507 14680 6508 14720
rect 6548 14680 6549 14720
rect 6507 14671 6549 14680
rect 6682 14720 6740 14721
rect 6682 14680 6691 14720
rect 6731 14680 6740 14720
rect 6682 14679 6740 14680
rect 6970 14720 7028 14721
rect 6970 14680 6979 14720
rect 7019 14680 7028 14720
rect 7387 14691 7388 14731
rect 7428 14691 7429 14731
rect 7387 14682 7429 14691
rect 7546 14720 7604 14721
rect 6970 14679 7028 14680
rect 7546 14680 7555 14720
rect 7595 14680 7604 14720
rect 7546 14679 7604 14680
rect 7671 14720 7713 14729
rect 7671 14680 7672 14720
rect 7712 14680 7713 14720
rect 7671 14671 7713 14680
rect 7834 14720 7892 14721
rect 7834 14680 7843 14720
rect 7883 14680 7892 14720
rect 7834 14679 7892 14680
rect 7956 14720 8014 14721
rect 7956 14680 7965 14720
rect 8005 14680 8014 14720
rect 7956 14679 8014 14680
rect 8139 14720 8181 14729
rect 8139 14680 8140 14720
rect 8180 14680 8181 14720
rect 8139 14671 8181 14680
rect 8331 14720 8373 14729
rect 8331 14680 8332 14720
rect 8372 14680 8373 14720
rect 8331 14671 8373 14680
rect 9178 14720 9236 14721
rect 9178 14680 9187 14720
rect 9227 14680 9236 14720
rect 9178 14679 9236 14680
rect 9483 14720 9525 14729
rect 9483 14680 9484 14720
rect 9524 14680 9525 14720
rect 9483 14671 9525 14680
rect 9675 14720 9717 14729
rect 9675 14680 9676 14720
rect 9716 14680 9717 14720
rect 9675 14671 9717 14680
rect 9850 14720 9908 14721
rect 9850 14680 9859 14720
rect 9899 14680 9908 14720
rect 9850 14679 9908 14680
rect 10107 14720 10149 14729
rect 10107 14680 10108 14720
rect 10148 14680 10149 14720
rect 10107 14671 10149 14680
rect 10422 14720 10464 14729
rect 10422 14680 10423 14720
rect 10463 14680 10464 14720
rect 10422 14671 10464 14680
rect 10570 14720 10628 14721
rect 10570 14680 10579 14720
rect 10619 14680 10628 14720
rect 10570 14679 10628 14680
rect 11215 14720 11273 14721
rect 11215 14680 11224 14720
rect 11264 14680 11273 14720
rect 11215 14679 11273 14680
rect 11403 14720 11445 14729
rect 11403 14680 11404 14720
rect 11444 14680 11445 14720
rect 11403 14671 11445 14680
rect 12843 14720 12885 14729
rect 12843 14680 12844 14720
rect 12884 14680 12885 14720
rect 12843 14671 12885 14680
rect 13114 14720 13172 14721
rect 13114 14680 13123 14720
rect 13163 14680 13172 14720
rect 13114 14679 13172 14680
rect 13232 14720 13290 14721
rect 13232 14680 13241 14720
rect 13281 14680 13290 14720
rect 13232 14679 13290 14680
rect 13398 14720 13456 14721
rect 13398 14680 13407 14720
rect 13447 14680 13456 14720
rect 13398 14679 13456 14680
rect 13498 14720 13556 14721
rect 13498 14680 13507 14720
rect 13547 14680 13556 14720
rect 13498 14679 13556 14680
rect 13675 14720 13733 14721
rect 13675 14680 13684 14720
rect 13724 14680 13733 14720
rect 13675 14679 13733 14680
rect 13995 14720 14037 14729
rect 13995 14680 13996 14720
rect 14036 14680 14037 14720
rect 13995 14671 14037 14680
rect 14224 14720 14282 14721
rect 14224 14680 14233 14720
rect 14273 14680 14282 14720
rect 14224 14679 14282 14680
rect 14667 14720 14709 14729
rect 14667 14680 14668 14720
rect 14708 14680 14709 14720
rect 14667 14671 14709 14680
rect 14896 14720 14954 14721
rect 14896 14680 14905 14720
rect 14945 14680 14954 14720
rect 14896 14679 14954 14680
rect 16207 14720 16265 14721
rect 16207 14680 16216 14720
rect 16256 14680 16265 14720
rect 16207 14679 16265 14680
rect 16491 14720 16533 14729
rect 16491 14680 16492 14720
rect 16532 14680 16533 14720
rect 16491 14671 16533 14680
rect 16708 14720 16750 14729
rect 16708 14680 16709 14720
rect 16749 14680 16750 14720
rect 16708 14671 16750 14680
rect 16875 14720 16917 14729
rect 16875 14680 16876 14720
rect 16916 14680 16917 14720
rect 16875 14671 16917 14680
rect 17067 14720 17109 14729
rect 17067 14680 17068 14720
rect 17108 14680 17109 14720
rect 17067 14671 17109 14680
rect 17234 14720 17292 14721
rect 17234 14680 17243 14720
rect 17283 14680 17292 14720
rect 17234 14679 17292 14680
rect 17360 14720 17418 14721
rect 17634 14720 17692 14721
rect 17360 14680 17369 14720
rect 17409 14680 17418 14720
rect 17360 14679 17418 14680
rect 17538 14711 17584 14720
rect 17538 14671 17539 14711
rect 17579 14671 17584 14711
rect 17634 14680 17643 14720
rect 17683 14680 17692 14720
rect 17634 14679 17692 14680
rect 17803 14720 17861 14721
rect 17803 14680 17812 14720
rect 17852 14680 17861 14720
rect 17803 14679 17861 14680
rect 18313 14720 18371 14721
rect 18313 14680 18322 14720
rect 18362 14680 18371 14720
rect 18313 14679 18371 14680
rect 18699 14720 18741 14729
rect 18699 14680 18700 14720
rect 18740 14680 18741 14720
rect 18699 14671 18741 14680
rect 18793 14720 18851 14721
rect 18793 14680 18802 14720
rect 18842 14680 18851 14720
rect 18793 14679 18851 14680
rect 19371 14720 19413 14729
rect 19371 14680 19372 14720
rect 19412 14680 19413 14720
rect 19371 14671 19413 14680
rect 19618 14720 19676 14721
rect 19618 14680 19627 14720
rect 19667 14680 19676 14720
rect 19618 14679 19676 14680
rect 19738 14720 19796 14721
rect 19738 14680 19747 14720
rect 19787 14680 19796 14720
rect 19738 14679 19796 14680
rect 20986 14720 21044 14721
rect 20986 14680 20995 14720
rect 21035 14680 21044 14720
rect 20986 14679 21044 14680
rect 21099 14720 21141 14729
rect 21099 14680 21100 14720
rect 21140 14680 21141 14720
rect 21099 14671 21141 14680
rect 21579 14720 21621 14729
rect 21579 14680 21580 14720
rect 21620 14680 21621 14720
rect 21579 14671 21621 14680
rect 22051 14720 22109 14721
rect 22051 14680 22060 14720
rect 22100 14680 22109 14720
rect 22051 14679 22109 14680
rect 22539 14720 22597 14721
rect 22539 14680 22548 14720
rect 22588 14680 22597 14720
rect 22539 14679 22597 14680
rect 23307 14720 23349 14729
rect 23307 14680 23308 14720
rect 23348 14680 23349 14720
rect 23307 14671 23349 14680
rect 23979 14720 24021 14729
rect 23979 14680 23980 14720
rect 24020 14680 24021 14720
rect 23979 14671 24021 14680
rect 24093 14720 24151 14721
rect 24093 14680 24102 14720
rect 24142 14680 24151 14720
rect 24211 14713 24212 14753
rect 24252 14713 24253 14753
rect 25554 14746 25600 14755
rect 24211 14704 24253 14713
rect 24555 14720 24597 14729
rect 24093 14679 24151 14680
rect 24555 14680 24556 14720
rect 24596 14680 24597 14720
rect 24555 14671 24597 14680
rect 24768 14720 24826 14721
rect 24768 14680 24777 14720
rect 24817 14680 24826 14720
rect 24768 14679 24826 14680
rect 24886 14720 24944 14721
rect 24886 14680 24895 14720
rect 24935 14680 24944 14720
rect 24886 14679 24944 14680
rect 25419 14720 25461 14729
rect 25419 14680 25420 14720
rect 25460 14680 25461 14720
rect 25419 14671 25461 14680
rect 25650 14720 25692 14729
rect 25650 14680 25651 14720
rect 25691 14680 25692 14720
rect 25650 14671 25692 14680
rect 26710 14720 26752 14729
rect 26955 14720 26997 14729
rect 26710 14680 26711 14720
rect 26751 14680 26752 14720
rect 26710 14671 26752 14680
rect 26850 14711 26896 14720
rect 26850 14671 26851 14711
rect 26891 14671 26896 14711
rect 26955 14680 26956 14720
rect 26996 14680 26997 14720
rect 26955 14671 26997 14680
rect 27243 14720 27285 14729
rect 27243 14680 27244 14720
rect 27284 14680 27285 14720
rect 27243 14671 27285 14680
rect 27435 14720 27477 14729
rect 27435 14680 27436 14720
rect 27476 14680 27477 14720
rect 27435 14671 27477 14680
rect 27819 14720 27861 14729
rect 27819 14680 27820 14720
rect 27860 14680 27861 14720
rect 27819 14671 27861 14680
rect 27994 14720 28052 14721
rect 27994 14680 28003 14720
rect 28043 14680 28052 14720
rect 27994 14679 28052 14680
rect 28491 14720 28533 14729
rect 28491 14680 28492 14720
rect 28532 14680 28533 14720
rect 28491 14671 28533 14680
rect 28971 14720 29013 14729
rect 28971 14680 28972 14720
rect 29012 14680 29013 14720
rect 28971 14671 29013 14680
rect 30507 14720 30549 14729
rect 30507 14680 30508 14720
rect 30548 14680 30549 14720
rect 30507 14671 30549 14680
rect 30699 14720 30741 14729
rect 30699 14680 30700 14720
rect 30740 14680 30741 14720
rect 30699 14671 30741 14680
rect 30891 14720 30933 14729
rect 30891 14680 30892 14720
rect 30932 14680 30933 14720
rect 30891 14671 30933 14680
rect 17538 14662 17584 14671
rect 26850 14662 26896 14671
rect 4774 14652 4816 14661
rect 1018 14636 1076 14637
rect 1018 14596 1027 14636
rect 1067 14596 1076 14636
rect 1018 14595 1076 14596
rect 2554 14636 2612 14637
rect 2554 14596 2563 14636
rect 2603 14596 2612 14636
rect 2554 14595 2612 14596
rect 2859 14636 2901 14645
rect 2859 14596 2860 14636
rect 2900 14596 2901 14636
rect 2859 14587 2901 14596
rect 4299 14636 4341 14645
rect 4299 14596 4300 14636
rect 4340 14596 4341 14636
rect 4299 14587 4341 14596
rect 8235 14636 8277 14645
rect 8235 14596 8236 14636
rect 8276 14596 8277 14636
rect 8235 14587 8277 14596
rect 9003 14636 9045 14645
rect 9003 14596 9004 14636
rect 9044 14596 9045 14636
rect 9003 14587 9045 14596
rect 18016 14636 18058 14645
rect 18016 14596 18017 14636
rect 18057 14596 18058 14636
rect 18016 14587 18058 14596
rect 18493 14636 18535 14645
rect 18493 14596 18494 14636
rect 18534 14596 18535 14636
rect 18493 14587 18535 14596
rect 29643 14636 29685 14645
rect 29643 14596 29644 14636
rect 29684 14596 29685 14636
rect 29643 14587 29685 14596
rect 1323 14552 1365 14561
rect 1323 14512 1324 14552
rect 1364 14512 1365 14552
rect 1323 14503 1365 14512
rect 1707 14552 1749 14561
rect 1707 14512 1708 14552
rect 1748 14512 1749 14552
rect 1707 14503 1749 14512
rect 2955 14552 2997 14561
rect 2955 14512 2956 14552
rect 2996 14512 2997 14552
rect 2955 14503 2997 14512
rect 5818 14552 5876 14553
rect 5818 14512 5827 14552
rect 5867 14512 5876 14552
rect 5818 14511 5876 14512
rect 13498 14552 13556 14553
rect 13498 14512 13507 14552
rect 13547 14512 13556 14552
rect 13498 14511 13556 14512
rect 13899 14552 13941 14561
rect 13899 14512 13900 14552
rect 13940 14512 13941 14552
rect 13899 14503 13941 14512
rect 14571 14552 14613 14561
rect 14571 14512 14572 14552
rect 14612 14512 14613 14552
rect 14571 14503 14613 14512
rect 16042 14552 16100 14553
rect 16042 14512 16051 14552
rect 16091 14512 16100 14552
rect 16042 14511 16100 14512
rect 16395 14552 16437 14561
rect 16395 14512 16396 14552
rect 16436 14512 16437 14552
rect 16395 14503 16437 14512
rect 16971 14552 17013 14561
rect 16971 14512 16972 14552
rect 17012 14512 17013 14552
rect 16971 14503 17013 14512
rect 17722 14552 17780 14553
rect 17722 14512 17731 14552
rect 17771 14512 17780 14552
rect 17722 14511 17780 14512
rect 18219 14552 18261 14561
rect 18219 14512 18220 14552
rect 18260 14512 18261 14552
rect 18219 14503 18261 14512
rect 22731 14552 22773 14561
rect 22731 14512 22732 14552
rect 22772 14512 22773 14552
rect 22731 14503 22773 14512
rect 23451 14552 23493 14561
rect 23451 14512 23452 14552
rect 23492 14512 23493 14552
rect 23451 14503 23493 14512
rect 29835 14552 29877 14561
rect 29835 14512 29836 14552
rect 29876 14512 29877 14552
rect 29835 14503 29877 14512
rect 576 14384 31392 14408
rect 576 14344 4352 14384
rect 4720 14344 12126 14384
rect 12494 14344 19900 14384
rect 20268 14344 27674 14384
rect 28042 14344 31392 14384
rect 576 14320 31392 14344
rect 1786 14216 1844 14217
rect 1786 14176 1795 14216
rect 1835 14176 1844 14216
rect 1786 14175 1844 14176
rect 1899 14216 1941 14225
rect 1899 14176 1900 14216
rect 1940 14176 1941 14216
rect 1899 14167 1941 14176
rect 3706 14216 3764 14217
rect 3706 14176 3715 14216
rect 3755 14176 3764 14216
rect 3706 14175 3764 14176
rect 4875 14216 4917 14225
rect 4875 14176 4876 14216
rect 4916 14176 4917 14216
rect 4875 14167 4917 14176
rect 5626 14216 5684 14217
rect 5626 14176 5635 14216
rect 5675 14176 5684 14216
rect 5626 14175 5684 14176
rect 9963 14216 10005 14225
rect 9963 14176 9964 14216
rect 10004 14176 10005 14216
rect 9963 14167 10005 14176
rect 10635 14216 10677 14225
rect 10635 14176 10636 14216
rect 10676 14176 10677 14216
rect 10635 14167 10677 14176
rect 14187 14216 14229 14225
rect 14187 14176 14188 14216
rect 14228 14176 14229 14216
rect 14187 14167 14229 14176
rect 14746 14216 14804 14217
rect 14746 14176 14755 14216
rect 14795 14176 14804 14216
rect 14746 14175 14804 14176
rect 15339 14216 15381 14225
rect 15339 14176 15340 14216
rect 15380 14176 15381 14216
rect 15339 14167 15381 14176
rect 16474 14216 16532 14217
rect 16474 14176 16483 14216
rect 16523 14176 16532 14216
rect 16474 14175 16532 14176
rect 19371 14216 19413 14225
rect 19371 14176 19372 14216
rect 19412 14176 19413 14216
rect 19371 14167 19413 14176
rect 22234 14216 22292 14217
rect 22234 14176 22243 14216
rect 22283 14176 22292 14216
rect 22234 14175 22292 14176
rect 24939 14216 24981 14225
rect 24939 14176 24940 14216
rect 24980 14176 24981 14216
rect 24939 14167 24981 14176
rect 25611 14216 25653 14225
rect 25611 14176 25612 14216
rect 25652 14176 25653 14216
rect 25611 14167 25653 14176
rect 26091 14216 26133 14225
rect 26091 14176 26092 14216
rect 26132 14176 26133 14216
rect 26091 14167 26133 14176
rect 26955 14216 26997 14225
rect 26955 14176 26956 14216
rect 26996 14176 26997 14216
rect 26955 14167 26997 14176
rect 27243 14216 27285 14225
rect 27243 14176 27244 14216
rect 27284 14176 27285 14216
rect 27243 14167 27285 14176
rect 1114 14132 1172 14133
rect 1114 14092 1123 14132
rect 1163 14092 1172 14132
rect 1114 14091 1172 14092
rect 2009 14132 2051 14141
rect 2009 14092 2010 14132
rect 2050 14092 2051 14132
rect 2009 14083 2051 14092
rect 2650 14132 2708 14133
rect 2650 14092 2659 14132
rect 2699 14092 2708 14132
rect 2650 14091 2708 14092
rect 14859 14132 14901 14141
rect 14859 14092 14860 14132
rect 14900 14092 14901 14132
rect 14859 14083 14901 14092
rect 15446 14132 15488 14141
rect 20139 14132 20181 14141
rect 15446 14092 15447 14132
rect 15487 14092 15488 14132
rect 15446 14083 15488 14092
rect 16770 14123 16816 14132
rect 16770 14083 16771 14123
rect 16811 14083 16816 14123
rect 20139 14092 20140 14132
rect 20180 14092 20181 14132
rect 20139 14083 20181 14092
rect 21483 14132 21525 14141
rect 21483 14092 21484 14132
rect 21524 14092 21525 14132
rect 21483 14083 21525 14092
rect 23883 14132 23925 14141
rect 23883 14092 23884 14132
rect 23924 14092 23925 14132
rect 23883 14083 23925 14092
rect 24555 14132 24597 14141
rect 24555 14092 24556 14132
rect 24596 14092 24597 14132
rect 24555 14083 24597 14092
rect 24662 14132 24704 14141
rect 24662 14092 24663 14132
rect 24703 14092 24704 14132
rect 24662 14083 24704 14092
rect 16770 14074 16816 14083
rect 1035 14048 1077 14057
rect 1035 14008 1036 14048
rect 1076 14008 1077 14048
rect 1035 13999 1077 14008
rect 1207 14048 1249 14057
rect 1207 14008 1208 14048
rect 1248 14008 1249 14048
rect 1207 13999 1249 14008
rect 1323 14048 1365 14057
rect 1323 14008 1324 14048
rect 1364 14008 1365 14048
rect 1323 13999 1365 14008
rect 1690 14048 1748 14049
rect 1690 14008 1699 14048
rect 1739 14008 1748 14048
rect 1690 14007 1748 14008
rect 2314 14048 2372 14049
rect 2314 14008 2323 14048
rect 2363 14008 2372 14048
rect 2314 14007 2372 14008
rect 2509 14048 2567 14049
rect 2509 14008 2518 14048
rect 2558 14008 2567 14048
rect 2509 14007 2567 14008
rect 3291 14048 3333 14057
rect 3291 14008 3292 14048
rect 3332 14008 3333 14048
rect 3291 13999 3333 14008
rect 3521 14048 3579 14049
rect 3521 14008 3530 14048
rect 3570 14008 3579 14048
rect 3521 14007 3579 14008
rect 3723 14048 3765 14057
rect 3723 14008 3724 14048
rect 3764 14008 3765 14048
rect 3723 13999 3765 14008
rect 4971 14048 5013 14057
rect 4971 14008 4972 14048
rect 5012 14008 5013 14048
rect 4971 13999 5013 14008
rect 5090 14048 5132 14057
rect 5090 14008 5091 14048
rect 5131 14008 5132 14048
rect 5090 13999 5132 14008
rect 5200 14048 5258 14049
rect 5200 14008 5209 14048
rect 5249 14008 5258 14048
rect 5200 14007 5258 14008
rect 5547 14048 5589 14057
rect 5547 14008 5548 14048
rect 5588 14008 5589 14048
rect 5547 13999 5589 14008
rect 5931 14048 5973 14057
rect 5931 14008 5932 14048
rect 5972 14008 5973 14048
rect 5931 13999 5973 14008
rect 6160 14048 6218 14049
rect 6160 14008 6169 14048
rect 6209 14008 6218 14048
rect 6160 14007 6218 14008
rect 6315 14048 6357 14057
rect 6315 14008 6316 14048
rect 6356 14008 6357 14048
rect 6315 13999 6357 14008
rect 6507 14048 6549 14057
rect 6507 14008 6508 14048
rect 6548 14008 6549 14048
rect 6507 13999 6549 14008
rect 10059 14048 10101 14057
rect 10059 14008 10060 14048
rect 10100 14008 10101 14048
rect 10059 13999 10101 14008
rect 10288 14048 10346 14049
rect 10288 14008 10297 14048
rect 10337 14008 10346 14048
rect 10288 14007 10346 14008
rect 10731 14048 10773 14057
rect 10731 14008 10732 14048
rect 10772 14008 10773 14048
rect 10731 13999 10773 14008
rect 10960 14048 11018 14049
rect 10960 14008 10969 14048
rect 11009 14008 11018 14048
rect 10960 14007 11018 14008
rect 11194 14048 11252 14049
rect 11194 14008 11203 14048
rect 11243 14008 11252 14048
rect 11194 14007 11252 14008
rect 12651 14048 12693 14057
rect 12651 14008 12652 14048
rect 12692 14008 12693 14048
rect 12651 13999 12693 14008
rect 12843 14048 12885 14057
rect 12843 14008 12844 14048
rect 12884 14008 12885 14048
rect 12843 13999 12885 14008
rect 14230 14048 14272 14057
rect 14475 14048 14517 14057
rect 14230 14008 14231 14048
rect 14271 14008 14272 14048
rect 14230 13999 14272 14008
rect 14370 14039 14416 14048
rect 14370 13999 14371 14039
rect 14411 13999 14416 14039
rect 14475 14008 14476 14048
rect 14516 14008 14517 14048
rect 14475 13999 14517 14008
rect 14656 14048 14698 14057
rect 15130 14048 15188 14049
rect 14656 14008 14657 14048
rect 14697 14008 14698 14048
rect 14656 13999 14698 14008
rect 14955 14039 14997 14048
rect 14955 13999 14956 14039
rect 14996 13999 14997 14039
rect 15130 14008 15139 14048
rect 15179 14008 15188 14048
rect 15130 14007 15188 14008
rect 15243 14048 15285 14057
rect 15243 14008 15244 14048
rect 15284 14008 15285 14048
rect 15243 13999 15285 14008
rect 16474 14048 16532 14049
rect 16858 14048 16916 14049
rect 16474 14008 16483 14048
rect 16523 14008 16532 14048
rect 16474 14007 16532 14008
rect 16587 14039 16629 14048
rect 16587 13999 16588 14039
rect 16628 13999 16629 14039
rect 16858 14008 16867 14048
rect 16907 14008 16916 14048
rect 16858 14007 16916 14008
rect 17035 14048 17093 14049
rect 17035 14008 17044 14048
rect 17084 14008 17093 14048
rect 17035 14007 17093 14008
rect 18891 14048 18933 14057
rect 18891 14008 18892 14048
rect 18932 14008 18933 14048
rect 18891 13999 18933 14008
rect 19083 14048 19125 14057
rect 19083 14008 19084 14048
rect 19124 14008 19125 14048
rect 19083 13999 19125 14008
rect 19275 14048 19317 14057
rect 19275 14008 19276 14048
rect 19316 14008 19317 14048
rect 19275 13999 19317 14008
rect 19467 14048 19509 14057
rect 19467 14008 19468 14048
rect 19508 14008 19509 14048
rect 19467 13999 19509 14008
rect 20240 14048 20298 14049
rect 20240 14008 20249 14048
rect 20289 14008 20298 14048
rect 20240 14007 20298 14008
rect 20523 14048 20565 14057
rect 20523 14008 20524 14048
rect 20564 14008 20565 14048
rect 20523 13999 20565 14008
rect 20811 14048 20853 14057
rect 20811 14008 20812 14048
rect 20852 14008 20853 14048
rect 20811 13999 20853 14008
rect 20986 14048 21044 14049
rect 20986 14008 20995 14048
rect 21035 14008 21044 14048
rect 20986 14007 21044 14008
rect 21147 14048 21189 14057
rect 21147 14008 21148 14048
rect 21188 14008 21189 14048
rect 21147 13999 21189 14008
rect 21584 14048 21642 14049
rect 21584 14008 21593 14048
rect 21633 14008 21642 14048
rect 21584 14007 21642 14008
rect 21867 14048 21909 14057
rect 21867 14008 21868 14048
rect 21908 14008 21909 14048
rect 21867 13999 21909 14008
rect 22522 14048 22580 14049
rect 22522 14008 22531 14048
rect 22571 14008 22580 14048
rect 22522 14007 22580 14008
rect 23268 14048 23326 14049
rect 23268 14008 23277 14048
rect 23317 14008 23326 14048
rect 23722 14048 23780 14049
rect 23268 14007 23326 14008
rect 23431 14006 23473 14015
rect 23722 14008 23731 14048
rect 23771 14008 23780 14048
rect 23722 14007 23780 14008
rect 23979 14048 24021 14057
rect 23979 14008 23980 14048
rect 24020 14008 24021 14048
rect 14370 13990 14416 13999
rect 14955 13990 14997 13999
rect 16587 13990 16629 13999
rect 5835 13964 5877 13973
rect 5835 13924 5836 13964
rect 5876 13924 5877 13964
rect 5835 13915 5877 13924
rect 6050 13964 6092 13973
rect 6050 13924 6051 13964
rect 6091 13924 6092 13964
rect 6050 13915 6092 13924
rect 10178 13964 10220 13973
rect 10178 13924 10179 13964
rect 10219 13924 10220 13964
rect 10178 13915 10220 13924
rect 10850 13964 10892 13973
rect 10850 13924 10851 13964
rect 10891 13924 10892 13964
rect 10850 13915 10892 13924
rect 11691 13964 11733 13973
rect 11691 13924 11692 13964
rect 11732 13924 11733 13964
rect 11691 13915 11733 13924
rect 12939 13964 12981 13973
rect 23431 13966 23432 14006
rect 23472 13966 23473 14006
rect 23979 13999 24021 14008
rect 24196 14048 24238 14057
rect 24196 14008 24197 14048
rect 24237 14008 24238 14048
rect 24196 13999 24238 14008
rect 24346 14048 24404 14049
rect 24346 14008 24355 14048
rect 24395 14008 24404 14048
rect 24346 14007 24404 14008
rect 24459 14048 24501 14057
rect 24459 14008 24460 14048
rect 24500 14008 24501 14048
rect 24459 13999 24501 14008
rect 24939 14048 24981 14057
rect 24939 14008 24940 14048
rect 24980 14008 24981 14048
rect 24939 13999 24981 14008
rect 25136 14048 25178 14057
rect 25136 14008 25137 14048
rect 25177 14008 25178 14048
rect 25136 13999 25178 14008
rect 25275 14048 25317 14057
rect 25275 14008 25276 14048
rect 25316 14008 25317 14048
rect 25803 14048 25845 14057
rect 25275 13999 25317 14008
rect 25457 14024 25515 14025
rect 25457 13984 25466 14024
rect 25506 13984 25515 14024
rect 25803 14008 25804 14048
rect 25844 14008 25845 14048
rect 25803 13999 25845 14008
rect 26134 14048 26192 14049
rect 26134 14008 26143 14048
rect 26183 14008 26192 14048
rect 26134 14007 26192 14008
rect 26667 14048 26709 14057
rect 26667 14008 26668 14048
rect 26708 14008 26709 14048
rect 26667 13999 26709 14008
rect 26998 14048 27056 14049
rect 27623 14048 27681 14049
rect 26998 14008 27007 14048
rect 27047 14008 27056 14048
rect 27522 14039 27568 14048
rect 26998 14007 27056 14008
rect 27404 14027 27446 14036
rect 25457 13983 25515 13984
rect 27404 13987 27405 14027
rect 27445 13987 27446 14027
rect 27522 13999 27523 14039
rect 27563 13999 27568 14039
rect 27623 14008 27632 14048
rect 27672 14008 27681 14048
rect 27623 14007 27681 14008
rect 28203 14048 28245 14057
rect 28203 14008 28204 14048
rect 28244 14008 28245 14048
rect 28203 13999 28245 14008
rect 28587 14048 28629 14057
rect 28587 14008 28588 14048
rect 28628 14008 28629 14048
rect 28587 13999 28629 14008
rect 30874 14048 30932 14049
rect 30874 14008 30883 14048
rect 30923 14008 30932 14048
rect 30874 14007 30932 14008
rect 27522 13990 27568 13999
rect 27404 13978 27446 13987
rect 12939 13924 12940 13964
rect 12980 13924 12981 13964
rect 12939 13915 12981 13924
rect 22138 13964 22196 13965
rect 22138 13924 22147 13964
rect 22187 13924 22196 13964
rect 22138 13923 22196 13924
rect 22714 13964 22772 13965
rect 22714 13924 22723 13964
rect 22763 13924 22772 13964
rect 23431 13957 23473 13966
rect 23595 13964 23637 13973
rect 22714 13923 22772 13924
rect 23595 13924 23596 13964
rect 23636 13924 23637 13964
rect 23595 13915 23637 13924
rect 24098 13964 24140 13973
rect 24098 13924 24099 13964
rect 24139 13924 24140 13964
rect 24098 13915 24140 13924
rect 26025 13964 26067 13973
rect 26025 13924 26026 13964
rect 26066 13924 26067 13964
rect 26025 13915 26067 13924
rect 26889 13964 26931 13973
rect 26889 13924 26890 13964
rect 26930 13924 26931 13964
rect 26889 13915 26931 13924
rect 29338 13964 29396 13965
rect 29338 13924 29347 13964
rect 29387 13924 29396 13964
rect 29338 13923 29396 13924
rect 31258 13964 31316 13965
rect 31258 13924 31267 13964
rect 31307 13924 31316 13964
rect 31258 13923 31316 13924
rect 843 13880 885 13889
rect 843 13840 844 13880
rect 884 13840 885 13880
rect 843 13831 885 13840
rect 6315 13880 6357 13889
rect 6315 13840 6316 13880
rect 6356 13840 6357 13880
rect 6315 13831 6357 13840
rect 11174 13880 11216 13889
rect 11174 13840 11175 13880
rect 11215 13840 11216 13880
rect 11174 13831 11216 13840
rect 20986 13880 21044 13881
rect 20986 13840 20995 13880
rect 21035 13840 21044 13880
rect 20986 13839 21044 13840
rect 23499 13880 23541 13889
rect 23499 13840 23500 13880
rect 23540 13840 23541 13880
rect 23499 13831 23541 13840
rect 26763 13880 26805 13889
rect 26763 13840 26764 13880
rect 26804 13840 26805 13880
rect 26763 13831 26805 13840
rect 28827 13880 28869 13889
rect 28827 13840 28828 13880
rect 28868 13840 28869 13880
rect 28827 13831 28869 13840
rect 5355 13796 5397 13805
rect 5355 13756 5356 13796
rect 5396 13756 5397 13796
rect 5355 13747 5397 13756
rect 11386 13796 11444 13797
rect 11386 13756 11395 13796
rect 11435 13756 11444 13796
rect 11386 13755 11444 13756
rect 11931 13796 11973 13805
rect 11931 13756 11932 13796
rect 11972 13756 11973 13796
rect 11931 13747 11973 13756
rect 18891 13796 18933 13805
rect 18891 13756 18892 13796
rect 18932 13756 18933 13796
rect 18891 13747 18933 13756
rect 19851 13796 19893 13805
rect 19851 13756 19852 13796
rect 19892 13756 19893 13796
rect 19851 13747 19893 13756
rect 25899 13796 25941 13805
rect 25899 13756 25900 13796
rect 25940 13756 25941 13796
rect 25899 13747 25941 13756
rect 28971 13796 29013 13805
rect 28971 13756 28972 13796
rect 29012 13756 29013 13796
rect 28971 13747 29013 13756
rect 576 13628 31392 13652
rect 576 13588 3112 13628
rect 3480 13588 10886 13628
rect 11254 13588 18660 13628
rect 19028 13588 26434 13628
rect 26802 13588 31392 13628
rect 576 13564 31392 13588
rect 2955 13460 2997 13469
rect 2955 13420 2956 13460
rect 2996 13420 2997 13460
rect 2955 13411 2997 13420
rect 3819 13460 3861 13469
rect 3819 13420 3820 13460
rect 3860 13420 3861 13460
rect 3819 13411 3861 13420
rect 14475 13460 14517 13469
rect 14475 13420 14476 13460
rect 14516 13420 14517 13460
rect 14475 13411 14517 13420
rect 16474 13460 16532 13461
rect 16474 13420 16483 13460
rect 16523 13420 16532 13460
rect 16474 13419 16532 13420
rect 17050 13460 17108 13461
rect 17050 13420 17059 13460
rect 17099 13420 17108 13460
rect 17050 13419 17108 13420
rect 20715 13460 20757 13469
rect 20715 13420 20716 13460
rect 20756 13420 20757 13460
rect 20715 13411 20757 13420
rect 21963 13460 22005 13469
rect 21963 13420 21964 13460
rect 22004 13420 22005 13460
rect 21963 13411 22005 13420
rect 23674 13460 23732 13461
rect 23674 13420 23683 13460
rect 23723 13420 23732 13460
rect 23674 13419 23732 13420
rect 24459 13460 24501 13469
rect 24459 13420 24460 13460
rect 24500 13420 24501 13460
rect 24459 13411 24501 13420
rect 25803 13460 25845 13469
rect 25803 13420 25804 13460
rect 25844 13420 25845 13460
rect 25803 13411 25845 13420
rect 26955 13460 26997 13469
rect 26955 13420 26956 13460
rect 26996 13420 26997 13460
rect 26955 13411 26997 13420
rect 5547 13376 5589 13385
rect 5547 13336 5548 13376
rect 5588 13336 5589 13376
rect 5547 13327 5589 13336
rect 6123 13376 6165 13385
rect 6123 13336 6124 13376
rect 6164 13336 6165 13376
rect 6123 13327 6165 13336
rect 6795 13376 6837 13385
rect 6795 13336 6796 13376
rect 6836 13336 6837 13376
rect 6795 13327 6837 13336
rect 8811 13376 8853 13385
rect 8811 13336 8812 13376
rect 8852 13336 8853 13376
rect 8811 13327 8853 13336
rect 9274 13376 9332 13377
rect 9274 13336 9283 13376
rect 9323 13336 9332 13376
rect 9274 13335 9332 13336
rect 10827 13376 10869 13385
rect 10827 13336 10828 13376
rect 10868 13336 10869 13376
rect 10827 13327 10869 13336
rect 13131 13376 13173 13385
rect 13131 13336 13132 13376
rect 13172 13336 13173 13376
rect 13131 13327 13173 13336
rect 13702 13376 13744 13385
rect 13702 13336 13703 13376
rect 13743 13336 13744 13376
rect 13702 13327 13744 13336
rect 15531 13376 15573 13385
rect 15531 13336 15532 13376
rect 15572 13336 15573 13376
rect 15531 13327 15573 13336
rect 19659 13376 19701 13385
rect 19659 13336 19660 13376
rect 19700 13336 19701 13376
rect 19659 13327 19701 13336
rect 27243 13376 27285 13385
rect 27243 13336 27244 13376
rect 27284 13336 27285 13376
rect 27243 13327 27285 13336
rect 29931 13376 29973 13385
rect 29931 13336 29932 13376
rect 29972 13336 29973 13376
rect 29931 13327 29973 13336
rect 651 13292 693 13301
rect 651 13252 652 13292
rect 692 13252 693 13292
rect 651 13243 693 13252
rect 2571 13292 2613 13301
rect 2571 13252 2572 13292
rect 2612 13252 2613 13292
rect 2571 13243 2613 13252
rect 4762 13292 4820 13293
rect 4762 13252 4771 13292
rect 4811 13252 4820 13292
rect 4762 13251 4820 13252
rect 4971 13292 5013 13301
rect 4971 13252 4972 13292
rect 5012 13252 5013 13292
rect 4971 13243 5013 13252
rect 5643 13292 5685 13301
rect 5643 13252 5644 13292
rect 5684 13252 5685 13292
rect 5643 13243 5685 13252
rect 6027 13292 6069 13301
rect 6027 13252 6028 13292
rect 6068 13252 6069 13292
rect 6027 13243 6069 13252
rect 6891 13292 6933 13301
rect 6891 13252 6892 13292
rect 6932 13252 6933 13292
rect 6891 13243 6933 13252
rect 8218 13292 8276 13293
rect 8218 13252 8227 13292
rect 8267 13252 8276 13292
rect 8218 13251 8276 13252
rect 8715 13292 8757 13301
rect 8715 13252 8716 13292
rect 8756 13252 8757 13292
rect 8715 13243 8757 13252
rect 10370 13292 10412 13301
rect 10370 13252 10371 13292
rect 10411 13252 10412 13292
rect 10370 13243 10412 13252
rect 10731 13292 10773 13301
rect 10731 13252 10732 13292
rect 10772 13252 10773 13292
rect 10731 13243 10773 13252
rect 12106 13292 12164 13293
rect 12106 13252 12115 13292
rect 12155 13252 12164 13292
rect 12106 13251 12164 13252
rect 12674 13292 12716 13301
rect 12674 13252 12675 13292
rect 12715 13252 12716 13292
rect 12674 13243 12716 13252
rect 13035 13292 13077 13301
rect 13035 13252 13036 13292
rect 13076 13252 13077 13292
rect 13805 13292 13847 13301
rect 13035 13243 13077 13252
rect 13611 13250 13653 13259
rect 7792 13219 7834 13228
rect 1018 13208 1076 13209
rect 1018 13168 1027 13208
rect 1067 13168 1076 13208
rect 1018 13167 1076 13168
rect 3610 13208 3668 13209
rect 3610 13168 3619 13208
rect 3659 13168 3668 13208
rect 3610 13167 3668 13168
rect 3723 13208 3765 13217
rect 3723 13168 3724 13208
rect 3764 13168 3765 13208
rect 3723 13159 3765 13168
rect 4642 13208 4700 13209
rect 4642 13168 4651 13208
rect 4691 13168 4700 13208
rect 4642 13167 4700 13168
rect 4875 13208 4917 13217
rect 4875 13168 4876 13208
rect 4916 13168 4917 13208
rect 4875 13159 4917 13168
rect 5486 13208 5528 13217
rect 5486 13168 5487 13208
rect 5527 13168 5528 13208
rect 5338 13166 5396 13167
rect 5338 13126 5347 13166
rect 5387 13126 5396 13166
rect 5486 13159 5528 13168
rect 5770 13208 5828 13209
rect 5770 13168 5779 13208
rect 5819 13168 5828 13208
rect 5770 13167 5828 13168
rect 5883 13208 5925 13217
rect 5883 13168 5884 13208
rect 5924 13168 5925 13208
rect 5883 13159 5925 13168
rect 6184 13208 6226 13217
rect 6184 13168 6185 13208
rect 6225 13168 6226 13208
rect 6184 13159 6226 13168
rect 6555 13208 6597 13217
rect 6555 13168 6556 13208
rect 6596 13168 6597 13208
rect 6298 13166 6356 13167
rect 5338 13125 5396 13126
rect 6298 13126 6307 13166
rect 6347 13126 6356 13166
rect 6555 13159 6597 13168
rect 6720 13208 6762 13217
rect 6720 13168 6721 13208
rect 6761 13168 6762 13208
rect 6720 13159 6762 13168
rect 7018 13208 7076 13209
rect 7018 13168 7027 13208
rect 7067 13168 7076 13208
rect 7018 13167 7076 13168
rect 7430 13208 7488 13209
rect 7430 13168 7439 13208
rect 7479 13168 7488 13208
rect 7430 13167 7488 13168
rect 7568 13208 7610 13217
rect 7568 13168 7569 13208
rect 7609 13168 7610 13208
rect 7568 13159 7610 13168
rect 7671 13208 7713 13217
rect 7671 13168 7672 13208
rect 7712 13168 7713 13208
rect 7792 13179 7793 13219
rect 7833 13179 7834 13219
rect 7792 13170 7834 13179
rect 7936 13208 7994 13209
rect 7671 13159 7713 13168
rect 7936 13168 7945 13208
rect 7985 13168 7994 13208
rect 7936 13167 7994 13168
rect 8086 13208 8128 13217
rect 8086 13168 8087 13208
rect 8127 13168 8128 13208
rect 8086 13159 8128 13168
rect 8331 13208 8373 13217
rect 8331 13168 8332 13208
rect 8372 13168 8373 13208
rect 9034 13208 9092 13209
rect 8331 13159 8373 13168
rect 8554 13166 8612 13167
rect 6298 13125 6356 13126
rect 8554 13126 8563 13166
rect 8603 13126 8612 13166
rect 8554 13125 8612 13126
rect 8879 13166 8921 13175
rect 9034 13168 9043 13208
rect 9083 13168 9092 13208
rect 9034 13167 9092 13168
rect 9291 13208 9333 13217
rect 9291 13168 9292 13208
rect 9332 13168 9333 13208
rect 8879 13126 8880 13166
rect 8920 13126 8921 13166
rect 9291 13159 9333 13168
rect 9483 13208 9525 13217
rect 9483 13168 9484 13208
rect 9524 13168 9525 13208
rect 9483 13159 9525 13168
rect 10251 13208 10293 13217
rect 10251 13168 10252 13208
rect 10292 13168 10293 13208
rect 10251 13159 10293 13168
rect 10468 13208 10510 13217
rect 10468 13168 10469 13208
rect 10509 13168 10510 13208
rect 10468 13159 10510 13168
rect 10587 13208 10629 13217
rect 10587 13168 10588 13208
rect 10628 13168 10629 13208
rect 10587 13159 10629 13168
rect 10902 13208 10944 13217
rect 10902 13168 10903 13208
rect 10943 13168 10944 13208
rect 10902 13159 10944 13168
rect 11042 13208 11084 13217
rect 11042 13168 11043 13208
rect 11083 13168 11084 13208
rect 11042 13159 11084 13168
rect 11307 13208 11349 13217
rect 11307 13168 11308 13208
rect 11348 13168 11349 13208
rect 11307 13159 11349 13168
rect 11595 13208 11637 13217
rect 11595 13168 11596 13208
rect 11636 13168 11637 13208
rect 11595 13159 11637 13168
rect 12271 13208 12329 13209
rect 12271 13168 12280 13208
rect 12320 13168 12329 13208
rect 12271 13167 12329 13168
rect 12555 13208 12597 13217
rect 12555 13168 12556 13208
rect 12596 13168 12597 13208
rect 12555 13159 12597 13168
rect 12772 13208 12814 13217
rect 12772 13168 12773 13208
rect 12813 13168 12814 13208
rect 12772 13159 12814 13168
rect 12891 13208 12933 13217
rect 12891 13168 12892 13208
rect 12932 13168 12933 13208
rect 12891 13159 12933 13168
rect 13192 13208 13234 13217
rect 13192 13168 13193 13208
rect 13233 13168 13234 13208
rect 13192 13159 13234 13168
rect 13467 13208 13509 13217
rect 13467 13168 13468 13208
rect 13508 13168 13509 13208
rect 13611 13210 13612 13250
rect 13652 13210 13653 13250
rect 13805 13252 13806 13292
rect 13846 13252 13847 13292
rect 13805 13243 13847 13252
rect 14859 13292 14901 13301
rect 14859 13252 14860 13292
rect 14900 13252 14901 13292
rect 14859 13243 14901 13252
rect 15627 13292 15669 13301
rect 15627 13252 15628 13292
rect 15668 13252 15669 13292
rect 15627 13243 15669 13252
rect 22658 13292 22700 13301
rect 22658 13252 22659 13292
rect 22699 13252 22700 13292
rect 22658 13243 22700 13252
rect 27108 13292 27150 13301
rect 27108 13252 27109 13292
rect 27149 13252 27150 13292
rect 27108 13243 27150 13252
rect 27675 13292 27717 13301
rect 27675 13252 27676 13292
rect 27716 13252 27717 13292
rect 27675 13243 27717 13252
rect 30795 13292 30837 13301
rect 30795 13252 30796 13292
rect 30836 13252 30837 13292
rect 30795 13243 30837 13252
rect 13611 13201 13653 13210
rect 14379 13208 14421 13217
rect 13306 13166 13364 13167
rect 8879 13117 8921 13126
rect 10155 13124 10197 13133
rect 10155 13084 10156 13124
rect 10196 13084 10197 13124
rect 10155 13075 10197 13084
rect 11403 13124 11445 13133
rect 11403 13084 11404 13124
rect 11444 13084 11445 13124
rect 11403 13075 11445 13084
rect 12459 13124 12501 13133
rect 13306 13126 13315 13166
rect 13355 13126 13364 13166
rect 13467 13159 13509 13168
rect 14379 13168 14380 13208
rect 14420 13168 14421 13208
rect 13930 13166 13988 13167
rect 13306 13125 13364 13126
rect 13930 13126 13939 13166
rect 13979 13126 13988 13166
rect 14379 13159 14421 13168
rect 14571 13208 14613 13217
rect 14571 13168 14572 13208
rect 14612 13168 14613 13208
rect 14571 13159 14613 13168
rect 14722 13208 14780 13209
rect 14722 13168 14731 13208
rect 14771 13168 14780 13208
rect 14722 13167 14780 13168
rect 15030 13208 15072 13217
rect 15030 13168 15031 13208
rect 15071 13168 15072 13208
rect 15030 13159 15072 13168
rect 15470 13208 15512 13217
rect 15470 13168 15471 13208
rect 15511 13168 15512 13208
rect 15130 13166 15188 13167
rect 13930 13125 13988 13126
rect 15130 13126 15139 13166
rect 15179 13126 15188 13166
rect 15130 13125 15188 13126
rect 15322 13166 15380 13167
rect 15322 13126 15331 13166
rect 15371 13126 15380 13166
rect 15470 13159 15512 13168
rect 15748 13208 15790 13217
rect 15748 13168 15749 13208
rect 15789 13168 15790 13208
rect 15748 13159 15790 13168
rect 16299 13208 16341 13217
rect 16299 13168 16300 13208
rect 16340 13168 16341 13208
rect 16299 13159 16341 13168
rect 16474 13208 16532 13209
rect 16474 13168 16483 13208
rect 16523 13168 16532 13208
rect 16474 13167 16532 13168
rect 16683 13208 16725 13217
rect 16683 13168 16684 13208
rect 16724 13168 16725 13208
rect 16683 13159 16725 13168
rect 16875 13208 16917 13217
rect 16875 13168 16876 13208
rect 16916 13168 16917 13208
rect 16875 13159 16917 13168
rect 17050 13208 17108 13209
rect 17050 13168 17059 13208
rect 17099 13168 17108 13208
rect 17050 13167 17108 13168
rect 17168 13208 17226 13209
rect 17168 13168 17177 13208
rect 17217 13168 17226 13208
rect 17168 13167 17226 13168
rect 17336 13208 17378 13217
rect 17336 13168 17337 13208
rect 17377 13168 17378 13208
rect 17336 13159 17378 13168
rect 17434 13208 17492 13209
rect 17434 13168 17443 13208
rect 17483 13168 17492 13208
rect 17434 13167 17492 13168
rect 17580 13208 17638 13209
rect 17580 13168 17589 13208
rect 17629 13168 17638 13208
rect 17580 13167 17638 13168
rect 17818 13208 17876 13209
rect 17818 13168 17827 13208
rect 17867 13168 17876 13208
rect 17818 13167 17876 13168
rect 17973 13208 18031 13209
rect 17973 13168 17982 13208
rect 18022 13168 18031 13208
rect 17973 13167 18031 13168
rect 18076 13208 18134 13209
rect 18076 13168 18085 13208
rect 18125 13168 18134 13208
rect 18076 13167 18134 13168
rect 18202 13208 18260 13209
rect 18202 13168 18211 13208
rect 18251 13168 18260 13208
rect 18202 13167 18260 13168
rect 18336 13208 18394 13209
rect 18336 13168 18345 13208
rect 18385 13168 18394 13208
rect 18336 13167 18394 13168
rect 18979 13208 19037 13209
rect 20331 13208 20373 13217
rect 18979 13168 18988 13208
rect 19028 13168 19037 13208
rect 18979 13167 19037 13168
rect 20043 13199 20085 13208
rect 20043 13159 20044 13199
rect 20084 13159 20085 13199
rect 20331 13168 20332 13208
rect 20372 13168 20373 13208
rect 20331 13159 20373 13168
rect 21003 13208 21045 13217
rect 21387 13208 21429 13217
rect 21003 13168 21004 13208
rect 21044 13168 21045 13208
rect 21003 13159 21045 13168
rect 21099 13199 21141 13208
rect 21099 13159 21100 13199
rect 21140 13159 21141 13199
rect 21387 13168 21388 13208
rect 21428 13168 21429 13208
rect 21387 13159 21429 13168
rect 21963 13208 22005 13217
rect 21963 13168 21964 13208
rect 22004 13168 22005 13208
rect 21963 13159 22005 13168
rect 22251 13208 22293 13217
rect 22251 13168 22252 13208
rect 22292 13168 22293 13208
rect 22251 13159 22293 13168
rect 22539 13208 22581 13217
rect 22539 13168 22540 13208
rect 22580 13168 22581 13208
rect 22539 13159 22581 13168
rect 22756 13208 22798 13217
rect 22756 13168 22757 13208
rect 22797 13168 22798 13208
rect 22756 13159 22798 13168
rect 23194 13208 23252 13209
rect 23194 13168 23203 13208
rect 23243 13168 23252 13208
rect 23194 13167 23252 13168
rect 23677 13208 23719 13217
rect 23677 13168 23678 13208
rect 23718 13168 23719 13208
rect 23677 13159 23719 13168
rect 23971 13208 24029 13209
rect 23971 13168 23980 13208
rect 24020 13168 24029 13208
rect 23971 13167 24029 13168
rect 24163 13208 24221 13209
rect 24163 13168 24172 13208
rect 24212 13168 24221 13208
rect 24163 13167 24221 13168
rect 24298 13208 24356 13209
rect 24298 13168 24307 13208
rect 24347 13168 24356 13208
rect 24298 13167 24356 13168
rect 24412 13208 24470 13209
rect 24412 13168 24421 13208
rect 24461 13168 24470 13208
rect 24412 13167 24470 13168
rect 25227 13208 25269 13217
rect 25227 13168 25228 13208
rect 25268 13168 25269 13208
rect 25227 13159 25269 13168
rect 25402 13208 25460 13209
rect 25402 13168 25411 13208
rect 25451 13168 25460 13208
rect 25402 13167 25460 13168
rect 25515 13208 25557 13217
rect 25515 13168 25516 13208
rect 25556 13168 25557 13208
rect 25515 13159 25557 13168
rect 25707 13208 25749 13217
rect 25707 13168 25708 13208
rect 25748 13168 25749 13208
rect 25707 13159 25749 13168
rect 25899 13208 25941 13217
rect 25899 13168 25900 13208
rect 25940 13168 25941 13208
rect 25899 13159 25941 13168
rect 27008 13208 27066 13209
rect 27008 13168 27017 13208
rect 27057 13168 27066 13208
rect 27008 13167 27066 13168
rect 27339 13208 27381 13217
rect 27339 13168 27340 13208
rect 27380 13168 27381 13208
rect 27339 13159 27381 13168
rect 27562 13208 27620 13209
rect 27562 13168 27571 13208
rect 27611 13168 27620 13208
rect 27562 13167 27620 13168
rect 28779 13208 28821 13217
rect 28779 13168 28780 13208
rect 28820 13168 28821 13208
rect 28779 13159 28821 13168
rect 28971 13208 29013 13217
rect 28971 13168 28972 13208
rect 29012 13168 29013 13208
rect 28971 13159 29013 13168
rect 30123 13208 30165 13217
rect 30123 13168 30124 13208
rect 30164 13168 30165 13208
rect 30123 13159 30165 13168
rect 20043 13150 20085 13159
rect 21099 13150 21141 13159
rect 15322 13125 15380 13126
rect 12459 13084 12460 13124
rect 12500 13084 12501 13124
rect 12459 13075 12501 13084
rect 16779 13124 16821 13133
rect 16779 13084 16780 13124
rect 16820 13084 16821 13124
rect 14938 13082 14996 13083
rect 7450 13040 7508 13041
rect 7450 13000 7459 13040
rect 7499 13000 7508 13040
rect 7450 12999 7508 13000
rect 8410 13040 8468 13041
rect 8410 13000 8419 13040
rect 8459 13000 8468 13040
rect 8410 12999 8468 13000
rect 9483 13040 9525 13049
rect 14938 13042 14947 13082
rect 14987 13042 14996 13082
rect 16779 13075 16821 13084
rect 18688 13124 18730 13133
rect 18688 13084 18689 13124
rect 18729 13084 18730 13124
rect 18688 13075 18730 13084
rect 19947 13124 19989 13133
rect 19947 13084 19948 13124
rect 19988 13084 19989 13124
rect 19947 13075 19989 13084
rect 22443 13124 22485 13133
rect 22443 13084 22444 13124
rect 22484 13084 22485 13124
rect 22443 13075 22485 13084
rect 23403 13124 23445 13133
rect 23403 13084 23404 13124
rect 23444 13084 23445 13124
rect 23403 13075 23445 13084
rect 23513 13124 23555 13133
rect 23513 13084 23514 13124
rect 23554 13084 23555 13124
rect 23513 13075 23555 13084
rect 25306 13124 25364 13125
rect 25306 13084 25315 13124
rect 25355 13084 25364 13124
rect 25306 13083 25364 13084
rect 28875 13124 28917 13133
rect 28875 13084 28876 13124
rect 28916 13084 28917 13124
rect 28875 13075 28917 13084
rect 14938 13041 14996 13042
rect 9483 13000 9484 13040
rect 9524 13000 9525 13040
rect 9483 12991 9525 13000
rect 18106 13040 18164 13041
rect 18106 13000 18115 13040
rect 18155 13000 18164 13040
rect 18106 12999 18164 13000
rect 18778 13040 18836 13041
rect 18778 13000 18787 13040
rect 18827 13000 18836 13040
rect 18778 12999 18836 13000
rect 18891 13040 18933 13049
rect 18891 13000 18892 13040
rect 18932 13000 18933 13040
rect 18891 12991 18933 13000
rect 23290 13040 23348 13041
rect 23290 13000 23299 13040
rect 23339 13000 23348 13040
rect 23290 12999 23348 13000
rect 23883 13040 23925 13049
rect 23883 13000 23884 13040
rect 23924 13000 23925 13040
rect 23883 12991 23925 13000
rect 30555 13040 30597 13049
rect 30555 13000 30556 13040
rect 30596 13000 30597 13040
rect 30555 12991 30597 13000
rect 576 12872 31392 12896
rect 576 12832 4352 12872
rect 4720 12832 12126 12872
rect 12494 12832 19900 12872
rect 20268 12832 27674 12872
rect 28042 12832 31392 12872
rect 576 12808 31392 12832
rect 3339 12704 3381 12713
rect 3339 12664 3340 12704
rect 3380 12664 3381 12704
rect 3339 12655 3381 12664
rect 4203 12704 4245 12713
rect 4203 12664 4204 12704
rect 4244 12664 4245 12704
rect 4203 12655 4245 12664
rect 4875 12704 4917 12713
rect 4875 12664 4876 12704
rect 4916 12664 4917 12704
rect 4875 12655 4917 12664
rect 5739 12704 5781 12713
rect 5739 12664 5740 12704
rect 5780 12664 5781 12704
rect 5739 12655 5781 12664
rect 6891 12704 6933 12713
rect 6891 12664 6892 12704
rect 6932 12664 6933 12704
rect 6891 12655 6933 12664
rect 7467 12704 7509 12713
rect 7467 12664 7468 12704
rect 7508 12664 7509 12704
rect 7467 12655 7509 12664
rect 9003 12704 9045 12713
rect 9003 12664 9004 12704
rect 9044 12664 9045 12704
rect 9003 12655 9045 12664
rect 11403 12704 11445 12713
rect 11403 12664 11404 12704
rect 11444 12664 11445 12704
rect 11403 12655 11445 12664
rect 13018 12704 13076 12705
rect 13018 12664 13027 12704
rect 13067 12664 13076 12704
rect 13018 12663 13076 12664
rect 14554 12704 14612 12705
rect 14554 12664 14563 12704
rect 14603 12664 14612 12704
rect 14554 12663 14612 12664
rect 14938 12704 14996 12705
rect 14938 12664 14947 12704
rect 14987 12664 14996 12704
rect 14938 12663 14996 12664
rect 17067 12704 17109 12713
rect 17067 12664 17068 12704
rect 17108 12664 17109 12704
rect 17067 12655 17109 12664
rect 19066 12704 19124 12705
rect 19066 12664 19075 12704
rect 19115 12664 19124 12704
rect 19066 12663 19124 12664
rect 22042 12704 22100 12705
rect 22042 12664 22051 12704
rect 22091 12664 22100 12704
rect 22042 12663 22100 12664
rect 23835 12704 23877 12713
rect 23835 12664 23836 12704
rect 23876 12664 23877 12704
rect 23835 12655 23877 12664
rect 24250 12704 24308 12705
rect 24250 12664 24259 12704
rect 24299 12664 24308 12704
rect 24250 12663 24308 12664
rect 25419 12704 25461 12713
rect 25419 12664 25420 12704
rect 25460 12664 25461 12704
rect 25419 12655 25461 12664
rect 25803 12704 25845 12713
rect 25803 12664 25804 12704
rect 25844 12664 25845 12704
rect 25803 12655 25845 12664
rect 26475 12704 26517 12713
rect 26475 12664 26476 12704
rect 26516 12664 26517 12704
rect 26475 12655 26517 12664
rect 26619 12704 26661 12713
rect 26619 12664 26620 12704
rect 26660 12664 26661 12704
rect 26619 12655 26661 12664
rect 26938 12704 26996 12705
rect 26938 12664 26947 12704
rect 26987 12664 26996 12704
rect 26938 12663 26996 12664
rect 27723 12704 27765 12713
rect 27723 12664 27724 12704
rect 27764 12664 27765 12704
rect 27723 12655 27765 12664
rect 28491 12704 28533 12713
rect 28491 12664 28492 12704
rect 28532 12664 28533 12704
rect 28491 12655 28533 12664
rect 23019 12620 23061 12629
rect 18479 12578 18521 12587
rect 1323 12536 1365 12545
rect 1323 12496 1324 12536
rect 1364 12496 1365 12536
rect 1323 12487 1365 12496
rect 1515 12536 1557 12545
rect 1515 12496 1516 12536
rect 1556 12496 1557 12536
rect 1515 12487 1557 12496
rect 2859 12536 2901 12545
rect 2859 12496 2860 12536
rect 2900 12496 2901 12536
rect 2859 12487 2901 12496
rect 3147 12536 3189 12545
rect 3147 12496 3148 12536
rect 3188 12496 3189 12536
rect 3147 12487 3189 12496
rect 4299 12536 4341 12545
rect 4299 12496 4300 12536
rect 4340 12496 4341 12536
rect 4299 12487 4341 12496
rect 4516 12536 4558 12545
rect 4516 12496 4517 12536
rect 4557 12496 4558 12536
rect 4516 12487 4558 12496
rect 4672 12536 4714 12545
rect 5835 12536 5877 12545
rect 4672 12496 4673 12536
rect 4713 12496 4714 12536
rect 4672 12487 4714 12496
rect 4971 12527 5013 12536
rect 4971 12487 4972 12527
rect 5012 12487 5013 12527
rect 5835 12496 5836 12536
rect 5876 12496 5877 12536
rect 5835 12487 5877 12496
rect 6052 12536 6094 12545
rect 6052 12496 6053 12536
rect 6093 12496 6094 12536
rect 6052 12487 6094 12496
rect 6987 12536 7029 12545
rect 6987 12496 6988 12536
rect 7028 12496 7029 12536
rect 7371 12536 7413 12545
rect 6987 12487 7029 12496
rect 7227 12494 7269 12503
rect 4971 12478 5013 12487
rect 4418 12452 4460 12461
rect 7106 12452 7148 12461
rect 4418 12412 4419 12452
rect 4459 12412 4460 12452
rect 4418 12403 4460 12412
rect 5970 12443 6016 12452
rect 5970 12403 5971 12443
rect 6011 12403 6016 12443
rect 7106 12412 7107 12452
rect 7147 12412 7148 12452
rect 7227 12454 7228 12494
rect 7268 12454 7269 12494
rect 7371 12496 7372 12536
rect 7412 12496 7413 12536
rect 7371 12487 7413 12496
rect 7562 12536 7604 12545
rect 7562 12496 7563 12536
rect 7603 12496 7604 12536
rect 7562 12487 7604 12496
rect 7755 12536 7797 12545
rect 7755 12496 7756 12536
rect 7796 12496 7797 12536
rect 7755 12487 7797 12496
rect 7952 12531 7994 12540
rect 7952 12491 7953 12531
rect 7993 12491 7994 12531
rect 8098 12536 8156 12537
rect 8098 12496 8107 12536
rect 8147 12496 8156 12536
rect 8098 12495 8156 12496
rect 8392 12536 8434 12545
rect 8392 12496 8393 12536
rect 8433 12496 8434 12536
rect 7952 12482 7994 12491
rect 8392 12487 8434 12496
rect 8546 12536 8588 12545
rect 8546 12496 8547 12536
rect 8587 12496 8588 12536
rect 8546 12487 8588 12496
rect 9099 12536 9141 12545
rect 9099 12496 9100 12536
rect 9140 12496 9141 12536
rect 9099 12487 9141 12496
rect 9328 12536 9386 12537
rect 9328 12496 9337 12536
rect 9377 12496 9386 12536
rect 9328 12495 9386 12496
rect 10491 12536 10533 12545
rect 10491 12496 10492 12536
rect 10532 12496 10533 12536
rect 10491 12487 10533 12496
rect 10656 12536 10698 12545
rect 10656 12496 10657 12536
rect 10697 12496 10698 12536
rect 10656 12487 10698 12496
rect 10954 12536 11012 12537
rect 10954 12496 10963 12536
rect 11003 12496 11012 12536
rect 10954 12495 11012 12496
rect 11115 12536 11157 12545
rect 11115 12496 11116 12536
rect 11156 12496 11157 12536
rect 12706 12536 12764 12537
rect 11115 12487 11157 12496
rect 11248 12504 11306 12505
rect 11248 12464 11257 12504
rect 11297 12464 11306 12504
rect 12706 12496 12715 12536
rect 12755 12496 12764 12536
rect 12706 12495 12764 12496
rect 12939 12536 12981 12545
rect 12939 12496 12940 12536
rect 12980 12496 12981 12536
rect 12939 12487 12981 12496
rect 13690 12536 13748 12537
rect 13690 12496 13699 12536
rect 13739 12496 13748 12536
rect 13690 12495 13748 12496
rect 14379 12536 14421 12545
rect 14379 12496 14380 12536
rect 14420 12496 14421 12536
rect 14379 12487 14421 12496
rect 14571 12536 14613 12545
rect 14571 12496 14572 12536
rect 14612 12496 14613 12536
rect 14571 12487 14613 12496
rect 14763 12536 14805 12545
rect 14763 12496 14764 12536
rect 14804 12496 14805 12536
rect 14763 12487 14805 12496
rect 14955 12536 14997 12545
rect 14955 12496 14956 12536
rect 14996 12496 14997 12536
rect 14955 12487 14997 12496
rect 16587 12536 16629 12545
rect 16587 12496 16588 12536
rect 16628 12496 16629 12536
rect 16587 12487 16629 12496
rect 16779 12536 16821 12545
rect 16779 12496 16780 12536
rect 16820 12496 16821 12536
rect 16779 12487 16821 12496
rect 16971 12536 17013 12545
rect 16971 12496 16972 12536
rect 17012 12496 17013 12536
rect 16971 12487 17013 12496
rect 17163 12536 17205 12545
rect 17163 12496 17164 12536
rect 17204 12496 17205 12536
rect 18479 12538 18480 12578
rect 18520 12538 18521 12578
rect 23019 12580 23020 12620
rect 23060 12580 23061 12620
rect 23019 12571 23061 12580
rect 18479 12529 18521 12538
rect 18626 12536 18668 12545
rect 17163 12487 17205 12496
rect 18171 12494 18213 12503
rect 11248 12463 11306 12464
rect 7227 12445 7269 12454
rect 8235 12452 8277 12461
rect 7106 12403 7148 12412
rect 8235 12412 8236 12452
rect 8276 12412 8277 12452
rect 8235 12403 8277 12412
rect 9218 12452 9260 12461
rect 9218 12412 9219 12452
rect 9259 12412 9260 12452
rect 9218 12403 9260 12412
rect 10827 12452 10869 12461
rect 18171 12454 18172 12494
rect 18212 12454 18213 12494
rect 18626 12496 18627 12536
rect 18667 12496 18668 12536
rect 18626 12487 18668 12496
rect 18754 12536 18812 12537
rect 18754 12496 18763 12536
rect 18803 12496 18812 12536
rect 18754 12495 18812 12496
rect 18987 12536 19029 12545
rect 18987 12496 18988 12536
rect 19028 12496 19029 12536
rect 18987 12487 19029 12496
rect 21099 12536 21141 12545
rect 21099 12496 21100 12536
rect 21140 12496 21141 12536
rect 21099 12487 21141 12496
rect 21200 12536 21258 12537
rect 21200 12496 21209 12536
rect 21249 12496 21258 12536
rect 21200 12495 21258 12496
rect 21483 12536 21525 12545
rect 21483 12496 21484 12536
rect 21524 12496 21525 12536
rect 21483 12487 21525 12496
rect 21867 12536 21909 12545
rect 21867 12496 21868 12536
rect 21908 12496 21909 12536
rect 21867 12487 21909 12496
rect 22059 12536 22101 12545
rect 22059 12496 22060 12536
rect 22100 12496 22101 12536
rect 22059 12487 22101 12496
rect 23115 12536 23157 12545
rect 23115 12496 23116 12536
rect 23156 12496 23157 12536
rect 23499 12536 23541 12545
rect 23115 12487 23157 12496
rect 23355 12494 23397 12503
rect 10827 12412 10828 12452
rect 10868 12412 10869 12452
rect 10827 12403 10869 12412
rect 12826 12452 12884 12453
rect 12826 12412 12835 12452
rect 12875 12412 12884 12452
rect 18171 12445 18213 12454
rect 18315 12452 18357 12461
rect 12826 12411 12884 12412
rect 18315 12412 18316 12452
rect 18356 12412 18357 12452
rect 18315 12403 18357 12412
rect 18874 12452 18932 12453
rect 18874 12412 18883 12452
rect 18923 12412 18932 12452
rect 18874 12411 18932 12412
rect 23234 12452 23276 12461
rect 23234 12412 23235 12452
rect 23275 12412 23276 12452
rect 23355 12454 23356 12494
rect 23396 12454 23397 12494
rect 23499 12496 23500 12536
rect 23540 12496 23541 12536
rect 23499 12487 23541 12496
rect 23691 12536 23733 12545
rect 23691 12496 23692 12536
rect 23732 12496 23733 12536
rect 23691 12487 23733 12496
rect 23979 12536 24021 12545
rect 23979 12496 23980 12536
rect 24020 12496 24021 12536
rect 23979 12487 24021 12496
rect 24171 12536 24213 12545
rect 24171 12496 24172 12536
rect 24212 12496 24213 12536
rect 24171 12487 24213 12496
rect 24459 12536 24501 12545
rect 24459 12496 24460 12536
rect 24500 12496 24501 12536
rect 24459 12487 24501 12496
rect 25323 12536 25365 12545
rect 25323 12496 25324 12536
rect 25364 12496 25365 12536
rect 25323 12487 25365 12496
rect 25515 12536 25557 12545
rect 25515 12496 25516 12536
rect 25556 12496 25557 12536
rect 25515 12487 25557 12496
rect 25707 12536 25749 12545
rect 25707 12496 25708 12536
rect 25748 12496 25749 12536
rect 25707 12487 25749 12496
rect 25899 12536 25941 12545
rect 25899 12496 25900 12536
rect 25940 12496 25941 12536
rect 25899 12487 25941 12496
rect 26091 12536 26133 12545
rect 26091 12496 26092 12536
rect 26132 12496 26133 12536
rect 26091 12487 26133 12496
rect 26205 12536 26263 12537
rect 26205 12496 26214 12536
rect 26254 12496 26263 12536
rect 26205 12495 26263 12496
rect 26316 12536 26374 12537
rect 26763 12536 26805 12545
rect 26316 12496 26325 12536
rect 26365 12496 26374 12536
rect 26316 12495 26374 12496
rect 26430 12527 26472 12536
rect 26430 12487 26431 12527
rect 26471 12487 26472 12527
rect 26763 12496 26764 12536
rect 26804 12496 26805 12536
rect 26763 12487 26805 12496
rect 27099 12536 27141 12545
rect 27099 12496 27100 12536
rect 27140 12496 27141 12536
rect 27099 12487 27141 12496
rect 27250 12536 27292 12545
rect 27250 12496 27251 12536
rect 27291 12496 27292 12536
rect 27250 12487 27292 12496
rect 27766 12536 27808 12545
rect 28011 12536 28053 12545
rect 27766 12496 27767 12536
rect 27807 12496 27808 12536
rect 27766 12487 27808 12496
rect 27906 12527 27952 12536
rect 27906 12487 27907 12527
rect 27947 12487 27952 12527
rect 28011 12496 28012 12536
rect 28052 12496 28053 12536
rect 28011 12487 28053 12496
rect 28200 12536 28242 12545
rect 28200 12496 28201 12536
rect 28241 12496 28242 12536
rect 28200 12487 28242 12496
rect 28317 12536 28375 12537
rect 28317 12496 28326 12536
rect 28366 12496 28375 12536
rect 30586 12536 30644 12537
rect 28317 12495 28375 12496
rect 28443 12518 28485 12527
rect 26430 12478 26472 12487
rect 27906 12478 27952 12487
rect 28443 12478 28444 12518
rect 28484 12478 28485 12518
rect 30586 12496 30595 12536
rect 30635 12496 30644 12536
rect 30586 12495 30644 12496
rect 28443 12469 28485 12478
rect 23355 12445 23397 12454
rect 29050 12452 29108 12453
rect 23234 12403 23276 12412
rect 29050 12412 29059 12452
rect 29099 12412 29108 12452
rect 29050 12411 29108 12412
rect 30970 12452 31028 12453
rect 30970 12412 30979 12452
rect 31019 12412 31028 12452
rect 30970 12411 31028 12412
rect 5970 12394 6016 12403
rect 1899 12368 1941 12377
rect 1899 12328 1900 12368
rect 1940 12328 1941 12368
rect 1899 12319 1941 12328
rect 8331 12368 8373 12377
rect 8331 12328 8332 12368
rect 8372 12328 8373 12368
rect 8331 12319 8373 12328
rect 10731 12368 10773 12377
rect 10731 12328 10732 12368
rect 10772 12328 10773 12368
rect 10731 12319 10773 12328
rect 13743 12368 13785 12377
rect 13743 12328 13744 12368
rect 13784 12328 13785 12368
rect 13743 12319 13785 12328
rect 18411 12368 18453 12377
rect 18411 12328 18412 12368
rect 18452 12328 18453 12368
rect 18411 12319 18453 12328
rect 20811 12368 20853 12377
rect 20811 12328 20812 12368
rect 20852 12328 20853 12368
rect 20811 12319 20853 12328
rect 27723 12368 27765 12377
rect 27723 12328 27724 12368
rect 27764 12328 27765 12368
rect 27723 12319 27765 12328
rect 1323 12284 1365 12293
rect 1323 12244 1324 12284
rect 1364 12244 1365 12284
rect 1323 12235 1365 12244
rect 4666 12284 4724 12285
rect 4666 12244 4675 12284
rect 4715 12244 4724 12284
rect 4666 12243 4724 12244
rect 7851 12284 7893 12293
rect 7851 12244 7852 12284
rect 7892 12244 7893 12284
rect 7851 12235 7893 12244
rect 13515 12284 13557 12293
rect 13515 12244 13516 12284
rect 13556 12244 13557 12284
rect 13515 12235 13557 12244
rect 16587 12284 16629 12293
rect 16587 12244 16588 12284
rect 16628 12244 16629 12284
rect 16587 12235 16629 12244
rect 23499 12284 23541 12293
rect 23499 12244 23500 12284
rect 23540 12244 23541 12284
rect 23499 12235 23541 12244
rect 24171 12284 24213 12293
rect 24171 12244 24172 12284
rect 24212 12244 24213 12284
rect 24171 12235 24213 12244
rect 28683 12284 28725 12293
rect 28683 12244 28684 12284
rect 28724 12244 28725 12284
rect 28683 12235 28725 12244
rect 576 12116 31392 12140
rect 576 12076 3112 12116
rect 3480 12076 10886 12116
rect 11254 12076 18660 12116
rect 19028 12076 26434 12116
rect 26802 12076 31392 12116
rect 576 12052 31392 12076
rect 4474 11948 4532 11949
rect 4474 11908 4483 11948
rect 4523 11908 4532 11948
rect 9466 11948 9524 11949
rect 4474 11907 4532 11908
rect 7563 11906 7605 11915
rect 9466 11908 9475 11948
rect 9515 11908 9524 11948
rect 9466 11907 9524 11908
rect 12171 11948 12213 11957
rect 12171 11908 12172 11948
rect 12212 11908 12213 11948
rect 3243 11864 3285 11873
rect 3243 11824 3244 11864
rect 3284 11824 3285 11864
rect 7563 11866 7564 11906
rect 7604 11866 7605 11906
rect 12171 11899 12213 11908
rect 13018 11948 13076 11949
rect 13018 11908 13027 11948
rect 13067 11908 13076 11948
rect 13018 11907 13076 11908
rect 16762 11948 16820 11949
rect 16762 11908 16771 11948
rect 16811 11908 16820 11948
rect 16762 11907 16820 11908
rect 18298 11948 18356 11949
rect 18298 11908 18307 11948
rect 18347 11908 18356 11948
rect 18298 11907 18356 11908
rect 23307 11948 23349 11957
rect 23307 11908 23308 11948
rect 23348 11908 23349 11948
rect 23307 11899 23349 11908
rect 25611 11948 25653 11957
rect 25611 11908 25612 11948
rect 25652 11908 25653 11948
rect 25611 11899 25653 11908
rect 26187 11948 26229 11957
rect 26187 11908 26188 11948
rect 26228 11908 26229 11948
rect 26187 11899 26229 11908
rect 26379 11948 26421 11957
rect 26379 11908 26380 11948
rect 26420 11908 26421 11948
rect 26379 11899 26421 11908
rect 28011 11948 28053 11957
rect 28011 11908 28012 11948
rect 28052 11908 28053 11948
rect 28011 11899 28053 11908
rect 29739 11948 29781 11957
rect 29739 11908 29740 11948
rect 29780 11908 29781 11948
rect 29739 11899 29781 11908
rect 7563 11857 7605 11866
rect 8139 11864 8181 11873
rect 3243 11815 3285 11824
rect 8139 11824 8140 11864
rect 8180 11824 8181 11864
rect 8139 11815 8181 11824
rect 10155 11864 10197 11873
rect 10155 11824 10156 11864
rect 10196 11824 10197 11864
rect 10155 11815 10197 11824
rect 11403 11864 11445 11873
rect 11403 11824 11404 11864
rect 11444 11824 11445 11864
rect 11403 11815 11445 11824
rect 13995 11864 14037 11873
rect 13995 11824 13996 11864
rect 14036 11824 14037 11864
rect 13995 11815 14037 11824
rect 14763 11864 14805 11873
rect 14763 11824 14764 11864
rect 14804 11824 14805 11864
rect 14763 11815 14805 11824
rect 16395 11864 16437 11873
rect 16395 11824 16396 11864
rect 16436 11824 16437 11864
rect 16395 11815 16437 11824
rect 18075 11855 18117 11864
rect 18075 11815 18076 11855
rect 18116 11815 18117 11855
rect 18075 11806 18117 11815
rect 2859 11780 2901 11789
rect 2859 11740 2860 11780
rect 2900 11740 2901 11780
rect 2859 11731 2901 11740
rect 4497 11780 4539 11789
rect 4497 11740 4498 11780
rect 4538 11740 4539 11780
rect 4497 11731 4539 11740
rect 5242 11780 5300 11781
rect 5242 11740 5251 11780
rect 5291 11740 5300 11780
rect 6970 11780 7028 11781
rect 5242 11739 5300 11740
rect 6843 11738 6885 11747
rect 6970 11740 6979 11780
rect 7019 11740 7028 11780
rect 6970 11739 7028 11740
rect 7467 11780 7509 11789
rect 7467 11740 7468 11780
rect 7508 11740 7509 11780
rect 5691 11707 5733 11716
rect 1306 11696 1364 11697
rect 1306 11656 1315 11696
rect 1355 11656 1364 11696
rect 1306 11655 1364 11656
rect 4107 11696 4149 11705
rect 4107 11656 4108 11696
rect 4148 11656 4149 11696
rect 4107 11647 4149 11656
rect 4587 11696 4629 11705
rect 4587 11656 4588 11696
rect 4628 11656 4629 11696
rect 4587 11647 4629 11656
rect 5110 11696 5152 11705
rect 5110 11656 5111 11696
rect 5151 11656 5152 11696
rect 5110 11647 5152 11656
rect 5355 11696 5397 11705
rect 5355 11656 5356 11696
rect 5396 11656 5397 11696
rect 5691 11667 5692 11707
rect 5732 11667 5733 11707
rect 5691 11658 5733 11667
rect 5818 11696 5876 11697
rect 5355 11647 5397 11656
rect 5818 11656 5827 11696
rect 5867 11656 5876 11696
rect 5818 11655 5876 11656
rect 5962 11696 6020 11697
rect 5962 11656 5971 11696
rect 6011 11656 6020 11696
rect 5962 11655 6020 11656
rect 6067 11696 6125 11697
rect 6067 11656 6076 11696
rect 6116 11656 6125 11696
rect 6067 11655 6125 11656
rect 6202 11696 6260 11697
rect 6202 11656 6211 11696
rect 6251 11656 6260 11696
rect 6202 11655 6260 11656
rect 6406 11696 6448 11705
rect 6406 11656 6407 11696
rect 6447 11656 6448 11696
rect 6406 11647 6448 11656
rect 6597 11696 6639 11705
rect 6597 11656 6598 11696
rect 6638 11656 6639 11696
rect 6843 11698 6844 11738
rect 6884 11698 6885 11738
rect 7467 11731 7509 11740
rect 8043 11780 8085 11789
rect 8043 11740 8044 11780
rect 8084 11740 8085 11780
rect 8043 11731 8085 11740
rect 10923 11780 10965 11789
rect 10923 11740 10924 11780
rect 10964 11740 10965 11780
rect 10923 11731 10965 11740
rect 11499 11780 11541 11789
rect 11499 11740 11500 11780
rect 11540 11740 11541 11780
rect 11499 11731 11541 11740
rect 13899 11780 13941 11789
rect 13899 11740 13900 11780
rect 13940 11740 13941 11780
rect 13899 11731 13941 11740
rect 15723 11780 15765 11789
rect 15723 11740 15724 11780
rect 15764 11740 15765 11780
rect 15723 11731 15765 11740
rect 16484 11780 16526 11789
rect 16484 11740 16485 11780
rect 16525 11740 16526 11780
rect 16484 11731 16526 11740
rect 20331 11780 20373 11789
rect 20331 11740 20332 11780
rect 20372 11740 20373 11780
rect 22539 11780 22581 11789
rect 20331 11731 20373 11740
rect 22375 11738 22417 11747
rect 6843 11689 6885 11698
rect 7083 11696 7125 11705
rect 6597 11647 6639 11656
rect 7083 11656 7084 11696
rect 7124 11656 7125 11696
rect 7083 11647 7125 11656
rect 7323 11696 7365 11705
rect 7323 11656 7324 11696
rect 7364 11656 7365 11696
rect 7323 11647 7365 11656
rect 7624 11696 7666 11705
rect 7624 11656 7625 11696
rect 7665 11656 7666 11696
rect 7624 11647 7666 11656
rect 7906 11696 7964 11697
rect 7906 11656 7915 11696
rect 7955 11656 7964 11696
rect 8362 11696 8420 11697
rect 7906 11655 7964 11656
rect 7738 11654 7796 11655
rect 922 11612 980 11613
rect 922 11572 931 11612
rect 971 11572 980 11612
rect 922 11571 980 11572
rect 6507 11612 6549 11621
rect 7738 11614 7747 11654
rect 7787 11614 7796 11654
rect 7738 11613 7796 11614
rect 8207 11654 8249 11663
rect 8362 11656 8371 11696
rect 8411 11656 8420 11696
rect 8362 11655 8420 11656
rect 9133 11696 9191 11697
rect 9133 11656 9142 11696
rect 9182 11656 9191 11696
rect 9133 11655 9191 11656
rect 9483 11696 9525 11705
rect 9483 11656 9484 11696
rect 9524 11656 9525 11696
rect 8207 11614 8208 11654
rect 8248 11614 8249 11654
rect 9483 11647 9525 11656
rect 9590 11696 9632 11705
rect 9590 11656 9591 11696
rect 9631 11656 9632 11696
rect 9590 11647 9632 11656
rect 10155 11696 10197 11705
rect 10155 11656 10156 11696
rect 10196 11656 10197 11696
rect 10155 11647 10197 11656
rect 10474 11696 10532 11697
rect 10474 11656 10483 11696
rect 10523 11656 10532 11696
rect 10474 11655 10532 11656
rect 11098 11696 11156 11697
rect 11098 11656 11107 11696
rect 11147 11656 11156 11696
rect 11098 11655 11156 11656
rect 11771 11696 11829 11697
rect 11771 11656 11780 11696
rect 11820 11656 11829 11696
rect 11771 11655 11829 11656
rect 12651 11696 12693 11705
rect 12651 11656 12652 11696
rect 12692 11656 12693 11696
rect 12651 11647 12693 11656
rect 12826 11696 12884 11697
rect 12826 11656 12835 11696
rect 12875 11656 12884 11696
rect 12826 11655 12884 11656
rect 13018 11696 13076 11697
rect 13018 11656 13027 11696
rect 13067 11656 13076 11696
rect 13018 11655 13076 11656
rect 13174 11696 13232 11697
rect 13174 11656 13183 11696
rect 13223 11656 13232 11696
rect 13174 11655 13232 11656
rect 13276 11696 13334 11697
rect 13276 11656 13285 11696
rect 13325 11656 13334 11696
rect 13276 11655 13334 11656
rect 13405 11696 13447 11705
rect 13405 11656 13406 11696
rect 13446 11656 13447 11696
rect 13405 11647 13447 11656
rect 13536 11696 13594 11697
rect 13536 11656 13545 11696
rect 13585 11656 13594 11696
rect 13536 11655 13594 11656
rect 13755 11696 13797 11705
rect 13755 11656 13756 11696
rect 13796 11656 13797 11696
rect 13755 11647 13797 11656
rect 14070 11696 14112 11705
rect 14070 11656 14071 11696
rect 14111 11656 14112 11696
rect 14070 11647 14112 11656
rect 14218 11696 14276 11697
rect 14218 11656 14227 11696
rect 14267 11656 14276 11696
rect 14218 11655 14276 11656
rect 14571 11696 14613 11705
rect 14571 11656 14572 11696
rect 14612 11656 14613 11696
rect 14571 11647 14613 11656
rect 14938 11696 14996 11697
rect 14938 11656 14947 11696
rect 14987 11656 14996 11696
rect 14938 11655 14996 11656
rect 15056 11696 15114 11697
rect 15056 11656 15065 11696
rect 15105 11656 15114 11696
rect 15056 11655 15114 11656
rect 15188 11696 15246 11697
rect 15188 11656 15197 11696
rect 15237 11656 15246 11696
rect 15188 11655 15246 11656
rect 15322 11696 15380 11697
rect 15322 11656 15331 11696
rect 15371 11656 15380 11696
rect 15322 11655 15380 11656
rect 15456 11696 15514 11697
rect 15456 11656 15465 11696
rect 15505 11656 15514 11696
rect 15456 11655 15514 11656
rect 15819 11696 15861 11705
rect 16059 11696 16101 11705
rect 15819 11656 15820 11696
rect 15860 11656 15861 11696
rect 15819 11647 15861 11656
rect 15954 11687 16000 11696
rect 15954 11647 15955 11687
rect 15995 11647 16000 11687
rect 16059 11656 16060 11696
rect 16100 11656 16101 11696
rect 16059 11647 16101 11656
rect 16162 11696 16204 11705
rect 16162 11656 16163 11696
rect 16203 11656 16204 11696
rect 16162 11647 16204 11656
rect 16334 11696 16376 11705
rect 16334 11656 16335 11696
rect 16375 11656 16376 11696
rect 16334 11647 16376 11656
rect 16612 11696 16654 11705
rect 16612 11656 16613 11696
rect 16653 11656 16654 11696
rect 16612 11647 16654 11656
rect 16762 11696 16820 11697
rect 16762 11656 16771 11696
rect 16811 11656 16820 11696
rect 16762 11655 16820 11656
rect 16906 11696 16964 11697
rect 16906 11656 16915 11696
rect 16955 11656 16964 11696
rect 16906 11655 16964 11656
rect 17154 11696 17212 11697
rect 17154 11656 17163 11696
rect 17203 11656 17212 11696
rect 17154 11655 17212 11656
rect 17323 11696 17381 11697
rect 17323 11656 17332 11696
rect 17372 11656 17381 11696
rect 17323 11655 17381 11656
rect 18106 11696 18164 11697
rect 18106 11656 18115 11696
rect 18155 11656 18164 11696
rect 18106 11655 18164 11656
rect 19354 11696 19412 11697
rect 19354 11656 19363 11696
rect 19403 11656 19412 11696
rect 19354 11655 19412 11656
rect 19843 11696 19901 11697
rect 19843 11656 19852 11696
rect 19892 11656 19901 11696
rect 19843 11655 19901 11656
rect 20427 11696 20469 11705
rect 20427 11656 20428 11696
rect 20468 11656 20469 11696
rect 15954 11638 16000 11647
rect 17058 11645 17104 11654
rect 20427 11647 20469 11656
rect 20811 11696 20853 11705
rect 20811 11656 20812 11696
rect 20852 11656 20853 11696
rect 20811 11647 20853 11656
rect 20921 11696 20979 11697
rect 20921 11656 20930 11696
rect 20970 11656 20979 11696
rect 20921 11655 20979 11656
rect 21867 11696 21909 11705
rect 21867 11656 21868 11696
rect 21908 11656 21909 11696
rect 21867 11647 21909 11656
rect 22042 11696 22100 11697
rect 22042 11656 22051 11696
rect 22091 11656 22100 11696
rect 22042 11655 22100 11656
rect 22203 11696 22245 11705
rect 22203 11656 22204 11696
rect 22244 11656 22245 11696
rect 22375 11698 22376 11738
rect 22416 11698 22417 11738
rect 22539 11740 22540 11780
rect 22580 11740 22581 11780
rect 22539 11731 22581 11740
rect 23115 11780 23157 11789
rect 23115 11740 23116 11780
rect 23156 11740 23157 11780
rect 23115 11731 23157 11740
rect 28418 11780 28460 11789
rect 28418 11740 28419 11780
rect 28459 11740 28460 11780
rect 28418 11731 28460 11740
rect 22375 11689 22417 11698
rect 22660 11696 22702 11705
rect 22203 11647 22245 11656
rect 22660 11656 22661 11696
rect 22701 11656 22702 11696
rect 22660 11647 22702 11656
rect 22802 11696 22844 11705
rect 22802 11656 22803 11696
rect 22843 11656 22844 11696
rect 22802 11647 22844 11656
rect 22906 11696 22964 11697
rect 22906 11656 22915 11696
rect 22955 11656 22964 11696
rect 22906 11655 22964 11656
rect 23019 11696 23061 11705
rect 23019 11656 23020 11696
rect 23060 11656 23061 11696
rect 23019 11647 23061 11656
rect 23307 11696 23349 11705
rect 23307 11656 23308 11696
rect 23348 11656 23349 11696
rect 23307 11647 23349 11656
rect 23600 11696 23658 11697
rect 23600 11656 23609 11696
rect 23649 11656 23658 11696
rect 23600 11655 23658 11656
rect 24459 11696 24501 11705
rect 24459 11656 24460 11696
rect 24500 11656 24501 11696
rect 24459 11647 24501 11656
rect 25323 11696 25365 11705
rect 25323 11656 25324 11696
rect 25364 11656 25365 11696
rect 25323 11647 25365 11656
rect 25437 11696 25495 11697
rect 25437 11656 25446 11696
rect 25486 11656 25495 11696
rect 25437 11655 25495 11656
rect 25563 11696 25605 11705
rect 25563 11656 25564 11696
rect 25604 11656 25605 11696
rect 25563 11647 25605 11656
rect 25995 11696 26037 11705
rect 25995 11656 25996 11696
rect 26036 11656 26037 11696
rect 25995 11647 26037 11656
rect 26379 11696 26421 11705
rect 26379 11656 26380 11696
rect 26420 11656 26421 11696
rect 26379 11647 26421 11656
rect 26576 11696 26618 11705
rect 26576 11656 26577 11696
rect 26617 11656 26618 11696
rect 26576 11647 26618 11656
rect 26859 11696 26901 11705
rect 26859 11656 26860 11696
rect 26900 11656 26901 11696
rect 26859 11647 26901 11656
rect 27706 11696 27764 11697
rect 27706 11656 27715 11696
rect 27755 11656 27764 11696
rect 27706 11655 27764 11656
rect 27819 11696 27861 11705
rect 27819 11656 27820 11696
rect 27860 11656 27861 11696
rect 27819 11647 27861 11656
rect 28299 11696 28341 11705
rect 28299 11656 28300 11696
rect 28340 11656 28341 11696
rect 28299 11647 28341 11656
rect 28516 11696 28558 11705
rect 28516 11656 28517 11696
rect 28557 11656 28558 11696
rect 28516 11647 28558 11656
rect 28875 11696 28917 11705
rect 28875 11656 28876 11696
rect 28916 11656 28917 11696
rect 28875 11647 28917 11656
rect 29547 11696 29589 11705
rect 29547 11656 29548 11696
rect 29588 11656 29589 11696
rect 29547 11647 29589 11656
rect 29739 11696 29781 11705
rect 29739 11656 29740 11696
rect 29780 11656 29781 11696
rect 29739 11647 29781 11656
rect 29931 11696 29973 11705
rect 29931 11656 29932 11696
rect 29972 11656 29973 11696
rect 29931 11647 29973 11656
rect 30123 11696 30165 11705
rect 30123 11656 30124 11696
rect 30164 11656 30165 11696
rect 30123 11647 30165 11656
rect 30315 11696 30357 11705
rect 30315 11656 30316 11696
rect 30356 11656 30357 11696
rect 30315 11647 30357 11656
rect 30682 11696 30740 11697
rect 30682 11656 30691 11696
rect 30731 11656 30740 11696
rect 30682 11655 30740 11656
rect 6507 11572 6508 11612
rect 6548 11572 6549 11612
rect 8207 11605 8249 11614
rect 8938 11612 8996 11613
rect 6507 11563 6549 11572
rect 8938 11572 8947 11612
rect 8987 11572 8996 11612
rect 8938 11571 8996 11572
rect 11403 11612 11445 11621
rect 11403 11572 11404 11612
rect 11444 11572 11445 11612
rect 11403 11563 11445 11572
rect 12747 11612 12789 11621
rect 12747 11572 12748 11612
rect 12788 11572 12789 11612
rect 17058 11605 17059 11645
rect 17099 11605 17104 11645
rect 17058 11596 17104 11605
rect 21963 11612 22005 11621
rect 12747 11563 12789 11572
rect 21963 11572 21964 11612
rect 22004 11572 22005 11612
rect 26475 11612 26517 11621
rect 21963 11563 22005 11572
rect 22457 11570 22499 11579
rect 3435 11528 3477 11537
rect 3435 11488 3436 11528
rect 3476 11488 3477 11528
rect 3435 11479 3477 11488
rect 5434 11528 5492 11529
rect 5434 11488 5443 11528
rect 5483 11488 5492 11528
rect 5434 11487 5492 11488
rect 5722 11528 5780 11529
rect 5722 11488 5731 11528
rect 5771 11488 5780 11528
rect 5722 11487 5780 11488
rect 7162 11528 7220 11529
rect 7162 11488 7171 11528
rect 7211 11488 7220 11528
rect 7162 11487 7220 11488
rect 13498 11528 13556 11529
rect 13498 11488 13507 11528
rect 13547 11488 13556 11528
rect 13498 11487 13556 11488
rect 14458 11528 14516 11529
rect 14458 11488 14467 11528
rect 14507 11488 14516 11528
rect 14458 11487 14516 11488
rect 15418 11528 15476 11529
rect 15418 11488 15427 11528
rect 15467 11488 15476 11528
rect 15418 11487 15476 11488
rect 19179 11528 19221 11537
rect 19179 11488 19180 11528
rect 19220 11488 19221 11528
rect 22457 11530 22458 11570
rect 22498 11530 22499 11570
rect 26475 11572 26476 11612
rect 26516 11572 26517 11612
rect 26475 11563 26517 11572
rect 28025 11612 28067 11621
rect 28025 11572 28026 11612
rect 28066 11572 28067 11612
rect 28025 11563 28067 11572
rect 28203 11612 28245 11621
rect 28203 11572 28204 11612
rect 28244 11572 28245 11612
rect 28203 11563 28245 11572
rect 30219 11612 30261 11621
rect 30219 11572 30220 11612
rect 30260 11572 30261 11612
rect 30219 11563 30261 11572
rect 22457 11521 22499 11530
rect 23787 11528 23829 11537
rect 19179 11479 19221 11488
rect 23787 11488 23788 11528
rect 23828 11488 23829 11528
rect 23787 11479 23829 11488
rect 25882 11528 25940 11529
rect 25882 11488 25891 11528
rect 25931 11488 25940 11528
rect 25882 11487 25940 11488
rect 27531 11528 27573 11537
rect 27531 11488 27532 11528
rect 27572 11488 27573 11528
rect 27531 11479 27573 11488
rect 30891 11528 30933 11537
rect 30891 11488 30892 11528
rect 30932 11488 30933 11528
rect 30891 11479 30933 11488
rect 576 11360 31392 11384
rect 576 11320 4352 11360
rect 4720 11320 12126 11360
rect 12494 11320 19900 11360
rect 20268 11320 27674 11360
rect 28042 11320 31392 11360
rect 576 11296 31392 11320
rect 4186 11192 4244 11193
rect 4186 11152 4195 11192
rect 4235 11152 4244 11192
rect 4186 11151 4244 11152
rect 4762 11192 4820 11193
rect 4762 11152 4771 11192
rect 4811 11152 4820 11192
rect 4762 11151 4820 11152
rect 5163 11192 5205 11201
rect 5163 11152 5164 11192
rect 5204 11152 5205 11192
rect 5163 11143 5205 11152
rect 6939 11192 6981 11201
rect 6939 11152 6940 11192
rect 6980 11152 6981 11192
rect 6939 11143 6981 11152
rect 7275 11192 7317 11201
rect 7275 11152 7276 11192
rect 7316 11152 7317 11192
rect 7275 11143 7317 11152
rect 8043 11192 8085 11201
rect 8043 11152 8044 11192
rect 8084 11152 8085 11192
rect 8043 11143 8085 11152
rect 8907 11192 8949 11201
rect 8907 11152 8908 11192
rect 8948 11152 8949 11192
rect 8907 11143 8949 11152
rect 10546 11192 10604 11193
rect 10546 11152 10555 11192
rect 10595 11152 10604 11192
rect 10546 11151 10604 11152
rect 11386 11192 11444 11193
rect 11386 11152 11395 11192
rect 11435 11152 11444 11192
rect 11386 11151 11444 11152
rect 11691 11192 11733 11201
rect 11691 11152 11692 11192
rect 11732 11152 11733 11192
rect 11691 11143 11733 11152
rect 12603 11192 12645 11201
rect 12603 11152 12604 11192
rect 12644 11152 12645 11192
rect 12603 11143 12645 11152
rect 13515 11192 13557 11201
rect 13515 11152 13516 11192
rect 13556 11152 13557 11192
rect 13515 11143 13557 11152
rect 14362 11192 14420 11193
rect 14362 11152 14371 11192
rect 14411 11152 14420 11192
rect 14362 11151 14420 11152
rect 15610 11192 15668 11193
rect 15610 11152 15619 11192
rect 15659 11152 15668 11192
rect 15610 11151 15668 11152
rect 16683 11192 16725 11201
rect 16683 11152 16684 11192
rect 16724 11152 16725 11192
rect 16683 11143 16725 11152
rect 17835 11192 17877 11201
rect 17835 11152 17836 11192
rect 17876 11152 17877 11192
rect 17835 11143 17877 11152
rect 19179 11192 19221 11201
rect 19179 11152 19180 11192
rect 19220 11152 19221 11192
rect 19179 11143 19221 11152
rect 19467 11192 19509 11201
rect 19467 11152 19468 11192
rect 19508 11152 19509 11192
rect 19467 11143 19509 11152
rect 21867 11192 21909 11201
rect 21867 11152 21868 11192
rect 21908 11152 21909 11192
rect 21867 11143 21909 11152
rect 26667 11192 26709 11201
rect 26667 11152 26668 11192
rect 26708 11152 26709 11192
rect 26667 11143 26709 11152
rect 26986 11192 27044 11193
rect 26986 11152 26995 11192
rect 27035 11152 27044 11192
rect 26986 11151 27044 11152
rect 27915 11192 27957 11201
rect 27915 11152 27916 11192
rect 27956 11152 27957 11192
rect 27915 11143 27957 11152
rect 3898 11108 3956 11109
rect 3898 11068 3907 11108
rect 3947 11068 3956 11108
rect 3898 11067 3956 11068
rect 14859 11108 14901 11117
rect 14859 11068 14860 11108
rect 14900 11068 14901 11108
rect 14859 11059 14901 11068
rect 17259 11108 17301 11117
rect 17259 11068 17260 11108
rect 17300 11068 17301 11108
rect 17259 11059 17301 11068
rect 22251 11108 22293 11117
rect 22251 11068 22252 11108
rect 22292 11068 22293 11108
rect 22251 11059 22293 11068
rect 23403 11108 23445 11117
rect 23403 11068 23404 11108
rect 23444 11068 23445 11108
rect 23403 11059 23445 11068
rect 31258 11108 31316 11109
rect 31258 11068 31267 11108
rect 31307 11068 31316 11108
rect 31258 11067 31316 11068
rect 1131 11024 1173 11033
rect 1131 10984 1132 11024
rect 1172 10984 1173 11024
rect 1131 10975 1173 10984
rect 1248 11024 1306 11025
rect 1248 10984 1257 11024
rect 1297 10984 1306 11024
rect 1248 10983 1306 10984
rect 1419 11024 1461 11033
rect 1419 10984 1420 11024
rect 1460 10984 1461 11024
rect 1419 10975 1461 10984
rect 2955 11024 2997 11033
rect 2955 10984 2956 11024
rect 2996 10984 2997 11024
rect 2955 10975 2997 10984
rect 3439 11024 3497 11025
rect 3439 10984 3448 11024
rect 3488 10984 3497 11024
rect 3439 10983 3497 10984
rect 4107 11024 4149 11033
rect 4107 10984 4108 11024
rect 4148 10984 4149 11024
rect 4107 10975 4149 10984
rect 4411 11024 4469 11025
rect 4411 10984 4420 11024
rect 4460 10984 4469 11024
rect 4411 10983 4469 10984
rect 4548 11024 4606 11025
rect 4548 10984 4557 11024
rect 4597 10984 4606 11024
rect 4548 10983 4606 10984
rect 4695 11024 4737 11033
rect 4695 10984 4696 11024
rect 4736 10984 4737 11024
rect 4695 10975 4737 10984
rect 4853 11024 4911 11025
rect 4853 10984 4862 11024
rect 4902 10984 4911 11024
rect 4853 10983 4911 10984
rect 4954 11024 5012 11025
rect 4954 10984 4963 11024
rect 5003 10984 5012 11024
rect 4954 10983 5012 10984
rect 5259 11024 5301 11033
rect 5259 10984 5260 11024
rect 5300 10984 5301 11024
rect 5259 10975 5301 10984
rect 5488 11024 5546 11025
rect 5488 10984 5497 11024
rect 5537 10984 5546 11024
rect 5488 10983 5546 10984
rect 6411 11024 6453 11033
rect 6411 10984 6412 11024
rect 6452 10984 6453 11024
rect 6411 10975 6453 10984
rect 6586 11024 6644 11025
rect 6586 10984 6595 11024
rect 6635 10984 6644 11024
rect 6586 10983 6644 10984
rect 7083 11024 7125 11033
rect 7083 10984 7084 11024
rect 7124 10984 7125 11024
rect 7083 10975 7125 10984
rect 7371 11024 7413 11033
rect 7371 10984 7372 11024
rect 7412 10984 7413 11024
rect 7371 10975 7413 10984
rect 7600 11024 7658 11025
rect 7600 10984 7609 11024
rect 7649 10984 7658 11024
rect 7600 10983 7658 10984
rect 8139 11024 8181 11033
rect 8139 10984 8140 11024
rect 8180 10984 8181 11024
rect 8139 10975 8181 10984
rect 8356 11024 8398 11033
rect 8356 10984 8357 11024
rect 8397 10984 8398 11024
rect 8356 10975 8398 10984
rect 8619 11024 8661 11033
rect 8619 10984 8620 11024
rect 8660 10984 8661 11024
rect 8619 10975 8661 10984
rect 8733 11024 8791 11025
rect 8733 10984 8742 11024
rect 8782 10984 8791 11024
rect 8733 10983 8791 10984
rect 8860 11024 8918 11025
rect 9480 11024 9538 11025
rect 10426 11024 10484 11025
rect 8860 10984 8869 11024
rect 8909 10984 8918 11024
rect 8860 10983 8918 10984
rect 9260 11015 9302 11024
rect 9260 10975 9261 11015
rect 9301 10975 9302 11015
rect 9260 10966 9302 10975
rect 9378 11015 9424 11024
rect 9378 10975 9379 11015
rect 9419 10975 9424 11015
rect 9480 10984 9489 11024
rect 9529 10984 9538 11024
rect 9480 10983 9538 10984
rect 10335 11015 10377 11024
rect 9378 10966 9424 10975
rect 10335 10975 10336 11015
rect 10376 10975 10377 11015
rect 10426 10984 10435 11024
rect 10475 10984 10484 11024
rect 10426 10983 10484 10984
rect 11062 11024 11104 11033
rect 11062 10984 11063 11024
rect 11103 10984 11104 11024
rect 11062 10975 11104 10984
rect 11305 11024 11347 11033
rect 11305 10984 11306 11024
rect 11346 10984 11347 11024
rect 11305 10975 11347 10984
rect 11595 11024 11637 11033
rect 11595 10984 11596 11024
rect 11636 10984 11637 11024
rect 11595 10975 11637 10984
rect 11787 11024 11829 11033
rect 11787 10984 11788 11024
rect 11828 10984 11829 11024
rect 11787 10975 11829 10984
rect 13131 11024 13173 11033
rect 13131 10984 13132 11024
rect 13172 10984 13173 11024
rect 13131 10975 13173 10984
rect 13300 11024 13342 11033
rect 13300 10984 13301 11024
rect 13341 10984 13342 11024
rect 13828 11024 13870 11033
rect 13300 10975 13342 10984
rect 13611 10982 13653 10991
rect 10335 10966 10377 10975
rect 3274 10940 3332 10941
rect 8258 10940 8300 10949
rect 3274 10900 3283 10940
rect 3323 10900 3332 10940
rect 3274 10899 3332 10900
rect 5394 10931 5440 10940
rect 5394 10891 5395 10931
rect 5435 10891 5440 10931
rect 5394 10882 5440 10891
rect 7506 10931 7552 10940
rect 7506 10891 7507 10931
rect 7547 10891 7552 10931
rect 8258 10900 8259 10940
rect 8299 10900 8300 10940
rect 8258 10891 8300 10900
rect 11194 10940 11252 10941
rect 11194 10900 11203 10940
rect 11243 10900 11252 10940
rect 11194 10899 11252 10900
rect 12363 10940 12405 10949
rect 12363 10900 12364 10940
rect 12404 10900 12405 10940
rect 13611 10942 13612 10982
rect 13652 10942 13653 10982
rect 13828 10984 13829 11024
rect 13869 10984 13870 11024
rect 13828 10975 13870 10984
rect 14269 11024 14311 11033
rect 14269 10984 14270 11024
rect 14310 10984 14311 11024
rect 14269 10975 14311 10984
rect 14475 11024 14517 11033
rect 14955 11024 14997 11033
rect 14475 10984 14476 11024
rect 14516 10984 14517 11024
rect 14475 10975 14517 10984
rect 14571 11015 14613 11024
rect 14571 10975 14572 11015
rect 14612 10975 14613 11015
rect 14955 10984 14956 11024
rect 14996 10984 14997 11024
rect 14955 10975 14997 10984
rect 15184 11024 15242 11025
rect 15184 10984 15193 11024
rect 15233 10984 15242 11024
rect 15184 10983 15242 10984
rect 15418 11024 15476 11025
rect 15418 10984 15427 11024
rect 15467 10984 15476 11024
rect 15418 10983 15476 10984
rect 15771 11024 15813 11033
rect 15771 10984 15772 11024
rect 15812 10984 15813 11024
rect 15771 10975 15813 10984
rect 16234 11024 16292 11025
rect 16234 10984 16243 11024
rect 16283 10984 16292 11024
rect 16234 10983 16292 10984
rect 16779 11024 16821 11033
rect 16779 10984 16780 11024
rect 16820 10984 16821 11024
rect 16090 10982 16148 10983
rect 14571 10966 14613 10975
rect 13611 10933 13653 10942
rect 13730 10940 13772 10949
rect 15915 10940 15957 10949
rect 16090 10942 16099 10982
rect 16139 10942 16148 10982
rect 16779 10975 16821 10984
rect 17008 11024 17066 11025
rect 17008 10984 17017 11024
rect 17057 10984 17066 11024
rect 17008 10983 17066 10984
rect 17355 11024 17397 11033
rect 17355 10984 17356 11024
rect 17396 10984 17397 11024
rect 17355 10975 17397 10984
rect 17584 11024 17642 11025
rect 17584 10984 17593 11024
rect 17633 10984 17642 11024
rect 17584 10983 17642 10984
rect 17739 11024 17781 11033
rect 17739 10984 17740 11024
rect 17780 10984 17781 11024
rect 17739 10975 17781 10984
rect 17931 11024 17973 11033
rect 17931 10984 17932 11024
rect 17972 10984 17973 11024
rect 17931 10975 17973 10984
rect 18682 11024 18740 11025
rect 18682 10984 18691 11024
rect 18731 10984 18740 11024
rect 18682 10983 18740 10984
rect 19083 11024 19125 11033
rect 19083 10984 19084 11024
rect 19124 10984 19125 11024
rect 19083 10975 19125 10984
rect 19275 11024 19317 11033
rect 19275 10984 19276 11024
rect 19316 10984 19317 11024
rect 19275 10975 19317 10984
rect 19642 11024 19700 11025
rect 20619 11024 20661 11033
rect 19642 10984 19651 11024
rect 19691 10984 19700 11024
rect 19642 10983 19700 10984
rect 20139 11015 20181 11024
rect 20139 10975 20140 11015
rect 20180 10975 20181 11015
rect 20619 10984 20620 11024
rect 20660 10984 20661 11024
rect 20619 10975 20661 10984
rect 21099 11024 21141 11033
rect 21099 10984 21100 11024
rect 21140 10984 21141 11024
rect 21099 10975 21141 10984
rect 21209 11024 21267 11025
rect 21209 10984 21218 11024
rect 21258 10984 21267 11024
rect 21209 10983 21267 10984
rect 21771 11024 21813 11033
rect 21771 10984 21772 11024
rect 21812 10984 21813 11024
rect 21771 10975 21813 10984
rect 21946 11024 22004 11025
rect 21946 10984 21955 11024
rect 21995 10984 22004 11024
rect 21946 10983 22004 10984
rect 22155 11024 22197 11033
rect 22155 10984 22156 11024
rect 22196 10984 22197 11024
rect 22155 10975 22197 10984
rect 22347 11024 22389 11033
rect 22347 10984 22348 11024
rect 22388 10984 22389 11024
rect 22347 10975 22389 10984
rect 22714 11024 22772 11025
rect 22714 10984 22723 11024
rect 22763 10984 22772 11024
rect 22714 10983 22772 10984
rect 22827 11024 22869 11033
rect 22827 10984 22828 11024
rect 22868 10984 22869 11024
rect 22827 10975 22869 10984
rect 23307 11024 23349 11033
rect 23307 10984 23308 11024
rect 23348 10984 23349 11024
rect 23307 10975 23349 10984
rect 23482 11024 23540 11025
rect 23482 10984 23491 11024
rect 23531 10984 23540 11024
rect 23482 10983 23540 10984
rect 23883 11024 23925 11033
rect 23883 10984 23884 11024
rect 23924 10984 23925 11024
rect 23883 10975 23925 10984
rect 24058 11024 24116 11025
rect 24058 10984 24067 11024
rect 24107 10984 24116 11024
rect 24730 11024 24788 11025
rect 24058 10983 24116 10984
rect 24169 11012 24227 11013
rect 20139 10966 20181 10975
rect 24169 10972 24178 11012
rect 24218 10972 24227 11012
rect 24730 10984 24739 11024
rect 24779 10984 24788 11024
rect 24730 10983 24788 10984
rect 27181 11024 27239 11025
rect 27181 10984 27190 11024
rect 27230 10984 27239 11024
rect 27181 10983 27239 10984
rect 27514 11024 27572 11025
rect 27514 10984 27523 11024
rect 27563 10984 27572 11024
rect 27514 10983 27572 10984
rect 27627 11024 27669 11033
rect 27627 10984 27628 11024
rect 27668 10984 27669 11024
rect 27627 10975 27669 10984
rect 28107 11024 28149 11033
rect 28107 10984 28108 11024
rect 28148 10984 28149 11024
rect 28107 10975 28149 10984
rect 30874 11024 30932 11025
rect 30874 10984 30883 11024
rect 30923 10984 30932 11024
rect 30874 10983 30932 10984
rect 24169 10971 24227 10972
rect 16090 10941 16148 10942
rect 18298 10940 18356 10941
rect 12363 10891 12405 10900
rect 13730 10900 13731 10940
rect 13771 10900 13772 10940
rect 13730 10891 13772 10900
rect 15090 10931 15136 10940
rect 15090 10891 15091 10931
rect 15131 10891 15136 10931
rect 15915 10900 15916 10940
rect 15956 10900 15957 10940
rect 15915 10891 15957 10900
rect 16914 10931 16960 10940
rect 16914 10891 16915 10931
rect 16955 10891 16960 10931
rect 7506 10882 7552 10891
rect 15090 10882 15136 10891
rect 16914 10882 16960 10891
rect 17490 10931 17536 10940
rect 17490 10891 17491 10931
rect 17531 10891 17536 10931
rect 18298 10900 18307 10940
rect 18347 10900 18356 10940
rect 18298 10899 18356 10900
rect 18874 10940 18932 10941
rect 18874 10900 18883 10940
rect 18923 10900 18932 10940
rect 18874 10899 18932 10900
rect 20715 10940 20757 10949
rect 20715 10900 20716 10940
rect 20756 10900 20757 10940
rect 20715 10891 20757 10900
rect 24363 10940 24405 10949
rect 24363 10900 24364 10940
rect 24404 10900 24405 10940
rect 24363 10891 24405 10900
rect 26283 10940 26325 10949
rect 26283 10900 26284 10940
rect 26324 10900 26325 10940
rect 26283 10891 26325 10900
rect 17490 10882 17536 10891
rect 1131 10856 1173 10865
rect 1131 10816 1132 10856
rect 1172 10816 1173 10856
rect 1131 10807 1173 10816
rect 9099 10856 9141 10865
rect 9099 10816 9100 10856
rect 9140 10816 9141 10856
rect 9099 10807 9141 10816
rect 10042 10856 10100 10857
rect 10042 10816 10051 10856
rect 10091 10816 10100 10856
rect 10042 10815 10100 10816
rect 15398 10856 15440 10865
rect 15398 10816 15399 10856
rect 15439 10816 15440 10856
rect 15398 10807 15440 10816
rect 16011 10856 16053 10865
rect 16011 10816 16012 10856
rect 16052 10816 16053 10856
rect 16011 10807 16053 10816
rect 18394 10856 18452 10857
rect 18394 10816 18403 10856
rect 18443 10816 18452 10856
rect 18394 10815 18452 10816
rect 24171 10856 24213 10865
rect 24171 10816 24172 10856
rect 24212 10816 24213 10856
rect 24171 10807 24213 10816
rect 2283 10772 2325 10781
rect 2283 10732 2284 10772
rect 2324 10732 2325 10772
rect 2283 10723 2325 10732
rect 6586 10772 6644 10773
rect 6586 10732 6595 10772
rect 6635 10732 6644 10772
rect 6586 10731 6644 10732
rect 13306 10772 13364 10773
rect 13306 10732 13315 10772
rect 13355 10732 13364 10772
rect 13306 10731 13364 10732
rect 23002 10772 23060 10773
rect 23002 10732 23011 10772
rect 23051 10732 23060 10772
rect 23002 10731 23060 10732
rect 28779 10772 28821 10781
rect 28779 10732 28780 10772
rect 28820 10732 28821 10772
rect 28779 10723 28821 10732
rect 28971 10772 29013 10781
rect 28971 10732 28972 10772
rect 29012 10732 29013 10772
rect 28971 10723 29013 10732
rect 29355 10772 29397 10781
rect 29355 10732 29356 10772
rect 29396 10732 29397 10772
rect 29355 10723 29397 10732
rect 576 10604 31392 10628
rect 576 10564 3112 10604
rect 3480 10564 10886 10604
rect 11254 10564 18660 10604
rect 19028 10564 26434 10604
rect 26802 10564 31392 10604
rect 576 10540 31392 10564
rect 651 10436 693 10445
rect 651 10396 652 10436
rect 692 10396 693 10436
rect 651 10387 693 10396
rect 4875 10436 4917 10445
rect 4875 10396 4876 10436
rect 4916 10396 4917 10436
rect 4875 10387 4917 10396
rect 5722 10436 5780 10437
rect 5722 10396 5731 10436
rect 5771 10396 5780 10436
rect 5722 10395 5780 10396
rect 9466 10436 9524 10437
rect 9466 10396 9475 10436
rect 9515 10396 9524 10436
rect 9466 10395 9524 10396
rect 14938 10436 14996 10437
rect 14938 10396 14947 10436
rect 14987 10396 14996 10436
rect 14938 10395 14996 10396
rect 21099 10436 21141 10445
rect 21099 10396 21100 10436
rect 21140 10396 21141 10436
rect 21099 10387 21141 10396
rect 22443 10436 22485 10445
rect 22443 10396 22444 10436
rect 22484 10396 22485 10436
rect 22443 10387 22485 10396
rect 24747 10436 24789 10445
rect 24747 10396 24748 10436
rect 24788 10396 24789 10436
rect 24747 10387 24789 10396
rect 27147 10436 27189 10445
rect 27147 10396 27148 10436
rect 27188 10396 27189 10436
rect 27147 10387 27189 10396
rect 29931 10436 29973 10445
rect 29931 10396 29932 10436
rect 29972 10396 29973 10436
rect 29931 10387 29973 10396
rect 2362 10352 2420 10353
rect 2362 10312 2371 10352
rect 2411 10312 2420 10352
rect 2362 10311 2420 10312
rect 7179 10352 7221 10361
rect 7179 10312 7180 10352
rect 7220 10312 7221 10352
rect 7179 10303 7221 10312
rect 12267 10352 12309 10361
rect 12267 10312 12268 10352
rect 12308 10312 12309 10352
rect 12267 10303 12309 10312
rect 18795 10352 18837 10361
rect 18795 10312 18796 10352
rect 18836 10312 18837 10352
rect 18795 10303 18837 10312
rect 25035 10352 25077 10361
rect 25035 10312 25036 10352
rect 25076 10312 25077 10352
rect 25035 10303 25077 10312
rect 25419 10352 25461 10361
rect 25419 10312 25420 10352
rect 25460 10312 25461 10352
rect 25419 10303 25461 10312
rect 28378 10352 28436 10353
rect 28378 10312 28387 10352
rect 28427 10312 28436 10352
rect 28378 10311 28436 10312
rect 3051 10268 3093 10277
rect 3051 10228 3052 10268
rect 3092 10228 3093 10268
rect 3051 10219 3093 10228
rect 6219 10268 6261 10277
rect 6914 10268 6956 10277
rect 6219 10228 6220 10268
rect 6260 10228 6261 10268
rect 6219 10219 6261 10228
rect 6450 10259 6496 10268
rect 6450 10219 6451 10259
rect 6491 10219 6496 10259
rect 6914 10228 6915 10268
rect 6955 10228 6956 10268
rect 6914 10219 6956 10228
rect 7642 10268 7700 10269
rect 7642 10228 7651 10268
rect 7691 10228 7700 10268
rect 7642 10227 7700 10228
rect 7851 10268 7893 10277
rect 7851 10228 7852 10268
rect 7892 10228 7893 10268
rect 7851 10219 7893 10228
rect 8427 10268 8469 10277
rect 8427 10228 8428 10268
rect 8468 10228 8469 10268
rect 8427 10219 8469 10228
rect 10754 10268 10796 10277
rect 10754 10228 10755 10268
rect 10795 10228 10796 10268
rect 11092 10268 11134 10277
rect 10754 10219 10796 10228
rect 10971 10226 11013 10235
rect 6450 10210 6496 10219
rect 4315 10195 4357 10204
rect 843 10184 885 10193
rect 843 10144 844 10184
rect 884 10144 885 10184
rect 843 10135 885 10144
rect 1419 10184 1461 10193
rect 1419 10144 1420 10184
rect 1460 10144 1461 10184
rect 1419 10135 1461 10144
rect 1546 10184 1604 10185
rect 1546 10144 1555 10184
rect 1595 10144 1604 10184
rect 1546 10143 1604 10144
rect 2074 10184 2132 10185
rect 2074 10144 2083 10184
rect 2123 10144 2132 10184
rect 2074 10143 2132 10144
rect 2187 10184 2229 10193
rect 2187 10144 2188 10184
rect 2228 10144 2229 10184
rect 2187 10135 2229 10144
rect 2710 10184 2752 10193
rect 2710 10144 2711 10184
rect 2751 10144 2752 10184
rect 2710 10135 2752 10144
rect 2842 10184 2900 10185
rect 2842 10144 2851 10184
rect 2891 10144 2900 10184
rect 2842 10143 2900 10144
rect 2955 10184 2997 10193
rect 2955 10144 2956 10184
rect 2996 10144 2997 10184
rect 2955 10135 2997 10144
rect 3531 10184 3573 10193
rect 3531 10144 3532 10184
rect 3572 10144 3573 10184
rect 3531 10135 3573 10144
rect 3915 10184 3957 10193
rect 3915 10144 3916 10184
rect 3956 10144 3957 10184
rect 4315 10155 4316 10195
rect 4356 10155 4357 10195
rect 4315 10146 4357 10155
rect 4498 10184 4556 10185
rect 3915 10135 3957 10144
rect 4498 10144 4507 10184
rect 4547 10144 4556 10184
rect 4498 10143 4556 10144
rect 4618 10184 4676 10185
rect 4618 10144 4627 10184
rect 4667 10144 4676 10184
rect 4618 10143 4676 10144
rect 4757 10184 4815 10185
rect 4757 10144 4766 10184
rect 4806 10144 4815 10184
rect 4757 10143 4815 10144
rect 4858 10184 4916 10185
rect 4858 10144 4867 10184
rect 4907 10144 4916 10184
rect 4858 10143 4916 10144
rect 5434 10184 5492 10185
rect 5434 10144 5443 10184
rect 5483 10144 5492 10184
rect 5434 10143 5492 10144
rect 5547 10184 5589 10193
rect 5547 10144 5548 10184
rect 5588 10144 5589 10184
rect 5547 10135 5589 10144
rect 6315 10184 6357 10193
rect 6315 10144 6316 10184
rect 6356 10144 6357 10184
rect 6315 10135 6357 10144
rect 6546 10184 6588 10193
rect 6546 10144 6547 10184
rect 6587 10144 6588 10184
rect 6546 10135 6588 10144
rect 6795 10184 6837 10193
rect 6795 10144 6796 10184
rect 6836 10144 6837 10184
rect 6795 10135 6837 10144
rect 7024 10184 7082 10185
rect 7024 10144 7033 10184
rect 7073 10144 7082 10184
rect 7024 10143 7082 10144
rect 7179 10184 7221 10193
rect 7179 10144 7180 10184
rect 7220 10144 7221 10184
rect 7179 10135 7221 10144
rect 7376 10184 7418 10193
rect 7376 10144 7377 10184
rect 7417 10144 7418 10184
rect 7376 10135 7418 10144
rect 7522 10184 7580 10185
rect 7522 10144 7531 10184
rect 7571 10144 7580 10184
rect 7522 10143 7580 10144
rect 7755 10184 7797 10193
rect 7755 10144 7756 10184
rect 7796 10144 7797 10184
rect 7755 10135 7797 10144
rect 8043 10184 8085 10193
rect 8043 10144 8044 10184
rect 8084 10144 8085 10184
rect 8043 10135 8085 10144
rect 8235 10184 8277 10193
rect 8235 10144 8236 10184
rect 8276 10144 8277 10184
rect 8235 10135 8277 10144
rect 8523 10184 8565 10193
rect 8523 10144 8524 10184
rect 8564 10144 8565 10184
rect 8523 10135 8565 10144
rect 8642 10184 8684 10193
rect 8642 10144 8643 10184
rect 8683 10144 8684 10184
rect 8642 10135 8684 10144
rect 8752 10184 8810 10185
rect 8752 10144 8761 10184
rect 8801 10144 8810 10184
rect 8752 10143 8810 10144
rect 9229 10184 9287 10185
rect 9229 10144 9238 10184
rect 9278 10144 9287 10184
rect 9229 10143 9287 10144
rect 9867 10184 9909 10193
rect 9867 10144 9868 10184
rect 9908 10144 9909 10184
rect 9867 10135 9909 10144
rect 10635 10184 10677 10193
rect 10635 10144 10636 10184
rect 10676 10144 10677 10184
rect 10635 10135 10677 10144
rect 10866 10184 10908 10193
rect 10866 10144 10867 10184
rect 10907 10144 10908 10184
rect 10971 10186 10972 10226
rect 11012 10186 11013 10226
rect 11092 10228 11093 10268
rect 11133 10228 11134 10268
rect 11092 10219 11134 10228
rect 11307 10268 11349 10277
rect 11307 10228 11308 10268
rect 11348 10228 11349 10268
rect 11307 10219 11349 10228
rect 11883 10268 11925 10277
rect 11883 10228 11884 10268
rect 11924 10228 11925 10268
rect 11883 10219 11925 10228
rect 12363 10268 12405 10277
rect 12363 10228 12364 10268
rect 12404 10228 12405 10268
rect 12363 10219 12405 10228
rect 13306 10268 13364 10269
rect 13306 10228 13315 10268
rect 13355 10228 13364 10268
rect 13306 10227 13364 10228
rect 13515 10268 13557 10277
rect 13515 10228 13516 10268
rect 13556 10228 13557 10268
rect 12490 10226 12548 10227
rect 10971 10177 11013 10186
rect 11196 10184 11254 10185
rect 10866 10135 10908 10144
rect 11196 10144 11205 10184
rect 11245 10144 11254 10184
rect 11196 10143 11254 10144
rect 11542 10184 11584 10193
rect 11542 10144 11543 10184
rect 11583 10144 11584 10184
rect 11542 10135 11584 10144
rect 11674 10184 11732 10185
rect 11674 10144 11683 10184
rect 11723 10144 11732 10184
rect 11674 10143 11732 10144
rect 11787 10184 11829 10193
rect 11787 10144 11788 10184
rect 11828 10144 11829 10184
rect 11787 10135 11829 10144
rect 12036 10184 12094 10185
rect 12036 10144 12045 10184
rect 12085 10144 12094 10184
rect 12036 10143 12094 10144
rect 12192 10184 12234 10193
rect 12490 10186 12499 10226
rect 12539 10186 12548 10226
rect 13515 10219 13557 10228
rect 14410 10268 14468 10269
rect 14410 10228 14419 10268
rect 14459 10228 14468 10268
rect 14410 10227 14468 10228
rect 15435 10268 15477 10277
rect 16491 10268 16533 10277
rect 17186 10268 17228 10277
rect 15435 10228 15436 10268
rect 15476 10228 15477 10268
rect 15435 10219 15477 10228
rect 15666 10259 15712 10268
rect 15666 10219 15667 10259
rect 15707 10219 15712 10259
rect 16491 10228 16492 10268
rect 16532 10228 16533 10268
rect 16491 10219 16533 10228
rect 16722 10259 16768 10268
rect 16722 10219 16723 10259
rect 16763 10219 16768 10259
rect 17186 10228 17187 10268
rect 17227 10228 17228 10268
rect 17186 10219 17228 10228
rect 31035 10268 31077 10277
rect 31035 10228 31036 10268
rect 31076 10228 31077 10268
rect 31035 10219 31077 10228
rect 15666 10210 15712 10219
rect 16722 10210 16768 10219
rect 12490 10185 12548 10186
rect 12192 10144 12193 10184
rect 12233 10144 12234 10184
rect 12192 10135 12234 10144
rect 13202 10184 13244 10193
rect 13202 10144 13203 10184
rect 13243 10144 13244 10184
rect 13202 10135 13244 10144
rect 13419 10184 13461 10193
rect 13419 10144 13420 10184
rect 13460 10144 13461 10184
rect 13419 10135 13461 10144
rect 14605 10184 14663 10185
rect 15147 10184 15189 10193
rect 14605 10144 14614 10184
rect 14654 10144 14663 10184
rect 14605 10143 14663 10144
rect 14850 10175 14896 10184
rect 14850 10135 14851 10175
rect 14891 10135 14896 10175
rect 15147 10144 15148 10184
rect 15188 10144 15189 10184
rect 15147 10135 15189 10144
rect 15531 10184 15573 10193
rect 15531 10144 15532 10184
rect 15572 10144 15573 10184
rect 15531 10135 15573 10144
rect 15760 10184 15818 10185
rect 15760 10144 15769 10184
rect 15809 10144 15818 10184
rect 15760 10143 15818 10144
rect 16587 10184 16629 10193
rect 16587 10144 16588 10184
rect 16628 10144 16629 10184
rect 16587 10135 16629 10144
rect 16816 10184 16874 10185
rect 16816 10144 16825 10184
rect 16865 10144 16874 10184
rect 16816 10143 16874 10144
rect 17067 10184 17109 10193
rect 17067 10144 17068 10184
rect 17108 10144 17109 10184
rect 17067 10135 17109 10144
rect 17296 10184 17354 10185
rect 17296 10144 17305 10184
rect 17345 10144 17354 10184
rect 17296 10143 17354 10144
rect 17446 10184 17488 10193
rect 17446 10144 17447 10184
rect 17487 10144 17488 10184
rect 17446 10135 17488 10144
rect 17626 10184 17684 10185
rect 17626 10144 17635 10184
rect 17675 10144 17684 10184
rect 17626 10143 17684 10144
rect 18603 10184 18645 10193
rect 18603 10144 18604 10184
rect 18644 10144 18645 10184
rect 18603 10135 18645 10144
rect 18718 10184 18760 10193
rect 18718 10144 18719 10184
rect 18759 10144 18760 10184
rect 18718 10135 18760 10144
rect 18891 10184 18933 10193
rect 18891 10144 18892 10184
rect 18932 10144 18933 10184
rect 18891 10135 18933 10144
rect 19083 10184 19125 10193
rect 19083 10144 19084 10184
rect 19124 10144 19125 10184
rect 19083 10135 19125 10144
rect 19275 10184 19317 10193
rect 19275 10144 19276 10184
rect 19316 10144 19317 10184
rect 19275 10135 19317 10144
rect 19947 10184 19989 10193
rect 19947 10144 19948 10184
rect 19988 10144 19989 10184
rect 19947 10135 19989 10144
rect 20035 10184 20093 10185
rect 20035 10144 20044 10184
rect 20084 10144 20093 10184
rect 20035 10143 20093 10144
rect 20311 10184 20369 10185
rect 20311 10144 20320 10184
rect 20360 10144 20369 10184
rect 20311 10143 20369 10144
rect 21147 10184 21189 10193
rect 21147 10144 21148 10184
rect 21188 10144 21189 10184
rect 21147 10135 21189 10144
rect 21291 10184 21333 10193
rect 21291 10144 21292 10184
rect 21332 10144 21333 10184
rect 21291 10135 21333 10144
rect 21771 10184 21813 10193
rect 21771 10144 21772 10184
rect 21812 10144 21813 10184
rect 21771 10135 21813 10144
rect 22635 10184 22677 10193
rect 22635 10144 22636 10184
rect 22676 10144 22677 10184
rect 22635 10135 22677 10144
rect 23499 10184 23541 10193
rect 23499 10144 23500 10184
rect 23540 10144 23541 10184
rect 23499 10135 23541 10144
rect 24555 10184 24597 10193
rect 24555 10144 24556 10184
rect 24596 10144 24597 10184
rect 24555 10135 24597 10144
rect 24939 10184 24981 10193
rect 24939 10144 24940 10184
rect 24980 10144 24981 10184
rect 24939 10135 24981 10144
rect 26667 10184 26709 10193
rect 26667 10144 26668 10184
rect 26708 10144 26709 10184
rect 26667 10135 26709 10144
rect 26859 10184 26901 10193
rect 26859 10144 26860 10184
rect 26900 10144 26901 10184
rect 26859 10135 26901 10144
rect 27051 10184 27093 10193
rect 27051 10144 27052 10184
rect 27092 10144 27093 10184
rect 27051 10135 27093 10144
rect 28107 10184 28149 10193
rect 28107 10144 28108 10184
rect 28148 10144 28149 10184
rect 28107 10135 28149 10144
rect 28395 10184 28437 10193
rect 28395 10144 28396 10184
rect 28436 10144 28437 10184
rect 28395 10135 28437 10144
rect 28587 10184 28629 10193
rect 28587 10144 28588 10184
rect 28628 10144 28629 10184
rect 28587 10135 28629 10144
rect 29067 10184 29109 10193
rect 29067 10144 29068 10184
rect 29108 10144 29109 10184
rect 29067 10135 29109 10144
rect 29931 10184 29973 10193
rect 29931 10144 29932 10184
rect 29972 10144 29973 10184
rect 29931 10135 29973 10144
rect 30046 10184 30088 10193
rect 30046 10144 30047 10184
rect 30087 10144 30088 10184
rect 30046 10135 30088 10144
rect 30219 10184 30261 10193
rect 30219 10144 30220 10184
rect 30260 10144 30261 10184
rect 30219 10135 30261 10144
rect 30346 10184 30404 10185
rect 30346 10144 30355 10184
rect 30395 10144 30404 10184
rect 30346 10143 30404 10144
rect 30841 10184 30899 10185
rect 30841 10144 30850 10184
rect 30890 10144 30899 10184
rect 30841 10143 30899 10144
rect 14850 10126 14896 10135
rect 4155 10100 4197 10109
rect 4155 10060 4156 10100
rect 4196 10060 4197 10100
rect 4155 10051 4197 10060
rect 9034 10100 9092 10101
rect 9034 10060 9043 10100
rect 9083 10060 9092 10100
rect 9034 10059 9092 10060
rect 10539 10100 10581 10109
rect 10539 10060 10540 10100
rect 10580 10060 10581 10100
rect 10539 10051 10581 10060
rect 16971 10100 17013 10109
rect 16971 10060 16972 10100
rect 17012 10060 17013 10100
rect 16971 10051 17013 10060
rect 19179 10100 19221 10109
rect 19179 10060 19180 10100
rect 19220 10060 19221 10100
rect 19179 10051 19221 10060
rect 19741 10100 19783 10109
rect 19741 10060 19742 10100
rect 19782 10060 19783 10100
rect 19741 10051 19783 10060
rect 20475 10100 20517 10109
rect 20475 10060 20476 10100
rect 20516 10060 20517 10100
rect 20475 10051 20517 10060
rect 26763 10100 26805 10109
rect 26763 10060 26764 10100
rect 26804 10060 26805 10100
rect 26763 10051 26805 10060
rect 29739 10100 29781 10109
rect 29739 10060 29740 10100
rect 29780 10060 29781 10100
rect 29739 10051 29781 10060
rect 30555 10100 30597 10109
rect 30555 10060 30556 10100
rect 30596 10060 30597 10100
rect 30555 10051 30597 10060
rect 922 10016 980 10017
rect 922 9976 931 10016
rect 971 9976 980 10016
rect 922 9975 980 9976
rect 1707 10016 1749 10025
rect 1707 9976 1708 10016
rect 1748 9976 1749 10016
rect 1707 9967 1749 9976
rect 5835 10016 5877 10025
rect 5835 9976 5836 10016
rect 5876 9976 5877 10016
rect 5835 9967 5877 9976
rect 6699 10016 6741 10025
rect 6699 9976 6700 10016
rect 6740 9976 6741 10016
rect 6699 9967 6741 9976
rect 8218 10016 8276 10017
rect 8218 9976 8227 10016
rect 8267 9976 8276 10016
rect 8218 9975 8276 9976
rect 17547 10016 17589 10025
rect 17547 9976 17548 10016
rect 17588 9976 17589 10016
rect 17547 9967 17589 9976
rect 19834 10016 19892 10017
rect 19834 9976 19843 10016
rect 19883 9976 19892 10016
rect 19834 9975 19892 9976
rect 23307 10016 23349 10025
rect 23307 9976 23308 10016
rect 23348 9976 23349 10016
rect 23307 9967 23349 9976
rect 24171 10016 24213 10025
rect 24171 9976 24172 10016
rect 24212 9976 24213 10016
rect 24171 9967 24213 9976
rect 24442 10016 24500 10017
rect 24442 9976 24451 10016
rect 24491 9976 24500 10016
rect 24442 9975 24500 9976
rect 27435 10016 27477 10025
rect 27435 9976 27436 10016
rect 27476 9976 27477 10016
rect 27435 9967 27477 9976
rect 576 9848 31392 9872
rect 576 9808 4352 9848
rect 4720 9808 12126 9848
rect 12494 9808 19900 9848
rect 20268 9808 27674 9848
rect 28042 9808 31392 9848
rect 576 9784 31392 9808
rect 1594 9680 1652 9681
rect 1594 9640 1603 9680
rect 1643 9640 1652 9680
rect 1594 9639 1652 9640
rect 1899 9680 1941 9689
rect 1899 9640 1900 9680
rect 1940 9640 1941 9680
rect 1899 9631 1941 9640
rect 2842 9680 2900 9681
rect 2842 9640 2851 9680
rect 2891 9640 2900 9680
rect 2842 9639 2900 9640
rect 5835 9680 5877 9689
rect 5835 9640 5836 9680
rect 5876 9640 5877 9680
rect 5835 9631 5877 9640
rect 6394 9680 6452 9681
rect 6394 9640 6403 9680
rect 6443 9640 6452 9680
rect 6394 9639 6452 9640
rect 7450 9680 7508 9681
rect 7450 9640 7459 9680
rect 7499 9640 7508 9680
rect 7450 9639 7508 9640
rect 8410 9680 8468 9681
rect 8410 9640 8419 9680
rect 8459 9640 8468 9680
rect 8410 9639 8468 9640
rect 8523 9680 8565 9689
rect 8523 9640 8524 9680
rect 8564 9640 8565 9680
rect 8523 9631 8565 9640
rect 8907 9680 8949 9689
rect 8907 9640 8908 9680
rect 8948 9640 8949 9680
rect 8907 9631 8949 9640
rect 10474 9680 10532 9681
rect 10474 9640 10483 9680
rect 10523 9640 10532 9680
rect 10474 9639 10532 9640
rect 11098 9680 11156 9681
rect 11098 9640 11107 9680
rect 11147 9640 11156 9680
rect 11098 9639 11156 9640
rect 11770 9680 11828 9681
rect 11770 9640 11779 9680
rect 11819 9640 11828 9680
rect 11770 9639 11828 9640
rect 13588 9680 13646 9681
rect 13588 9640 13597 9680
rect 13637 9640 13646 9680
rect 13588 9639 13646 9640
rect 14427 9680 14469 9689
rect 14427 9640 14428 9680
rect 14468 9640 14469 9680
rect 14427 9631 14469 9640
rect 15531 9680 15573 9689
rect 15531 9640 15532 9680
rect 15572 9640 15573 9680
rect 15531 9631 15573 9640
rect 15963 9680 16005 9689
rect 15963 9640 15964 9680
rect 16004 9640 16005 9680
rect 15963 9631 16005 9640
rect 18826 9680 18884 9681
rect 18826 9640 18835 9680
rect 18875 9640 18884 9680
rect 18826 9639 18884 9640
rect 19371 9680 19413 9689
rect 19371 9640 19372 9680
rect 19412 9640 19413 9680
rect 19371 9631 19413 9640
rect 20523 9680 20565 9689
rect 20523 9640 20524 9680
rect 20564 9640 20565 9680
rect 20523 9631 20565 9640
rect 25611 9680 25653 9689
rect 25611 9640 25612 9680
rect 25652 9640 25653 9680
rect 25611 9631 25653 9640
rect 27610 9680 27668 9681
rect 27610 9640 27619 9680
rect 27659 9640 27668 9680
rect 27610 9639 27668 9640
rect 27723 9680 27765 9689
rect 27723 9640 27724 9680
rect 27764 9640 27765 9680
rect 27723 9631 27765 9640
rect 28779 9680 28821 9689
rect 28779 9640 28780 9680
rect 28820 9640 28821 9680
rect 28779 9631 28821 9640
rect 28971 9680 29013 9689
rect 28971 9640 28972 9680
rect 29012 9640 29013 9680
rect 28971 9631 29013 9640
rect 2955 9596 2997 9605
rect 2955 9556 2956 9596
rect 2996 9556 2997 9596
rect 2955 9547 2997 9556
rect 6617 9596 6659 9605
rect 6617 9556 6618 9596
rect 6658 9556 6659 9596
rect 6617 9547 6659 9556
rect 6891 9596 6933 9605
rect 6891 9556 6892 9596
rect 6932 9556 6933 9596
rect 6891 9547 6933 9556
rect 7851 9596 7893 9605
rect 7851 9556 7852 9596
rect 7892 9556 7893 9596
rect 7851 9547 7893 9556
rect 8320 9596 8362 9605
rect 8320 9556 8321 9596
rect 8361 9556 8362 9596
rect 8320 9547 8362 9556
rect 11211 9596 11253 9605
rect 11211 9556 11212 9596
rect 11252 9556 11253 9596
rect 11211 9547 11253 9556
rect 11931 9596 11973 9605
rect 11931 9556 11932 9596
rect 11972 9556 11973 9596
rect 11931 9547 11973 9556
rect 20122 9596 20180 9597
rect 20122 9556 20131 9596
rect 20171 9556 20180 9596
rect 20122 9555 20180 9556
rect 24202 9596 24260 9597
rect 24202 9556 24211 9596
rect 24251 9556 24260 9596
rect 24202 9555 24260 9556
rect 31258 9596 31316 9597
rect 31258 9556 31267 9596
rect 31307 9556 31316 9596
rect 31258 9555 31316 9556
rect 1114 9512 1172 9513
rect 1114 9472 1123 9512
rect 1163 9472 1172 9512
rect 1114 9471 1172 9472
rect 1419 9512 1461 9521
rect 1419 9472 1420 9512
rect 1460 9472 1461 9512
rect 1419 9463 1461 9472
rect 1707 9512 1749 9521
rect 1707 9472 1708 9512
rect 1748 9472 1749 9512
rect 1707 9463 1749 9472
rect 2050 9512 2108 9513
rect 2050 9472 2059 9512
rect 2099 9472 2108 9512
rect 2050 9471 2108 9472
rect 2344 9512 2386 9521
rect 2344 9472 2345 9512
rect 2385 9472 2386 9512
rect 2344 9463 2386 9472
rect 2506 9512 2564 9513
rect 2506 9472 2515 9512
rect 2555 9472 2564 9512
rect 2506 9471 2564 9472
rect 2746 9512 2804 9513
rect 2746 9472 2755 9512
rect 2795 9472 2804 9512
rect 2746 9471 2804 9472
rect 3062 9512 3104 9521
rect 3062 9472 3063 9512
rect 3103 9472 3104 9512
rect 3062 9463 3104 9472
rect 5931 9512 5973 9521
rect 5931 9472 5932 9512
rect 5972 9472 5973 9512
rect 5931 9463 5973 9472
rect 6148 9512 6190 9521
rect 6148 9472 6149 9512
rect 6189 9472 6190 9512
rect 6148 9463 6190 9472
rect 6298 9512 6356 9513
rect 6298 9472 6307 9512
rect 6347 9472 6356 9512
rect 6298 9471 6356 9472
rect 6411 9512 6453 9521
rect 6411 9472 6412 9512
rect 6452 9472 6453 9512
rect 6411 9463 6453 9472
rect 6795 9512 6837 9521
rect 6795 9472 6796 9512
rect 6836 9472 6837 9512
rect 6795 9463 6837 9472
rect 6970 9512 7028 9513
rect 6970 9472 6979 9512
rect 7019 9472 7028 9512
rect 6970 9471 7028 9472
rect 7126 9512 7168 9521
rect 7126 9472 7127 9512
rect 7167 9472 7168 9512
rect 7126 9463 7168 9472
rect 7371 9512 7413 9521
rect 7371 9472 7372 9512
rect 7412 9472 7413 9512
rect 7371 9463 7413 9472
rect 7947 9512 7989 9521
rect 7947 9472 7948 9512
rect 7988 9472 7989 9512
rect 7947 9463 7989 9472
rect 8181 9512 8223 9521
rect 8811 9512 8853 9521
rect 8181 9472 8182 9512
rect 8222 9472 8223 9512
rect 8181 9463 8223 9472
rect 8619 9503 8661 9512
rect 8619 9463 8620 9503
rect 8660 9463 8661 9503
rect 8811 9472 8812 9512
rect 8852 9472 8853 9512
rect 8811 9463 8853 9472
rect 9003 9512 9045 9521
rect 9003 9472 9004 9512
rect 9044 9472 9045 9512
rect 9003 9463 9045 9472
rect 10639 9512 10697 9513
rect 10639 9472 10648 9512
rect 10688 9472 10697 9512
rect 10639 9471 10697 9472
rect 11005 9512 11047 9521
rect 11446 9512 11488 9521
rect 11005 9472 11006 9512
rect 11046 9472 11047 9512
rect 11005 9463 11047 9472
rect 11307 9503 11349 9512
rect 11307 9463 11308 9503
rect 11348 9463 11349 9503
rect 11446 9472 11447 9512
rect 11487 9472 11488 9512
rect 11446 9463 11488 9472
rect 11691 9512 11733 9521
rect 11691 9472 11692 9512
rect 11732 9472 11733 9512
rect 11691 9463 11733 9472
rect 12075 9512 12117 9521
rect 12075 9472 12076 9512
rect 12116 9472 12117 9512
rect 12075 9463 12117 9472
rect 12843 9512 12885 9521
rect 12843 9472 12844 9512
rect 12884 9472 12885 9512
rect 12843 9463 12885 9472
rect 13227 9512 13269 9521
rect 13227 9472 13228 9512
rect 13268 9472 13269 9512
rect 13227 9463 13269 9472
rect 13690 9512 13748 9513
rect 15435 9512 15477 9521
rect 13690 9472 13699 9512
rect 13739 9472 13748 9512
rect 13690 9471 13748 9472
rect 13803 9503 13845 9512
rect 13803 9463 13804 9503
rect 13844 9463 13845 9503
rect 8619 9454 8661 9463
rect 11307 9454 11349 9463
rect 13803 9454 13845 9463
rect 14274 9503 14320 9512
rect 14274 9463 14275 9503
rect 14315 9463 14320 9503
rect 14274 9454 14320 9463
rect 14754 9503 14800 9512
rect 14754 9463 14755 9503
rect 14795 9463 14800 9503
rect 15435 9472 15436 9512
rect 15476 9472 15477 9512
rect 15435 9463 15477 9472
rect 15610 9512 15668 9513
rect 16587 9512 16629 9521
rect 15610 9472 15619 9512
rect 15659 9472 15668 9512
rect 15610 9471 15668 9472
rect 15810 9503 15856 9512
rect 15810 9463 15811 9503
rect 15851 9463 15856 9503
rect 16587 9472 16588 9512
rect 16628 9472 16629 9512
rect 16587 9463 16629 9472
rect 16702 9512 16744 9521
rect 16702 9472 16703 9512
rect 16743 9472 16744 9512
rect 16702 9463 16744 9472
rect 16875 9512 16917 9521
rect 16875 9472 16876 9512
rect 16916 9472 16917 9512
rect 16875 9463 16917 9472
rect 17590 9512 17632 9521
rect 17590 9472 17591 9512
rect 17631 9472 17632 9512
rect 17590 9463 17632 9472
rect 17835 9512 17877 9521
rect 17835 9472 17836 9512
rect 17876 9472 17877 9512
rect 17835 9463 17877 9472
rect 19021 9512 19079 9513
rect 19021 9472 19030 9512
rect 19070 9472 19079 9512
rect 19021 9471 19079 9472
rect 19467 9512 19509 9521
rect 19467 9472 19468 9512
rect 19508 9472 19509 9512
rect 19810 9512 19868 9513
rect 19467 9463 19509 9472
rect 19707 9470 19749 9479
rect 19810 9472 19819 9512
rect 19859 9472 19868 9512
rect 19810 9471 19868 9472
rect 20028 9512 20086 9513
rect 20028 9472 20037 9512
rect 20077 9472 20086 9512
rect 20028 9471 20086 9472
rect 22426 9512 22484 9513
rect 22426 9472 22435 9512
rect 22475 9472 22484 9512
rect 22426 9471 22484 9472
rect 23407 9512 23465 9513
rect 23407 9472 23416 9512
rect 23456 9472 23465 9512
rect 23407 9471 23465 9472
rect 23595 9512 23637 9521
rect 23595 9472 23596 9512
rect 23636 9472 23637 9512
rect 14754 9454 14800 9463
rect 15810 9454 15856 9463
rect 2187 9428 2229 9437
rect 2187 9388 2188 9428
rect 2228 9388 2229 9428
rect 2187 9379 2229 9388
rect 6050 9428 6092 9437
rect 6050 9388 6051 9428
rect 6091 9388 6092 9428
rect 6050 9379 6092 9388
rect 7258 9428 7316 9429
rect 11578 9428 11636 9429
rect 7258 9388 7267 9428
rect 7307 9388 7316 9428
rect 7258 9387 7316 9388
rect 8082 9419 8128 9428
rect 8082 9379 8083 9419
rect 8123 9379 8128 9419
rect 11578 9388 11587 9428
rect 11627 9388 11636 9428
rect 11578 9387 11636 9388
rect 14907 9428 14949 9437
rect 14907 9388 14908 9428
rect 14948 9388 14949 9428
rect 14907 9379 14949 9388
rect 17722 9428 17780 9429
rect 17722 9388 17731 9428
rect 17771 9388 17780 9428
rect 17722 9387 17780 9388
rect 17931 9428 17973 9437
rect 17931 9388 17932 9428
rect 17972 9388 17973 9428
rect 17931 9379 17973 9388
rect 19586 9428 19628 9437
rect 19586 9388 19587 9428
rect 19627 9388 19628 9428
rect 19707 9430 19708 9470
rect 19748 9430 19749 9470
rect 23595 9463 23637 9472
rect 23770 9512 23828 9513
rect 23770 9472 23779 9512
rect 23819 9472 23828 9512
rect 23770 9471 23828 9472
rect 24367 9512 24425 9513
rect 24367 9472 24376 9512
rect 24416 9472 24425 9512
rect 25803 9512 25845 9521
rect 24367 9471 24425 9472
rect 24854 9485 24896 9494
rect 24854 9445 24855 9485
rect 24895 9445 24896 9485
rect 25803 9472 25804 9512
rect 25844 9472 25845 9512
rect 25803 9463 25845 9472
rect 26091 9512 26133 9521
rect 26091 9472 26092 9512
rect 26132 9472 26133 9512
rect 26091 9463 26133 9472
rect 26205 9512 26263 9513
rect 26205 9472 26214 9512
rect 26254 9472 26263 9512
rect 26205 9471 26263 9472
rect 26332 9512 26390 9513
rect 26332 9472 26341 9512
rect 26381 9472 26390 9512
rect 26332 9471 26390 9472
rect 26571 9512 26613 9521
rect 26571 9472 26572 9512
rect 26612 9472 26613 9512
rect 26571 9463 26613 9472
rect 26746 9512 26804 9513
rect 26746 9472 26755 9512
rect 26795 9472 26804 9512
rect 26746 9471 26804 9472
rect 26859 9512 26901 9521
rect 26859 9472 26860 9512
rect 26900 9472 26901 9512
rect 26859 9463 26901 9472
rect 27370 9512 27428 9513
rect 27370 9472 27379 9512
rect 27419 9472 27428 9512
rect 27370 9471 27428 9472
rect 27514 9512 27572 9513
rect 27514 9472 27523 9512
rect 27563 9472 27572 9512
rect 27514 9471 27572 9472
rect 27833 9512 27875 9521
rect 27833 9472 27834 9512
rect 27874 9472 27875 9512
rect 28618 9512 28676 9513
rect 27833 9463 27875 9472
rect 28480 9485 28522 9494
rect 19707 9421 19749 9430
rect 19924 9428 19966 9437
rect 19586 9379 19628 9388
rect 19924 9388 19925 9428
rect 19965 9388 19966 9428
rect 19924 9379 19966 9388
rect 20890 9428 20948 9429
rect 20890 9388 20899 9428
rect 20939 9388 20948 9428
rect 20890 9387 20948 9388
rect 22810 9428 22868 9429
rect 22810 9388 22819 9428
rect 22859 9388 22868 9428
rect 22810 9387 22868 9388
rect 23242 9428 23300 9429
rect 23242 9388 23251 9428
rect 23291 9388 23300 9428
rect 23242 9387 23300 9388
rect 24753 9428 24795 9437
rect 24854 9436 24896 9445
rect 28480 9445 28481 9485
rect 28521 9445 28522 9485
rect 28618 9472 28627 9512
rect 28667 9472 28676 9512
rect 28618 9471 28676 9472
rect 30874 9512 30932 9513
rect 30874 9472 30883 9512
rect 30923 9472 30932 9512
rect 30874 9471 30932 9472
rect 28480 9436 28522 9445
rect 24753 9388 24754 9428
rect 24794 9388 24795 9428
rect 24753 9379 24795 9388
rect 27178 9428 27236 9429
rect 27178 9388 27187 9428
rect 27227 9388 27236 9428
rect 27178 9387 27236 9388
rect 29338 9428 29396 9429
rect 29338 9388 29347 9428
rect 29387 9388 29396 9428
rect 29338 9387 29396 9388
rect 8082 9370 8128 9379
rect 2283 9344 2325 9353
rect 2283 9304 2284 9344
rect 2324 9304 2325 9344
rect 2283 9295 2325 9304
rect 16587 9344 16629 9353
rect 16587 9304 16588 9344
rect 16628 9304 16629 9344
rect 16587 9295 16629 9304
rect 26379 9344 26421 9353
rect 26379 9304 26380 9344
rect 26420 9304 26421 9344
rect 26379 9295 26421 9304
rect 1419 9260 1461 9269
rect 1419 9220 1420 9260
rect 1460 9220 1461 9260
rect 1419 9211 1461 9220
rect 6603 9260 6645 9269
rect 6603 9220 6604 9260
rect 6644 9220 6645 9260
rect 6603 9211 6645 9220
rect 13467 9260 13509 9269
rect 13467 9220 13468 9260
rect 13508 9220 13509 9260
rect 13467 9211 13509 9220
rect 14091 9260 14133 9269
rect 14091 9220 14092 9260
rect 14132 9220 14133 9260
rect 14091 9211 14133 9220
rect 23770 9260 23828 9261
rect 23770 9220 23779 9260
rect 23819 9220 23828 9260
rect 23770 9219 23828 9220
rect 24651 9260 24693 9269
rect 24651 9220 24652 9260
rect 24692 9220 24693 9260
rect 24651 9211 24693 9220
rect 26859 9260 26901 9269
rect 26859 9220 26860 9260
rect 26900 9220 26901 9260
rect 26859 9211 26901 9220
rect 576 9092 31392 9116
rect 576 9052 3112 9092
rect 3480 9052 10886 9092
rect 11254 9052 18660 9092
rect 19028 9052 26434 9092
rect 26802 9052 31392 9092
rect 576 9028 31392 9052
rect 1210 8924 1268 8925
rect 1210 8884 1219 8924
rect 1259 8884 1268 8924
rect 1210 8883 1268 8884
rect 3898 8924 3956 8925
rect 3898 8884 3907 8924
rect 3947 8884 3956 8924
rect 3898 8883 3956 8884
rect 4875 8924 4917 8933
rect 4875 8884 4876 8924
rect 4916 8884 4917 8924
rect 4875 8875 4917 8884
rect 5626 8924 5684 8925
rect 5626 8884 5635 8924
rect 5675 8884 5684 8924
rect 5626 8883 5684 8884
rect 8314 8924 8372 8925
rect 8314 8884 8323 8924
rect 8363 8884 8372 8924
rect 8314 8883 8372 8884
rect 12651 8924 12693 8933
rect 12651 8884 12652 8924
rect 12692 8884 12693 8924
rect 12651 8875 12693 8884
rect 13899 8924 13941 8933
rect 13899 8884 13900 8924
rect 13940 8884 13941 8924
rect 13899 8875 13941 8884
rect 14458 8924 14516 8925
rect 14458 8884 14467 8924
rect 14507 8884 14516 8924
rect 14458 8883 14516 8884
rect 20026 8924 20084 8925
rect 20026 8884 20035 8924
rect 20075 8884 20084 8924
rect 20026 8883 20084 8884
rect 23451 8924 23493 8933
rect 23451 8884 23452 8924
rect 23492 8884 23493 8924
rect 23451 8875 23493 8884
rect 27099 8924 27141 8933
rect 27099 8884 27100 8924
rect 27140 8884 27141 8924
rect 27099 8875 27141 8884
rect 28971 8924 29013 8933
rect 28971 8884 28972 8924
rect 29012 8884 29013 8924
rect 28971 8875 29013 8884
rect 29931 8924 29973 8933
rect 29931 8884 29932 8924
rect 29972 8884 29973 8924
rect 29931 8875 29973 8884
rect 11194 8840 11252 8841
rect 19851 8840 19893 8849
rect 11194 8800 11203 8840
rect 11243 8800 11252 8840
rect 11194 8799 11252 8800
rect 17787 8831 17829 8840
rect 17787 8791 17788 8831
rect 17828 8791 17829 8831
rect 19851 8800 19852 8840
rect 19892 8800 19893 8840
rect 19851 8791 19893 8800
rect 21771 8840 21813 8849
rect 21771 8800 21772 8840
rect 21812 8800 21813 8840
rect 21771 8791 21813 8800
rect 26571 8840 26613 8849
rect 26571 8800 26572 8840
rect 26612 8800 26613 8840
rect 26571 8791 26613 8800
rect 31083 8840 31125 8849
rect 31083 8800 31084 8840
rect 31124 8800 31125 8840
rect 31083 8791 31125 8800
rect 17787 8782 17829 8791
rect 2554 8756 2612 8757
rect 2554 8716 2563 8756
rect 2603 8716 2612 8756
rect 2554 8715 2612 8716
rect 2763 8756 2805 8765
rect 2763 8716 2764 8756
rect 2804 8716 2805 8756
rect 2763 8707 2805 8716
rect 4977 8756 5019 8765
rect 4977 8716 4978 8756
rect 5018 8716 5019 8756
rect 4977 8707 5019 8716
rect 9195 8756 9237 8765
rect 9195 8716 9196 8756
rect 9236 8716 9237 8756
rect 9195 8707 9237 8716
rect 11578 8756 11636 8757
rect 11578 8716 11587 8756
rect 11627 8716 11636 8756
rect 11578 8715 11636 8716
rect 11787 8756 11829 8765
rect 11787 8716 11788 8756
rect 11828 8716 11829 8756
rect 11787 8707 11829 8716
rect 15531 8756 15573 8765
rect 15531 8716 15532 8756
rect 15572 8716 15573 8756
rect 12367 8705 12409 8714
rect 15531 8707 15573 8716
rect 15746 8756 15788 8765
rect 18219 8756 18261 8765
rect 30033 8756 30075 8765
rect 15746 8716 15747 8756
rect 15787 8716 15788 8756
rect 15746 8707 15788 8716
rect 17202 8747 17248 8756
rect 17202 8707 17203 8747
rect 17243 8707 17248 8747
rect 18219 8716 18220 8756
rect 18260 8716 18261 8756
rect 18219 8707 18261 8716
rect 18450 8747 18496 8756
rect 18450 8707 18451 8747
rect 18491 8707 18496 8747
rect 30033 8716 30034 8756
rect 30074 8716 30075 8756
rect 1611 8672 1653 8681
rect 1611 8632 1612 8672
rect 1652 8632 1653 8672
rect 1611 8623 1653 8632
rect 2091 8672 2133 8681
rect 2091 8632 2092 8672
rect 2132 8632 2133 8672
rect 2091 8623 2133 8632
rect 2283 8672 2325 8681
rect 2283 8632 2284 8672
rect 2324 8632 2325 8672
rect 2283 8623 2325 8632
rect 2422 8672 2464 8681
rect 2422 8632 2423 8672
rect 2463 8632 2464 8672
rect 2422 8623 2464 8632
rect 2667 8672 2709 8681
rect 2667 8632 2668 8672
rect 2708 8632 2709 8672
rect 2667 8623 2709 8632
rect 2938 8672 2996 8673
rect 2938 8632 2947 8672
rect 2987 8632 2996 8672
rect 2938 8631 2996 8632
rect 3243 8672 3285 8681
rect 3243 8632 3244 8672
rect 3284 8632 3285 8672
rect 3243 8623 3285 8632
rect 3610 8672 3668 8673
rect 3610 8632 3619 8672
rect 3659 8632 3668 8672
rect 3610 8631 3668 8632
rect 3723 8672 3765 8681
rect 3723 8632 3724 8672
rect 3764 8632 3765 8672
rect 3723 8623 3765 8632
rect 4186 8672 4244 8673
rect 4186 8632 4195 8672
rect 4235 8632 4244 8672
rect 4186 8631 4244 8632
rect 4299 8672 4341 8681
rect 4299 8632 4300 8672
rect 4340 8632 4341 8672
rect 4299 8623 4341 8632
rect 5067 8672 5109 8681
rect 5067 8632 5068 8672
rect 5108 8632 5109 8672
rect 5067 8623 5109 8632
rect 6027 8672 6069 8681
rect 6027 8632 6028 8672
rect 6068 8632 6069 8672
rect 6027 8623 6069 8632
rect 6874 8672 6932 8673
rect 6874 8632 6883 8672
rect 6923 8632 6932 8672
rect 6874 8631 6932 8632
rect 6987 8672 7029 8681
rect 6987 8632 6988 8672
rect 7028 8632 7029 8672
rect 6987 8623 7029 8632
rect 8026 8672 8084 8673
rect 8026 8632 8035 8672
rect 8075 8632 8084 8672
rect 8026 8631 8084 8632
rect 8139 8672 8181 8681
rect 8139 8632 8140 8672
rect 8180 8632 8181 8672
rect 8139 8623 8181 8632
rect 8698 8672 8756 8673
rect 8698 8632 8707 8672
rect 8747 8632 8756 8672
rect 8698 8631 8756 8632
rect 8811 8672 8853 8681
rect 8811 8632 8812 8672
rect 8852 8632 8853 8672
rect 8811 8623 8853 8632
rect 9291 8672 9333 8681
rect 9291 8632 9292 8672
rect 9332 8632 9333 8672
rect 9291 8623 9333 8632
rect 9763 8672 9821 8673
rect 9763 8632 9772 8672
rect 9812 8632 9821 8672
rect 9763 8631 9821 8632
rect 10282 8672 10340 8673
rect 10282 8632 10291 8672
rect 10331 8632 10340 8672
rect 10282 8631 10340 8632
rect 10906 8672 10964 8673
rect 10906 8632 10915 8672
rect 10955 8632 10964 8672
rect 10906 8631 10964 8632
rect 11019 8672 11061 8681
rect 11019 8632 11020 8672
rect 11060 8632 11061 8672
rect 11019 8623 11061 8632
rect 11458 8672 11516 8673
rect 11458 8632 11467 8672
rect 11507 8632 11516 8672
rect 11458 8631 11516 8632
rect 11691 8672 11733 8681
rect 11691 8632 11692 8672
rect 11732 8632 11733 8672
rect 11691 8623 11733 8632
rect 12250 8672 12308 8673
rect 12250 8632 12259 8672
rect 12299 8632 12308 8672
rect 12367 8665 12368 8705
rect 12408 8665 12409 8705
rect 17202 8698 17248 8707
rect 18450 8698 18496 8707
rect 24634 8714 24692 8715
rect 16299 8683 16341 8692
rect 12367 8656 12409 8665
rect 13594 8672 13652 8673
rect 12250 8631 12308 8632
rect 13594 8632 13603 8672
rect 13643 8632 13652 8672
rect 13594 8631 13652 8632
rect 13707 8672 13749 8681
rect 13707 8632 13708 8672
rect 13748 8632 13749 8672
rect 13707 8623 13749 8632
rect 14755 8672 14813 8673
rect 14755 8632 14764 8672
rect 14804 8632 14813 8672
rect 14755 8631 14813 8632
rect 15031 8672 15089 8673
rect 15031 8632 15040 8672
rect 15080 8632 15089 8672
rect 15031 8631 15089 8632
rect 15627 8672 15669 8681
rect 15627 8632 15628 8672
rect 15668 8632 15669 8672
rect 15627 8623 15669 8632
rect 15856 8672 15914 8673
rect 15856 8632 15865 8672
rect 15905 8632 15914 8672
rect 15856 8631 15914 8632
rect 16186 8672 16244 8673
rect 16186 8632 16195 8672
rect 16235 8632 16244 8672
rect 16299 8643 16300 8683
rect 16340 8643 16341 8683
rect 16299 8634 16341 8643
rect 16436 8672 16494 8673
rect 16186 8631 16244 8632
rect 16436 8632 16445 8672
rect 16485 8632 16494 8672
rect 16436 8631 16494 8632
rect 16566 8672 16624 8673
rect 16566 8632 16575 8672
rect 16615 8632 16624 8672
rect 16566 8631 16624 8632
rect 16704 8672 16762 8673
rect 16704 8632 16713 8672
rect 16753 8632 16762 8672
rect 16704 8631 16762 8632
rect 17067 8672 17109 8681
rect 17067 8632 17068 8672
rect 17108 8632 17109 8672
rect 17067 8623 17109 8632
rect 17296 8672 17354 8673
rect 17296 8632 17305 8672
rect 17345 8632 17354 8672
rect 17296 8631 17354 8632
rect 17818 8672 17876 8673
rect 17818 8632 17827 8672
rect 17867 8632 17876 8672
rect 17818 8631 17876 8632
rect 18314 8672 18356 8681
rect 18314 8632 18315 8672
rect 18355 8632 18356 8672
rect 18314 8623 18356 8632
rect 18544 8672 18602 8673
rect 18544 8632 18553 8672
rect 18593 8632 18602 8672
rect 18544 8631 18602 8632
rect 19179 8672 19221 8681
rect 19179 8632 19180 8672
rect 19220 8632 19221 8672
rect 19179 8623 19221 8632
rect 19450 8672 19508 8673
rect 19450 8632 19459 8672
rect 19499 8632 19508 8672
rect 19450 8631 19508 8632
rect 20235 8672 20277 8681
rect 20235 8632 20236 8672
rect 20276 8632 20277 8672
rect 20235 8623 20277 8632
rect 20329 8672 20387 8673
rect 20329 8632 20338 8672
rect 20378 8632 20387 8672
rect 20329 8631 20387 8632
rect 23787 8672 23829 8681
rect 23787 8632 23788 8672
rect 23828 8632 23829 8672
rect 23787 8623 23829 8632
rect 24075 8672 24117 8681
rect 24075 8632 24076 8672
rect 24116 8632 24117 8672
rect 24075 8623 24117 8632
rect 24454 8672 24496 8681
rect 24634 8674 24643 8714
rect 24683 8674 24692 8714
rect 30033 8707 30075 8716
rect 24634 8673 24692 8674
rect 24454 8632 24455 8672
rect 24495 8632 24496 8672
rect 24454 8623 24496 8632
rect 24843 8672 24885 8681
rect 24843 8632 24844 8672
rect 24884 8632 24885 8672
rect 24843 8623 24885 8632
rect 26955 8672 26997 8681
rect 26955 8632 26956 8672
rect 26996 8632 26997 8672
rect 26955 8623 26997 8632
rect 28107 8672 28149 8681
rect 28107 8632 28108 8672
rect 28148 8632 28149 8672
rect 28107 8623 28149 8632
rect 29643 8672 29685 8681
rect 29643 8632 29644 8672
rect 29684 8632 29685 8672
rect 29643 8623 29685 8632
rect 30123 8672 30165 8681
rect 30123 8632 30124 8672
rect 30164 8632 30165 8672
rect 30123 8623 30165 8632
rect 30538 8672 30596 8673
rect 30538 8632 30547 8672
rect 30587 8632 30596 8672
rect 30538 8631 30596 8632
rect 4502 8588 4544 8597
rect 4502 8548 4503 8588
rect 4543 8548 4544 8588
rect 4502 8539 4544 8548
rect 5722 8588 5780 8589
rect 5722 8548 5731 8588
rect 5771 8548 5780 8588
rect 5722 8547 5780 8548
rect 13913 8588 13955 8597
rect 13913 8548 13914 8588
rect 13954 8548 13955 8588
rect 13913 8539 13955 8548
rect 14464 8588 14506 8597
rect 14464 8548 14465 8588
rect 14505 8548 14506 8588
rect 14464 8539 14506 8548
rect 18027 8588 18069 8597
rect 18027 8548 18028 8588
rect 18068 8548 18069 8588
rect 18027 8539 18069 8548
rect 19563 8588 19605 8597
rect 19563 8548 19564 8588
rect 19604 8548 19605 8588
rect 19563 8539 19605 8548
rect 20029 8588 20071 8597
rect 20029 8548 20030 8588
rect 20070 8548 20071 8588
rect 20029 8539 20071 8548
rect 24555 8588 24597 8597
rect 24555 8548 24556 8588
rect 24596 8548 24597 8588
rect 24555 8539 24597 8548
rect 2266 8504 2324 8505
rect 2266 8464 2275 8504
rect 2315 8464 2324 8504
rect 2266 8463 2324 8464
rect 3147 8504 3189 8513
rect 3147 8464 3148 8504
rect 3188 8464 3189 8504
rect 3147 8455 3189 8464
rect 4395 8504 4437 8513
rect 4395 8464 4396 8504
rect 4436 8464 4437 8504
rect 4395 8455 4437 8464
rect 7275 8504 7317 8513
rect 7275 8464 7276 8504
rect 7316 8464 7317 8504
rect 7275 8455 7317 8464
rect 10443 8504 10485 8513
rect 14667 8504 14709 8513
rect 10443 8464 10444 8504
rect 10484 8464 10485 8504
rect 10443 8455 10485 8464
rect 12162 8495 12208 8504
rect 12162 8455 12163 8495
rect 12203 8455 12208 8495
rect 14667 8464 14668 8504
rect 14708 8464 14709 8504
rect 14667 8455 14709 8464
rect 15195 8504 15237 8513
rect 15195 8464 15196 8504
rect 15236 8464 15237 8504
rect 15195 8455 15237 8464
rect 16666 8504 16724 8505
rect 16666 8464 16675 8504
rect 16715 8464 16724 8504
rect 16666 8463 16724 8464
rect 16971 8504 17013 8513
rect 16971 8464 16972 8504
rect 17012 8464 17013 8504
rect 16971 8455 17013 8464
rect 28779 8504 28821 8513
rect 28779 8464 28780 8504
rect 28820 8464 28821 8504
rect 28779 8455 28821 8464
rect 30747 8504 30789 8513
rect 30747 8464 30748 8504
rect 30788 8464 30789 8504
rect 30747 8455 30789 8464
rect 12162 8446 12208 8455
rect 576 8336 31392 8360
rect 576 8296 4352 8336
rect 4720 8296 12126 8336
rect 12494 8296 19900 8336
rect 20268 8296 27674 8336
rect 28042 8296 31392 8336
rect 576 8272 31392 8296
rect 2475 8168 2517 8177
rect 2475 8128 2476 8168
rect 2516 8128 2517 8168
rect 2475 8119 2517 8128
rect 3226 8168 3284 8169
rect 3226 8128 3235 8168
rect 3275 8128 3284 8168
rect 3226 8127 3284 8128
rect 4186 8168 4244 8169
rect 4186 8128 4195 8168
rect 4235 8128 4244 8168
rect 4186 8127 4244 8128
rect 4491 8168 4533 8177
rect 4491 8128 4492 8168
rect 4532 8128 4533 8168
rect 4491 8119 4533 8128
rect 5163 8168 5205 8177
rect 5163 8128 5164 8168
rect 5204 8128 5205 8168
rect 5163 8119 5205 8128
rect 5386 8168 5444 8169
rect 5386 8128 5395 8168
rect 5435 8128 5444 8168
rect 5386 8127 5444 8128
rect 6987 8168 7029 8177
rect 6987 8128 6988 8168
rect 7028 8128 7029 8168
rect 6987 8119 7029 8128
rect 7450 8168 7508 8169
rect 7450 8128 7459 8168
rect 7499 8128 7508 8168
rect 7450 8127 7508 8128
rect 11866 8168 11924 8169
rect 11866 8128 11875 8168
rect 11915 8128 11924 8168
rect 11866 8127 11924 8128
rect 12250 8168 12308 8169
rect 12250 8128 12259 8168
rect 12299 8128 12308 8168
rect 12250 8127 12308 8128
rect 13323 8168 13365 8177
rect 13323 8128 13324 8168
rect 13364 8128 13365 8168
rect 13323 8119 13365 8128
rect 13899 8168 13941 8177
rect 13899 8128 13900 8168
rect 13940 8128 13941 8168
rect 13899 8119 13941 8128
rect 16587 8168 16629 8177
rect 16587 8128 16588 8168
rect 16628 8128 16629 8168
rect 16587 8119 16629 8128
rect 16875 8168 16917 8177
rect 16875 8128 16876 8168
rect 16916 8128 16917 8168
rect 16875 8119 16917 8128
rect 18010 8168 18068 8169
rect 18010 8128 18019 8168
rect 18059 8128 18068 8168
rect 18010 8127 18068 8128
rect 18123 8168 18165 8177
rect 18123 8128 18124 8168
rect 18164 8128 18165 8168
rect 18123 8119 18165 8128
rect 18411 8168 18453 8177
rect 18411 8128 18412 8168
rect 18452 8128 18453 8168
rect 18411 8119 18453 8128
rect 19354 8168 19412 8169
rect 19354 8128 19363 8168
rect 19403 8128 19412 8168
rect 19354 8127 19412 8128
rect 19467 8168 19509 8177
rect 19467 8128 19468 8168
rect 19508 8128 19509 8168
rect 19467 8119 19509 8128
rect 19738 8168 19796 8169
rect 19738 8128 19747 8168
rect 19787 8128 19796 8168
rect 19738 8127 19796 8128
rect 22059 8168 22101 8177
rect 22059 8128 22060 8168
rect 22100 8128 22101 8168
rect 22059 8119 22101 8128
rect 25419 8168 25461 8177
rect 25419 8128 25420 8168
rect 25460 8128 25461 8168
rect 25419 8119 25461 8128
rect 27915 8168 27957 8177
rect 27915 8128 27916 8168
rect 27956 8128 27957 8168
rect 27915 8119 27957 8128
rect 29163 8168 29205 8177
rect 29163 8128 29164 8168
rect 29204 8128 29205 8168
rect 29163 8119 29205 8128
rect 30123 8168 30165 8177
rect 30123 8128 30124 8168
rect 30164 8128 30165 8168
rect 30123 8119 30165 8128
rect 7755 8084 7797 8093
rect 7755 8044 7756 8084
rect 7796 8044 7797 8084
rect 7755 8035 7797 8044
rect 12089 8084 12131 8093
rect 12089 8044 12090 8084
rect 12130 8044 12131 8084
rect 12089 8035 12131 8044
rect 17355 8084 17397 8093
rect 17355 8044 17356 8084
rect 17396 8044 17397 8084
rect 17355 8035 17397 8044
rect 17920 8084 17962 8093
rect 17920 8044 17921 8084
rect 17961 8044 17962 8084
rect 17920 8035 17962 8044
rect 23098 8084 23156 8085
rect 23098 8044 23107 8084
rect 23147 8044 23156 8084
rect 23098 8043 23156 8044
rect 25594 8084 25652 8085
rect 25594 8044 25603 8084
rect 25643 8044 25652 8084
rect 25594 8043 25652 8044
rect 939 8000 981 8009
rect 939 7960 940 8000
rect 980 7960 981 8000
rect 939 7951 981 7960
rect 1131 8000 1173 8009
rect 1131 7960 1132 8000
rect 1172 7960 1173 8000
rect 1131 7951 1173 7960
rect 1498 8000 1556 8001
rect 1498 7960 1507 8000
rect 1547 7960 1556 8000
rect 1498 7959 1556 7960
rect 1611 8000 1653 8009
rect 1611 7960 1612 8000
rect 1652 7960 1653 8000
rect 1611 7951 1653 7960
rect 2379 8000 2421 8009
rect 2379 7960 2380 8000
rect 2420 7960 2421 8000
rect 2379 7951 2421 7960
rect 2902 8000 2944 8009
rect 2902 7960 2903 8000
rect 2943 7960 2944 8000
rect 2554 7958 2612 7959
rect 2554 7918 2563 7958
rect 2603 7918 2612 7958
rect 2902 7951 2944 7960
rect 3147 8000 3189 8009
rect 3147 7960 3148 8000
rect 3188 7960 3189 8000
rect 3147 7951 3189 7960
rect 4299 8000 4341 8009
rect 4299 7960 4300 8000
rect 4340 7960 4341 8000
rect 4299 7951 4341 7960
rect 4683 8000 4725 8009
rect 4683 7960 4684 8000
rect 4724 7960 4725 8000
rect 4683 7951 4725 7960
rect 5067 8000 5109 8009
rect 5067 7960 5068 8000
rect 5108 7960 5109 8000
rect 5067 7951 5109 7960
rect 5530 8000 5588 8001
rect 6586 8000 6644 8001
rect 5530 7960 5539 8000
rect 5579 7960 5588 8000
rect 5530 7959 5588 7960
rect 5643 7991 5685 8000
rect 5643 7951 5644 7991
rect 5684 7951 5685 7991
rect 6586 7960 6595 8000
rect 6635 7960 6644 8000
rect 6586 7959 6644 7960
rect 6699 8000 6741 8009
rect 6699 7960 6700 8000
rect 6740 7960 6741 8000
rect 6699 7951 6741 7960
rect 7126 8000 7168 8009
rect 7126 7960 7127 8000
rect 7167 7960 7168 8000
rect 7126 7951 7168 7960
rect 7371 8000 7413 8009
rect 7371 7960 7372 8000
rect 7412 7960 7413 8000
rect 7371 7951 7413 7960
rect 7659 8000 7701 8009
rect 7659 7960 7660 8000
rect 7700 7960 7701 8000
rect 7659 7951 7701 7960
rect 7851 8000 7893 8009
rect 7851 7960 7852 8000
rect 7892 7960 7893 8000
rect 7851 7951 7893 7960
rect 9579 8000 9621 8009
rect 9579 7960 9580 8000
rect 9620 7960 9621 8000
rect 9579 7951 9621 7960
rect 11770 8000 11828 8001
rect 11770 7960 11779 8000
rect 11819 7960 11828 8000
rect 11770 7959 11828 7960
rect 11883 8000 11925 8009
rect 11883 7960 11884 8000
rect 11924 7960 11925 8000
rect 11883 7951 11925 7960
rect 12444 8000 12486 8009
rect 12444 7960 12445 8000
rect 12485 7960 12486 8000
rect 12444 7951 12486 7960
rect 12555 8000 12597 8009
rect 12555 7960 12556 8000
rect 12596 7960 12597 8000
rect 12555 7951 12597 7960
rect 13035 8000 13077 8009
rect 13035 7960 13036 8000
rect 13076 7960 13077 8000
rect 14091 8000 14133 8009
rect 13035 7951 13077 7960
rect 13169 7968 13227 7969
rect 5643 7942 5685 7951
rect 13169 7928 13178 7968
rect 13218 7928 13227 7968
rect 14091 7960 14092 8000
rect 14132 7960 14133 8000
rect 14091 7951 14133 7960
rect 14667 8000 14709 8009
rect 14667 7960 14668 8000
rect 14708 7960 14709 8000
rect 14667 7951 14709 7960
rect 14859 8000 14901 8009
rect 14859 7960 14860 8000
rect 14900 7960 14901 8000
rect 14859 7951 14901 7960
rect 16491 8000 16533 8009
rect 16491 7960 16492 8000
rect 16532 7960 16533 8000
rect 16491 7951 16533 7960
rect 16666 8000 16724 8001
rect 16666 7960 16675 8000
rect 16715 7960 16724 8000
rect 16666 7959 16724 7960
rect 16875 8000 16917 8009
rect 16875 7960 16876 8000
rect 16916 7960 16917 8000
rect 16875 7951 16917 7960
rect 17067 8000 17109 8009
rect 17067 7960 17068 8000
rect 17108 7960 17109 8000
rect 17067 7951 17109 7960
rect 17259 8000 17301 8009
rect 17259 7960 17260 8000
rect 17300 7960 17301 8000
rect 17259 7951 17301 7960
rect 17451 8000 17493 8009
rect 18507 8000 18549 8009
rect 17451 7960 17452 8000
rect 17492 7960 17493 8000
rect 17451 7951 17493 7960
rect 18219 7991 18261 8000
rect 18219 7951 18220 7991
rect 18260 7951 18261 7991
rect 18507 7960 18508 8000
rect 18548 7960 18549 8000
rect 19264 8000 19306 8009
rect 20043 8000 20085 8009
rect 22330 8000 22388 8001
rect 18507 7951 18549 7960
rect 18747 7958 18789 7967
rect 18219 7942 18261 7951
rect 13169 7927 13227 7928
rect 2554 7917 2612 7918
rect 3034 7916 3092 7917
rect 3034 7876 3043 7916
rect 3083 7876 3092 7916
rect 3034 7875 3092 7876
rect 7258 7916 7316 7917
rect 7258 7876 7267 7916
rect 7307 7876 7316 7916
rect 7258 7875 7316 7876
rect 18626 7916 18668 7925
rect 18626 7876 18627 7916
rect 18667 7876 18668 7916
rect 18747 7918 18748 7958
rect 18788 7918 18789 7958
rect 19264 7960 19265 8000
rect 19305 7960 19306 8000
rect 19264 7951 19306 7960
rect 19563 7991 19605 8000
rect 19563 7951 19564 7991
rect 19604 7951 19605 7991
rect 20043 7960 20044 8000
rect 20084 7960 20085 8000
rect 20043 7951 20085 7960
rect 21675 7991 21717 8000
rect 21675 7951 21676 7991
rect 21716 7951 21717 7991
rect 19563 7942 19605 7951
rect 21675 7942 21717 7951
rect 21786 7991 21828 8000
rect 21786 7951 21787 7991
rect 21827 7951 21828 7991
rect 21786 7942 21828 7951
rect 21906 7991 21952 8000
rect 21906 7951 21907 7991
rect 21947 7951 21952 7991
rect 22330 7960 22339 8000
rect 22379 7960 22388 8000
rect 22330 7959 22388 7960
rect 22731 8000 22773 8009
rect 22731 7960 22732 8000
rect 22772 7960 22773 8000
rect 22731 7951 22773 7960
rect 23482 8000 23540 8001
rect 23482 7960 23491 8000
rect 23531 7960 23540 8000
rect 23482 7959 23540 7960
rect 25978 8000 26036 8001
rect 25978 7960 25987 8000
rect 26027 7960 26036 8000
rect 25978 7959 26036 7960
rect 28762 8000 28820 8001
rect 28762 7960 28771 8000
rect 28811 7960 28820 8000
rect 28762 7959 28820 7960
rect 28875 8000 28917 8009
rect 28875 7960 28876 8000
rect 28916 7960 28917 8000
rect 28875 7951 28917 7960
rect 29722 8000 29780 8001
rect 29722 7960 29731 8000
rect 29771 7960 29780 8000
rect 29722 7959 29780 7960
rect 29829 8000 29887 8001
rect 29829 7960 29838 8000
rect 29878 7960 29887 8000
rect 29829 7959 29887 7960
rect 30490 8000 30548 8001
rect 30490 7960 30499 8000
rect 30539 7960 30548 8000
rect 30490 7959 30548 7960
rect 30603 8000 30645 8009
rect 30603 7960 30604 8000
rect 30644 7960 30645 8000
rect 30603 7951 30645 7960
rect 21906 7942 21952 7951
rect 18747 7909 18789 7918
rect 19953 7916 19995 7925
rect 18626 7867 18668 7876
rect 19953 7876 19954 7916
rect 19994 7876 19995 7916
rect 19953 7867 19995 7876
rect 27531 7916 27573 7925
rect 27531 7876 27532 7916
rect 27572 7876 27573 7916
rect 27531 7867 27573 7876
rect 1035 7832 1077 7841
rect 1035 7792 1036 7832
rect 1076 7792 1077 7832
rect 1035 7783 1077 7792
rect 5931 7832 5973 7841
rect 5931 7792 5932 7832
rect 5972 7792 5973 7832
rect 5931 7783 5973 7792
rect 31083 7832 31125 7841
rect 31083 7792 31084 7832
rect 31124 7792 31125 7832
rect 31083 7783 31125 7792
rect 1786 7748 1844 7749
rect 1786 7708 1795 7748
rect 1835 7708 1844 7748
rect 1786 7707 1844 7708
rect 9435 7748 9477 7757
rect 9435 7708 9436 7748
rect 9476 7708 9477 7748
rect 9435 7699 9477 7708
rect 12075 7748 12117 7757
rect 12075 7708 12076 7748
rect 12116 7708 12117 7748
rect 12075 7699 12117 7708
rect 14763 7748 14805 7757
rect 14763 7708 14764 7748
rect 14804 7708 14805 7748
rect 14763 7699 14805 7708
rect 25035 7748 25077 7757
rect 25035 7708 25036 7748
rect 25076 7708 25077 7748
rect 25035 7699 25077 7708
rect 30699 7748 30741 7757
rect 30699 7708 30700 7748
rect 30740 7708 30741 7748
rect 30699 7699 30741 7708
rect 576 7580 31392 7604
rect 576 7540 3112 7580
rect 3480 7540 10886 7580
rect 11254 7540 18660 7580
rect 19028 7540 26434 7580
rect 26802 7540 31392 7580
rect 576 7516 31392 7540
rect 1498 7412 1556 7413
rect 1498 7372 1507 7412
rect 1547 7372 1556 7412
rect 1498 7371 1556 7372
rect 3147 7412 3189 7421
rect 3147 7372 3148 7412
rect 3188 7372 3189 7412
rect 3147 7363 3189 7372
rect 4971 7412 5013 7421
rect 4971 7372 4972 7412
rect 5012 7372 5013 7412
rect 4971 7363 5013 7372
rect 6874 7412 6932 7413
rect 6874 7372 6883 7412
rect 6923 7372 6932 7412
rect 6874 7371 6932 7372
rect 9963 7412 10005 7421
rect 9963 7372 9964 7412
rect 10004 7372 10005 7412
rect 9963 7363 10005 7372
rect 11979 7412 12021 7421
rect 11979 7372 11980 7412
rect 12020 7372 12021 7412
rect 11979 7363 12021 7372
rect 12730 7412 12788 7413
rect 12730 7372 12739 7412
rect 12779 7372 12788 7412
rect 12730 7371 12788 7372
rect 14746 7412 14804 7413
rect 14746 7372 14755 7412
rect 14795 7372 14804 7412
rect 14746 7371 14804 7372
rect 18219 7412 18261 7421
rect 18219 7372 18220 7412
rect 18260 7372 18261 7412
rect 18219 7363 18261 7372
rect 20410 7412 20468 7413
rect 20410 7372 20419 7412
rect 20459 7372 20468 7412
rect 20410 7371 20468 7372
rect 21291 7412 21333 7421
rect 21291 7372 21292 7412
rect 21332 7372 21333 7412
rect 21291 7363 21333 7372
rect 22059 7412 22101 7421
rect 22059 7372 22060 7412
rect 22100 7372 22101 7412
rect 22059 7363 22101 7372
rect 30507 7412 30549 7421
rect 30507 7372 30508 7412
rect 30548 7372 30549 7412
rect 30507 7363 30549 7372
rect 8122 7328 8180 7329
rect 8122 7288 8131 7328
rect 8171 7288 8180 7328
rect 8122 7287 8180 7288
rect 19450 7328 19508 7329
rect 19450 7288 19459 7328
rect 19499 7288 19508 7328
rect 19450 7287 19508 7288
rect 19611 7328 19653 7337
rect 19611 7288 19612 7328
rect 19652 7288 19653 7328
rect 19611 7279 19653 7288
rect 24651 7328 24693 7337
rect 24651 7288 24652 7328
rect 24692 7288 24693 7328
rect 24651 7279 24693 7288
rect 28875 7328 28917 7337
rect 28875 7288 28876 7328
rect 28916 7288 28917 7328
rect 28875 7279 28917 7288
rect 29643 7328 29685 7337
rect 29643 7288 29644 7328
rect 29684 7288 29685 7328
rect 29643 7279 29685 7288
rect 12490 7272 12548 7273
rect 1882 7244 1940 7245
rect 1882 7204 1891 7244
rect 1931 7204 1940 7244
rect 1882 7203 1940 7204
rect 2091 7244 2133 7253
rect 8907 7244 8949 7253
rect 2091 7204 2092 7244
rect 2132 7204 2133 7244
rect 2091 7195 2133 7204
rect 4434 7235 4480 7244
rect 4434 7195 4435 7235
rect 4475 7195 4480 7235
rect 8907 7204 8908 7244
rect 8948 7204 8949 7244
rect 8907 7195 8949 7204
rect 9483 7244 9525 7253
rect 9483 7204 9484 7244
rect 9524 7204 9525 7244
rect 12490 7232 12499 7272
rect 12539 7232 12548 7272
rect 12490 7231 12548 7232
rect 18490 7244 18548 7245
rect 9483 7195 9525 7204
rect 18490 7204 18499 7244
rect 18539 7204 18548 7244
rect 18490 7203 18548 7204
rect 18699 7244 18741 7253
rect 18699 7204 18700 7244
rect 18740 7204 18741 7244
rect 4434 7186 4480 7195
rect 4677 7193 4735 7194
rect 1210 7160 1268 7161
rect 1210 7120 1219 7160
rect 1259 7120 1268 7160
rect 1210 7119 1268 7120
rect 1323 7160 1365 7169
rect 1323 7120 1324 7160
rect 1364 7120 1365 7160
rect 1323 7111 1365 7120
rect 1750 7160 1792 7169
rect 1750 7120 1751 7160
rect 1791 7120 1792 7160
rect 1750 7111 1792 7120
rect 1995 7160 2037 7169
rect 1995 7120 1996 7160
rect 2036 7120 2037 7160
rect 1995 7111 2037 7120
rect 2283 7160 2325 7169
rect 2283 7120 2284 7160
rect 2324 7120 2325 7160
rect 2283 7111 2325 7120
rect 2475 7160 2517 7169
rect 2475 7120 2476 7160
rect 2516 7120 2517 7160
rect 2475 7111 2517 7120
rect 2842 7160 2900 7161
rect 2842 7120 2851 7160
rect 2891 7120 2900 7160
rect 2842 7119 2900 7120
rect 2955 7160 2997 7169
rect 2955 7120 2956 7160
rect 2996 7120 2997 7160
rect 2955 7111 2997 7120
rect 4299 7160 4341 7169
rect 4299 7120 4300 7160
rect 4340 7120 4341 7160
rect 4299 7111 4341 7120
rect 4533 7160 4575 7169
rect 4533 7120 4534 7160
rect 4574 7120 4575 7160
rect 4677 7153 4686 7193
rect 4726 7153 4735 7193
rect 10155 7193 10197 7202
rect 18699 7195 18741 7204
rect 27562 7244 27620 7245
rect 27562 7204 27571 7244
rect 27611 7204 27620 7244
rect 27562 7203 27620 7204
rect 29914 7244 29972 7245
rect 29914 7204 29923 7244
rect 29963 7204 29972 7244
rect 29914 7203 29972 7204
rect 30123 7244 30165 7253
rect 30123 7204 30124 7244
rect 30164 7204 30165 7244
rect 4677 7152 4735 7153
rect 4982 7160 5024 7169
rect 4533 7111 4575 7120
rect 4982 7120 4983 7160
rect 5023 7120 5024 7160
rect 4982 7111 5024 7120
rect 6699 7160 6741 7169
rect 6699 7120 6700 7160
rect 6740 7120 6741 7160
rect 6699 7111 6741 7120
rect 6874 7160 6932 7161
rect 6874 7120 6883 7160
rect 6923 7120 6932 7160
rect 6874 7119 6932 7120
rect 7834 7160 7892 7161
rect 7834 7120 7843 7160
rect 7883 7120 7892 7160
rect 7834 7119 7892 7120
rect 7947 7160 7989 7169
rect 7947 7120 7948 7160
rect 7988 7120 7989 7160
rect 7947 7111 7989 7120
rect 8374 7160 8416 7169
rect 8374 7120 8375 7160
rect 8415 7120 8416 7160
rect 8374 7111 8416 7120
rect 8506 7160 8564 7161
rect 8506 7120 8515 7160
rect 8555 7120 8564 7160
rect 8506 7119 8564 7120
rect 8619 7160 8661 7169
rect 8619 7120 8620 7160
rect 8660 7120 8661 7160
rect 8619 7111 8661 7120
rect 9082 7160 9140 7161
rect 9082 7120 9091 7160
rect 9131 7120 9140 7160
rect 9082 7119 9140 7120
rect 10044 7160 10086 7169
rect 10044 7120 10045 7160
rect 10085 7120 10086 7160
rect 10155 7153 10156 7193
rect 10196 7153 10197 7193
rect 29595 7193 29637 7202
rect 30123 7195 30165 7204
rect 30609 7244 30651 7253
rect 30609 7204 30610 7244
rect 30650 7204 30651 7244
rect 30609 7195 30651 7204
rect 10155 7144 10197 7153
rect 10966 7160 11008 7169
rect 10044 7111 10086 7120
rect 10966 7120 10967 7160
rect 11007 7120 11008 7160
rect 10966 7111 11008 7120
rect 11098 7160 11156 7161
rect 11098 7120 11107 7160
rect 11147 7120 11156 7160
rect 11098 7119 11156 7120
rect 11211 7160 11253 7169
rect 11211 7120 11212 7160
rect 11252 7120 11253 7160
rect 11211 7111 11253 7120
rect 12171 7160 12213 7169
rect 12171 7120 12172 7160
rect 12212 7120 12213 7160
rect 12171 7111 12213 7120
rect 12538 7160 12596 7161
rect 12538 7120 12547 7160
rect 12587 7120 12596 7160
rect 12538 7119 12596 7120
rect 13227 7160 13269 7169
rect 13227 7120 13228 7160
rect 13268 7120 13269 7160
rect 13227 7111 13269 7120
rect 13414 7160 13472 7161
rect 13414 7120 13423 7160
rect 13463 7120 13472 7160
rect 13414 7119 13472 7120
rect 14458 7160 14516 7161
rect 14458 7120 14467 7160
rect 14507 7120 14516 7160
rect 14458 7119 14516 7120
rect 14571 7160 14613 7169
rect 14571 7120 14572 7160
rect 14612 7120 14613 7160
rect 14571 7111 14613 7120
rect 15195 7160 15237 7169
rect 15195 7120 15196 7160
rect 15236 7120 15237 7160
rect 15195 7111 15237 7120
rect 15339 7160 15381 7169
rect 15339 7120 15340 7160
rect 15380 7120 15381 7160
rect 15339 7111 15381 7120
rect 18012 7160 18054 7169
rect 18012 7120 18013 7160
rect 18053 7120 18054 7160
rect 18012 7111 18054 7120
rect 18358 7160 18400 7169
rect 18358 7120 18359 7160
rect 18399 7120 18400 7160
rect 18358 7111 18400 7120
rect 18603 7160 18645 7169
rect 18603 7120 18604 7160
rect 18644 7120 18645 7160
rect 18603 7111 18645 7120
rect 19275 7160 19317 7169
rect 19275 7120 19276 7160
rect 19316 7120 19317 7160
rect 19275 7111 19317 7120
rect 19450 7160 19508 7161
rect 19450 7120 19459 7160
rect 19499 7120 19508 7160
rect 19450 7119 19508 7120
rect 19947 7160 19989 7169
rect 19947 7120 19948 7160
rect 19988 7120 19989 7160
rect 19947 7111 19989 7120
rect 20235 7160 20277 7169
rect 20235 7120 20236 7160
rect 20276 7120 20277 7160
rect 20235 7111 20277 7120
rect 20413 7160 20455 7169
rect 20413 7120 20414 7160
rect 20454 7120 20455 7160
rect 20413 7111 20455 7120
rect 20707 7160 20765 7161
rect 20707 7120 20716 7160
rect 20756 7120 20765 7160
rect 20707 7119 20765 7120
rect 21339 7160 21381 7169
rect 21339 7120 21340 7160
rect 21380 7120 21381 7160
rect 21339 7111 21381 7120
rect 21483 7160 21525 7169
rect 21483 7120 21484 7160
rect 21524 7120 21525 7160
rect 21483 7111 21525 7120
rect 22140 7160 22182 7169
rect 22140 7120 22141 7160
rect 22181 7120 22182 7160
rect 22140 7111 22182 7120
rect 22251 7160 22293 7169
rect 22251 7120 22252 7160
rect 22292 7120 22293 7160
rect 22251 7111 22293 7120
rect 23307 7160 23349 7169
rect 23307 7120 23308 7160
rect 23348 7120 23349 7160
rect 23307 7111 23349 7120
rect 23499 7160 23541 7169
rect 23499 7120 23500 7160
rect 23540 7120 23541 7160
rect 23499 7111 23541 7120
rect 23767 7160 23825 7161
rect 23767 7120 23776 7160
rect 23816 7120 23825 7160
rect 23767 7119 23825 7120
rect 24267 7160 24309 7169
rect 24267 7120 24268 7160
rect 24308 7120 24309 7160
rect 24267 7111 24309 7120
rect 25015 7160 25073 7161
rect 25015 7120 25024 7160
rect 25064 7120 25073 7160
rect 25015 7119 25073 7120
rect 25179 7160 25221 7169
rect 25179 7120 25180 7160
rect 25220 7120 25221 7160
rect 25179 7111 25221 7120
rect 27757 7160 27815 7161
rect 27757 7120 27766 7160
rect 27806 7120 27815 7160
rect 27757 7119 27815 7120
rect 28587 7160 28629 7169
rect 28587 7120 28588 7160
rect 28628 7120 28629 7160
rect 28587 7111 28629 7120
rect 28875 7160 28917 7169
rect 28875 7120 28876 7160
rect 28916 7120 28917 7160
rect 28875 7111 28917 7120
rect 28990 7160 29032 7169
rect 28990 7120 28991 7160
rect 29031 7120 29032 7160
rect 28990 7111 29032 7120
rect 29163 7160 29205 7169
rect 29163 7120 29164 7160
rect 29204 7120 29205 7160
rect 29163 7111 29205 7120
rect 29347 7160 29405 7161
rect 29347 7120 29356 7160
rect 29396 7120 29405 7160
rect 29347 7119 29405 7120
rect 29469 7160 29527 7161
rect 29469 7120 29478 7160
rect 29518 7120 29527 7160
rect 29595 7153 29596 7193
rect 29636 7153 29637 7193
rect 29595 7144 29637 7153
rect 29782 7160 29824 7169
rect 29469 7119 29527 7120
rect 29782 7120 29783 7160
rect 29823 7120 29824 7160
rect 29782 7111 29824 7120
rect 30027 7160 30069 7169
rect 30027 7120 30028 7160
rect 30068 7120 30069 7160
rect 30027 7111 30069 7120
rect 30699 7160 30741 7169
rect 30699 7120 30700 7160
rect 30740 7120 30741 7160
rect 30699 7111 30741 7120
rect 2379 7076 2421 7085
rect 2379 7036 2380 7076
rect 2420 7036 2421 7076
rect 2379 7027 2421 7036
rect 3158 7076 3200 7085
rect 3158 7036 3159 7076
rect 3199 7036 3200 7076
rect 3158 7027 3200 7036
rect 4203 7076 4245 7085
rect 4203 7036 4204 7076
rect 4244 7036 4245 7076
rect 4203 7027 4245 7036
rect 9387 7076 9429 7085
rect 9387 7036 9388 7076
rect 9428 7036 9429 7076
rect 9387 7027 9429 7036
rect 23194 7076 23252 7077
rect 23194 7036 23203 7076
rect 23243 7036 23252 7076
rect 23194 7035 23252 7036
rect 28186 7076 28244 7077
rect 28186 7036 28195 7076
rect 28235 7036 28244 7076
rect 28186 7035 28244 7036
rect 4762 6992 4820 6993
rect 4762 6952 4771 6992
rect 4811 6952 4820 6992
rect 4762 6951 4820 6952
rect 8698 6992 8756 6993
rect 8698 6952 8707 6992
rect 8747 6952 8756 6992
rect 8698 6951 8756 6952
rect 11290 6992 11348 6993
rect 11290 6952 11299 6992
rect 11339 6952 11348 6992
rect 11290 6951 11348 6952
rect 12250 6992 12308 6993
rect 12250 6952 12259 6992
rect 12299 6952 12308 6992
rect 12250 6951 12308 6952
rect 13402 6992 13460 6993
rect 13402 6952 13411 6992
rect 13451 6952 13460 6992
rect 13402 6951 13460 6952
rect 15034 6992 15092 6993
rect 15034 6952 15043 6992
rect 15083 6952 15092 6992
rect 15034 6951 15092 6952
rect 17914 6992 17972 6993
rect 17914 6952 17923 6992
rect 17963 6952 17972 6992
rect 17914 6951 17972 6952
rect 20619 6992 20661 7001
rect 20619 6952 20620 6992
rect 20660 6952 20661 6992
rect 20619 6943 20661 6952
rect 23499 6992 23541 7001
rect 23499 6952 23500 6992
rect 23540 6952 23541 6992
rect 23499 6943 23541 6952
rect 23931 6992 23973 7001
rect 23931 6952 23932 6992
rect 23972 6952 23973 6992
rect 23931 6943 23973 6952
rect 24363 6992 24405 7001
rect 24363 6952 24364 6992
rect 24404 6952 24405 6992
rect 24363 6943 24405 6952
rect 576 6824 31392 6848
rect 576 6784 4352 6824
rect 4720 6784 12126 6824
rect 12494 6784 19900 6824
rect 20268 6784 27674 6824
rect 28042 6784 31392 6824
rect 576 6760 31392 6784
rect 1899 6656 1941 6665
rect 1899 6616 1900 6656
rect 1940 6616 1941 6656
rect 1899 6607 1941 6616
rect 2667 6656 2709 6665
rect 2667 6616 2668 6656
rect 2708 6616 2709 6656
rect 2667 6607 2709 6616
rect 3915 6656 3957 6665
rect 3915 6616 3916 6656
rect 3956 6616 3957 6656
rect 3915 6607 3957 6616
rect 4683 6656 4725 6665
rect 4683 6616 4684 6656
rect 4724 6616 4725 6656
rect 4683 6607 4725 6616
rect 6202 6656 6260 6657
rect 6202 6616 6211 6656
rect 6251 6616 6260 6656
rect 6202 6615 6260 6616
rect 7467 6656 7509 6665
rect 7467 6616 7468 6656
rect 7508 6616 7509 6656
rect 7467 6607 7509 6616
rect 8026 6656 8084 6657
rect 8026 6616 8035 6656
rect 8075 6616 8084 6656
rect 8026 6615 8084 6616
rect 9291 6656 9333 6665
rect 9291 6616 9292 6656
rect 9332 6616 9333 6656
rect 9291 6607 9333 6616
rect 10155 6656 10197 6665
rect 10155 6616 10156 6656
rect 10196 6616 10197 6656
rect 10155 6607 10197 6616
rect 10827 6656 10869 6665
rect 10827 6616 10828 6656
rect 10868 6616 10869 6656
rect 10827 6607 10869 6616
rect 12538 6656 12596 6657
rect 12538 6616 12547 6656
rect 12587 6616 12596 6656
rect 12538 6615 12596 6616
rect 13515 6656 13557 6665
rect 13515 6616 13516 6656
rect 13556 6616 13557 6656
rect 13515 6607 13557 6616
rect 16971 6656 17013 6665
rect 16971 6616 16972 6656
rect 17012 6616 17013 6656
rect 16971 6607 17013 6616
rect 18202 6656 18260 6657
rect 18202 6616 18211 6656
rect 18251 6616 18260 6656
rect 18202 6615 18260 6616
rect 21562 6656 21620 6657
rect 21562 6616 21571 6656
rect 21611 6616 21620 6656
rect 21562 6615 21620 6616
rect 22491 6656 22533 6665
rect 22491 6616 22492 6656
rect 22532 6616 22533 6656
rect 22491 6607 22533 6616
rect 23499 6656 23541 6665
rect 23499 6616 23500 6656
rect 23540 6616 23541 6656
rect 23499 6607 23541 6616
rect 23674 6656 23732 6657
rect 23674 6616 23683 6656
rect 23723 6616 23732 6656
rect 23674 6615 23732 6616
rect 26746 6656 26804 6657
rect 26746 6616 26755 6656
rect 26795 6616 26804 6656
rect 26746 6615 26804 6616
rect 28779 6656 28821 6665
rect 28779 6616 28780 6656
rect 28820 6616 28821 6656
rect 28779 6607 28821 6616
rect 29530 6656 29588 6657
rect 29530 6616 29539 6656
rect 29579 6616 29588 6656
rect 29530 6615 29588 6616
rect 6603 6572 6645 6581
rect 6603 6532 6604 6572
rect 6644 6532 6645 6572
rect 6603 6523 6645 6532
rect 6710 6572 6752 6581
rect 6710 6532 6711 6572
rect 6751 6532 6752 6572
rect 6710 6523 6752 6532
rect 8139 6572 8181 6581
rect 8139 6532 8140 6572
rect 8180 6532 8181 6572
rect 8139 6523 8181 6532
rect 14091 6572 14133 6581
rect 14091 6532 14092 6572
rect 14132 6532 14133 6572
rect 14091 6523 14133 6532
rect 15034 6572 15092 6573
rect 15034 6532 15043 6572
rect 15083 6532 15092 6572
rect 15034 6531 15092 6532
rect 29242 6572 29300 6573
rect 29242 6532 29251 6572
rect 29291 6532 29300 6572
rect 29242 6531 29300 6532
rect 29750 6572 29792 6581
rect 29750 6532 29751 6572
rect 29791 6532 29792 6572
rect 29750 6523 29792 6532
rect 1498 6488 1556 6489
rect 1498 6448 1507 6488
rect 1547 6448 1556 6488
rect 1498 6447 1556 6448
rect 1611 6488 1653 6497
rect 1611 6448 1612 6488
rect 1652 6448 1653 6488
rect 1611 6439 1653 6448
rect 2187 6488 2229 6497
rect 2187 6448 2188 6488
rect 2228 6448 2229 6488
rect 2187 6439 2229 6448
rect 2475 6488 2517 6497
rect 2475 6448 2476 6488
rect 2516 6448 2517 6488
rect 2475 6439 2517 6448
rect 2955 6488 2997 6497
rect 2955 6448 2956 6488
rect 2996 6448 2997 6488
rect 2955 6439 2997 6448
rect 3147 6488 3189 6497
rect 3147 6448 3148 6488
rect 3188 6448 3189 6488
rect 3147 6439 3189 6448
rect 3514 6488 3572 6489
rect 3514 6448 3523 6488
rect 3563 6448 3572 6488
rect 3514 6447 3572 6448
rect 3627 6488 3669 6497
rect 3627 6448 3628 6488
rect 3668 6448 3669 6488
rect 3627 6439 3669 6448
rect 4282 6488 4340 6489
rect 4282 6448 4291 6488
rect 4331 6448 4340 6488
rect 4282 6447 4340 6448
rect 4395 6488 4437 6497
rect 4395 6448 4396 6488
rect 4436 6448 4437 6488
rect 4395 6439 4437 6448
rect 4875 6488 4917 6497
rect 4875 6448 4876 6488
rect 4916 6448 4917 6488
rect 4875 6439 4917 6448
rect 5067 6488 5109 6497
rect 5067 6448 5068 6488
rect 5108 6448 5109 6488
rect 6123 6488 6165 6497
rect 5067 6439 5109 6448
rect 5883 6446 5925 6455
rect 3051 6404 3093 6413
rect 3051 6364 3052 6404
rect 3092 6364 3093 6404
rect 5883 6406 5884 6446
rect 5924 6406 5925 6446
rect 6123 6448 6124 6488
rect 6164 6448 6165 6488
rect 6123 6439 6165 6448
rect 6394 6488 6452 6489
rect 6394 6448 6403 6488
rect 6443 6448 6452 6488
rect 6394 6447 6452 6448
rect 6507 6488 6549 6497
rect 6507 6448 6508 6488
rect 6548 6448 6549 6488
rect 6507 6439 6549 6448
rect 6987 6488 7029 6497
rect 6987 6448 6988 6488
rect 7028 6448 7029 6488
rect 6987 6439 7029 6448
rect 7275 6488 7317 6497
rect 7275 6448 7276 6488
rect 7316 6448 7317 6488
rect 7275 6439 7317 6448
rect 7933 6488 7975 6497
rect 9195 6488 9237 6497
rect 7933 6448 7934 6488
rect 7974 6448 7975 6488
rect 7933 6439 7975 6448
rect 8235 6479 8277 6488
rect 8235 6439 8236 6479
rect 8276 6439 8277 6479
rect 9195 6448 9196 6488
rect 9236 6448 9237 6488
rect 9195 6439 9237 6448
rect 9387 6488 9429 6497
rect 9387 6448 9388 6488
rect 9428 6448 9429 6488
rect 9387 6439 9429 6448
rect 9675 6488 9717 6497
rect 9675 6448 9676 6488
rect 9716 6448 9717 6488
rect 9675 6439 9717 6448
rect 9963 6488 10005 6497
rect 9963 6448 9964 6488
rect 10004 6448 10005 6488
rect 9963 6439 10005 6448
rect 10539 6488 10581 6497
rect 10539 6448 10540 6488
rect 10580 6448 10581 6488
rect 10539 6439 10581 6448
rect 10678 6488 10720 6497
rect 10678 6448 10679 6488
rect 10719 6448 10720 6488
rect 10678 6439 10720 6448
rect 11866 6488 11924 6489
rect 11866 6448 11875 6488
rect 11915 6448 11924 6488
rect 11866 6447 11924 6448
rect 11979 6488 12021 6497
rect 11979 6448 11980 6488
rect 12020 6448 12021 6488
rect 11979 6439 12021 6448
rect 12747 6488 12789 6497
rect 12747 6448 12748 6488
rect 12788 6448 12789 6488
rect 12747 6439 12789 6448
rect 13035 6488 13077 6497
rect 13035 6448 13036 6488
rect 13076 6448 13077 6488
rect 13035 6439 13077 6448
rect 13611 6488 13653 6497
rect 13611 6448 13612 6488
rect 13652 6448 13653 6488
rect 13611 6439 13653 6448
rect 13730 6488 13772 6497
rect 13730 6448 13731 6488
rect 13771 6448 13772 6488
rect 13730 6439 13772 6448
rect 13840 6488 13898 6489
rect 13840 6448 13849 6488
rect 13889 6448 13898 6488
rect 13840 6447 13898 6448
rect 13995 6488 14037 6497
rect 13995 6448 13996 6488
rect 14036 6448 14037 6488
rect 13995 6439 14037 6448
rect 14170 6488 14228 6489
rect 14170 6448 14179 6488
rect 14219 6448 14228 6488
rect 14170 6447 14228 6448
rect 14710 6488 14752 6497
rect 14710 6448 14711 6488
rect 14751 6448 14752 6488
rect 14710 6439 14752 6448
rect 14955 6488 14997 6497
rect 14955 6448 14956 6488
rect 14996 6448 14997 6488
rect 14955 6439 14997 6448
rect 15802 6488 15860 6489
rect 15802 6448 15811 6488
rect 15851 6448 15860 6488
rect 15802 6447 15860 6448
rect 15915 6488 15957 6497
rect 15915 6448 15916 6488
rect 15956 6448 15957 6488
rect 15915 6439 15957 6448
rect 16672 6488 16714 6497
rect 16672 6448 16673 6488
rect 16713 6448 16714 6488
rect 16672 6439 16714 6448
rect 16810 6488 16868 6489
rect 16810 6448 16819 6488
rect 16859 6448 16868 6488
rect 16810 6447 16868 6448
rect 17434 6488 17492 6489
rect 17434 6448 17443 6488
rect 17483 6448 17492 6488
rect 17434 6447 17492 6448
rect 17739 6488 17781 6497
rect 17739 6448 17740 6488
rect 17780 6448 17781 6488
rect 18124 6488 18166 6497
rect 17739 6439 17781 6448
rect 17883 6446 17925 6455
rect 8235 6430 8277 6439
rect 5883 6397 5925 6406
rect 17883 6406 17884 6446
rect 17924 6406 17925 6446
rect 18124 6448 18125 6488
rect 18165 6448 18166 6488
rect 18124 6439 18166 6448
rect 19083 6488 19125 6497
rect 19083 6448 19084 6488
rect 19124 6448 19125 6488
rect 19083 6439 19125 6448
rect 20314 6488 20372 6489
rect 20314 6448 20323 6488
rect 20363 6448 20372 6488
rect 20314 6447 20372 6448
rect 21771 6488 21813 6497
rect 21771 6448 21772 6488
rect 21812 6448 21813 6488
rect 21771 6439 21813 6448
rect 22059 6488 22101 6497
rect 22059 6448 22060 6488
rect 22100 6448 22101 6488
rect 22059 6439 22101 6448
rect 22347 6488 22389 6497
rect 22347 6448 22348 6488
rect 22388 6448 22389 6488
rect 22347 6439 22389 6448
rect 23098 6488 23156 6489
rect 23098 6448 23107 6488
rect 23147 6448 23156 6488
rect 23098 6447 23156 6448
rect 23211 6488 23253 6497
rect 23211 6448 23212 6488
rect 23252 6448 23253 6488
rect 23211 6439 23253 6448
rect 23979 6488 24021 6497
rect 23979 6448 23980 6488
rect 24020 6448 24021 6488
rect 23979 6439 24021 6448
rect 25210 6488 25268 6489
rect 25210 6448 25219 6488
rect 25259 6448 25268 6488
rect 25210 6447 25268 6448
rect 25947 6488 25989 6497
rect 25947 6448 25948 6488
rect 25988 6448 25989 6488
rect 25947 6439 25989 6448
rect 26091 6488 26133 6497
rect 26091 6448 26092 6488
rect 26132 6448 26133 6488
rect 26091 6439 26133 6448
rect 27051 6488 27093 6497
rect 27051 6448 27052 6488
rect 27092 6448 27093 6488
rect 27051 6439 27093 6448
rect 27819 6488 27861 6497
rect 27819 6448 27820 6488
rect 27860 6448 27861 6488
rect 27819 6439 27861 6448
rect 28059 6488 28101 6497
rect 28059 6448 28060 6488
rect 28100 6448 28101 6488
rect 28059 6439 28101 6448
rect 28299 6488 28341 6497
rect 28299 6448 28300 6488
rect 28340 6448 28341 6488
rect 28299 6439 28341 6448
rect 28443 6488 28485 6497
rect 28443 6448 28444 6488
rect 28484 6448 28485 6488
rect 28443 6439 28485 6448
rect 28587 6488 28629 6497
rect 28587 6448 28588 6488
rect 28628 6448 28629 6488
rect 28587 6439 28629 6448
rect 28918 6488 28960 6497
rect 28918 6448 28919 6488
rect 28959 6448 28960 6488
rect 28918 6439 28960 6448
rect 29163 6488 29205 6497
rect 29163 6448 29164 6488
rect 29204 6448 29205 6488
rect 29163 6439 29205 6448
rect 29434 6488 29492 6489
rect 29434 6448 29443 6488
rect 29483 6448 29492 6488
rect 29434 6447 29492 6448
rect 30603 6488 30645 6497
rect 30603 6448 30604 6488
rect 30644 6448 30645 6488
rect 30603 6439 30645 6448
rect 6010 6404 6068 6405
rect 3051 6355 3093 6364
rect 6010 6364 6019 6404
rect 6059 6364 6068 6404
rect 6010 6363 6068 6364
rect 14842 6404 14900 6405
rect 14842 6364 14851 6404
rect 14891 6364 14900 6404
rect 17883 6397 17925 6406
rect 18010 6404 18068 6405
rect 14842 6363 14900 6364
rect 18010 6364 18019 6404
rect 18059 6364 18068 6404
rect 18010 6363 18068 6364
rect 23889 6404 23931 6413
rect 23889 6364 23890 6404
rect 23930 6364 23931 6404
rect 23889 6355 23931 6364
rect 25035 6404 25077 6413
rect 25035 6364 25036 6404
rect 25076 6364 25077 6404
rect 25035 6355 25077 6364
rect 25611 6404 25653 6413
rect 25611 6364 25612 6404
rect 25652 6364 25653 6404
rect 25611 6355 25653 6364
rect 26961 6404 27003 6413
rect 26961 6364 26962 6404
rect 27002 6364 27003 6404
rect 26961 6355 27003 6364
rect 27466 6404 27524 6405
rect 27466 6364 27475 6404
rect 27515 6364 27524 6404
rect 27466 6363 27524 6364
rect 29050 6404 29108 6405
rect 29050 6364 29059 6404
rect 29099 6364 29108 6404
rect 29050 6363 29108 6364
rect 30513 6404 30555 6413
rect 30513 6364 30514 6404
rect 30554 6364 30555 6404
rect 30513 6355 30555 6364
rect 12154 6320 12212 6321
rect 12154 6280 12163 6320
rect 12203 6280 12212 6320
rect 12154 6279 12212 6280
rect 25515 6320 25557 6329
rect 25515 6280 25516 6320
rect 25556 6280 25557 6320
rect 25515 6271 25557 6280
rect 4971 6236 5013 6245
rect 4971 6196 4972 6236
rect 5012 6196 5013 6236
rect 4971 6187 5013 6196
rect 16090 6236 16148 6237
rect 16090 6196 16099 6236
rect 16139 6196 16148 6236
rect 16090 6195 16148 6196
rect 17739 6236 17781 6245
rect 17739 6196 17740 6236
rect 17780 6196 17781 6236
rect 17739 6187 17781 6196
rect 18682 6236 18740 6237
rect 18682 6196 18691 6236
rect 18731 6196 18740 6236
rect 18682 6195 18740 6196
rect 20715 6236 20757 6245
rect 20715 6196 20716 6236
rect 20756 6196 20757 6236
rect 20715 6187 20757 6196
rect 25978 6236 26036 6237
rect 25978 6196 25987 6236
rect 26027 6196 26036 6236
rect 25978 6195 26036 6196
rect 29739 6236 29781 6245
rect 29739 6196 29740 6236
rect 29780 6196 29781 6236
rect 29739 6187 29781 6196
rect 30411 6236 30453 6245
rect 30411 6196 30412 6236
rect 30452 6196 30453 6236
rect 30411 6187 30453 6196
rect 576 6068 31392 6092
rect 576 6028 3112 6068
rect 3480 6028 10886 6068
rect 11254 6028 18660 6068
rect 19028 6028 26434 6068
rect 26802 6028 31392 6068
rect 576 6004 31392 6028
rect 4347 5900 4389 5909
rect 4347 5860 4348 5900
rect 4388 5860 4389 5900
rect 4347 5851 4389 5860
rect 16474 5900 16532 5901
rect 16474 5860 16483 5900
rect 16523 5860 16532 5900
rect 16474 5859 16532 5860
rect 20907 5900 20949 5909
rect 20907 5860 20908 5900
rect 20948 5860 20949 5900
rect 20907 5851 20949 5860
rect 21466 5900 21524 5901
rect 21466 5860 21475 5900
rect 21515 5860 21524 5900
rect 21466 5859 21524 5860
rect 25402 5900 25460 5901
rect 25402 5860 25411 5900
rect 25451 5860 25460 5900
rect 25402 5859 25460 5860
rect 27898 5900 27956 5901
rect 27898 5860 27907 5900
rect 27947 5860 27956 5900
rect 27898 5859 27956 5860
rect 29259 5900 29301 5909
rect 29259 5860 29260 5900
rect 29300 5860 29301 5900
rect 29259 5851 29301 5860
rect 30586 5900 30644 5901
rect 30586 5860 30595 5900
rect 30635 5860 30644 5900
rect 30586 5859 30644 5860
rect 4683 5816 4725 5825
rect 7275 5816 7317 5825
rect 4683 5776 4684 5816
rect 4724 5776 4725 5816
rect 4683 5767 4725 5776
rect 6267 5807 6309 5816
rect 6267 5767 6268 5807
rect 6308 5767 6309 5807
rect 7275 5776 7276 5816
rect 7316 5776 7317 5816
rect 7275 5767 7317 5776
rect 9579 5816 9621 5825
rect 9579 5776 9580 5816
rect 9620 5776 9621 5816
rect 9579 5767 9621 5776
rect 22042 5816 22100 5817
rect 22042 5776 22051 5816
rect 22091 5776 22100 5816
rect 22042 5775 22100 5776
rect 6267 5758 6309 5767
rect 2458 5732 2516 5733
rect 2458 5692 2467 5732
rect 2507 5692 2516 5732
rect 2458 5691 2516 5692
rect 2667 5732 2709 5741
rect 2667 5692 2668 5732
rect 2708 5692 2709 5732
rect 2667 5683 2709 5692
rect 4587 5732 4629 5741
rect 4587 5692 4588 5732
rect 4628 5692 4629 5732
rect 4587 5683 4629 5692
rect 6778 5732 6836 5733
rect 6778 5692 6787 5732
rect 6827 5692 6836 5732
rect 6778 5691 6836 5692
rect 6987 5732 7029 5741
rect 6987 5692 6988 5732
rect 7028 5692 7029 5732
rect 9483 5732 9525 5741
rect 4762 5690 4820 5691
rect 651 5648 693 5657
rect 651 5608 652 5648
rect 692 5608 693 5648
rect 651 5599 693 5608
rect 1035 5648 1077 5657
rect 1035 5608 1036 5648
rect 1076 5608 1077 5648
rect 1035 5599 1077 5608
rect 1594 5648 1652 5649
rect 1594 5608 1603 5648
rect 1643 5608 1652 5648
rect 1594 5607 1652 5608
rect 1707 5648 1749 5657
rect 1707 5608 1708 5648
rect 1748 5608 1749 5648
rect 1707 5599 1749 5608
rect 2326 5648 2368 5657
rect 2326 5608 2327 5648
rect 2367 5608 2368 5648
rect 2326 5599 2368 5608
rect 2571 5648 2613 5657
rect 2571 5608 2572 5648
rect 2612 5608 2613 5648
rect 2571 5599 2613 5608
rect 2859 5648 2901 5657
rect 2859 5608 2860 5648
rect 2900 5608 2901 5648
rect 2859 5599 2901 5608
rect 3051 5648 3093 5657
rect 3051 5608 3052 5648
rect 3092 5608 3093 5648
rect 3051 5599 3093 5608
rect 3435 5648 3477 5657
rect 3435 5608 3436 5648
rect 3476 5608 3477 5648
rect 3435 5599 3477 5608
rect 3627 5648 3669 5657
rect 3627 5608 3628 5648
rect 3668 5608 3669 5648
rect 3627 5599 3669 5608
rect 4203 5648 4245 5657
rect 4762 5650 4771 5690
rect 4811 5650 4820 5690
rect 6987 5683 7029 5692
rect 9339 5690 9381 5699
rect 4762 5649 4820 5650
rect 4203 5608 4204 5648
rect 4244 5608 4245 5648
rect 4203 5599 4245 5608
rect 4898 5648 4940 5657
rect 4898 5608 4899 5648
rect 4939 5608 4940 5648
rect 4426 5606 4484 5607
rect 2955 5564 2997 5573
rect 4426 5566 4435 5606
rect 4475 5566 4484 5606
rect 4898 5599 4940 5608
rect 5451 5648 5493 5657
rect 5451 5608 5452 5648
rect 5492 5608 5493 5648
rect 5451 5599 5493 5608
rect 5739 5648 5781 5657
rect 5739 5608 5740 5648
rect 5780 5608 5781 5648
rect 5739 5599 5781 5608
rect 6298 5648 6356 5649
rect 6298 5608 6307 5648
rect 6347 5608 6356 5648
rect 6298 5607 6356 5608
rect 6646 5648 6688 5657
rect 6646 5608 6647 5648
rect 6687 5608 6688 5648
rect 6646 5599 6688 5608
rect 6891 5648 6933 5657
rect 6891 5608 6892 5648
rect 6932 5608 6933 5648
rect 6891 5599 6933 5608
rect 7179 5648 7221 5657
rect 7179 5608 7180 5648
rect 7220 5608 7221 5648
rect 7179 5599 7221 5608
rect 7851 5648 7893 5657
rect 7851 5608 7852 5648
rect 7892 5608 7893 5648
rect 7851 5599 7893 5608
rect 8235 5648 8277 5657
rect 8235 5608 8236 5648
rect 8276 5608 8277 5648
rect 8235 5599 8277 5608
rect 8763 5648 8805 5657
rect 8763 5608 8764 5648
rect 8804 5608 8805 5648
rect 8763 5599 8805 5608
rect 8907 5648 8949 5657
rect 8907 5608 8908 5648
rect 8948 5608 8949 5648
rect 9339 5650 9340 5690
rect 9380 5650 9381 5690
rect 9483 5692 9484 5732
rect 9524 5692 9525 5732
rect 9483 5683 9525 5692
rect 10858 5732 10916 5733
rect 10858 5692 10867 5732
rect 10907 5692 10916 5732
rect 10858 5691 10916 5692
rect 13227 5732 13269 5741
rect 13227 5692 13228 5732
rect 13268 5692 13269 5732
rect 13227 5683 13269 5692
rect 18682 5732 18740 5733
rect 18682 5692 18691 5732
rect 18731 5692 18740 5732
rect 18682 5691 18740 5692
rect 18891 5732 18933 5741
rect 18891 5692 18892 5732
rect 18932 5692 18933 5732
rect 16299 5681 16341 5690
rect 9339 5641 9381 5650
rect 9802 5648 9860 5649
rect 8907 5599 8949 5608
rect 9647 5606 9689 5615
rect 9802 5608 9811 5648
rect 9851 5608 9860 5648
rect 9802 5607 9860 5608
rect 11050 5648 11108 5649
rect 11050 5608 11059 5648
rect 11099 5608 11108 5648
rect 11050 5607 11108 5608
rect 11194 5648 11252 5649
rect 11194 5608 11203 5648
rect 11243 5608 11252 5648
rect 11194 5607 11252 5608
rect 12448 5648 12490 5657
rect 12448 5608 12449 5648
rect 12489 5608 12490 5648
rect 4426 5565 4484 5566
rect 2955 5524 2956 5564
rect 2996 5524 2997 5564
rect 2955 5515 2997 5524
rect 6507 5564 6549 5573
rect 6507 5524 6508 5564
rect 6548 5524 6549 5564
rect 9647 5566 9648 5606
rect 9688 5566 9689 5606
rect 12448 5599 12490 5608
rect 12739 5648 12797 5649
rect 12739 5608 12748 5648
rect 12788 5608 12797 5648
rect 12739 5607 12797 5608
rect 12891 5648 12933 5657
rect 12891 5608 12892 5648
rect 12932 5608 12933 5648
rect 12891 5599 12933 5608
rect 13018 5648 13076 5649
rect 13018 5608 13027 5648
rect 13067 5608 13076 5648
rect 13018 5607 13076 5608
rect 13131 5648 13173 5657
rect 13131 5608 13132 5648
rect 13172 5608 13173 5648
rect 13131 5599 13173 5608
rect 13995 5648 14037 5657
rect 13995 5608 13996 5648
rect 14036 5608 14037 5648
rect 13995 5599 14037 5608
rect 14283 5648 14325 5657
rect 14283 5608 14284 5648
rect 14324 5608 14325 5648
rect 14283 5599 14325 5608
rect 14619 5648 14661 5657
rect 14619 5608 14620 5648
rect 14660 5608 14661 5648
rect 14619 5599 14661 5608
rect 14763 5648 14805 5657
rect 14763 5608 14764 5648
rect 14804 5608 14805 5648
rect 14763 5599 14805 5608
rect 15226 5648 15284 5649
rect 15226 5608 15235 5648
rect 15275 5608 15284 5648
rect 15226 5607 15284 5608
rect 15339 5648 15381 5657
rect 15339 5608 15340 5648
rect 15380 5608 15381 5648
rect 15339 5599 15381 5608
rect 16186 5648 16244 5649
rect 16186 5608 16195 5648
rect 16235 5608 16244 5648
rect 16299 5641 16300 5681
rect 16340 5641 16341 5681
rect 17691 5681 17733 5690
rect 18891 5683 18933 5692
rect 21489 5732 21531 5741
rect 21489 5692 21490 5732
rect 21530 5692 21531 5732
rect 21489 5683 21531 5692
rect 29722 5732 29780 5733
rect 29722 5692 29731 5732
rect 29771 5692 29780 5732
rect 29722 5691 29780 5692
rect 29931 5732 29973 5741
rect 29931 5692 29932 5732
rect 29972 5692 29973 5732
rect 16299 5632 16341 5641
rect 17547 5648 17589 5657
rect 16186 5607 16244 5608
rect 17547 5608 17548 5648
rect 17588 5608 17589 5648
rect 17691 5641 17692 5681
rect 17732 5641 17733 5681
rect 22335 5681 22377 5690
rect 29931 5683 29973 5692
rect 17691 5632 17733 5641
rect 18123 5648 18165 5657
rect 17547 5599 17589 5608
rect 18123 5608 18124 5648
rect 18164 5608 18165 5648
rect 18123 5599 18165 5608
rect 18262 5648 18304 5657
rect 18262 5608 18263 5648
rect 18303 5608 18304 5648
rect 18262 5599 18304 5608
rect 18550 5648 18592 5657
rect 18550 5608 18551 5648
rect 18591 5608 18592 5648
rect 18550 5599 18592 5608
rect 18795 5648 18837 5657
rect 18795 5608 18796 5648
rect 18836 5608 18837 5648
rect 18795 5599 18837 5608
rect 20139 5648 20181 5657
rect 20139 5608 20140 5648
rect 20180 5608 20181 5648
rect 20139 5599 20181 5608
rect 20427 5648 20469 5657
rect 20427 5608 20428 5648
rect 20468 5608 20469 5648
rect 20427 5599 20469 5608
rect 20602 5648 20660 5649
rect 20602 5608 20611 5648
rect 20651 5608 20660 5648
rect 20602 5607 20660 5608
rect 20715 5648 20757 5657
rect 20715 5608 20716 5648
rect 20756 5608 20757 5648
rect 20715 5599 20757 5608
rect 21579 5648 21621 5657
rect 21579 5608 21580 5648
rect 21620 5608 21621 5648
rect 22335 5641 22336 5681
rect 22376 5641 22377 5681
rect 30262 5681 30304 5690
rect 22335 5632 22377 5641
rect 22426 5648 22484 5649
rect 21579 5599 21621 5608
rect 22426 5608 22435 5648
rect 22475 5608 22484 5648
rect 22426 5607 22484 5608
rect 24459 5648 24501 5657
rect 24459 5608 24460 5648
rect 24500 5608 24501 5648
rect 24459 5599 24501 5608
rect 24747 5648 24789 5657
rect 24747 5608 24748 5648
rect 24788 5608 24789 5648
rect 24747 5599 24789 5608
rect 25227 5648 25269 5657
rect 25227 5608 25228 5648
rect 25268 5608 25269 5648
rect 25227 5599 25269 5608
rect 25402 5648 25460 5649
rect 25402 5608 25411 5648
rect 25451 5608 25460 5648
rect 25402 5607 25460 5608
rect 25803 5648 25845 5657
rect 25803 5608 25804 5648
rect 25844 5608 25845 5648
rect 25803 5599 25845 5608
rect 25910 5648 25952 5657
rect 25910 5608 25911 5648
rect 25951 5608 25952 5648
rect 25910 5599 25952 5608
rect 27610 5648 27668 5649
rect 27610 5608 27619 5648
rect 27659 5608 27668 5648
rect 27610 5607 27668 5608
rect 27723 5648 27765 5657
rect 27723 5608 27724 5648
rect 27764 5608 27765 5648
rect 27723 5599 27765 5608
rect 28474 5648 28532 5649
rect 28474 5608 28483 5648
rect 28523 5608 28532 5648
rect 28474 5607 28532 5608
rect 28971 5648 29013 5657
rect 28971 5608 28972 5648
rect 29012 5608 29013 5648
rect 28971 5599 29013 5608
rect 29085 5648 29143 5649
rect 29085 5608 29094 5648
rect 29134 5608 29143 5648
rect 29085 5607 29143 5608
rect 29212 5648 29270 5649
rect 29212 5608 29221 5648
rect 29261 5608 29270 5648
rect 29212 5607 29270 5608
rect 29590 5648 29632 5657
rect 29590 5608 29591 5648
rect 29631 5608 29632 5648
rect 29590 5599 29632 5608
rect 29836 5648 29878 5657
rect 29836 5608 29837 5648
rect 29877 5608 29878 5648
rect 29836 5599 29878 5608
rect 30123 5648 30165 5657
rect 30123 5608 30124 5648
rect 30164 5608 30165 5648
rect 30262 5641 30263 5681
rect 30303 5641 30304 5681
rect 30262 5632 30304 5641
rect 30883 5648 30941 5649
rect 30123 5599 30165 5608
rect 30883 5608 30892 5648
rect 30932 5608 30941 5648
rect 30883 5607 30941 5608
rect 9647 5557 9689 5566
rect 11510 5564 11552 5573
rect 6507 5515 6549 5524
rect 11510 5524 11511 5564
rect 11551 5524 11552 5564
rect 11510 5515 11552 5524
rect 12538 5564 12596 5565
rect 12538 5524 12547 5564
rect 12587 5524 12596 5564
rect 12538 5523 12596 5524
rect 15435 5564 15477 5573
rect 15435 5524 15436 5564
rect 15476 5524 15477 5564
rect 15435 5515 15477 5524
rect 15542 5564 15584 5573
rect 15542 5524 15543 5564
rect 15583 5524 15584 5564
rect 15542 5515 15584 5524
rect 20918 5564 20960 5573
rect 20918 5524 20919 5564
rect 20959 5524 20960 5564
rect 20918 5515 20960 5524
rect 28793 5564 28835 5573
rect 28793 5524 28794 5564
rect 28834 5524 28835 5564
rect 28793 5515 28835 5524
rect 30589 5564 30631 5573
rect 30589 5524 30590 5564
rect 30630 5524 30631 5564
rect 30589 5515 30631 5524
rect 1131 5480 1173 5489
rect 1131 5440 1132 5480
rect 1172 5440 1173 5480
rect 1131 5431 1173 5440
rect 1995 5480 2037 5489
rect 1995 5440 1996 5480
rect 2036 5440 2037 5480
rect 1995 5431 2037 5440
rect 3610 5480 3668 5481
rect 3610 5440 3619 5480
rect 3659 5440 3668 5480
rect 3610 5439 3668 5440
rect 5931 5480 5973 5489
rect 5931 5440 5932 5480
rect 5972 5440 5973 5480
rect 5931 5431 5973 5440
rect 8331 5480 8373 5489
rect 8331 5440 8332 5480
rect 8372 5440 8373 5480
rect 8331 5431 8373 5440
rect 8602 5480 8660 5481
rect 8602 5440 8611 5480
rect 8651 5440 8660 5480
rect 8602 5439 8660 5440
rect 11290 5480 11348 5481
rect 11290 5440 11299 5480
rect 11339 5440 11348 5480
rect 11290 5439 11348 5440
rect 11403 5480 11445 5489
rect 11403 5440 11404 5480
rect 11444 5440 11445 5480
rect 11403 5431 11445 5440
rect 12651 5480 12693 5489
rect 12651 5440 12652 5480
rect 12692 5440 12693 5480
rect 12651 5431 12693 5440
rect 13786 5480 13844 5481
rect 13786 5440 13795 5480
rect 13835 5440 13844 5480
rect 13786 5439 13844 5440
rect 14458 5480 14516 5481
rect 14458 5440 14467 5480
rect 14507 5440 14516 5480
rect 14458 5439 14516 5440
rect 17835 5480 17877 5489
rect 17835 5440 17836 5480
rect 17876 5440 17877 5480
rect 17835 5431 17877 5440
rect 18411 5480 18453 5489
rect 18411 5440 18412 5480
rect 18452 5440 18453 5480
rect 18411 5431 18453 5440
rect 19930 5480 19988 5481
rect 19930 5440 19939 5480
rect 19979 5440 19988 5480
rect 19930 5439 19988 5440
rect 20698 5480 20756 5481
rect 20698 5440 20707 5480
rect 20747 5440 20756 5480
rect 20698 5439 20756 5440
rect 22546 5480 22604 5481
rect 22546 5440 22555 5480
rect 22595 5440 22604 5480
rect 22546 5439 22604 5440
rect 24939 5480 24981 5489
rect 24939 5440 24940 5480
rect 24980 5440 24981 5480
rect 24939 5431 24981 5440
rect 25594 5480 25652 5481
rect 25594 5440 25603 5480
rect 25643 5440 25652 5480
rect 25594 5439 25652 5440
rect 28570 5480 28628 5481
rect 28570 5440 28579 5480
rect 28619 5440 28628 5480
rect 28570 5439 28628 5440
rect 28683 5480 28725 5489
rect 28683 5440 28684 5480
rect 28724 5440 28725 5480
rect 28683 5431 28725 5440
rect 30411 5480 30453 5489
rect 30411 5440 30412 5480
rect 30452 5440 30453 5480
rect 30411 5431 30453 5440
rect 30795 5480 30837 5489
rect 30795 5440 30796 5480
rect 30836 5440 30837 5480
rect 30795 5431 30837 5440
rect 576 5312 31392 5336
rect 576 5272 4352 5312
rect 4720 5272 12126 5312
rect 12494 5272 19900 5312
rect 20268 5272 27674 5312
rect 28042 5272 31392 5312
rect 576 5248 31392 5272
rect 3243 5144 3285 5153
rect 3243 5104 3244 5144
rect 3284 5104 3285 5144
rect 3243 5095 3285 5104
rect 3915 5144 3957 5153
rect 3915 5104 3916 5144
rect 3956 5104 3957 5144
rect 3915 5095 3957 5104
rect 5739 5144 5781 5153
rect 5739 5104 5740 5144
rect 5780 5104 5781 5144
rect 5739 5095 5781 5104
rect 8043 5144 8085 5153
rect 8043 5104 8044 5144
rect 8084 5104 8085 5144
rect 8043 5095 8085 5104
rect 9771 5144 9813 5153
rect 9771 5104 9772 5144
rect 9812 5104 9813 5144
rect 9771 5095 9813 5104
rect 10539 5144 10581 5153
rect 10539 5104 10540 5144
rect 10580 5104 10581 5144
rect 10539 5095 10581 5104
rect 11002 5144 11060 5145
rect 11002 5104 11011 5144
rect 11051 5104 11060 5144
rect 11002 5103 11060 5104
rect 12267 5144 12309 5153
rect 12267 5104 12268 5144
rect 12308 5104 12309 5144
rect 12267 5095 12309 5104
rect 12442 5144 12500 5145
rect 12442 5104 12451 5144
rect 12491 5104 12500 5144
rect 12442 5103 12500 5104
rect 14458 5144 14516 5145
rect 14458 5104 14467 5144
rect 14507 5104 14516 5144
rect 14458 5103 14516 5104
rect 14763 5144 14805 5153
rect 14763 5104 14764 5144
rect 14804 5104 14805 5144
rect 14763 5095 14805 5104
rect 15723 5144 15765 5153
rect 15723 5104 15724 5144
rect 15764 5104 15765 5144
rect 15723 5095 15765 5104
rect 16491 5144 16533 5153
rect 16491 5104 16492 5144
rect 16532 5104 16533 5144
rect 16491 5095 16533 5104
rect 17355 5144 17397 5153
rect 17355 5104 17356 5144
rect 17396 5104 17397 5144
rect 17355 5095 17397 5104
rect 18411 5144 18453 5153
rect 18411 5104 18412 5144
rect 18452 5104 18453 5144
rect 18411 5095 18453 5104
rect 19275 5144 19317 5153
rect 19275 5104 19276 5144
rect 19316 5104 19317 5144
rect 19275 5095 19317 5104
rect 20139 5144 20181 5153
rect 20139 5104 20140 5144
rect 20180 5104 20181 5144
rect 20139 5095 20181 5104
rect 20410 5144 20468 5145
rect 20410 5104 20419 5144
rect 20459 5104 20468 5144
rect 20410 5103 20468 5104
rect 20715 5144 20757 5153
rect 20715 5104 20716 5144
rect 20756 5104 20757 5144
rect 20715 5095 20757 5104
rect 21562 5144 21620 5145
rect 21562 5104 21571 5144
rect 21611 5104 21620 5144
rect 21562 5103 21620 5104
rect 21867 5144 21909 5153
rect 21867 5104 21868 5144
rect 21908 5104 21909 5144
rect 21867 5095 21909 5104
rect 22906 5144 22964 5145
rect 22906 5104 22915 5144
rect 22955 5104 22964 5144
rect 22906 5103 22964 5104
rect 24171 5144 24213 5153
rect 24171 5104 24172 5144
rect 24212 5104 24213 5144
rect 24171 5095 24213 5104
rect 24346 5144 24404 5145
rect 24346 5104 24355 5144
rect 24395 5104 24404 5144
rect 24346 5103 24404 5104
rect 25786 5144 25844 5145
rect 25786 5104 25795 5144
rect 25835 5104 25844 5144
rect 25786 5103 25844 5104
rect 26650 5144 26708 5145
rect 26650 5104 26659 5144
rect 26699 5104 26708 5144
rect 26650 5103 26708 5104
rect 28011 5144 28053 5153
rect 28011 5104 28012 5144
rect 28052 5104 28053 5144
rect 28011 5095 28053 5104
rect 28378 5144 28436 5145
rect 28378 5104 28387 5144
rect 28427 5104 28436 5144
rect 28378 5103 28436 5104
rect 30315 5144 30357 5153
rect 30315 5104 30316 5144
rect 30356 5104 30357 5144
rect 30315 5095 30357 5104
rect 30490 5144 30548 5145
rect 30490 5104 30499 5144
rect 30539 5104 30548 5144
rect 30490 5103 30548 5104
rect 1707 5060 1749 5069
rect 1707 5020 1708 5060
rect 1748 5020 1749 5060
rect 1707 5011 1749 5020
rect 4474 5060 4532 5061
rect 4474 5020 4483 5060
rect 4523 5020 4532 5060
rect 4474 5019 4532 5020
rect 7642 5060 7700 5061
rect 7642 5020 7651 5060
rect 7691 5020 7700 5060
rect 7642 5019 7700 5020
rect 7837 5060 7879 5069
rect 7837 5020 7838 5060
rect 7878 5020 7879 5060
rect 7837 5011 7879 5020
rect 16683 5060 16725 5069
rect 16683 5020 16684 5060
rect 16724 5020 16725 5060
rect 16683 5011 16725 5020
rect 17242 5060 17300 5061
rect 17242 5020 17251 5060
rect 17291 5020 17300 5060
rect 17242 5019 17300 5020
rect 19162 5060 19220 5061
rect 19162 5020 19171 5060
rect 19211 5020 19220 5060
rect 19162 5019 19220 5020
rect 28491 5060 28533 5069
rect 28491 5020 28492 5060
rect 28532 5020 28533 5060
rect 28491 5011 28533 5020
rect 1611 4976 1653 4985
rect 1611 4936 1612 4976
rect 1652 4936 1653 4976
rect 1611 4927 1653 4936
rect 1803 4976 1845 4985
rect 1803 4936 1804 4976
rect 1844 4936 1845 4976
rect 1803 4927 1845 4936
rect 2842 4976 2900 4977
rect 2842 4936 2851 4976
rect 2891 4936 2900 4976
rect 2842 4935 2900 4936
rect 2955 4976 2997 4985
rect 2955 4936 2956 4976
rect 2996 4936 2997 4976
rect 2955 4927 2997 4936
rect 3435 4976 3477 4985
rect 3435 4936 3436 4976
rect 3476 4936 3477 4976
rect 3435 4927 3477 4936
rect 3723 4976 3765 4985
rect 3723 4936 3724 4976
rect 3764 4936 3765 4976
rect 3723 4927 3765 4936
rect 4150 4976 4192 4985
rect 4150 4936 4151 4976
rect 4191 4936 4192 4976
rect 4150 4927 4192 4936
rect 4395 4976 4437 4985
rect 4395 4936 4396 4976
rect 4436 4936 4437 4976
rect 4395 4927 4437 4936
rect 5338 4976 5396 4977
rect 5338 4936 5347 4976
rect 5387 4936 5396 4976
rect 5338 4935 5396 4936
rect 5451 4976 5493 4985
rect 5451 4936 5452 4976
rect 5492 4936 5493 4976
rect 5451 4927 5493 4936
rect 7330 4976 7388 4977
rect 7330 4936 7339 4976
rect 7379 4936 7388 4976
rect 7330 4935 7388 4936
rect 7563 4976 7605 4985
rect 8811 4976 8853 4985
rect 7563 4936 7564 4976
rect 7604 4936 7605 4976
rect 7563 4927 7605 4936
rect 8139 4967 8181 4976
rect 8139 4927 8140 4967
rect 8180 4927 8181 4967
rect 8811 4936 8812 4976
rect 8852 4936 8853 4976
rect 8811 4927 8853 4936
rect 9370 4976 9428 4977
rect 9370 4936 9379 4976
rect 9419 4936 9428 4976
rect 9370 4935 9428 4936
rect 9483 4976 9525 4985
rect 9483 4936 9484 4976
rect 9524 4936 9525 4976
rect 9483 4927 9525 4936
rect 10138 4976 10196 4977
rect 10138 4936 10147 4976
rect 10187 4936 10196 4976
rect 10138 4935 10196 4936
rect 10251 4976 10293 4985
rect 10251 4936 10252 4976
rect 10292 4936 10293 4976
rect 10251 4927 10293 4936
rect 10690 4976 10748 4977
rect 10690 4936 10699 4976
rect 10739 4936 10748 4976
rect 10690 4935 10748 4936
rect 10923 4976 10965 4985
rect 10923 4936 10924 4976
rect 10964 4936 10965 4976
rect 10923 4927 10965 4936
rect 11866 4976 11924 4977
rect 11866 4936 11875 4976
rect 11915 4936 11924 4976
rect 11866 4935 11924 4936
rect 11985 4976 12027 4985
rect 11985 4936 11986 4976
rect 12026 4936 12027 4976
rect 11985 4927 12027 4936
rect 12603 4976 12645 4985
rect 12603 4936 12604 4976
rect 12644 4936 12645 4976
rect 12603 4927 12645 4936
rect 12747 4976 12789 4985
rect 12747 4936 12748 4976
rect 12788 4936 12789 4976
rect 12747 4927 12789 4936
rect 13174 4976 13216 4985
rect 13174 4936 13175 4976
rect 13215 4936 13216 4976
rect 13174 4927 13216 4936
rect 13419 4976 13461 4985
rect 13419 4936 13420 4976
rect 13460 4936 13461 4976
rect 13419 4927 13461 4936
rect 14571 4976 14613 4985
rect 14571 4936 14572 4976
rect 14612 4936 14613 4976
rect 14571 4927 14613 4936
rect 15322 4976 15380 4977
rect 15322 4936 15331 4976
rect 15371 4936 15380 4976
rect 15322 4935 15380 4936
rect 15435 4976 15477 4985
rect 15435 4936 15436 4976
rect 15476 4936 15477 4976
rect 15435 4927 15477 4936
rect 16090 4976 16148 4977
rect 16090 4936 16099 4976
rect 16139 4936 16148 4976
rect 16090 4935 16148 4936
rect 16203 4976 16245 4985
rect 16203 4936 16204 4976
rect 16244 4936 16245 4976
rect 16203 4927 16245 4936
rect 16779 4976 16821 4985
rect 16779 4936 16780 4976
rect 16820 4936 16821 4976
rect 16779 4927 16821 4936
rect 17010 4976 17052 4985
rect 17010 4936 17011 4976
rect 17051 4936 17052 4976
rect 17010 4927 17052 4936
rect 17152 4976 17194 4985
rect 17152 4936 17153 4976
rect 17193 4936 17194 4976
rect 17152 4927 17194 4936
rect 17449 4976 17507 4977
rect 17449 4936 17458 4976
rect 17498 4936 17507 4976
rect 17449 4935 17507 4936
rect 18010 4976 18068 4977
rect 18010 4936 18019 4976
rect 18059 4936 18068 4976
rect 18010 4935 18068 4936
rect 18123 4976 18165 4985
rect 18123 4936 18124 4976
rect 18164 4936 18165 4976
rect 18123 4927 18165 4936
rect 18699 4976 18741 4985
rect 18699 4936 18700 4976
rect 18740 4936 18741 4976
rect 18699 4927 18741 4936
rect 18916 4976 18958 4985
rect 18916 4936 18917 4976
rect 18957 4936 18958 4976
rect 18916 4927 18958 4936
rect 19072 4976 19114 4985
rect 19659 4976 19701 4985
rect 19072 4936 19073 4976
rect 19113 4936 19114 4976
rect 19072 4927 19114 4936
rect 19371 4967 19413 4976
rect 19371 4927 19372 4967
rect 19412 4927 19413 4967
rect 19659 4936 19660 4976
rect 19700 4936 19701 4976
rect 19659 4927 19701 4936
rect 20043 4976 20085 4985
rect 20043 4936 20044 4976
rect 20084 4936 20085 4976
rect 20043 4927 20085 4936
rect 20523 4976 20565 4985
rect 20523 4936 20524 4976
rect 20564 4936 20565 4976
rect 20523 4927 20565 4936
rect 21675 4976 21717 4985
rect 21675 4936 21676 4976
rect 21716 4936 21717 4976
rect 21675 4927 21717 4936
rect 23115 4976 23157 4985
rect 23115 4936 23116 4976
rect 23156 4936 23157 4976
rect 23115 4927 23157 4936
rect 23434 4976 23492 4977
rect 23434 4936 23443 4976
rect 23483 4936 23492 4976
rect 23434 4935 23492 4936
rect 23770 4976 23828 4977
rect 23770 4936 23779 4976
rect 23819 4936 23828 4976
rect 23770 4935 23828 4936
rect 23883 4976 23925 4985
rect 23883 4936 23884 4976
rect 23924 4936 23925 4976
rect 23883 4927 23925 4936
rect 24540 4976 24582 4985
rect 24540 4936 24541 4976
rect 24581 4936 24582 4976
rect 24540 4927 24582 4936
rect 24651 4976 24693 4985
rect 24651 4936 24652 4976
rect 24692 4936 24693 4976
rect 24651 4927 24693 4936
rect 25980 4976 26022 4985
rect 25980 4936 25981 4976
rect 26021 4936 26022 4976
rect 25980 4927 26022 4936
rect 26091 4976 26133 4985
rect 26091 4936 26092 4976
rect 26132 4936 26133 4976
rect 26091 4927 26133 4936
rect 26859 4976 26901 4985
rect 26859 4936 26860 4976
rect 26900 4936 26901 4976
rect 26859 4927 26901 4936
rect 27147 4976 27189 4985
rect 27147 4936 27148 4976
rect 27188 4936 27189 4976
rect 27147 4927 27189 4936
rect 27802 4976 27860 4977
rect 27802 4936 27811 4976
rect 27851 4936 27860 4976
rect 27802 4935 27860 4936
rect 28107 4976 28149 4985
rect 28107 4936 28108 4976
rect 28148 4936 28149 4976
rect 28107 4927 28149 4936
rect 28288 4976 28330 4985
rect 29071 4976 29129 4977
rect 28288 4936 28289 4976
rect 28329 4936 28330 4976
rect 28288 4927 28330 4936
rect 28587 4967 28629 4976
rect 28587 4927 28588 4967
rect 28628 4927 28629 4967
rect 29071 4936 29080 4976
rect 29120 4936 29129 4976
rect 29071 4935 29129 4936
rect 29355 4976 29397 4985
rect 29355 4936 29356 4976
rect 29396 4936 29397 4976
rect 29355 4927 29397 4936
rect 29530 4976 29588 4977
rect 29530 4936 29539 4976
rect 29579 4936 29588 4976
rect 29530 4935 29588 4936
rect 29914 4976 29972 4977
rect 29914 4936 29923 4976
rect 29963 4936 29972 4976
rect 29914 4935 29972 4936
rect 30027 4976 30069 4985
rect 30027 4936 30028 4976
rect 30068 4936 30069 4976
rect 30027 4927 30069 4936
rect 30651 4976 30693 4985
rect 30651 4936 30652 4976
rect 30692 4936 30693 4976
rect 30651 4927 30693 4936
rect 30795 4976 30837 4985
rect 30795 4936 30796 4976
rect 30836 4936 30837 4976
rect 30795 4927 30837 4936
rect 8139 4918 8181 4927
rect 19371 4918 19413 4927
rect 28587 4918 28629 4927
rect 4282 4892 4340 4893
rect 4282 4852 4291 4892
rect 4331 4852 4340 4892
rect 4282 4851 4340 4852
rect 7450 4892 7508 4893
rect 7450 4852 7459 4892
rect 7499 4852 7508 4892
rect 7450 4851 7508 4852
rect 10810 4892 10868 4893
rect 10810 4852 10819 4892
rect 10859 4852 10868 4892
rect 10810 4851 10868 4852
rect 13306 4892 13364 4893
rect 13306 4852 13315 4892
rect 13355 4852 13364 4892
rect 13306 4851 13364 4852
rect 13515 4892 13557 4901
rect 18603 4892 18645 4901
rect 13515 4852 13516 4892
rect 13556 4852 13557 4892
rect 13515 4843 13557 4852
rect 16914 4883 16960 4892
rect 16914 4843 16915 4883
rect 16955 4843 16960 4883
rect 18603 4852 18604 4892
rect 18644 4852 18645 4892
rect 18603 4843 18645 4852
rect 18818 4892 18860 4901
rect 18818 4852 18819 4892
rect 18859 4852 18860 4892
rect 18818 4843 18860 4852
rect 28906 4892 28964 4893
rect 28906 4852 28915 4892
rect 28955 4852 28964 4892
rect 28906 4851 28964 4852
rect 16914 4834 16960 4843
rect 7834 4724 7892 4725
rect 7834 4684 7843 4724
rect 7883 4684 7892 4724
rect 7834 4683 7892 4684
rect 8955 4724 8997 4733
rect 8955 4684 8956 4724
rect 8996 4684 8997 4724
rect 8955 4675 8997 4684
rect 29530 4724 29588 4725
rect 29530 4684 29539 4724
rect 29579 4684 29588 4724
rect 29530 4683 29588 4684
rect 576 4556 31392 4580
rect 576 4516 3112 4556
rect 3480 4516 10886 4556
rect 11254 4516 18660 4556
rect 19028 4516 26434 4556
rect 26802 4516 31392 4556
rect 576 4492 31392 4516
rect 3435 4388 3477 4397
rect 3435 4348 3436 4388
rect 3476 4348 3477 4388
rect 3435 4339 3477 4348
rect 7371 4388 7413 4397
rect 7371 4348 7372 4388
rect 7412 4348 7413 4388
rect 7371 4339 7413 4348
rect 9099 4388 9141 4397
rect 9099 4348 9100 4388
rect 9140 4348 9141 4388
rect 9099 4339 9141 4348
rect 13131 4388 13173 4397
rect 13131 4348 13132 4388
rect 13172 4348 13173 4388
rect 13131 4339 13173 4348
rect 16299 4388 16341 4397
rect 16299 4348 16300 4388
rect 16340 4348 16341 4388
rect 16299 4339 16341 4348
rect 18411 4388 18453 4397
rect 18411 4348 18412 4388
rect 18452 4348 18453 4388
rect 18411 4339 18453 4348
rect 21675 4388 21717 4397
rect 21675 4348 21676 4388
rect 21716 4348 21717 4388
rect 21675 4339 21717 4348
rect 25882 4388 25940 4389
rect 25882 4348 25891 4388
rect 25931 4348 25940 4388
rect 25882 4347 25940 4348
rect 26650 4388 26708 4389
rect 26650 4348 26659 4388
rect 26699 4348 26708 4388
rect 26650 4347 26708 4348
rect 27322 4388 27380 4389
rect 27322 4348 27331 4388
rect 27371 4348 27380 4388
rect 27322 4347 27380 4348
rect 5067 4304 5109 4313
rect 5067 4264 5068 4304
rect 5108 4264 5109 4304
rect 5067 4255 5109 4264
rect 5338 4304 5396 4305
rect 5338 4264 5347 4304
rect 5387 4264 5396 4304
rect 5338 4263 5396 4264
rect 10635 4304 10677 4313
rect 10635 4264 10636 4304
rect 10676 4264 10677 4304
rect 10635 4255 10677 4264
rect 21274 4304 21332 4305
rect 21274 4264 21283 4304
rect 21323 4264 21332 4304
rect 21274 4263 21332 4264
rect 28203 4304 28245 4313
rect 28203 4264 28204 4304
rect 28244 4264 28245 4304
rect 28203 4255 28245 4264
rect 30219 4304 30261 4313
rect 30219 4264 30220 4304
rect 30260 4264 30261 4304
rect 30219 4255 30261 4264
rect 5242 4220 5300 4221
rect 5242 4180 5251 4220
rect 5291 4180 5300 4220
rect 5242 4179 5300 4180
rect 5499 4220 5541 4229
rect 5499 4180 5500 4220
rect 5540 4180 5541 4220
rect 5499 4171 5541 4180
rect 7834 4220 7892 4221
rect 7834 4180 7843 4220
rect 7883 4180 7892 4220
rect 7834 4179 7892 4180
rect 9201 4220 9243 4229
rect 9201 4180 9202 4220
rect 9242 4180 9243 4220
rect 9201 4171 9243 4180
rect 10906 4220 10964 4221
rect 10906 4180 10915 4220
rect 10955 4180 10964 4220
rect 10906 4179 10964 4180
rect 17626 4220 17684 4221
rect 17626 4180 17635 4220
rect 17675 4180 17684 4220
rect 17626 4179 17684 4180
rect 19665 4220 19707 4229
rect 19665 4180 19666 4220
rect 19706 4180 19707 4220
rect 19665 4171 19707 4180
rect 21777 4220 21819 4229
rect 21777 4180 21778 4220
rect 21818 4180 21819 4220
rect 29626 4220 29684 4221
rect 21777 4171 21819 4180
rect 29499 4178 29541 4187
rect 29626 4180 29635 4220
rect 29675 4180 29684 4220
rect 29626 4179 29684 4180
rect 30699 4220 30741 4229
rect 30699 4180 30700 4220
rect 30740 4180 30741 4220
rect 25874 4147 25916 4156
rect 747 4136 789 4145
rect 747 4096 748 4136
rect 788 4096 789 4136
rect 747 4087 789 4096
rect 922 4136 980 4137
rect 922 4096 931 4136
rect 971 4096 980 4136
rect 922 4095 980 4096
rect 1423 4136 1481 4137
rect 1423 4096 1432 4136
rect 1472 4096 1481 4136
rect 1423 4095 1481 4096
rect 1654 4136 1696 4145
rect 1654 4096 1655 4136
rect 1695 4096 1696 4136
rect 1654 4087 1696 4096
rect 1786 4136 1844 4137
rect 1786 4096 1795 4136
rect 1835 4096 1844 4136
rect 1786 4095 1844 4096
rect 1899 4136 1941 4145
rect 1899 4096 1900 4136
rect 1940 4096 1941 4136
rect 1899 4087 1941 4096
rect 2187 4136 2229 4145
rect 2187 4096 2188 4136
rect 2228 4096 2229 4136
rect 2187 4087 2229 4096
rect 2379 4136 2421 4145
rect 2379 4096 2380 4136
rect 2420 4096 2421 4136
rect 2379 4087 2421 4096
rect 3339 4136 3381 4145
rect 3339 4096 3340 4136
rect 3380 4096 3381 4136
rect 3339 4087 3381 4096
rect 3531 4136 3573 4145
rect 3531 4096 3532 4136
rect 3572 4096 3573 4136
rect 3531 4087 3573 4096
rect 4875 4136 4917 4145
rect 4875 4096 4876 4136
rect 4916 4096 4917 4136
rect 4875 4087 4917 4096
rect 5626 4136 5684 4137
rect 5626 4096 5635 4136
rect 5675 4096 5684 4136
rect 5626 4095 5684 4096
rect 6219 4136 6261 4145
rect 6219 4096 6220 4136
rect 6260 4096 6261 4136
rect 6219 4087 6261 4096
rect 6603 4136 6645 4145
rect 6603 4096 6604 4136
rect 6644 4096 6645 4136
rect 6603 4087 6645 4096
rect 7162 4136 7220 4137
rect 7162 4096 7171 4136
rect 7211 4096 7220 4136
rect 7162 4095 7220 4096
rect 7275 4136 7317 4145
rect 7275 4096 7276 4136
rect 7316 4096 7317 4136
rect 7275 4087 7317 4096
rect 7702 4136 7744 4145
rect 7702 4096 7703 4136
rect 7743 4096 7744 4136
rect 7702 4087 7744 4096
rect 7947 4136 7989 4145
rect 7947 4096 7948 4136
rect 7988 4096 7989 4136
rect 7947 4087 7989 4096
rect 8506 4136 8564 4137
rect 8506 4096 8515 4136
rect 8555 4096 8564 4136
rect 8506 4095 8564 4096
rect 9291 4136 9333 4145
rect 9291 4096 9292 4136
rect 9332 4096 9333 4136
rect 9291 4087 9333 4096
rect 9963 4136 10005 4145
rect 9963 4096 9964 4136
rect 10004 4096 10005 4136
rect 9963 4087 10005 4096
rect 10330 4136 10388 4137
rect 10330 4096 10339 4136
rect 10379 4096 10388 4136
rect 10330 4095 10388 4096
rect 10635 4136 10677 4145
rect 10635 4096 10636 4136
rect 10676 4096 10677 4136
rect 10635 4087 10677 4096
rect 10774 4136 10816 4145
rect 10774 4096 10775 4136
rect 10815 4096 10816 4136
rect 10774 4087 10816 4096
rect 11019 4136 11061 4145
rect 11019 4096 11020 4136
rect 11060 4096 11061 4136
rect 11019 4087 11061 4096
rect 11451 4136 11493 4145
rect 11451 4096 11452 4136
rect 11492 4096 11493 4136
rect 11451 4087 11493 4096
rect 11595 4136 11637 4145
rect 11595 4096 11596 4136
rect 11636 4096 11637 4136
rect 11595 4087 11637 4096
rect 12363 4136 12405 4145
rect 12363 4096 12364 4136
rect 12404 4096 12405 4136
rect 12363 4087 12405 4096
rect 12497 4136 12555 4137
rect 12497 4096 12506 4136
rect 12546 4096 12555 4136
rect 12497 4095 12555 4096
rect 13035 4136 13077 4145
rect 13035 4096 13036 4136
rect 13076 4096 13077 4136
rect 13035 4087 13077 4096
rect 13227 4136 13269 4145
rect 13227 4096 13228 4136
rect 13268 4096 13269 4136
rect 13227 4087 13269 4096
rect 14091 4136 14133 4145
rect 14091 4096 14092 4136
rect 14132 4096 14133 4136
rect 14091 4087 14133 4096
rect 14475 4136 14517 4145
rect 14475 4096 14476 4136
rect 14516 4096 14517 4136
rect 14475 4087 14517 4096
rect 15994 4136 16052 4137
rect 15994 4096 16003 4136
rect 16043 4096 16052 4136
rect 15994 4095 16052 4096
rect 16491 4136 16533 4145
rect 16491 4096 16492 4136
rect 16532 4096 16533 4136
rect 16491 4087 16533 4096
rect 16683 4136 16725 4145
rect 16683 4096 16684 4136
rect 16724 4096 16725 4136
rect 16683 4087 16725 4096
rect 17506 4136 17564 4137
rect 17506 4096 17515 4136
rect 17555 4096 17564 4136
rect 17506 4095 17564 4096
rect 17739 4136 17781 4145
rect 17739 4096 17740 4136
rect 17780 4096 17781 4136
rect 17739 4087 17781 4096
rect 18202 4136 18260 4137
rect 18202 4096 18211 4136
rect 18251 4096 18260 4136
rect 18202 4095 18260 4096
rect 18315 4136 18357 4145
rect 18315 4096 18316 4136
rect 18356 4096 18357 4136
rect 18315 4087 18357 4096
rect 19755 4136 19797 4145
rect 19755 4096 19756 4136
rect 19796 4096 19797 4136
rect 19755 4087 19797 4096
rect 20986 4136 21044 4137
rect 20986 4096 20995 4136
rect 21035 4096 21044 4136
rect 20986 4095 21044 4096
rect 21099 4136 21141 4145
rect 21099 4096 21100 4136
rect 21140 4096 21141 4136
rect 21099 4087 21141 4096
rect 21867 4136 21909 4145
rect 21867 4096 21868 4136
rect 21908 4096 21909 4136
rect 21867 4087 21909 4096
rect 23499 4136 23541 4145
rect 23499 4096 23500 4136
rect 23540 4096 23541 4136
rect 23499 4087 23541 4096
rect 23691 4136 23733 4145
rect 23691 4096 23692 4136
rect 23732 4096 23733 4136
rect 23691 4087 23733 4096
rect 24939 4136 24981 4145
rect 24939 4096 24940 4136
rect 24980 4096 24981 4136
rect 24939 4087 24981 4096
rect 25323 4136 25365 4145
rect 25323 4096 25324 4136
rect 25364 4096 25365 4136
rect 25874 4107 25875 4147
rect 25915 4107 25916 4147
rect 25874 4098 25916 4107
rect 26010 4136 26068 4137
rect 25323 4087 25365 4096
rect 26010 4096 26019 4136
rect 26059 4096 26068 4136
rect 26010 4095 26068 4096
rect 26306 4136 26364 4137
rect 26306 4096 26315 4136
rect 26355 4096 26364 4136
rect 26306 4095 26364 4096
rect 26443 4136 26501 4137
rect 26443 4096 26452 4136
rect 26492 4096 26501 4136
rect 26443 4095 26501 4096
rect 26947 4136 27005 4137
rect 26947 4096 26956 4136
rect 26996 4096 27005 4136
rect 26947 4095 27005 4096
rect 27159 4136 27201 4145
rect 27159 4096 27160 4136
rect 27200 4096 27201 4136
rect 26178 4085 26224 4094
rect 27159 4087 27201 4096
rect 27338 4136 27380 4145
rect 27338 4096 27339 4136
rect 27379 4096 27380 4136
rect 27338 4087 27380 4096
rect 27675 4136 27733 4137
rect 27675 4096 27684 4136
rect 27724 4096 27733 4136
rect 27675 4095 27733 4096
rect 27819 4136 27861 4145
rect 27819 4096 27820 4136
rect 27860 4096 27861 4136
rect 27819 4087 27861 4096
rect 27997 4136 28039 4145
rect 27997 4096 27998 4136
rect 28038 4096 28039 4136
rect 27997 4087 28039 4096
rect 28128 4136 28186 4137
rect 28128 4096 28137 4136
rect 28177 4096 28186 4136
rect 28128 4095 28186 4096
rect 28299 4136 28341 4145
rect 28299 4096 28300 4136
rect 28340 4096 28341 4136
rect 28299 4087 28341 4096
rect 29355 4136 29397 4145
rect 29355 4096 29356 4136
rect 29396 4096 29397 4136
rect 29499 4138 29500 4178
rect 29540 4138 29541 4178
rect 30699 4171 30741 4180
rect 29499 4129 29541 4138
rect 29739 4136 29781 4145
rect 29355 4087 29397 4096
rect 29739 4096 29740 4136
rect 29780 4096 29781 4136
rect 29739 4087 29781 4096
rect 30358 4136 30400 4145
rect 30358 4096 30359 4136
rect 30399 4096 30400 4136
rect 30358 4087 30400 4096
rect 30490 4136 30548 4137
rect 30490 4096 30499 4136
rect 30539 4096 30548 4136
rect 30490 4095 30548 4096
rect 30603 4136 30645 4145
rect 30603 4096 30604 4136
rect 30644 4096 30645 4136
rect 30603 4087 30645 4096
rect 30891 4136 30933 4145
rect 30891 4096 30892 4136
rect 30932 4096 30933 4136
rect 30891 4087 30933 4096
rect 31083 4136 31125 4145
rect 31083 4096 31084 4136
rect 31124 4096 31125 4136
rect 31083 4087 31125 4096
rect 843 4052 885 4061
rect 843 4012 844 4052
rect 884 4012 885 4052
rect 843 4003 885 4012
rect 2283 4052 2325 4061
rect 2283 4012 2284 4052
rect 2324 4012 2325 4052
rect 2283 4003 2325 4012
rect 8825 4052 8867 4061
rect 8825 4012 8826 4052
rect 8866 4012 8867 4052
rect 8825 4003 8867 4012
rect 9754 4052 9812 4053
rect 9754 4012 9763 4052
rect 9803 4012 9812 4052
rect 9754 4011 9812 4012
rect 16313 4052 16355 4061
rect 16313 4012 16314 4052
rect 16354 4012 16355 4052
rect 16313 4003 16355 4012
rect 16587 4052 16629 4061
rect 16587 4012 16588 4052
rect 16628 4012 16629 4052
rect 16587 4003 16629 4012
rect 17818 4052 17876 4053
rect 17818 4012 17827 4052
rect 17867 4012 17876 4052
rect 26178 4045 26179 4085
rect 26219 4045 26224 4085
rect 26178 4036 26224 4045
rect 26653 4052 26695 4061
rect 17818 4011 17876 4012
rect 26653 4012 26654 4052
rect 26694 4012 26695 4052
rect 26653 4003 26695 4012
rect 29818 4052 29876 4053
rect 29818 4012 29827 4052
rect 29867 4012 29876 4052
rect 29818 4011 29876 4012
rect 30987 4052 31029 4061
rect 30987 4012 30988 4052
rect 31028 4012 31029 4052
rect 30987 4003 31029 4012
rect 1258 3968 1316 3969
rect 1258 3928 1267 3968
rect 1307 3928 1316 3968
rect 1258 3927 1316 3928
rect 1978 3968 2036 3969
rect 1978 3928 1987 3968
rect 2027 3928 2036 3968
rect 1978 3927 2036 3928
rect 4762 3968 4820 3969
rect 4762 3928 4771 3968
rect 4811 3928 4820 3968
rect 4762 3927 4820 3928
rect 6699 3968 6741 3977
rect 6699 3928 6700 3968
rect 6740 3928 6741 3968
rect 6699 3919 6741 3928
rect 8026 3968 8084 3969
rect 8026 3928 8035 3968
rect 8075 3928 8084 3968
rect 8026 3927 8084 3928
rect 8602 3968 8660 3969
rect 8602 3928 8611 3968
rect 8651 3928 8660 3968
rect 8602 3927 8660 3928
rect 8715 3968 8757 3977
rect 8715 3928 8716 3968
rect 8756 3928 8757 3968
rect 8715 3919 8757 3928
rect 10042 3968 10100 3969
rect 10042 3928 10051 3968
rect 10091 3928 10100 3968
rect 10042 3927 10100 3928
rect 11098 3968 11156 3969
rect 11098 3928 11107 3968
rect 11147 3928 11156 3968
rect 11098 3927 11156 3928
rect 11290 3968 11348 3969
rect 11290 3928 11299 3968
rect 11339 3928 11348 3968
rect 11290 3927 11348 3928
rect 12651 3968 12693 3977
rect 12651 3928 12652 3968
rect 12692 3928 12693 3968
rect 12651 3919 12693 3928
rect 14571 3968 14613 3977
rect 14571 3928 14572 3968
rect 14612 3928 14613 3968
rect 14571 3919 14613 3928
rect 16090 3968 16148 3969
rect 16090 3928 16099 3968
rect 16139 3928 16148 3968
rect 16090 3927 16148 3928
rect 19450 3968 19508 3969
rect 19450 3928 19459 3968
rect 19499 3928 19508 3968
rect 19450 3927 19508 3928
rect 23595 3968 23637 3977
rect 23595 3928 23596 3968
rect 23636 3928 23637 3968
rect 23595 3919 23637 3928
rect 24826 3968 24884 3969
rect 24826 3928 24835 3968
rect 24875 3928 24884 3968
rect 24826 3927 24884 3928
rect 26859 3968 26901 3977
rect 26859 3928 26860 3968
rect 26900 3928 26901 3968
rect 26859 3919 26901 3928
rect 27514 3968 27572 3969
rect 27514 3928 27523 3968
rect 27563 3928 27572 3968
rect 27514 3927 27572 3928
rect 28683 3968 28725 3977
rect 28683 3928 28684 3968
rect 28724 3928 28725 3968
rect 28683 3919 28725 3928
rect 576 3800 31392 3824
rect 576 3760 4352 3800
rect 4720 3760 12126 3800
rect 12494 3760 19900 3800
rect 20268 3760 27674 3800
rect 28042 3760 31392 3800
rect 576 3736 31392 3760
rect 4875 3632 4917 3641
rect 4875 3592 4876 3632
rect 4916 3592 4917 3632
rect 4875 3583 4917 3592
rect 5643 3632 5685 3641
rect 5643 3592 5644 3632
rect 5684 3592 5685 3632
rect 5643 3583 5685 3592
rect 5914 3632 5972 3633
rect 5914 3592 5923 3632
rect 5963 3592 5972 3632
rect 5914 3591 5972 3592
rect 7738 3632 7796 3633
rect 7738 3592 7747 3632
rect 7787 3592 7796 3632
rect 7738 3591 7796 3592
rect 9867 3632 9909 3641
rect 9867 3592 9868 3632
rect 9908 3592 9909 3632
rect 9867 3583 9909 3592
rect 11019 3632 11061 3641
rect 11019 3592 11020 3632
rect 11060 3592 11061 3632
rect 11019 3583 11061 3592
rect 11979 3632 12021 3641
rect 11979 3592 11980 3632
rect 12020 3592 12021 3632
rect 11979 3583 12021 3592
rect 12651 3632 12693 3641
rect 12651 3592 12652 3632
rect 12692 3592 12693 3632
rect 12651 3583 12693 3592
rect 13306 3632 13364 3633
rect 13306 3592 13315 3632
rect 13355 3592 13364 3632
rect 13306 3591 13364 3592
rect 13995 3632 14037 3641
rect 13995 3592 13996 3632
rect 14036 3592 14037 3632
rect 13995 3583 14037 3592
rect 14266 3632 14324 3633
rect 14266 3592 14275 3632
rect 14315 3592 14324 3632
rect 14266 3591 14324 3592
rect 16587 3632 16629 3641
rect 16587 3592 16588 3632
rect 16628 3592 16629 3632
rect 16587 3583 16629 3592
rect 17355 3632 17397 3641
rect 17355 3592 17356 3632
rect 17396 3592 17397 3632
rect 17355 3583 17397 3592
rect 17962 3632 18020 3633
rect 17962 3592 17971 3632
rect 18011 3592 18020 3632
rect 17962 3591 18020 3592
rect 19162 3632 19220 3633
rect 19162 3592 19171 3632
rect 19211 3592 19220 3632
rect 19162 3591 19220 3592
rect 19738 3632 19796 3633
rect 19738 3592 19747 3632
rect 19787 3592 19796 3632
rect 19738 3591 19796 3592
rect 20506 3632 20564 3633
rect 20506 3592 20515 3632
rect 20555 3592 20564 3632
rect 20506 3591 20564 3592
rect 21466 3632 21524 3633
rect 21466 3592 21475 3632
rect 21515 3592 21524 3632
rect 21466 3591 21524 3592
rect 22234 3632 22292 3633
rect 22234 3592 22243 3632
rect 22283 3592 22292 3632
rect 22234 3591 22292 3592
rect 22906 3632 22964 3633
rect 22906 3592 22915 3632
rect 22955 3592 22964 3632
rect 22906 3591 22964 3592
rect 23674 3632 23732 3633
rect 23674 3592 23683 3632
rect 23723 3592 23732 3632
rect 23674 3591 23732 3592
rect 25419 3632 25461 3641
rect 25419 3592 25420 3632
rect 25460 3592 25461 3632
rect 25419 3583 25461 3592
rect 25690 3632 25748 3633
rect 25690 3592 25699 3632
rect 25739 3592 25748 3632
rect 25690 3591 25748 3592
rect 25995 3632 26037 3641
rect 25995 3592 25996 3632
rect 26036 3592 26037 3632
rect 25995 3583 26037 3592
rect 27819 3632 27861 3641
rect 27819 3592 27820 3632
rect 27860 3592 27861 3632
rect 27819 3583 27861 3592
rect 28971 3632 29013 3641
rect 28971 3592 28972 3632
rect 29012 3592 29013 3632
rect 28971 3583 29013 3592
rect 31258 3548 31316 3549
rect 15311 3506 15353 3515
rect 31258 3508 31267 3548
rect 31307 3508 31316 3548
rect 31258 3507 31316 3508
rect 1131 3464 1173 3473
rect 1131 3424 1132 3464
rect 1172 3424 1173 3464
rect 1131 3415 1173 3424
rect 1786 3464 1844 3465
rect 1786 3424 1795 3464
rect 1835 3424 1844 3464
rect 1786 3423 1844 3424
rect 4395 3464 4437 3473
rect 4395 3424 4396 3464
rect 4436 3424 4437 3464
rect 4395 3415 4437 3424
rect 4683 3464 4725 3473
rect 4683 3424 4684 3464
rect 4724 3424 4725 3464
rect 4683 3415 4725 3424
rect 5163 3464 5205 3473
rect 5163 3424 5164 3464
rect 5204 3424 5205 3464
rect 5163 3415 5205 3424
rect 5547 3464 5589 3473
rect 5547 3424 5548 3464
rect 5588 3424 5589 3464
rect 5547 3415 5589 3424
rect 6027 3464 6069 3473
rect 6027 3424 6028 3464
rect 6068 3424 6069 3464
rect 6027 3415 6069 3424
rect 7546 3464 7604 3465
rect 7546 3424 7555 3464
rect 7595 3424 7604 3464
rect 7546 3423 7604 3424
rect 9466 3464 9524 3465
rect 9466 3424 9475 3464
rect 9515 3424 9524 3464
rect 9466 3423 9524 3424
rect 9579 3464 9621 3473
rect 9579 3424 9580 3464
rect 9620 3424 9621 3464
rect 9579 3415 9621 3424
rect 10618 3464 10676 3465
rect 10618 3424 10627 3464
rect 10667 3424 10676 3464
rect 10618 3423 10676 3424
rect 10731 3464 10773 3473
rect 10731 3424 10732 3464
rect 10772 3424 10773 3464
rect 10731 3415 10773 3424
rect 11578 3464 11636 3465
rect 11578 3424 11587 3464
rect 11627 3424 11636 3464
rect 11578 3423 11636 3424
rect 11691 3464 11733 3473
rect 11691 3424 11692 3464
rect 11732 3424 11733 3464
rect 11691 3415 11733 3424
rect 12171 3464 12213 3473
rect 12171 3424 12172 3464
rect 12212 3424 12213 3464
rect 12171 3415 12213 3424
rect 12459 3464 12501 3473
rect 12459 3424 12460 3464
rect 12500 3424 12501 3464
rect 12459 3415 12501 3424
rect 12994 3464 13052 3465
rect 12994 3424 13003 3464
rect 13043 3424 13052 3464
rect 12994 3423 13052 3424
rect 13227 3464 13269 3473
rect 13227 3424 13228 3464
rect 13268 3424 13269 3464
rect 13227 3415 13269 3424
rect 13792 3464 13834 3473
rect 14460 3464 14502 3473
rect 13792 3424 13793 3464
rect 13833 3424 13834 3464
rect 13792 3415 13834 3424
rect 14091 3455 14133 3464
rect 14091 3415 14092 3455
rect 14132 3415 14133 3455
rect 14460 3424 14461 3464
rect 14501 3424 14502 3464
rect 14460 3415 14502 3424
rect 14571 3464 14613 3473
rect 15311 3466 15312 3506
rect 15352 3466 15353 3506
rect 14571 3424 14572 3464
rect 14612 3424 14613 3464
rect 14571 3415 14613 3424
rect 15010 3464 15068 3465
rect 15010 3424 15019 3464
rect 15059 3424 15068 3464
rect 15311 3457 15353 3466
rect 15466 3464 15524 3465
rect 15010 3423 15068 3424
rect 15466 3424 15475 3464
rect 15515 3424 15524 3464
rect 15466 3423 15524 3424
rect 16107 3464 16149 3473
rect 16107 3424 16108 3464
rect 16148 3424 16149 3464
rect 16107 3415 16149 3424
rect 16491 3464 16533 3473
rect 16491 3424 16492 3464
rect 16532 3424 16533 3464
rect 16491 3415 16533 3424
rect 16875 3464 16917 3473
rect 16875 3424 16876 3464
rect 16916 3424 16917 3464
rect 16875 3415 16917 3424
rect 17163 3464 17205 3473
rect 17163 3424 17164 3464
rect 17204 3424 17205 3464
rect 17163 3415 17205 3424
rect 18127 3464 18185 3465
rect 18127 3424 18136 3464
rect 18176 3424 18185 3464
rect 18127 3423 18185 3424
rect 18298 3464 18356 3465
rect 18298 3424 18307 3464
rect 18347 3424 18356 3464
rect 18298 3423 18356 3424
rect 18603 3464 18645 3473
rect 18603 3424 18604 3464
rect 18644 3424 18645 3464
rect 18603 3415 18645 3424
rect 19275 3464 19317 3473
rect 19275 3424 19276 3464
rect 19316 3424 19317 3464
rect 19275 3415 19317 3424
rect 19851 3464 19893 3473
rect 19851 3424 19852 3464
rect 19892 3424 19893 3464
rect 19851 3415 19893 3424
rect 20235 3464 20277 3473
rect 20235 3424 20236 3464
rect 20276 3424 20277 3464
rect 20235 3415 20277 3424
rect 20619 3464 20661 3473
rect 20619 3424 20620 3464
rect 20660 3424 20661 3464
rect 20619 3415 20661 3424
rect 21003 3464 21045 3473
rect 21003 3424 21004 3464
rect 21044 3424 21045 3464
rect 21003 3415 21045 3424
rect 21675 3464 21717 3473
rect 21675 3424 21676 3464
rect 21716 3424 21717 3464
rect 21675 3415 21717 3424
rect 21963 3464 22005 3473
rect 21963 3424 21964 3464
rect 22004 3424 22005 3464
rect 21963 3415 22005 3424
rect 22347 3464 22389 3473
rect 22347 3424 22348 3464
rect 22388 3424 22389 3464
rect 22347 3415 22389 3424
rect 22731 3464 22773 3473
rect 22731 3424 22732 3464
rect 22772 3424 22773 3464
rect 22731 3415 22773 3424
rect 23211 3464 23253 3473
rect 23211 3424 23212 3464
rect 23252 3424 23253 3464
rect 23211 3415 23253 3424
rect 23979 3464 24021 3473
rect 23979 3424 23980 3464
rect 24020 3424 24021 3464
rect 23979 3415 24021 3424
rect 24459 3464 24501 3473
rect 24459 3424 24460 3464
rect 24500 3424 24501 3464
rect 24459 3415 24501 3424
rect 24651 3464 24693 3473
rect 24651 3424 24652 3464
rect 24692 3424 24693 3464
rect 24651 3415 24693 3424
rect 24939 3464 24981 3473
rect 24939 3424 24940 3464
rect 24980 3424 24981 3464
rect 24939 3415 24981 3424
rect 25323 3464 25365 3473
rect 25323 3424 25324 3464
rect 25364 3424 25365 3464
rect 25323 3415 25365 3424
rect 25803 3464 25845 3473
rect 25803 3424 25804 3464
rect 25844 3424 25845 3464
rect 25803 3415 25845 3424
rect 27418 3464 27476 3465
rect 27418 3424 27427 3464
rect 27467 3424 27476 3464
rect 27418 3423 27476 3424
rect 27531 3464 27573 3473
rect 27531 3424 27532 3464
rect 27572 3424 27573 3464
rect 27531 3415 27573 3424
rect 28395 3464 28437 3473
rect 28395 3424 28396 3464
rect 28436 3424 28437 3464
rect 28395 3415 28437 3424
rect 28779 3464 28821 3473
rect 28779 3424 28780 3464
rect 28820 3424 28821 3464
rect 28779 3415 28821 3424
rect 30874 3464 30932 3465
rect 30874 3424 30883 3464
rect 30923 3424 30932 3464
rect 30874 3423 30932 3424
rect 14091 3406 14133 3415
rect 1275 3380 1317 3389
rect 1275 3340 1276 3380
rect 1316 3340 1317 3380
rect 1275 3331 1317 3340
rect 1419 3380 1461 3389
rect 1419 3340 1420 3380
rect 1460 3340 1461 3380
rect 1419 3331 1461 3340
rect 13114 3380 13172 3381
rect 13114 3340 13123 3380
rect 13163 3340 13172 3380
rect 13114 3339 13172 3340
rect 15147 3380 15189 3389
rect 15147 3340 15148 3380
rect 15188 3340 15189 3380
rect 15147 3331 15189 3340
rect 23121 3380 23163 3389
rect 23121 3340 23122 3380
rect 23162 3340 23163 3380
rect 23121 3331 23163 3340
rect 23889 3380 23931 3389
rect 23889 3340 23890 3380
rect 23930 3340 23931 3380
rect 23889 3331 23931 3340
rect 7526 3296 7568 3305
rect 7526 3256 7527 3296
rect 7567 3256 7568 3296
rect 7526 3247 7568 3256
rect 15243 3296 15285 3305
rect 15243 3256 15244 3296
rect 15284 3256 15285 3296
rect 15243 3247 15285 3256
rect 3339 3212 3381 3221
rect 3339 3172 3340 3212
rect 3380 3172 3381 3212
rect 3339 3163 3381 3172
rect 3723 3212 3765 3221
rect 3723 3172 3724 3212
rect 3764 3172 3765 3212
rect 3723 3163 3765 3172
rect 6219 3212 6261 3221
rect 6219 3172 6220 3212
rect 6260 3172 6261 3212
rect 6219 3163 6261 3172
rect 13786 3212 13844 3213
rect 13786 3172 13795 3212
rect 13835 3172 13844 3212
rect 13786 3171 13844 3172
rect 14458 3212 14516 3213
rect 14458 3172 14467 3212
rect 14507 3172 14516 3212
rect 14458 3171 14516 3172
rect 18603 3212 18645 3221
rect 18603 3172 18604 3212
rect 18644 3172 18645 3212
rect 18603 3163 18645 3172
rect 19467 3212 19509 3221
rect 19467 3172 19468 3212
rect 19508 3172 19509 3212
rect 19467 3163 19509 3172
rect 24555 3212 24597 3221
rect 24555 3172 24556 3212
rect 24596 3172 24597 3212
rect 24555 3163 24597 3172
rect 28155 3212 28197 3221
rect 28155 3172 28156 3212
rect 28196 3172 28197 3212
rect 28155 3163 28197 3172
rect 29355 3212 29397 3221
rect 29355 3172 29356 3212
rect 29396 3172 29397 3212
rect 29355 3163 29397 3172
rect 576 3044 31392 3068
rect 576 3004 3112 3044
rect 3480 3004 10886 3044
rect 11254 3004 18660 3044
rect 19028 3004 26434 3044
rect 26802 3004 31392 3044
rect 576 2980 31392 3004
rect 1899 2876 1941 2885
rect 1899 2836 1900 2876
rect 1940 2836 1941 2876
rect 1899 2827 1941 2836
rect 3915 2876 3957 2885
rect 3915 2836 3916 2876
rect 3956 2836 3957 2876
rect 3915 2827 3957 2836
rect 7354 2876 7412 2877
rect 7354 2836 7363 2876
rect 7403 2836 7412 2876
rect 7354 2835 7412 2836
rect 9466 2876 9524 2877
rect 9466 2836 9475 2876
rect 9515 2836 9524 2876
rect 9466 2835 9524 2836
rect 13419 2876 13461 2885
rect 13419 2836 13420 2876
rect 13460 2836 13461 2876
rect 13419 2827 13461 2836
rect 18507 2876 18549 2885
rect 18507 2836 18508 2876
rect 18548 2836 18549 2876
rect 18507 2827 18549 2836
rect 20235 2876 20277 2885
rect 20235 2836 20236 2876
rect 20276 2836 20277 2876
rect 20235 2827 20277 2836
rect 21178 2876 21236 2877
rect 21178 2836 21187 2876
rect 21227 2836 21236 2876
rect 21178 2835 21236 2836
rect 23163 2876 23205 2885
rect 23163 2836 23164 2876
rect 23204 2836 23205 2876
rect 23163 2827 23205 2836
rect 24843 2876 24885 2885
rect 24843 2836 24844 2876
rect 24884 2836 24885 2876
rect 24843 2827 24885 2836
rect 28762 2876 28820 2877
rect 28762 2836 28771 2876
rect 28811 2836 28820 2876
rect 28762 2835 28820 2836
rect 2475 2792 2517 2801
rect 2475 2752 2476 2792
rect 2516 2752 2517 2792
rect 2475 2743 2517 2752
rect 6699 2792 6741 2801
rect 6699 2752 6700 2792
rect 6740 2752 6741 2792
rect 6699 2743 6741 2752
rect 22827 2792 22869 2801
rect 22827 2752 22828 2792
rect 22868 2752 22869 2792
rect 22827 2743 22869 2752
rect 25563 2792 25605 2801
rect 25563 2752 25564 2792
rect 25604 2752 25605 2792
rect 25563 2743 25605 2752
rect 26859 2792 26901 2801
rect 26859 2752 26860 2792
rect 26900 2752 26901 2792
rect 26859 2743 26901 2752
rect 30315 2792 30357 2801
rect 30315 2752 30316 2792
rect 30356 2752 30357 2792
rect 30315 2743 30357 2752
rect 1131 2708 1173 2717
rect 1131 2668 1132 2708
rect 1172 2668 1173 2708
rect 1131 2659 1173 2668
rect 1346 2708 1388 2717
rect 1346 2668 1347 2708
rect 1387 2668 1388 2708
rect 1346 2659 1388 2668
rect 9850 2708 9908 2709
rect 9850 2668 9859 2708
rect 9899 2668 9908 2708
rect 9850 2667 9908 2668
rect 12442 2708 12500 2709
rect 12442 2668 12451 2708
rect 12491 2668 12500 2708
rect 12442 2667 12500 2668
rect 12651 2708 12693 2717
rect 12651 2668 12652 2708
rect 12692 2668 12693 2708
rect 6423 2657 6465 2666
rect 1227 2624 1269 2633
rect 1227 2584 1228 2624
rect 1268 2584 1269 2624
rect 1227 2575 1269 2584
rect 1456 2624 1514 2625
rect 1456 2584 1465 2624
rect 1505 2584 1514 2624
rect 1456 2583 1514 2584
rect 1594 2624 1652 2625
rect 1594 2584 1603 2624
rect 1643 2584 1652 2624
rect 1594 2583 1652 2584
rect 1707 2624 1749 2633
rect 1707 2584 1708 2624
rect 1748 2584 1749 2624
rect 1707 2575 1749 2584
rect 3051 2624 3093 2633
rect 3051 2584 3052 2624
rect 3092 2584 3093 2624
rect 3051 2575 3093 2584
rect 3243 2624 3285 2633
rect 3243 2584 3244 2624
rect 3284 2584 3285 2624
rect 3243 2575 3285 2584
rect 3514 2624 3572 2625
rect 3514 2584 3523 2624
rect 3563 2584 3572 2624
rect 3514 2583 3572 2584
rect 4587 2624 4629 2633
rect 4587 2584 4588 2624
rect 4628 2584 4629 2624
rect 4587 2575 4629 2584
rect 4893 2624 4935 2633
rect 4893 2584 4894 2624
rect 4934 2584 4935 2624
rect 4893 2575 4935 2584
rect 6027 2624 6069 2633
rect 6027 2584 6028 2624
rect 6068 2584 6069 2624
rect 6027 2575 6069 2584
rect 6298 2624 6356 2625
rect 6298 2584 6307 2624
rect 6347 2584 6356 2624
rect 6423 2617 6424 2657
rect 6464 2617 6465 2657
rect 7798 2657 7840 2666
rect 12651 2659 12693 2668
rect 14955 2708 14997 2717
rect 14955 2668 14956 2708
rect 14996 2668 14997 2708
rect 14955 2659 14997 2668
rect 15915 2708 15957 2717
rect 15915 2668 15916 2708
rect 15956 2668 15957 2708
rect 17745 2708 17787 2717
rect 15915 2659 15957 2668
rect 16251 2666 16293 2675
rect 6423 2608 6465 2617
rect 7066 2624 7124 2625
rect 6298 2583 6356 2584
rect 7066 2584 7075 2624
rect 7115 2584 7124 2624
rect 7066 2583 7124 2584
rect 7179 2624 7221 2633
rect 7179 2584 7180 2624
rect 7220 2584 7221 2624
rect 7179 2575 7221 2584
rect 7659 2624 7701 2633
rect 7659 2584 7660 2624
rect 7700 2584 7701 2624
rect 7798 2617 7799 2657
rect 7839 2617 7840 2657
rect 7798 2608 7840 2617
rect 8410 2624 8468 2625
rect 7659 2575 7701 2584
rect 8410 2584 8419 2624
rect 8459 2584 8468 2624
rect 8410 2583 8468 2584
rect 8523 2624 8565 2633
rect 8523 2584 8524 2624
rect 8564 2584 8565 2624
rect 8523 2575 8565 2584
rect 9178 2624 9236 2625
rect 9178 2584 9187 2624
rect 9227 2584 9236 2624
rect 9178 2583 9236 2584
rect 9291 2624 9333 2633
rect 9291 2584 9292 2624
rect 9332 2584 9333 2624
rect 9291 2575 9333 2584
rect 9718 2624 9760 2633
rect 9718 2584 9719 2624
rect 9759 2584 9760 2624
rect 9718 2575 9760 2584
rect 9963 2624 10005 2633
rect 9963 2584 9964 2624
rect 10004 2584 10005 2624
rect 9963 2575 10005 2584
rect 10731 2624 10773 2633
rect 10731 2584 10732 2624
rect 10772 2584 10773 2624
rect 10731 2575 10773 2584
rect 12310 2624 12352 2633
rect 12310 2584 12311 2624
rect 12351 2584 12352 2624
rect 12310 2575 12352 2584
rect 12555 2624 12597 2633
rect 12555 2584 12556 2624
rect 12596 2584 12597 2624
rect 12555 2575 12597 2584
rect 13114 2624 13172 2625
rect 13114 2584 13123 2624
rect 13163 2584 13172 2624
rect 13114 2583 13172 2584
rect 13433 2624 13475 2633
rect 13433 2584 13434 2624
rect 13474 2584 13475 2624
rect 13433 2575 13475 2584
rect 14614 2624 14656 2633
rect 14614 2584 14615 2624
rect 14655 2584 14656 2624
rect 14614 2575 14656 2584
rect 14746 2624 14804 2625
rect 14746 2584 14755 2624
rect 14795 2584 14804 2624
rect 14746 2583 14804 2584
rect 14859 2624 14901 2633
rect 14859 2584 14860 2624
rect 14900 2584 14901 2624
rect 14859 2575 14901 2584
rect 16011 2624 16053 2633
rect 16011 2584 16012 2624
rect 16052 2584 16053 2624
rect 16011 2575 16053 2584
rect 16130 2624 16172 2633
rect 16130 2584 16131 2624
rect 16171 2584 16172 2624
rect 16251 2626 16252 2666
rect 16292 2626 16293 2666
rect 17745 2668 17746 2708
rect 17786 2668 17787 2708
rect 17745 2659 17787 2668
rect 18609 2708 18651 2717
rect 18609 2668 18610 2708
rect 18650 2668 18651 2708
rect 18609 2659 18651 2668
rect 23578 2708 23636 2709
rect 23578 2668 23587 2708
rect 23627 2668 23636 2708
rect 23578 2667 23636 2668
rect 23787 2708 23829 2717
rect 23787 2668 23788 2708
rect 23828 2668 23829 2708
rect 23787 2659 23829 2668
rect 16251 2617 16293 2626
rect 16426 2624 16484 2625
rect 16130 2575 16172 2584
rect 16426 2584 16435 2624
rect 16475 2584 16484 2624
rect 16426 2583 16484 2584
rect 16529 2624 16587 2625
rect 16529 2584 16538 2624
rect 16578 2584 16587 2624
rect 16529 2583 16587 2584
rect 17155 2624 17213 2625
rect 17155 2584 17164 2624
rect 17204 2584 17213 2624
rect 17155 2583 17213 2584
rect 17835 2624 17877 2633
rect 17835 2584 17836 2624
rect 17876 2584 17877 2624
rect 17835 2575 17877 2584
rect 18699 2624 18741 2633
rect 18699 2584 18700 2624
rect 18740 2584 18741 2624
rect 18699 2575 18741 2584
rect 19930 2624 19988 2625
rect 19930 2584 19939 2624
rect 19979 2584 19988 2624
rect 19930 2583 19988 2584
rect 20246 2624 20288 2633
rect 20246 2584 20247 2624
rect 20287 2584 20288 2624
rect 20246 2575 20288 2584
rect 21475 2624 21533 2625
rect 21475 2584 21484 2624
rect 21524 2584 21533 2624
rect 21475 2583 21533 2584
rect 21675 2624 21717 2633
rect 21675 2584 21676 2624
rect 21716 2584 21717 2624
rect 21675 2575 21717 2584
rect 22539 2624 22581 2633
rect 22539 2584 22540 2624
rect 22580 2584 22581 2624
rect 22539 2575 22581 2584
rect 22653 2624 22711 2625
rect 22653 2584 22662 2624
rect 22702 2584 22711 2624
rect 22653 2583 22711 2584
rect 22780 2624 22838 2625
rect 22780 2584 22789 2624
rect 22829 2584 22838 2624
rect 22780 2583 22838 2584
rect 23307 2624 23349 2633
rect 23307 2584 23308 2624
rect 23348 2584 23349 2624
rect 23307 2575 23349 2584
rect 23458 2624 23516 2625
rect 23458 2584 23467 2624
rect 23507 2584 23516 2624
rect 23458 2583 23516 2584
rect 23691 2624 23733 2633
rect 23691 2584 23692 2624
rect 23732 2584 23733 2624
rect 23691 2575 23733 2584
rect 23979 2624 24021 2633
rect 23979 2584 23980 2624
rect 24020 2584 24021 2624
rect 23979 2575 24021 2584
rect 24154 2624 24212 2625
rect 24154 2584 24163 2624
rect 24203 2584 24212 2624
rect 24154 2583 24212 2584
rect 24363 2624 24405 2633
rect 24363 2584 24364 2624
rect 24404 2584 24405 2624
rect 24363 2575 24405 2584
rect 24507 2624 24549 2633
rect 24507 2584 24508 2624
rect 24548 2584 24549 2624
rect 24507 2575 24549 2584
rect 24651 2624 24693 2633
rect 24651 2584 24652 2624
rect 24692 2584 24693 2624
rect 24651 2575 24693 2584
rect 25323 2624 25365 2633
rect 25323 2584 25324 2624
rect 25364 2584 25365 2624
rect 25323 2575 25365 2584
rect 25411 2624 25469 2625
rect 25411 2584 25420 2624
rect 25460 2584 25469 2624
rect 25411 2583 25469 2584
rect 25755 2624 25797 2633
rect 25755 2584 25756 2624
rect 25796 2584 25797 2624
rect 25755 2575 25797 2584
rect 28203 2624 28245 2633
rect 28203 2584 28204 2624
rect 28244 2584 28245 2624
rect 28203 2575 28245 2584
rect 28395 2624 28437 2633
rect 28395 2584 28396 2624
rect 28436 2584 28437 2624
rect 28395 2575 28437 2584
rect 28587 2624 28629 2633
rect 28587 2584 28588 2624
rect 28628 2584 28629 2624
rect 28587 2575 28629 2584
rect 28762 2624 28820 2625
rect 28762 2584 28771 2624
rect 28811 2584 28820 2624
rect 28762 2583 28820 2584
rect 28954 2624 29012 2625
rect 28954 2584 28963 2624
rect 29003 2584 29012 2624
rect 28954 2583 29012 2584
rect 29259 2624 29301 2633
rect 29259 2584 29260 2624
rect 29300 2584 29301 2624
rect 29259 2575 29301 2584
rect 29434 2624 29492 2625
rect 29434 2584 29443 2624
rect 29483 2584 29492 2624
rect 29434 2583 29492 2584
rect 30123 2624 30165 2633
rect 30123 2584 30124 2624
rect 30164 2584 30165 2624
rect 30123 2575 30165 2584
rect 1913 2540 1955 2549
rect 1913 2500 1914 2540
rect 1954 2500 1955 2540
rect 1913 2491 1955 2500
rect 4683 2540 4725 2549
rect 4683 2500 4684 2540
rect 4724 2500 4725 2540
rect 4683 2491 4725 2500
rect 13227 2540 13269 2549
rect 13227 2500 13228 2540
rect 13268 2500 13269 2540
rect 13227 2491 13269 2500
rect 16864 2540 16906 2549
rect 16864 2500 16865 2540
rect 16905 2500 16906 2540
rect 16864 2491 16906 2500
rect 20043 2540 20085 2549
rect 20043 2500 20044 2540
rect 20084 2500 20085 2540
rect 20043 2491 20085 2500
rect 21181 2540 21223 2549
rect 21181 2500 21182 2540
rect 21222 2500 21223 2540
rect 21181 2491 21223 2500
rect 24075 2540 24117 2549
rect 24075 2500 24076 2540
rect 24116 2500 24117 2540
rect 24075 2491 24117 2500
rect 25120 2540 25162 2549
rect 25120 2500 25121 2540
rect 25161 2500 25162 2540
rect 25120 2491 25162 2500
rect 3226 2456 3284 2457
rect 3226 2416 3235 2456
rect 3275 2416 3284 2456
rect 3226 2415 3284 2416
rect 4779 2456 4821 2465
rect 4779 2416 4780 2456
rect 4820 2416 4821 2456
rect 4779 2407 4821 2416
rect 5067 2456 5109 2465
rect 5067 2416 5068 2456
rect 5108 2416 5109 2456
rect 5067 2407 5109 2416
rect 5355 2456 5397 2465
rect 7947 2456 7989 2465
rect 5355 2416 5356 2456
rect 5396 2416 5397 2456
rect 5355 2407 5397 2416
rect 6210 2447 6256 2456
rect 6210 2407 6211 2447
rect 6251 2407 6256 2447
rect 7947 2416 7948 2456
rect 7988 2416 7989 2456
rect 7947 2407 7989 2416
rect 8811 2456 8853 2465
rect 8811 2416 8812 2456
rect 8852 2416 8853 2456
rect 8811 2407 8853 2416
rect 10042 2456 10100 2457
rect 10042 2416 10051 2456
rect 10091 2416 10100 2456
rect 10042 2415 10100 2416
rect 10618 2456 10676 2457
rect 10618 2416 10627 2456
rect 10667 2416 10676 2456
rect 10618 2415 10676 2416
rect 10923 2456 10965 2465
rect 10923 2416 10924 2456
rect 10964 2416 10965 2456
rect 10923 2407 10965 2416
rect 16683 2456 16725 2465
rect 16683 2416 16684 2456
rect 16724 2416 16725 2456
rect 16683 2407 16725 2416
rect 16954 2456 17012 2457
rect 16954 2416 16963 2456
rect 17003 2416 17012 2456
rect 16954 2415 17012 2416
rect 17067 2456 17109 2465
rect 17067 2416 17068 2456
rect 17108 2416 17109 2456
rect 17067 2407 17109 2416
rect 17530 2456 17588 2457
rect 17530 2416 17539 2456
rect 17579 2416 17588 2456
rect 17530 2415 17588 2416
rect 21387 2456 21429 2465
rect 21387 2416 21388 2456
rect 21428 2416 21429 2456
rect 21387 2407 21429 2416
rect 22347 2456 22389 2465
rect 22347 2416 22348 2456
rect 22388 2416 22389 2456
rect 22347 2407 22389 2416
rect 22827 2456 22869 2465
rect 22827 2416 22828 2456
rect 22868 2416 22869 2456
rect 22827 2407 22869 2416
rect 25210 2456 25268 2457
rect 25210 2416 25219 2456
rect 25259 2416 25268 2456
rect 25210 2415 25268 2416
rect 28299 2456 28341 2465
rect 28299 2416 28300 2456
rect 28340 2416 28341 2456
rect 28299 2407 28341 2416
rect 29163 2456 29205 2465
rect 29163 2416 29164 2456
rect 29204 2416 29205 2456
rect 29163 2407 29205 2416
rect 6210 2398 6256 2407
rect 576 2288 31392 2312
rect 576 2248 4352 2288
rect 4720 2248 12126 2288
rect 12494 2248 19900 2288
rect 20268 2248 27674 2288
rect 28042 2248 31392 2288
rect 576 2224 31392 2248
rect 4186 2120 4244 2121
rect 4186 2080 4195 2120
rect 4235 2080 4244 2120
rect 4186 2079 4244 2080
rect 5259 2120 5301 2129
rect 5259 2080 5260 2120
rect 5300 2080 5301 2120
rect 5259 2071 5301 2080
rect 6795 2120 6837 2129
rect 6795 2080 6796 2120
rect 6836 2080 6837 2120
rect 6795 2071 6837 2080
rect 9003 2120 9045 2129
rect 9003 2080 9004 2120
rect 9044 2080 9045 2120
rect 9003 2071 9045 2080
rect 10347 2120 10389 2129
rect 10347 2080 10348 2120
rect 10388 2080 10389 2120
rect 10347 2071 10389 2080
rect 10714 2120 10772 2121
rect 10714 2080 10723 2120
rect 10763 2080 10772 2120
rect 10714 2079 10772 2080
rect 12267 2120 12309 2129
rect 12267 2080 12268 2120
rect 12308 2080 12309 2120
rect 12267 2071 12309 2080
rect 13131 2120 13173 2129
rect 13131 2080 13132 2120
rect 13172 2080 13173 2120
rect 13131 2071 13173 2080
rect 13738 2120 13796 2121
rect 13738 2080 13747 2120
rect 13787 2080 13796 2120
rect 13738 2079 13796 2080
rect 13995 2120 14037 2129
rect 13995 2080 13996 2120
rect 14036 2080 14037 2120
rect 13995 2071 14037 2080
rect 14266 2120 14324 2121
rect 14266 2080 14275 2120
rect 14315 2080 14324 2120
rect 14266 2079 14324 2080
rect 14890 2120 14948 2121
rect 14890 2080 14899 2120
rect 14939 2080 14948 2120
rect 14890 2079 14948 2080
rect 16203 2120 16245 2129
rect 16203 2080 16204 2120
rect 16244 2080 16245 2120
rect 16203 2071 16245 2080
rect 18010 2120 18068 2121
rect 18010 2080 18019 2120
rect 18059 2080 18068 2120
rect 18010 2079 18068 2080
rect 18603 2120 18645 2129
rect 18603 2080 18604 2120
rect 18644 2080 18645 2120
rect 18603 2071 18645 2080
rect 21483 2120 21525 2129
rect 21483 2080 21484 2120
rect 21524 2080 21525 2120
rect 21483 2071 21525 2080
rect 24651 2120 24693 2129
rect 24651 2080 24652 2120
rect 24692 2080 24693 2120
rect 24651 2071 24693 2080
rect 28107 2120 28149 2129
rect 28107 2080 28108 2120
rect 28148 2080 28149 2120
rect 28107 2071 28149 2080
rect 28570 2120 28628 2121
rect 28570 2080 28579 2120
rect 28619 2080 28628 2120
rect 28570 2079 28628 2080
rect 31083 2120 31125 2129
rect 31083 2080 31084 2120
rect 31124 2080 31125 2120
rect 31083 2071 31125 2080
rect 1323 2036 1365 2045
rect 1323 1996 1324 2036
rect 1364 1996 1365 2036
rect 1323 1987 1365 1996
rect 1594 2036 1652 2037
rect 1594 1996 1603 2036
rect 1643 1996 1652 2036
rect 1594 1995 1652 1996
rect 18233 2036 18275 2045
rect 18233 1996 18234 2036
rect 18274 1996 18275 2036
rect 18233 1987 18275 1996
rect 28683 2036 28725 2045
rect 28683 1996 28684 2036
rect 28724 1996 28725 2036
rect 28683 1987 28725 1996
rect 1227 1952 1269 1961
rect 1227 1912 1228 1952
rect 1268 1912 1269 1952
rect 1227 1903 1269 1912
rect 1402 1952 1460 1953
rect 1402 1912 1411 1952
rect 1451 1912 1460 1952
rect 1402 1911 1460 1912
rect 1978 1952 2036 1953
rect 1978 1912 1987 1952
rect 2027 1912 2036 1952
rect 1978 1911 2036 1912
rect 4299 1952 4341 1961
rect 4299 1912 4300 1952
rect 4340 1912 4341 1952
rect 4299 1903 4341 1912
rect 4683 1952 4725 1961
rect 4683 1912 4684 1952
rect 4724 1912 4725 1952
rect 4683 1903 4725 1912
rect 5451 1952 5493 1961
rect 5451 1912 5452 1952
rect 5492 1912 5493 1952
rect 5451 1903 5493 1912
rect 6411 1952 6453 1961
rect 6411 1912 6412 1952
rect 6452 1912 6453 1952
rect 6411 1903 6453 1912
rect 6970 1952 7028 1953
rect 6970 1912 6979 1952
rect 7019 1912 7028 1952
rect 6970 1911 7028 1912
rect 9003 1952 9045 1961
rect 9003 1912 9004 1952
rect 9044 1912 9045 1952
rect 9003 1903 9045 1912
rect 9195 1952 9237 1961
rect 9195 1912 9196 1952
rect 9236 1912 9237 1952
rect 9195 1903 9237 1912
rect 9867 1952 9909 1961
rect 9867 1912 9868 1952
rect 9908 1912 9909 1952
rect 9867 1903 9909 1912
rect 10251 1952 10293 1961
rect 10251 1912 10252 1952
rect 10292 1912 10293 1952
rect 10251 1903 10293 1912
rect 10827 1952 10869 1961
rect 10827 1912 10828 1952
rect 10868 1912 10869 1952
rect 10827 1903 10869 1912
rect 11211 1952 11253 1961
rect 11211 1912 11212 1952
rect 11252 1912 11253 1952
rect 11211 1903 11253 1912
rect 11787 1952 11829 1961
rect 11787 1912 11788 1952
rect 11828 1912 11829 1952
rect 11787 1903 11829 1912
rect 12171 1952 12213 1961
rect 12171 1912 12172 1952
rect 12212 1912 12213 1952
rect 12171 1903 12213 1912
rect 12730 1952 12788 1953
rect 12730 1912 12739 1952
rect 12779 1912 12788 1952
rect 12730 1911 12788 1912
rect 12843 1952 12885 1961
rect 12843 1912 12844 1952
rect 12884 1912 12885 1952
rect 12843 1903 12885 1912
rect 13323 1952 13365 1961
rect 13323 1912 13324 1952
rect 13364 1912 13365 1952
rect 13323 1903 13365 1912
rect 13515 1952 13557 1961
rect 13515 1912 13516 1952
rect 13556 1912 13557 1952
rect 13515 1903 13557 1912
rect 13803 1952 13845 1961
rect 13803 1912 13804 1952
rect 13844 1912 13845 1952
rect 13803 1903 13845 1912
rect 14379 1952 14421 1961
rect 14379 1912 14380 1952
rect 14420 1912 14421 1952
rect 14379 1903 14421 1912
rect 14763 1952 14805 1961
rect 14763 1912 14764 1952
rect 14804 1912 14805 1952
rect 14763 1903 14805 1912
rect 15034 1952 15092 1953
rect 16299 1952 16341 1961
rect 15034 1912 15043 1952
rect 15083 1912 15092 1952
rect 15034 1911 15092 1912
rect 15147 1943 15189 1952
rect 15147 1903 15148 1943
rect 15188 1903 15189 1943
rect 16299 1912 16300 1952
rect 16340 1912 16341 1952
rect 16299 1903 16341 1912
rect 17914 1952 17972 1953
rect 17914 1912 17923 1952
rect 17963 1912 17972 1952
rect 17914 1911 17972 1912
rect 18027 1952 18069 1961
rect 18027 1912 18028 1952
rect 18068 1912 18069 1952
rect 18027 1903 18069 1912
rect 18586 1952 18644 1953
rect 18586 1912 18595 1952
rect 18635 1912 18644 1952
rect 18586 1911 18644 1912
rect 18699 1952 18741 1961
rect 22826 1954 22868 1963
rect 18699 1912 18700 1952
rect 18740 1912 18741 1952
rect 18699 1903 18741 1912
rect 19546 1952 19604 1953
rect 19546 1912 19555 1952
rect 19595 1912 19604 1952
rect 19546 1911 19604 1912
rect 21802 1952 21860 1953
rect 21802 1912 21811 1952
rect 21851 1912 21860 1952
rect 21802 1911 21860 1912
rect 21997 1952 22055 1953
rect 21997 1912 22006 1952
rect 22046 1912 22055 1952
rect 21997 1911 22055 1912
rect 22714 1952 22772 1953
rect 22714 1912 22723 1952
rect 22763 1912 22772 1952
rect 22714 1911 22772 1912
rect 22826 1914 22827 1954
rect 22867 1914 22868 1954
rect 22826 1905 22868 1914
rect 23307 1952 23349 1961
rect 23307 1912 23308 1952
rect 23348 1912 23349 1952
rect 23307 1903 23349 1912
rect 23499 1952 23541 1961
rect 23499 1912 23500 1952
rect 23540 1912 23541 1952
rect 23499 1903 23541 1912
rect 24154 1952 24212 1953
rect 24154 1912 24163 1952
rect 24203 1912 24212 1952
rect 24154 1911 24212 1912
rect 24459 1952 24501 1961
rect 24459 1912 24460 1952
rect 24500 1912 24501 1952
rect 24459 1903 24501 1912
rect 25323 1952 25365 1961
rect 25323 1912 25324 1952
rect 25364 1912 25365 1952
rect 25323 1903 25365 1912
rect 26170 1952 26228 1953
rect 26170 1912 26179 1952
rect 26219 1912 26228 1952
rect 26170 1911 26228 1912
rect 28477 1952 28519 1961
rect 29835 1952 29877 1961
rect 28477 1912 28478 1952
rect 28518 1912 28519 1952
rect 28477 1903 28519 1912
rect 28779 1943 28821 1952
rect 28779 1903 28780 1943
rect 28820 1903 28821 1943
rect 29835 1912 29836 1952
rect 29876 1912 29877 1952
rect 29835 1903 29877 1912
rect 30123 1952 30165 1961
rect 30123 1912 30124 1952
rect 30164 1912 30165 1952
rect 30123 1903 30165 1912
rect 30987 1952 31029 1961
rect 30987 1912 30988 1952
rect 31028 1912 31029 1952
rect 30987 1903 31029 1912
rect 31179 1952 31221 1961
rect 31179 1912 31180 1952
rect 31220 1912 31221 1952
rect 31179 1903 31221 1912
rect 15147 1894 15189 1903
rect 28779 1894 28821 1903
rect 3531 1868 3573 1877
rect 3531 1828 3532 1868
rect 3572 1828 3573 1868
rect 3531 1819 3573 1828
rect 19179 1868 19221 1877
rect 19179 1828 19180 1868
rect 19220 1828 19221 1868
rect 19179 1819 19221 1828
rect 25803 1868 25845 1877
rect 25803 1828 25804 1868
rect 25844 1828 25845 1868
rect 25803 1819 25845 1828
rect 27723 1868 27765 1877
rect 27723 1828 27724 1868
rect 27764 1828 27765 1868
rect 27723 1819 27765 1828
rect 29146 1868 29204 1869
rect 29146 1828 29155 1868
rect 29195 1828 29204 1868
rect 29146 1827 29204 1828
rect 3915 1784 3957 1793
rect 3915 1744 3916 1784
rect 3956 1744 3957 1784
rect 3915 1735 3957 1744
rect 7023 1784 7065 1793
rect 7023 1744 7024 1784
rect 7064 1744 7065 1784
rect 7023 1735 7065 1744
rect 7563 1784 7605 1793
rect 7563 1744 7564 1784
rect 7604 1744 7605 1784
rect 7563 1735 7605 1744
rect 15435 1784 15477 1793
rect 15435 1744 15436 1784
rect 15476 1744 15477 1784
rect 15435 1735 15477 1744
rect 16779 1784 16821 1793
rect 16779 1744 16780 1784
rect 16820 1744 16821 1784
rect 16779 1735 16821 1744
rect 21099 1784 21141 1793
rect 21099 1744 21100 1784
rect 21140 1744 21141 1784
rect 21099 1735 21141 1744
rect 23002 1784 23060 1785
rect 23002 1744 23011 1784
rect 23051 1744 23060 1784
rect 23002 1743 23060 1744
rect 23787 1784 23829 1793
rect 23787 1744 23788 1784
rect 23828 1744 23829 1784
rect 23787 1735 23829 1744
rect 24459 1784 24501 1793
rect 24459 1744 24460 1784
rect 24500 1744 24501 1784
rect 24459 1735 24501 1744
rect 5050 1700 5108 1701
rect 5050 1660 5059 1700
rect 5099 1660 5108 1700
rect 5050 1659 5108 1660
rect 5739 1700 5781 1709
rect 5739 1660 5740 1700
rect 5780 1660 5781 1700
rect 5739 1651 5781 1660
rect 13419 1700 13461 1709
rect 13419 1660 13420 1700
rect 13460 1660 13461 1700
rect 13419 1651 13461 1660
rect 18219 1700 18261 1709
rect 18219 1660 18220 1700
rect 18260 1660 18261 1700
rect 18219 1651 18261 1660
rect 18891 1700 18933 1709
rect 18891 1660 18892 1700
rect 18932 1660 18933 1700
rect 18891 1651 18933 1660
rect 23307 1700 23349 1709
rect 23307 1660 23308 1700
rect 23348 1660 23349 1700
rect 23307 1651 23349 1660
rect 30795 1700 30837 1709
rect 30795 1660 30796 1700
rect 30836 1660 30837 1700
rect 30795 1651 30837 1660
rect 576 1532 31392 1556
rect 576 1492 3112 1532
rect 3480 1492 10886 1532
rect 11254 1492 18660 1532
rect 19028 1492 26434 1532
rect 26802 1492 31392 1532
rect 576 1468 31392 1492
rect 8427 1364 8469 1373
rect 8427 1324 8428 1364
rect 8468 1324 8469 1364
rect 8427 1315 8469 1324
rect 10347 1364 10389 1373
rect 10347 1324 10348 1364
rect 10388 1324 10389 1364
rect 10347 1315 10389 1324
rect 11211 1364 11253 1373
rect 11211 1324 11212 1364
rect 11252 1324 11253 1364
rect 11211 1315 11253 1324
rect 12843 1364 12885 1373
rect 12843 1324 12844 1364
rect 12884 1324 12885 1364
rect 12843 1315 12885 1324
rect 17643 1364 17685 1373
rect 17643 1324 17644 1364
rect 17684 1324 17685 1364
rect 17643 1315 17685 1324
rect 25227 1364 25269 1373
rect 25227 1324 25228 1364
rect 25268 1324 25269 1364
rect 25227 1315 25269 1324
rect 28491 1364 28533 1373
rect 28491 1324 28492 1364
rect 28532 1324 28533 1364
rect 28491 1315 28533 1324
rect 2667 1280 2709 1289
rect 2667 1240 2668 1280
rect 2708 1240 2709 1280
rect 2667 1231 2709 1240
rect 4378 1280 4436 1281
rect 4378 1240 4387 1280
rect 4427 1240 4436 1280
rect 4378 1239 4436 1240
rect 4827 1280 4869 1289
rect 4827 1240 4828 1280
rect 4868 1240 4869 1280
rect 4827 1231 4869 1240
rect 10539 1280 10581 1289
rect 10539 1240 10540 1280
rect 10580 1240 10581 1280
rect 10539 1231 10581 1240
rect 18987 1280 19029 1289
rect 18987 1240 18988 1280
rect 19028 1240 19029 1280
rect 18987 1231 19029 1240
rect 20907 1280 20949 1289
rect 20907 1240 20908 1280
rect 20948 1240 20949 1280
rect 20907 1231 20949 1240
rect 21675 1280 21717 1289
rect 21675 1240 21676 1280
rect 21716 1240 21717 1280
rect 21675 1231 21717 1240
rect 25035 1280 25077 1289
rect 25035 1240 25036 1280
rect 25076 1240 25077 1280
rect 25035 1231 25077 1240
rect 5050 1196 5108 1197
rect 5050 1156 5059 1196
rect 5099 1156 5108 1196
rect 5050 1155 5108 1156
rect 6507 1196 6549 1205
rect 6507 1156 6508 1196
rect 6548 1156 6549 1196
rect 5922 1145 5968 1154
rect 6507 1147 6549 1156
rect 24651 1196 24693 1205
rect 24651 1156 24652 1196
rect 24692 1156 24693 1196
rect 24651 1147 24693 1156
rect 26842 1196 26900 1197
rect 26842 1156 26851 1196
rect 26891 1156 26900 1196
rect 26842 1155 26900 1156
rect 30778 1196 30836 1197
rect 30778 1156 30787 1196
rect 30827 1156 30836 1196
rect 30778 1155 30836 1156
rect 4203 1112 4245 1121
rect 4203 1072 4204 1112
rect 4244 1072 4245 1112
rect 4203 1063 4245 1072
rect 4378 1112 4436 1113
rect 4378 1072 4387 1112
rect 4427 1072 4436 1112
rect 4378 1071 4436 1072
rect 4683 1112 4725 1121
rect 4683 1072 4684 1112
rect 4724 1072 4725 1112
rect 4683 1063 4725 1072
rect 4918 1112 4960 1121
rect 4918 1072 4919 1112
rect 4959 1072 4960 1112
rect 4918 1063 4960 1072
rect 5164 1112 5206 1121
rect 5164 1072 5165 1112
rect 5205 1072 5206 1112
rect 5164 1063 5206 1072
rect 5434 1112 5492 1113
rect 5434 1072 5443 1112
rect 5483 1072 5492 1112
rect 5922 1105 5923 1145
rect 5963 1105 5968 1145
rect 5922 1096 5968 1105
rect 6874 1112 6932 1113
rect 5434 1071 5492 1072
rect 6874 1072 6883 1112
rect 6923 1072 6932 1112
rect 6874 1071 6932 1072
rect 9195 1112 9237 1121
rect 9195 1072 9196 1112
rect 9236 1072 9237 1112
rect 9195 1063 9237 1072
rect 9867 1112 9909 1121
rect 9867 1072 9868 1112
rect 9908 1072 9909 1112
rect 9867 1063 9909 1072
rect 10138 1112 10196 1113
rect 10138 1072 10147 1112
rect 10187 1072 10196 1112
rect 10138 1071 10196 1072
rect 10906 1112 10964 1113
rect 10906 1072 10915 1112
rect 10955 1072 10964 1112
rect 10906 1071 10964 1072
rect 11383 1112 11441 1113
rect 11383 1072 11392 1112
rect 11432 1072 11441 1112
rect 11383 1071 11441 1072
rect 11547 1112 11589 1121
rect 11547 1072 11548 1112
rect 11588 1072 11589 1112
rect 11547 1063 11589 1072
rect 12634 1112 12692 1113
rect 12634 1072 12643 1112
rect 12683 1072 12692 1112
rect 12634 1071 12692 1072
rect 12747 1112 12789 1121
rect 12747 1072 12748 1112
rect 12788 1072 12789 1112
rect 12747 1063 12789 1072
rect 13174 1112 13216 1121
rect 13174 1072 13175 1112
rect 13215 1072 13216 1112
rect 13174 1063 13216 1072
rect 13306 1112 13364 1113
rect 13306 1072 13315 1112
rect 13355 1072 13364 1112
rect 13306 1071 13364 1072
rect 13419 1112 13461 1121
rect 13419 1072 13420 1112
rect 13460 1072 13461 1112
rect 13419 1063 13461 1072
rect 14283 1112 14325 1121
rect 14283 1072 14284 1112
rect 14324 1072 14325 1112
rect 14283 1063 14325 1072
rect 14458 1112 14516 1113
rect 14458 1072 14467 1112
rect 14507 1072 14516 1112
rect 14458 1071 14516 1072
rect 14811 1112 14853 1121
rect 14811 1072 14812 1112
rect 14852 1072 14853 1112
rect 14811 1063 14853 1072
rect 14955 1112 14997 1121
rect 14955 1072 14956 1112
rect 14996 1072 14997 1112
rect 14955 1063 14997 1072
rect 16090 1112 16148 1113
rect 16090 1072 16099 1112
rect 16139 1072 16148 1112
rect 16090 1071 16148 1072
rect 18795 1112 18837 1121
rect 18795 1072 18796 1112
rect 18836 1072 18837 1112
rect 18795 1063 18837 1072
rect 18910 1112 18952 1121
rect 18910 1072 18911 1112
rect 18951 1072 18952 1112
rect 18910 1063 18952 1072
rect 19083 1112 19125 1121
rect 19083 1072 19084 1112
rect 19124 1072 19125 1112
rect 19083 1063 19125 1072
rect 20043 1112 20085 1121
rect 20043 1072 20044 1112
rect 20084 1072 20085 1112
rect 20043 1063 20085 1072
rect 20715 1112 20757 1121
rect 20715 1072 20716 1112
rect 20756 1072 20757 1112
rect 20715 1063 20757 1072
rect 21466 1112 21524 1113
rect 21466 1072 21475 1112
rect 21515 1072 21524 1112
rect 21466 1071 21524 1072
rect 23098 1112 23156 1113
rect 23098 1072 23107 1112
rect 23147 1072 23156 1112
rect 23098 1071 23156 1072
rect 25851 1112 25893 1121
rect 25851 1072 25852 1112
rect 25892 1072 25893 1112
rect 25851 1063 25893 1072
rect 26091 1112 26133 1121
rect 26091 1072 26092 1112
rect 26132 1072 26133 1112
rect 26091 1063 26133 1072
rect 26283 1112 26325 1121
rect 26283 1072 26284 1112
rect 26324 1072 26325 1112
rect 26283 1063 26325 1072
rect 27531 1112 27573 1121
rect 27531 1072 27532 1112
rect 27572 1072 27573 1112
rect 27531 1063 27573 1072
rect 30394 1112 30452 1113
rect 30394 1072 30403 1112
rect 30443 1072 30452 1112
rect 30394 1071 30452 1072
rect 5643 1028 5685 1037
rect 5643 988 5644 1028
rect 5684 988 5685 1028
rect 5643 979 5685 988
rect 5753 1028 5795 1037
rect 5753 988 5754 1028
rect 5794 988 5795 1028
rect 5753 979 5795 988
rect 11019 1028 11061 1037
rect 11019 988 11020 1028
rect 11060 988 11061 1028
rect 11019 979 11061 988
rect 11225 1028 11267 1037
rect 11225 988 11226 1028
rect 11266 988 11267 1028
rect 11225 979 11267 988
rect 13498 1028 13556 1029
rect 13498 988 13507 1028
rect 13547 988 13556 1028
rect 13498 987 13556 988
rect 15706 1028 15764 1029
rect 15706 988 15715 1028
rect 15755 988 15764 1028
rect 15706 987 15764 988
rect 22714 1028 22772 1029
rect 22714 988 22723 1028
rect 22763 988 22772 1028
rect 22714 987 22772 988
rect 26187 1028 26229 1037
rect 26187 988 26188 1028
rect 26228 988 26229 1028
rect 26187 979 26229 988
rect 5242 944 5300 945
rect 5242 904 5251 944
rect 5291 904 5300 944
rect 5242 903 5300 904
rect 5530 944 5588 945
rect 5530 904 5539 944
rect 5579 904 5588 944
rect 5530 903 5588 904
rect 6075 944 6117 953
rect 6075 904 6076 944
rect 6116 904 6117 944
rect 6075 895 6117 904
rect 8811 944 8853 953
rect 8811 904 8812 944
rect 8852 904 8853 944
rect 8811 895 8853 904
rect 13035 944 13077 953
rect 13035 904 13036 944
rect 13076 904 13077 944
rect 13035 895 13077 904
rect 14379 944 14421 953
rect 14379 904 14380 944
rect 14420 904 14421 944
rect 14379 895 14421 904
rect 14650 944 14708 945
rect 14650 904 14659 944
rect 14699 904 14708 944
rect 14650 903 14708 904
rect 18027 944 18069 953
rect 18027 904 18028 944
rect 18068 904 18069 944
rect 18027 895 18069 904
rect 21675 944 21717 953
rect 21675 904 21676 944
rect 21716 904 21717 944
rect 21675 895 21717 904
rect 576 776 31392 800
rect 576 736 4352 776
rect 4720 736 12126 776
rect 12494 736 19900 776
rect 20268 736 27674 776
rect 28042 736 31392 776
rect 576 712 31392 736
<< via1 >>
rect 4352 27952 4720 27992
rect 12126 27952 12494 27992
rect 19900 27952 20268 27992
rect 27674 27952 28042 27992
rect 11203 27700 11243 27740
rect 22339 27700 22379 27740
rect 25123 27700 25163 27740
rect 25507 27700 25547 27740
rect 3619 27616 3659 27656
rect 6115 27616 6155 27656
rect 8611 27616 8651 27656
rect 11587 27616 11627 27656
rect 14188 27616 14228 27656
rect 16387 27616 16427 27656
rect 17068 27616 17108 27656
rect 18115 27616 18155 27656
rect 22723 27616 22763 27656
rect 25036 27616 25076 27656
rect 25219 27616 25259 27656
rect 25324 27616 25364 27656
rect 25891 27616 25931 27656
rect 28012 27616 28052 27656
rect 28867 27607 28907 27647
rect 29347 27607 29387 27647
rect 29827 27607 29867 27647
rect 3244 27532 3284 27572
rect 5740 27532 5780 27572
rect 8236 27532 8276 27572
rect 16771 27532 16811 27572
rect 17740 27532 17780 27572
rect 29020 27532 29060 27572
rect 29500 27532 29540 27572
rect 29980 27532 30020 27572
rect 30892 27532 30932 27572
rect 3052 27448 3092 27488
rect 13708 27448 13748 27488
rect 20236 27448 20276 27488
rect 20812 27448 20852 27488
rect 30316 27448 30356 27488
rect 31084 27448 31124 27488
rect 5548 27364 5588 27404
rect 8044 27364 8084 27404
rect 10540 27364 10580 27404
rect 13516 27364 13556 27404
rect 14044 27364 14084 27404
rect 14476 27364 14516 27404
rect 16924 27364 16964 27404
rect 20044 27364 20084 27404
rect 24652 27364 24692 27404
rect 27820 27364 27860 27404
rect 28684 27364 28724 27404
rect 30652 27364 30692 27404
rect 3112 27196 3480 27236
rect 10886 27196 11254 27236
rect 18660 27196 19028 27236
rect 26434 27196 26802 27236
rect 11692 27028 11732 27068
rect 14083 27028 14123 27068
rect 16780 27028 16820 27068
rect 17932 27028 17972 27068
rect 26851 27028 26891 27068
rect 2764 26944 2804 26984
rect 3148 26944 3188 26984
rect 3532 26944 3572 26984
rect 3724 26944 3764 26984
rect 5452 26944 5492 26984
rect 6700 26944 6740 26984
rect 9292 26944 9332 26984
rect 11884 26944 11924 26984
rect 13708 26944 13748 26984
rect 15724 26944 15764 26984
rect 17740 26944 17780 26984
rect 24460 26944 24500 26984
rect 27820 26944 27860 26984
rect 8476 26860 8516 26900
rect 15244 26860 15284 26900
rect 23308 26860 23348 26900
rect 24835 26860 24875 26900
rect 28963 26860 29003 26900
rect 3724 26776 3764 26816
rect 3916 26776 3956 26816
rect 6316 26776 6356 26816
rect 7468 26776 7508 26816
rect 8320 26776 8360 26816
rect 10252 26776 10292 26816
rect 10396 26776 10436 26816
rect 10732 26776 10772 26816
rect 10828 26776 10868 26816
rect 11020 26776 11060 26816
rect 12556 26776 12596 26816
rect 12748 26776 12788 26816
rect 14380 26776 14420 26816
rect 14572 26776 14612 26816
rect 16108 26776 16148 26816
rect 17068 26776 17108 26816
rect 17347 26776 17387 26816
rect 18604 26776 18644 26816
rect 19468 26776 19508 26816
rect 20131 26776 20171 26816
rect 23800 26776 23840 26816
rect 23968 26776 24008 26816
rect 25516 26776 25556 26816
rect 25900 26776 25940 26816
rect 26021 26776 26061 26816
rect 26323 26776 26363 26816
rect 27052 26776 27092 26816
rect 27148 26776 27188 26816
rect 27283 26776 27323 26816
rect 28387 26776 28427 26816
rect 28492 26776 28532 26816
rect 30883 26776 30923 26816
rect 8140 26692 8180 26732
rect 10526 26692 10566 26732
rect 14078 26692 14118 26732
rect 17452 26692 17492 26732
rect 18787 26692 18827 26732
rect 19747 26692 19787 26732
rect 25699 26692 25739 26732
rect 26846 26692 26886 26732
rect 31267 26692 31307 26732
rect 4300 26608 4340 26648
rect 4684 26608 4724 26648
rect 5068 26608 5108 26648
rect 5644 26608 5684 26648
rect 7276 26608 7316 26648
rect 8812 26608 8852 26648
rect 10627 26608 10667 26648
rect 13420 26608 13460 26648
rect 14284 26608 14324 26648
rect 22060 26608 22100 26648
rect 23068 26608 23108 26648
rect 23635 26608 23675 26648
rect 24124 26608 24164 26648
rect 26002 26608 26042 26648
rect 26524 26608 26564 26648
rect 27484 26608 27524 26648
rect 28780 26608 28820 26648
rect 4352 26440 4720 26480
rect 12126 26440 12494 26480
rect 19900 26440 20268 26480
rect 27674 26440 28042 26480
rect 4723 26272 4763 26312
rect 7948 26272 7988 26312
rect 8284 26272 8324 26312
rect 8716 26272 8756 26312
rect 9667 26272 9707 26312
rect 9964 26272 10004 26312
rect 11395 26272 11435 26312
rect 11923 26272 11963 26312
rect 15148 26272 15188 26312
rect 17443 26272 17483 26312
rect 18115 26272 18155 26312
rect 18796 26272 18836 26312
rect 19756 26272 19796 26312
rect 23971 26272 24011 26312
rect 26092 26272 26132 26312
rect 30508 26272 30548 26312
rect 5164 26188 5204 26228
rect 5635 26188 5675 26228
rect 10435 26179 10475 26219
rect 12835 26188 12875 26228
rect 15532 26188 15572 26228
rect 18590 26188 18630 26228
rect 18691 26188 18731 26228
rect 24076 26188 24116 26228
rect 27859 26188 27899 26228
rect 3619 26104 3659 26144
rect 4480 26095 4520 26135
rect 4579 26104 4619 26144
rect 5068 26104 5108 26144
rect 5260 26104 5300 26144
rect 6019 26104 6059 26144
rect 8140 26104 8180 26144
rect 8425 26104 8465 26144
rect 8551 26104 8591 26144
rect 8677 26104 8717 26144
rect 8908 26104 8948 26144
rect 9048 26104 9088 26144
rect 9157 26104 9197 26144
rect 9772 26104 9812 26144
rect 10147 26104 10187 26144
rect 10252 26095 10292 26135
rect 10531 26104 10571 26144
rect 10665 26104 10705 26144
rect 11068 26062 11108 26102
rect 11308 26104 11348 26144
rect 12088 26104 12128 26144
rect 12237 26104 12277 26144
rect 12399 26104 12439 26144
rect 12691 26104 12731 26144
rect 13219 26104 13259 26144
rect 15436 26104 15476 26144
rect 15628 26104 15668 26144
rect 16003 26104 16043 26144
rect 16108 26104 16148 26144
rect 16555 26104 16595 26144
rect 16780 26104 16820 26144
rect 17548 26104 17588 26144
rect 17932 26104 17972 26144
rect 18220 26104 18260 26144
rect 18892 26095 18932 26135
rect 19070 26104 19110 26144
rect 19276 26104 19316 26144
rect 19372 26095 19412 26135
rect 20428 26104 20468 26144
rect 20716 26104 20756 26144
rect 20953 26104 20993 26144
rect 21772 26104 21812 26144
rect 23873 26104 23913 26144
rect 24172 26095 24212 26135
rect 24739 26095 24779 26135
rect 25507 26095 25547 26135
rect 25996 26104 26036 26144
rect 26179 26104 26219 26144
rect 26872 26104 26912 26144
rect 27057 26104 27097 26144
rect 27244 26104 27284 26144
rect 27493 26104 27533 26144
rect 28054 26104 28094 26144
rect 28204 26104 28244 26144
rect 4003 26020 4043 26060
rect 11203 26020 11243 26060
rect 12559 26020 12599 26060
rect 16675 26020 16715 26060
rect 16876 26020 16916 26060
rect 20620 26020 20660 26060
rect 20835 26020 20875 26060
rect 24892 26020 24932 26060
rect 25660 26020 25700 26060
rect 27366 26062 27406 26102
rect 28387 26104 28427 26144
rect 28819 26104 28859 26144
rect 29014 26104 29054 26144
rect 29155 26104 29195 26144
rect 29836 26104 29876 26144
rect 30412 26104 30452 26144
rect 30604 26104 30644 26144
rect 26668 26020 26708 26060
rect 30988 26020 31028 26060
rect 1708 25936 1748 25976
rect 4195 25936 4235 25976
rect 9196 25936 9236 25976
rect 12460 25936 12500 25976
rect 16291 25936 16331 25976
rect 18412 25936 18452 25976
rect 22252 25936 22292 25976
rect 26428 25936 26468 25976
rect 27532 25936 27572 25976
rect 30028 25936 30068 25976
rect 30748 25936 30788 25976
rect 10147 25852 10187 25892
rect 19075 25852 19115 25892
rect 21100 25852 21140 25892
rect 26860 25852 26900 25892
rect 28387 25852 28427 25892
rect 3112 25684 3480 25724
rect 10886 25684 11254 25724
rect 18660 25684 19028 25724
rect 26434 25684 26802 25724
rect 5539 25516 5579 25556
rect 9283 25516 9323 25556
rect 10828 25516 10868 25556
rect 12652 25516 12692 25556
rect 16156 25516 16196 25556
rect 19900 25516 19940 25556
rect 25420 25516 25460 25556
rect 5155 25432 5195 25472
rect 6892 25432 6932 25472
rect 13036 25432 13076 25472
rect 14668 25432 14708 25472
rect 24844 25432 24884 25472
rect 26956 25432 26996 25472
rect 28099 25432 28139 25472
rect 11155 25348 11195 25388
rect 23884 25348 23924 25388
rect 3139 25264 3179 25304
rect 4481 25264 4521 25304
rect 4780 25289 4820 25329
rect 4972 25264 5012 25304
rect 5155 25264 5195 25304
rect 5356 25264 5396 25304
rect 5539 25264 5579 25304
rect 6508 25264 6548 25304
rect 8236 25264 8276 25304
rect 9283 25264 9323 25304
rect 9411 25264 9451 25304
rect 9533 25264 9573 25304
rect 9667 25264 9707 25304
rect 9844 25264 9884 25304
rect 11347 25306 11387 25346
rect 10540 25264 10580 25304
rect 10662 25264 10702 25304
rect 10789 25264 10829 25304
rect 11488 25264 11528 25304
rect 11980 25264 12020 25304
rect 12355 25264 12395 25304
rect 12663 25264 12703 25304
rect 14284 25264 14324 25304
rect 14476 25264 14516 25304
rect 15340 25264 15380 25304
rect 16492 25264 16532 25304
rect 16780 25264 16820 25304
rect 17347 25264 17387 25304
rect 17462 25264 17502 25304
rect 18109 25264 18149 25304
rect 18220 25264 18260 25304
rect 18700 25264 18740 25304
rect 18892 25264 18932 25304
rect 19372 25264 19412 25304
rect 19660 25264 19700 25304
rect 20044 25264 20084 25304
rect 20332 25264 20372 25304
rect 20611 25264 20651 25304
rect 21571 25264 21611 25304
rect 23980 25264 24020 25304
rect 24099 25264 24139 25304
rect 24220 25306 24260 25346
rect 24395 25297 24435 25337
rect 24547 25255 24587 25295
rect 24652 25264 24692 25304
rect 24844 25264 24884 25304
rect 24969 25264 25009 25304
rect 25137 25299 25177 25339
rect 25555 25339 25595 25379
rect 28579 25348 28619 25388
rect 25324 25264 25364 25304
rect 25663 25264 25703 25304
rect 25900 25264 25940 25304
rect 26371 25264 26411 25304
rect 26476 25264 26516 25304
rect 26860 25264 26900 25304
rect 26982 25264 27022 25304
rect 27109 25264 27149 25304
rect 27811 25264 27851 25304
rect 27918 25264 27958 25304
rect 28439 25264 28479 25304
rect 28684 25264 28724 25304
rect 29347 25264 29387 25304
rect 3523 25180 3563 25220
rect 11644 25180 11684 25220
rect 14380 25180 14420 25220
rect 20716 25180 20756 25220
rect 21187 25180 21227 25220
rect 26659 25180 26699 25220
rect 28771 25180 28811 25220
rect 28963 25180 29003 25220
rect 1228 25096 1268 25136
rect 4579 25096 4619 25136
rect 4684 25096 4724 25136
rect 5836 25096 5876 25136
rect 7276 25096 7316 25136
rect 8131 25096 8171 25136
rect 8428 25096 8468 25136
rect 12451 25096 12491 25136
rect 16012 25096 16052 25136
rect 17740 25096 17780 25136
rect 17923 25096 17963 25136
rect 18883 25096 18923 25136
rect 19171 25096 19211 25136
rect 21052 25096 21092 25136
rect 23500 25096 23540 25136
rect 24364 25096 24404 25136
rect 25420 25096 25460 25136
rect 26380 25096 26420 25136
rect 31276 25096 31316 25136
rect 4352 24928 4720 24968
rect 12126 24928 12494 24968
rect 19900 24928 20268 24968
rect 27674 24928 28042 24968
rect 4099 24760 4139 24800
rect 4972 24760 5012 24800
rect 5548 24760 5588 24800
rect 8140 24760 8180 24800
rect 8899 24760 8939 24800
rect 9196 24760 9236 24800
rect 10627 24760 10667 24800
rect 14755 24760 14795 24800
rect 16819 24760 16859 24800
rect 17827 24760 17867 24800
rect 17932 24760 17972 24800
rect 21196 24760 21236 24800
rect 23500 24760 23540 24800
rect 25324 24760 25364 24800
rect 26380 24760 26420 24800
rect 27052 24760 27092 24800
rect 28099 24760 28139 24800
rect 28876 24760 28916 24800
rect 10051 24667 10091 24707
rect 18039 24676 18079 24716
rect 19555 24667 19595 24707
rect 25219 24676 25259 24716
rect 2188 24592 2228 24632
rect 4204 24592 4244 24632
rect 4588 24592 4628 24632
rect 4780 24592 4820 24632
rect 5155 24592 5195 24632
rect 5452 24592 5492 24632
rect 5635 24592 5675 24632
rect 6211 24592 6251 24632
rect 8301 24592 8341 24632
rect 8449 24592 8489 24632
rect 8741 24592 8781 24632
rect 9004 24592 9044 24632
rect 9763 24592 9803 24632
rect 9868 24583 9908 24623
rect 10155 24592 10195 24632
rect 10324 24592 10364 24632
rect 10915 24592 10955 24632
rect 11447 24592 11487 24632
rect 11692 24592 11732 24632
rect 12355 24592 12395 24632
rect 14423 24592 14463 24632
rect 14563 24592 14603 24632
rect 14668 24592 14708 24632
rect 14947 24583 14987 24623
rect 16108 24592 16148 24632
rect 16984 24592 17024 24632
rect 17731 24592 17771 24632
rect 18215 24587 18255 24627
rect 18412 24592 18452 24632
rect 18700 24592 18740 24632
rect 18988 24592 19028 24632
rect 19132 24592 19172 24632
rect 19267 24592 19307 24632
rect 19372 24583 19412 24623
rect 19651 24592 19691 24632
rect 19785 24592 19825 24632
rect 19996 24592 20036 24632
rect 20297 24592 20337 24632
rect 20467 24592 20507 24632
rect 21868 24592 21908 24632
rect 22828 24592 22868 24632
rect 23596 24592 23636 24632
rect 24333 24592 24373 24632
rect 24495 24592 24535 24632
rect 24773 24592 24813 24632
rect 25118 24592 25158 24632
rect 25426 24589 25466 24629
rect 25849 24583 25889 24623
rect 25951 24592 25991 24632
rect 26083 24583 26123 24623
rect 26188 24592 26228 24632
rect 26369 24592 26409 24632
rect 26577 24592 26617 24632
rect 26956 24592 26996 24632
rect 27139 24592 27179 24632
rect 27436 24592 27476 24632
rect 27628 24592 27668 24632
rect 27916 24592 27956 24632
rect 28108 24592 28148 24632
rect 28298 24619 28338 24659
rect 28492 24592 28532 24632
rect 29548 24592 29588 24632
rect 30796 24592 30836 24632
rect 5836 24508 5876 24548
rect 8620 24508 8660 24548
rect 10531 24508 10571 24548
rect 11107 24508 11147 24548
rect 11587 24508 11627 24548
rect 11788 24508 11828 24548
rect 11980 24508 12020 24548
rect 15100 24508 15140 24548
rect 18316 24508 18356 24548
rect 20140 24508 20180 24548
rect 22147 24508 22187 24548
rect 23500 24508 23540 24548
rect 24652 24508 24692 24548
rect 27724 24508 27764 24548
rect 28396 24508 28436 24548
rect 1900 24424 1940 24464
rect 3052 24424 3092 24464
rect 4396 24424 4436 24464
rect 5200 24424 5240 24464
rect 8524 24424 8564 24464
rect 14284 24424 14324 24464
rect 17164 24424 17204 24464
rect 20236 24424 20276 24464
rect 23020 24424 23060 24464
rect 24556 24424 24596 24464
rect 29932 24424 29972 24464
rect 30988 24424 31028 24464
rect 2860 24340 2900 24380
rect 4588 24340 4628 24380
rect 9763 24340 9803 24380
rect 13900 24340 13940 24380
rect 15436 24340 15476 24380
rect 19267 24340 19307 24380
rect 25900 24340 25940 24380
rect 27139 24340 27179 24380
rect 30124 24340 30164 24380
rect 3112 24172 3480 24212
rect 10886 24172 11254 24212
rect 18660 24172 19028 24212
rect 26434 24172 26802 24212
rect 5251 24004 5291 24044
rect 7939 24004 7979 24044
rect 9292 24004 9332 24044
rect 9676 24004 9716 24044
rect 12268 24004 12308 24044
rect 18604 24004 18644 24044
rect 19459 24004 19499 24044
rect 28204 24004 28244 24044
rect 31276 24004 31316 24044
rect 3148 23920 3188 23960
rect 6220 23920 6260 23960
rect 7084 23920 7124 23960
rect 9100 23920 9140 23960
rect 11971 23920 12011 23960
rect 18860 23911 18900 23951
rect 27532 23920 27572 23960
rect 2947 23836 2987 23876
rect 4243 23836 4283 23876
rect 5011 23827 5051 23867
rect 12547 23836 12587 23876
rect 14515 23836 14555 23876
rect 15436 23836 15476 23876
rect 19804 23836 19844 23876
rect 23107 23836 23147 23876
rect 24700 23836 24740 23876
rect 28972 23836 29012 23876
rect 2563 23752 2603 23792
rect 3532 23743 3572 23783
rect 3820 23752 3860 23792
rect 4438 23752 4478 23792
rect 4875 23752 4915 23792
rect 5113 23752 5153 23792
rect 5548 23752 5588 23792
rect 6892 23752 6932 23792
rect 7937 23752 7977 23792
rect 8236 23752 8276 23792
rect 8524 23752 8564 23792
rect 8716 23752 8756 23792
rect 9292 23752 9332 23792
rect 9484 23752 9524 23792
rect 9676 23752 9716 23792
rect 9868 23752 9908 23792
rect 10684 23752 10724 23792
rect 10924 23752 10964 23792
rect 11788 23752 11828 23792
rect 11971 23752 12011 23792
rect 12155 23752 12195 23792
rect 12364 23752 12404 23792
rect 13228 23752 13268 23792
rect 14188 23752 14228 23792
rect 14680 23752 14720 23792
rect 15047 23752 15087 23792
rect 15244 23752 15284 23792
rect 15811 23752 15851 23792
rect 17932 23752 17972 23792
rect 18883 23752 18923 23792
rect 19276 23752 19316 23792
rect 19459 23752 19499 23792
rect 19648 23752 19688 23792
rect 22723 23752 22763 23792
rect 23452 23752 23492 23792
rect 23596 23752 23636 23792
rect 24268 23752 24308 23792
rect 24364 23752 24404 23792
rect 24499 23752 24539 23792
rect 24983 23752 25023 23792
rect 25123 23752 25163 23792
rect 25226 23752 25266 23792
rect 25516 23752 25556 23792
rect 25658 23752 25698 23792
rect 26188 23752 26228 23792
rect 26380 23752 26420 23792
rect 26668 23752 26708 23792
rect 27244 23752 27284 23792
rect 27427 23752 27467 23792
rect 27532 23752 27572 23792
rect 27868 23752 27908 23792
rect 28011 23752 28051 23792
rect 28387 23752 28427 23792
rect 28698 23752 28738 23792
rect 29347 23752 29387 23792
rect 643 23668 683 23708
rect 3436 23668 3476 23708
rect 4780 23668 4820 23708
rect 5249 23668 5289 23708
rect 10051 23668 10091 23708
rect 13507 23668 13547 23708
rect 24062 23668 24102 23708
rect 24163 23668 24203 23708
rect 28588 23668 28628 23708
rect 5452 23584 5492 23624
rect 8140 23584 8180 23624
rect 8707 23584 8747 23624
rect 11596 23584 11636 23624
rect 15235 23584 15275 23624
rect 17740 23584 17780 23624
rect 19075 23584 19115 23624
rect 20812 23584 20852 23624
rect 23299 23584 23339 23624
rect 24268 23584 24308 23624
rect 25315 23584 25355 23624
rect 25804 23584 25844 23624
rect 26188 23584 26228 23624
rect 26563 23584 26603 23624
rect 26860 23584 26900 23624
rect 27916 23584 27956 23624
rect 28483 23584 28523 23624
rect 4352 23416 4720 23456
rect 12126 23416 12494 23456
rect 19900 23416 20268 23456
rect 27674 23416 28042 23456
rect 4867 23248 4907 23288
rect 5068 23248 5108 23288
rect 11356 23248 11396 23288
rect 12556 23248 12596 23288
rect 15532 23248 15572 23288
rect 16531 23248 16571 23288
rect 20419 23248 20459 23288
rect 23596 23248 23636 23288
rect 27763 23248 27803 23288
rect 31276 23248 31316 23288
rect 5539 23164 5579 23204
rect 8419 23164 8459 23204
rect 11059 23164 11099 23204
rect 26563 23155 26603 23195
rect 2284 23080 2324 23120
rect 3148 23080 3188 23120
rect 3532 23080 3572 23120
rect 4684 23080 4724 23120
rect 4876 23080 4916 23120
rect 5164 23080 5204 23120
rect 5401 23080 5441 23120
rect 5923 23080 5963 23120
rect 8044 23080 8084 23120
rect 8803 23080 8843 23120
rect 11224 23080 11264 23120
rect 11774 23080 11814 23120
rect 11886 23080 11926 23120
rect 12076 23080 12116 23120
rect 12268 23080 12308 23120
rect 12412 23059 12452 23099
rect 12517 23080 12557 23120
rect 12748 23080 12788 23120
rect 12871 23080 12911 23120
rect 12988 23080 13028 23120
rect 13603 23080 13643 23120
rect 16726 23080 16766 23120
rect 17356 23080 17396 23120
rect 17635 23071 17675 23111
rect 17788 23080 17828 23120
rect 18307 23080 18347 23120
rect 18412 23080 18452 23120
rect 19036 23080 19076 23120
rect 19180 23080 19220 23120
rect 19843 23080 19883 23120
rect 19948 23080 19988 23120
rect 20572 23080 20612 23120
rect 20716 23080 20756 23120
rect 21292 23080 21332 23120
rect 21529 23080 21569 23120
rect 21671 23080 21711 23120
rect 21868 23080 21908 23120
rect 22252 23080 22292 23120
rect 22924 23080 22964 23120
rect 23500 23080 23540 23120
rect 23683 23080 23723 23120
rect 24172 23080 24212 23120
rect 24460 23080 24500 23120
rect 24643 23080 24683 23120
rect 25219 23080 25259 23120
rect 25507 23080 25547 23120
rect 25804 23080 25844 23120
rect 25996 23080 26036 23120
rect 26286 23080 26326 23120
rect 26380 23071 26420 23111
rect 26659 23080 26699 23120
rect 26836 23080 26876 23120
rect 27148 23080 27188 23120
rect 27340 23080 27380 23120
rect 27928 23080 27968 23120
rect 28108 23080 28148 23120
rect 28780 23080 28820 23120
rect 28972 23080 29012 23120
rect 29347 23080 29387 23120
rect 5283 22996 5323 23036
rect 7468 22996 7508 23036
rect 10348 22996 10388 23036
rect 11596 22996 11636 23036
rect 13228 22996 13268 23036
rect 21196 22996 21236 23036
rect 21411 22996 21451 23036
rect 24316 22996 24356 23036
rect 25036 22996 25076 23036
rect 25612 22996 25652 23036
rect 2092 22912 2132 22952
rect 7852 22912 7892 22952
rect 10732 22912 10772 22952
rect 11980 22912 12020 22952
rect 13036 22912 13076 22952
rect 18595 22912 18635 22952
rect 24643 22912 24683 22952
rect 2956 22828 2996 22868
rect 3772 22828 3812 22868
rect 8188 22828 8228 22868
rect 16963 22828 17003 22868
rect 19075 22828 19115 22868
rect 20131 22828 20171 22868
rect 21772 22828 21812 22868
rect 25804 22828 25844 22868
rect 26275 22828 26315 22868
rect 27244 22828 27284 22868
rect 30892 22828 30932 22868
rect 3112 22660 3480 22700
rect 10886 22660 11254 22700
rect 18660 22660 19028 22700
rect 26434 22660 26802 22700
rect 844 22492 884 22532
rect 14851 22492 14891 22532
rect 19372 22492 19412 22532
rect 24652 22492 24692 22532
rect 25603 22492 25643 22532
rect 4012 22408 4052 22448
rect 6508 22408 6548 22448
rect 11356 22408 11396 22448
rect 12940 22408 12980 22448
rect 24988 22399 25028 22439
rect 25219 22408 25259 22448
rect 27052 22408 27092 22448
rect 28483 22408 28523 22448
rect 7516 22324 7556 22364
rect 8515 22324 8555 22364
rect 22930 22324 22970 22364
rect 30691 22324 30731 22364
rect 30892 22324 30932 22364
rect 2755 22240 2795 22280
rect 3619 22240 3659 22280
rect 4291 22240 4331 22280
rect 4396 22240 4436 22280
rect 4972 22240 5012 22280
rect 5836 22240 5876 22280
rect 6028 22240 6068 22280
rect 7660 22240 7700 22280
rect 8375 22240 8415 22280
rect 8620 22240 8660 22280
rect 10156 22240 10196 22280
rect 10444 22240 10484 22280
rect 10813 22240 10853 22280
rect 10924 22240 10964 22280
rect 11500 22240 11540 22280
rect 12172 22240 12212 22280
rect 12316 22240 12356 22280
rect 12760 22240 12800 22280
rect 12926 22240 12966 22280
rect 13036 22240 13076 22280
rect 13238 22240 13278 22280
rect 15244 22240 15284 22280
rect 16099 22240 16139 22280
rect 18700 22240 18740 22280
rect 19075 22240 19115 22280
rect 19180 22240 19220 22280
rect 21100 22240 21140 22280
rect 21292 22240 21332 22280
rect 21431 22240 21471 22280
rect 21571 22240 21611 22280
rect 21676 22240 21716 22280
rect 22147 22240 22187 22280
rect 22252 22240 22292 22280
rect 23020 22240 23060 22280
rect 23500 22240 23540 22280
rect 23692 22240 23732 22280
rect 24460 22240 24500 22280
rect 24763 22240 24803 22280
rect 25027 22240 25067 22280
rect 25891 22273 25931 22313
rect 25996 22240 26036 22280
rect 26563 22240 26603 22280
rect 26755 22240 26795 22280
rect 27187 22240 27227 22280
rect 27383 22240 27423 22280
rect 27505 22240 27545 22280
rect 27628 22240 27668 22280
rect 28195 22240 28235 22280
rect 28300 22240 28340 22280
rect 29452 22240 29492 22280
rect 30412 22240 30452 22280
rect 30551 22240 30591 22280
rect 30796 22240 30836 22280
rect 31084 22240 31124 22280
rect 31276 22240 31316 22280
rect 3139 22156 3179 22196
rect 4492 22156 4532 22196
rect 4602 22156 4642 22196
rect 5932 22156 5972 22196
rect 8707 22156 8747 22196
rect 12595 22156 12635 22196
rect 16492 22156 16532 22196
rect 19386 22156 19426 22196
rect 29731 22156 29771 22196
rect 31180 22156 31220 22196
rect 5644 22072 5684 22112
rect 9955 22072 9995 22112
rect 10627 22072 10667 22112
rect 18595 22072 18635 22112
rect 18892 22072 18932 22112
rect 21283 22072 21323 22112
rect 21763 22072 21803 22112
rect 22540 22072 22580 22112
rect 22723 22072 22763 22112
rect 23683 22072 23723 22112
rect 26107 22072 26147 22112
rect 27340 22072 27380 22112
rect 28780 22072 28820 22112
rect 4352 21904 4720 21944
rect 12126 21904 12494 21944
rect 19900 21904 20268 21944
rect 27674 21904 28042 21944
rect 7756 21736 7796 21776
rect 16579 21736 16619 21776
rect 17347 21736 17387 21776
rect 18172 21736 18212 21776
rect 20035 21736 20075 21776
rect 20275 21736 20315 21776
rect 21964 21736 22004 21776
rect 22780 21736 22820 21776
rect 24940 21736 24980 21776
rect 25507 21736 25547 21776
rect 28972 21736 29012 21776
rect 29923 21736 29963 21776
rect 30460 21736 30500 21776
rect 4195 21652 4235 21692
rect 5443 21652 5483 21692
rect 21388 21652 21428 21692
rect 29822 21652 29862 21692
rect 30028 21652 30068 21692
rect 30931 21652 30971 21692
rect 1708 21568 1748 21608
rect 4108 21568 4148 21608
rect 4291 21568 4331 21608
rect 4402 21536 4442 21576
rect 4579 21568 4619 21608
rect 4869 21568 4909 21608
rect 5068 21568 5108 21608
rect 5260 21568 5300 21608
rect 5827 21568 5867 21608
rect 9196 21568 9236 21608
rect 9772 21568 9812 21608
rect 11587 21559 11627 21599
rect 11884 21568 11924 21608
rect 13324 21568 13364 21608
rect 13612 21568 13652 21608
rect 16867 21568 16907 21608
rect 17635 21568 17675 21608
rect 18019 21559 18059 21599
rect 19372 21568 19412 21608
rect 19948 21568 19988 21608
rect 20332 21568 20372 21608
rect 20995 21568 21035 21608
rect 21868 21568 21908 21608
rect 22051 21568 22091 21608
rect 22924 21568 22964 21608
rect 24652 21568 24692 21608
rect 24780 21565 24820 21605
rect 25612 21568 25652 21608
rect 25996 21568 26036 21608
rect 26188 21568 26228 21608
rect 26385 21568 26425 21608
rect 26515 21568 26555 21608
rect 26620 21568 26660 21608
rect 26719 21559 26759 21599
rect 27148 21568 27188 21608
rect 27331 21568 27371 21608
rect 27523 21568 27563 21608
rect 27820 21568 27860 21608
rect 28108 21568 28148 21608
rect 28299 21568 28339 21608
rect 28483 21568 28523 21608
rect 28588 21568 28628 21608
rect 29644 21568 29684 21608
rect 30124 21559 30164 21599
rect 30307 21559 30347 21599
rect 31096 21568 31136 21608
rect 9682 21484 9722 21524
rect 11779 21484 11819 21524
rect 12364 21484 12404 21524
rect 16060 21484 16100 21524
rect 16300 21484 16340 21524
rect 16483 21484 16523 21524
rect 17059 21484 17099 21524
rect 17251 21484 17291 21524
rect 17827 21484 17867 21524
rect 25132 21484 25172 21524
rect 2572 21400 2612 21440
rect 4876 21400 4916 21440
rect 14476 21400 14516 21440
rect 16579 21400 16619 21440
rect 19756 21400 19796 21440
rect 20524 21400 20564 21440
rect 22444 21400 22484 21440
rect 25372 21400 25412 21440
rect 27820 21400 27860 21440
rect 2380 21316 2420 21356
rect 5068 21316 5108 21356
rect 7372 21316 7412 21356
rect 7756 21316 7796 21356
rect 8803 21316 8843 21356
rect 9667 21316 9707 21356
rect 12124 21316 12164 21356
rect 12988 21316 13028 21356
rect 19180 21316 19220 21356
rect 21196 21316 21236 21356
rect 25804 21316 25844 21356
rect 25996 21316 26036 21356
rect 26668 21316 26708 21356
rect 27331 21316 27371 21356
rect 28588 21316 28628 21356
rect 3112 21148 3480 21188
rect 10886 21148 11254 21188
rect 18660 21148 19028 21188
rect 26434 21148 26802 21188
rect 652 20980 692 21020
rect 6220 20980 6260 21020
rect 15724 20980 15764 21020
rect 23692 20980 23732 21020
rect 25900 20980 25940 21020
rect 26860 20980 26900 21020
rect 28204 20980 28244 21020
rect 31276 20980 31316 21020
rect 3772 20896 3812 20936
rect 9244 20896 9284 20936
rect 11683 20896 11723 20936
rect 13228 20896 13268 20936
rect 25036 20896 25076 20936
rect 26668 20896 26708 20936
rect 4483 20812 4523 20852
rect 5443 20812 5483 20852
rect 8131 20812 8171 20852
rect 9004 20812 9044 20852
rect 10348 20812 10388 20852
rect 10819 20812 10859 20852
rect 11395 20812 11435 20852
rect 11587 20812 11627 20852
rect 12163 20812 12203 20852
rect 13420 20812 13460 20852
rect 15340 20812 15380 20852
rect 16300 20812 16340 20852
rect 17260 20812 17300 20852
rect 17836 20812 17876 20852
rect 19315 20812 19355 20852
rect 20643 20812 20683 20852
rect 20995 20812 21035 20852
rect 25612 20812 25652 20852
rect 25747 20803 25787 20843
rect 27427 20812 27467 20852
rect 28972 20812 29012 20852
rect 2563 20728 2603 20768
rect 3148 20728 3188 20768
rect 3532 20728 3572 20768
rect 4684 20728 4724 20768
rect 5303 20728 5343 20768
rect 5548 20728 5588 20768
rect 6892 20728 6932 20768
rect 8011 20728 8051 20768
rect 8236 20728 8276 20768
rect 10444 20728 10484 20768
rect 10563 20728 10603 20768
rect 10681 20728 10721 20768
rect 11203 20728 11243 20768
rect 11971 20728 12011 20768
rect 12556 20728 12596 20768
rect 12835 20728 12875 20768
rect 13795 20728 13835 20768
rect 15959 20728 15999 20768
rect 16099 20728 16139 20768
rect 16204 20728 16244 20768
rect 17443 20728 17483 20768
rect 17731 20728 17771 20768
rect 17971 20728 18011 20768
rect 19510 20728 19550 20768
rect 19660 20728 19700 20768
rect 19852 20728 19892 20768
rect 20524 20728 20564 20768
rect 20741 20728 20781 20768
rect 20875 20728 20915 20768
rect 21100 20728 21140 20768
rect 21763 20728 21803 20768
rect 23884 20728 23924 20768
rect 24556 20728 24596 20768
rect 24835 20728 24875 20768
rect 25516 20728 25556 20768
rect 25855 20728 25895 20768
rect 26092 20728 26132 20768
rect 26254 20728 26294 20768
rect 26372 20761 26412 20801
rect 26474 20728 26514 20768
rect 26903 20728 26943 20768
rect 27043 20719 27083 20759
rect 27148 20728 27188 20768
rect 27287 20728 27327 20768
rect 27532 20728 27572 20768
rect 27820 20728 27860 20768
rect 28021 20728 28061 20768
rect 28204 20728 28244 20768
rect 28492 20728 28532 20768
rect 29347 20728 29387 20768
rect 2947 20644 2987 20684
rect 4291 20644 4331 20684
rect 9244 20644 9284 20684
rect 12940 20644 12980 20684
rect 19756 20644 19796 20684
rect 20428 20644 20468 20684
rect 21187 20644 21227 20684
rect 21379 20644 21419 20684
rect 5635 20560 5675 20600
rect 8323 20560 8363 20600
rect 10915 20560 10955 20600
rect 18172 20560 18212 20600
rect 27619 20560 27659 20600
rect 27820 20560 27860 20600
rect 4352 20392 4720 20432
rect 12126 20392 12494 20432
rect 19900 20392 20268 20432
rect 27674 20392 28042 20432
rect 12739 20224 12779 20264
rect 13411 20224 13451 20264
rect 15715 20224 15755 20264
rect 16780 20224 16820 20264
rect 17539 20224 17579 20264
rect 17740 20224 17780 20264
rect 20380 20224 20420 20264
rect 25027 20224 25067 20264
rect 26860 20224 26900 20264
rect 27139 20224 27179 20264
rect 2668 20140 2708 20180
rect 6700 20140 6740 20180
rect 8707 20140 8747 20180
rect 14371 20140 14411 20180
rect 16492 20140 16532 20180
rect 29635 20140 29675 20180
rect 1804 20056 1844 20096
rect 2041 20056 2081 20096
rect 2284 20056 2324 20096
rect 2563 20056 2603 20096
rect 3379 20056 3419 20096
rect 3574 20056 3614 20096
rect 3820 20056 3860 20096
rect 4057 20056 4097 20096
rect 4300 20056 4340 20096
rect 4492 20056 4532 20096
rect 5155 20056 5195 20096
rect 5923 20056 5963 20096
rect 6494 20056 6534 20096
rect 6796 20047 6836 20087
rect 7084 20056 7124 20096
rect 7276 20056 7316 20096
rect 7747 20056 7787 20096
rect 8995 20056 9035 20096
rect 9379 20047 9419 20087
rect 10444 20056 10484 20096
rect 10636 20056 10676 20096
rect 11011 20056 11051 20096
rect 11299 20056 11339 20096
rect 13219 20056 13259 20096
rect 13795 20056 13835 20096
rect 15052 20056 15092 20096
rect 15820 20056 15860 20096
rect 1708 19972 1748 20012
rect 1939 19963 1979 20003
rect 3724 19972 3764 20012
rect 3955 19963 3995 20003
rect 4588 19972 4628 20012
rect 4972 19972 5012 20012
rect 5548 19972 5588 20012
rect 5740 19972 5780 20012
rect 6316 19972 6356 20012
rect 7564 19972 7604 20012
rect 8140 19972 8180 20012
rect 8611 19972 8651 20012
rect 9187 19972 9227 20012
rect 9532 19972 9572 20012
rect 10828 19972 10868 20012
rect 11404 19972 11444 20012
rect 13036 19972 13076 20012
rect 15571 20014 15611 20054
rect 16396 20056 16436 20096
rect 16579 20056 16619 20096
rect 16875 20056 16915 20096
rect 17107 20056 17147 20096
rect 17212 20056 17252 20096
rect 17452 20056 17492 20096
rect 17836 20056 17876 20096
rect 17955 20056 17995 20096
rect 18073 20056 18113 20096
rect 18499 20047 18539 20087
rect 19276 20056 19316 20096
rect 19468 20056 19508 20096
rect 19703 20056 19743 20096
rect 19948 20056 19988 20096
rect 20236 20056 20276 20096
rect 20707 20056 20747 20096
rect 20995 20056 21035 20096
rect 21283 20047 21323 20087
rect 24460 20056 24500 20096
rect 24643 20056 24683 20096
rect 24748 20056 24788 20096
rect 25027 20056 25067 20096
rect 25315 20056 25355 20096
rect 25507 20056 25547 20096
rect 25699 20056 25739 20096
rect 26572 20056 26612 20096
rect 27052 20056 27092 20096
rect 27307 20056 27347 20096
rect 27532 20056 27572 20096
rect 28195 20056 28235 20096
rect 28300 20056 28340 20096
rect 29452 20056 29492 20096
rect 30316 20056 30356 20096
rect 30499 20047 30539 20087
rect 30988 20056 31028 20096
rect 31180 20056 31220 20096
rect 13708 19972 13748 20012
rect 15379 19972 15419 20012
rect 16995 19972 17035 20012
rect 17347 19972 17387 20012
rect 18652 19972 18692 20012
rect 19843 19972 19883 20012
rect 20044 19972 20084 20012
rect 20524 19972 20564 20012
rect 21100 19972 21140 20012
rect 21436 19972 21476 20012
rect 26428 19972 26468 20012
rect 27427 19972 27467 20012
rect 27628 19972 27668 20012
rect 30652 19972 30692 20012
rect 2956 19888 2996 19928
rect 5452 19888 5492 19928
rect 6220 19888 6260 19928
rect 7075 19888 7115 19928
rect 8044 19888 8084 19928
rect 16012 19888 16052 19928
rect 21004 19888 21044 19928
rect 26284 19888 26324 19928
rect 28483 19888 28523 19928
rect 6499 19804 6539 19844
rect 10444 19804 10484 19844
rect 19276 19804 19316 19844
rect 24748 19804 24788 19844
rect 28780 19804 28820 19844
rect 30988 19804 31028 19844
rect 3112 19636 3480 19676
rect 10886 19636 11254 19676
rect 18660 19636 19028 19676
rect 26434 19636 26802 19676
rect 4156 19468 4196 19508
rect 16195 19468 16235 19508
rect 16675 19468 16715 19508
rect 17635 19468 17675 19508
rect 19468 19468 19508 19508
rect 26179 19468 26219 19508
rect 28972 19468 29012 19508
rect 8140 19384 8180 19424
rect 11980 19384 12020 19424
rect 15052 19384 15092 19424
rect 21292 19384 21332 19424
rect 23011 19384 23051 19424
rect 23395 19384 23435 19424
rect 24556 19384 24596 19424
rect 1132 19300 1172 19340
rect 1708 19300 1748 19340
rect 3171 19300 3211 19340
rect 4396 19300 4436 19340
rect 5836 19300 5876 19340
rect 1315 19216 1355 19256
rect 1894 19249 1934 19289
rect 2199 19216 2239 19256
rect 2462 19216 2502 19256
rect 2764 19216 2804 19256
rect 3052 19216 3092 19256
rect 3269 19216 3309 19256
rect 3436 19216 3476 19256
rect 3619 19216 3659 19256
rect 5515 19216 5555 19256
rect 5635 19216 5675 19256
rect 5740 19216 5780 19256
rect 6124 19216 6164 19256
rect 6308 19216 6348 19256
rect 6667 19216 6707 19256
rect 6787 19216 6827 19256
rect 6892 19216 6932 19256
rect 7132 19258 7172 19298
rect 7253 19300 7293 19340
rect 7468 19300 7508 19340
rect 7660 19300 7700 19340
rect 8236 19300 8276 19340
rect 8931 19300 8971 19340
rect 9859 19300 9899 19340
rect 10531 19300 10571 19340
rect 10924 19300 10964 19340
rect 11155 19291 11195 19331
rect 13420 19300 13460 19340
rect 19939 19300 19979 19340
rect 20419 19300 20459 19340
rect 20620 19300 20660 19340
rect 20812 19300 20852 19340
rect 21388 19300 21428 19340
rect 23299 19300 23339 19340
rect 23548 19300 23588 19340
rect 25036 19300 25076 19340
rect 31267 19300 31307 19340
rect 7372 19216 7412 19256
rect 7843 19216 7883 19256
rect 8812 19216 8852 19256
rect 9049 19216 9089 19256
rect 9280 19216 9320 19256
rect 9719 19216 9759 19256
rect 9964 19216 10004 19256
rect 10391 19216 10431 19256
rect 10636 19216 10676 19256
rect 11020 19216 11060 19256
rect 11257 19216 11297 19256
rect 11500 19216 11540 19256
rect 11619 19216 11659 19256
rect 11737 19216 11777 19256
rect 11884 19216 11924 19256
rect 12076 19216 12116 19256
rect 12268 19216 12308 19256
rect 12460 19216 12500 19256
rect 13132 19216 13172 19256
rect 13324 19216 13364 19256
rect 13804 19216 13844 19256
rect 14419 19216 14459 19256
rect 14614 19216 14654 19256
rect 14755 19207 14795 19247
rect 15052 19216 15092 19256
rect 15436 19216 15476 19256
rect 16012 19216 16052 19256
rect 16195 19216 16235 19256
rect 16972 19216 17012 19256
rect 17260 19216 17300 19256
rect 17379 19216 17419 19256
rect 17497 19216 17537 19256
rect 17938 19216 17978 19256
rect 19171 19216 19211 19256
rect 19479 19216 19519 19256
rect 19799 19216 19839 19256
rect 20044 19216 20084 19256
rect 20279 19216 20319 19256
rect 20524 19216 20564 19256
rect 20995 19216 21035 19256
rect 21523 19216 21563 19256
rect 22723 19216 22763 19256
rect 22828 19216 22868 19256
rect 23690 19216 23730 19256
rect 24163 19216 24203 19256
rect 24272 19249 24312 19289
rect 25219 19216 25259 19256
rect 25891 19216 25931 19256
rect 25996 19216 26036 19256
rect 26476 19216 26516 19256
rect 28108 19216 28148 19256
rect 28291 19216 28331 19256
rect 30883 19216 30923 19256
rect 1612 19132 1652 19172
rect 2563 19132 2603 19172
rect 6019 19132 6059 19172
rect 8716 19132 8756 19172
rect 11404 19132 11444 19172
rect 13603 19132 13643 19172
rect 16108 19132 16148 19172
rect 16670 19132 16710 19172
rect 17630 19132 17670 19172
rect 27148 19132 27188 19172
rect 28599 19132 28639 19172
rect 1987 19048 2027 19088
rect 2092 19048 2132 19088
rect 2668 19048 2708 19088
rect 2956 19048 2996 19088
rect 3532 19048 3572 19088
rect 6979 19048 7019 19088
rect 9436 19048 9476 19088
rect 10051 19048 10091 19088
rect 10723 19048 10763 19088
rect 12364 19048 12404 19088
rect 13891 19048 13931 19088
rect 15331 19048 15371 19088
rect 15619 19048 15659 19088
rect 16876 19048 16916 19088
rect 17164 19048 17204 19088
rect 17836 19048 17876 19088
rect 19267 19048 19307 19088
rect 20131 19048 20171 19088
rect 21724 19048 21764 19088
rect 23116 19048 23156 19088
rect 23395 19048 23435 19088
rect 24067 19039 24107 19079
rect 24739 19048 24779 19088
rect 27436 19048 27476 19088
rect 28387 19048 28427 19088
rect 28492 19048 28532 19088
rect 28972 19048 29012 19088
rect 4352 18880 4720 18920
rect 12126 18880 12494 18920
rect 19900 18880 20268 18920
rect 27674 18880 28042 18920
rect 1411 18712 1451 18752
rect 1891 18712 1931 18752
rect 3052 18712 3092 18752
rect 4204 18712 4244 18752
rect 5251 18712 5291 18752
rect 6412 18712 6452 18752
rect 7276 18712 7316 18752
rect 8899 18712 8939 18752
rect 9244 18712 9284 18752
rect 11020 18712 11060 18752
rect 11308 18712 11348 18752
rect 13891 18712 13931 18752
rect 16684 18712 16724 18752
rect 17923 18712 17963 18752
rect 18403 18712 18443 18752
rect 19363 18712 19403 18752
rect 22924 18712 22964 18752
rect 27763 18712 27803 18752
rect 28972 18712 29012 18752
rect 2092 18628 2132 18668
rect 2558 18628 2598 18668
rect 2659 18628 2699 18668
rect 3998 18628 4038 18668
rect 7660 18628 7700 18668
rect 8179 18628 8219 18668
rect 8798 18628 8838 18668
rect 9004 18628 9044 18668
rect 13603 18628 13643 18668
rect 16972 18628 17012 18668
rect 18508 18628 18548 18668
rect 19756 18628 19796 18668
rect 20323 18628 20363 18668
rect 21388 18628 21428 18668
rect 24451 18628 24491 18668
rect 27331 18628 27371 18668
rect 1079 18544 1119 18584
rect 1324 18544 1364 18584
rect 1564 18502 1604 18542
rect 1804 18544 1844 18584
rect 2188 18544 2228 18584
rect 2425 18544 2465 18584
rect 2764 18544 2804 18584
rect 2860 18535 2900 18575
rect 3148 18544 3188 18584
rect 3267 18544 3307 18584
rect 1219 18460 1259 18500
rect 1699 18460 1739 18500
rect 2092 18460 2132 18500
rect 2307 18460 2347 18500
rect 3388 18502 3428 18542
rect 4300 18535 4340 18575
rect 4939 18544 4979 18584
rect 5164 18544 5204 18584
rect 4819 18502 4859 18542
rect 5548 18544 5588 18584
rect 5765 18544 5805 18584
rect 5921 18544 5961 18584
rect 6124 18544 6164 18584
rect 6220 18535 6260 18575
rect 6508 18544 6548 18584
rect 6745 18544 6785 18584
rect 7180 18544 7220 18584
rect 7371 18544 7411 18584
rect 7555 18544 7595 18584
rect 7863 18544 7903 18584
rect 8374 18544 8414 18584
rect 8524 18544 8564 18584
rect 9100 18535 9140 18575
rect 10732 18544 10772 18584
rect 10874 18544 10914 18584
rect 11212 18544 11252 18584
rect 11395 18544 11435 18584
rect 12694 18544 12734 18584
rect 13324 18544 13364 18584
rect 13804 18544 13844 18584
rect 14668 18544 14708 18584
rect 14860 18544 14900 18584
rect 16204 18544 16244 18584
rect 16373 18544 16413 18584
rect 16492 18544 16532 18584
rect 16867 18544 16907 18584
rect 17175 18544 17215 18584
rect 17299 18544 17339 18584
rect 17827 18544 17867 18584
rect 18135 18544 18175 18584
rect 18302 18544 18342 18584
rect 18604 18535 18644 18575
rect 19031 18544 19071 18584
rect 19274 18544 19314 18584
rect 19555 18544 19595 18584
rect 19660 18544 19700 18584
rect 19863 18544 19903 18584
rect 19996 18544 20036 18584
rect 20131 18544 20171 18584
rect 20236 18544 20276 18584
rect 21091 18544 21131 18584
rect 22915 18544 22955 18584
rect 23020 18544 23060 18584
rect 24364 18544 24404 18584
rect 24556 18544 24596 18584
rect 26947 18544 26987 18584
rect 27955 18544 27995 18584
rect 28075 18544 28115 18584
rect 28531 18544 28571 18584
rect 28780 18544 28820 18584
rect 3820 18460 3860 18500
rect 4627 18460 4667 18500
rect 5059 18460 5099 18500
rect 5452 18460 5492 18500
rect 5683 18451 5723 18491
rect 6627 18460 6667 18500
rect 9484 18460 9524 18500
rect 12499 18460 12539 18500
rect 17500 18460 17540 18500
rect 19171 18460 19211 18500
rect 20908 18460 20948 18500
rect 21484 18460 21524 18500
rect 21868 18460 21908 18500
rect 28204 18460 28244 18500
rect 28368 18502 28408 18542
rect 30883 18544 30923 18584
rect 28636 18460 28676 18500
rect 31267 18460 31307 18500
rect 23212 18376 23252 18416
rect 25420 18376 25460 18416
rect 28300 18376 28340 18416
rect 3580 18292 3620 18332
rect 4003 18292 4043 18332
rect 5923 18292 5963 18332
rect 7852 18292 7892 18332
rect 13132 18292 13172 18332
rect 14764 18292 14804 18332
rect 17164 18292 17204 18332
rect 18124 18292 18164 18332
rect 21628 18292 21668 18332
rect 25036 18292 25076 18332
rect 3112 18124 3480 18164
rect 10886 18124 11254 18164
rect 18660 18124 19028 18164
rect 26434 18124 26802 18164
rect 1411 17956 1451 17996
rect 2179 17956 2219 17996
rect 5740 17956 5780 17996
rect 7555 17956 7595 17996
rect 8860 17956 8900 17996
rect 16300 17956 16340 17996
rect 18220 17956 18260 17996
rect 19756 17956 19796 17996
rect 22636 17956 22676 17996
rect 27724 17956 27764 17996
rect 30700 17956 30740 17996
rect 29836 17872 29876 17912
rect 30892 17872 30932 17912
rect 2995 17788 3035 17828
rect 4108 17788 4148 17828
rect 4531 17779 4571 17819
rect 9772 17788 9812 17828
rect 10828 17788 10868 17828
rect 11731 17788 11771 17828
rect 1708 17704 1748 17744
rect 2177 17704 2217 17744
rect 2476 17704 2516 17744
rect 3190 17704 3230 17744
rect 3628 17704 3668 17744
rect 3772 17704 3812 17744
rect 3907 17704 3947 17744
rect 4012 17704 4052 17744
rect 4396 17704 4436 17744
rect 4633 17704 4673 17744
rect 4876 17704 4916 17744
rect 4995 17704 5035 17744
rect 5113 17704 5153 17744
rect 5740 17704 5780 17744
rect 5932 17704 5972 17744
rect 6604 17704 6644 17744
rect 6795 17704 6835 17744
rect 6988 17704 7028 17744
rect 7171 17704 7211 17744
rect 7372 17704 7412 17744
rect 7555 17704 7595 17744
rect 8083 17704 8123 17744
rect 8278 17704 8318 17744
rect 9004 17704 9044 17744
rect 9292 17704 9332 17744
rect 9411 17704 9451 17744
rect 9529 17704 9569 17744
rect 9676 17704 9716 17744
rect 9868 17704 9908 17744
rect 10348 17704 10388 17744
rect 10540 17704 10580 17744
rect 10732 17704 10772 17744
rect 10924 17704 10964 17744
rect 11063 17704 11103 17744
rect 11203 17704 11243 17744
rect 11308 17704 11348 17744
rect 11926 17704 11966 17744
rect 13123 17704 13163 17744
rect 13420 17704 13460 17744
rect 14806 17704 14846 17744
rect 15148 17704 15188 17744
rect 15436 17704 15476 17744
rect 15628 17704 15668 17744
rect 16003 17704 16043 17744
rect 16492 17704 16532 17744
rect 16684 17704 16724 17744
rect 17548 17704 17588 17744
rect 17717 17704 17757 17744
rect 17923 17704 17963 17744
rect 18231 17704 18271 17744
rect 19459 17704 19499 17744
rect 19770 17704 19810 17744
rect 22636 17704 22676 17744
rect 22939 17704 22979 17744
rect 23107 17695 23147 17735
rect 23404 17704 23444 17744
rect 24172 17704 24212 17744
rect 24460 17704 24500 17744
rect 24844 17704 24884 17744
rect 24988 17704 25028 17744
rect 25900 17704 25940 17744
rect 26092 17704 26132 17744
rect 27628 17704 27668 17744
rect 27820 17704 27860 17744
rect 28396 17704 28436 17744
rect 28579 17704 28619 17744
rect 29260 17704 29300 17744
rect 30028 17704 30068 17744
rect 1409 17620 1449 17660
rect 3329 17620 3369 17660
rect 4300 17620 4340 17660
rect 6700 17620 6740 17660
rect 9196 17620 9236 17660
rect 11395 17620 11435 17660
rect 12940 17620 12980 17660
rect 15532 17620 15572 17660
rect 16314 17620 16354 17660
rect 16588 17620 16628 17660
rect 23212 17620 23252 17660
rect 24643 17620 24683 17660
rect 28492 17620 28532 17660
rect 1612 17536 1652 17576
rect 2380 17536 2420 17576
rect 3427 17536 3467 17576
rect 3532 17536 3572 17576
rect 4780 17536 4820 17576
rect 7084 17536 7124 17576
rect 10444 17536 10484 17576
rect 14611 17536 14651 17576
rect 14956 17536 14996 17576
rect 15235 17536 15275 17576
rect 16099 17536 16139 17576
rect 17644 17536 17684 17576
rect 18019 17536 18059 17576
rect 19555 17536 19595 17576
rect 23971 17536 24011 17576
rect 24940 17536 24980 17576
rect 25996 17536 26036 17576
rect 29155 17536 29195 17576
rect 29452 17536 29492 17576
rect 4352 17368 4720 17408
rect 12126 17368 12494 17408
rect 19900 17368 20268 17408
rect 27674 17368 28042 17408
rect 5164 17200 5204 17240
rect 6172 17200 6212 17240
rect 9100 17200 9140 17240
rect 11107 17200 11147 17240
rect 11587 17200 11627 17240
rect 13420 17200 13460 17240
rect 16867 17200 16907 17240
rect 18979 17200 19019 17240
rect 25747 17200 25787 17240
rect 29356 17200 29396 17240
rect 641 17116 681 17156
rect 1900 17116 1940 17156
rect 4867 17116 4907 17156
rect 6595 17116 6635 17156
rect 8332 17116 8372 17156
rect 9187 17107 9227 17147
rect 10819 17116 10859 17156
rect 11006 17116 11046 17156
rect 11212 17116 11252 17156
rect 11692 17116 11732 17156
rect 18115 17107 18155 17147
rect 20419 17116 20459 17156
rect 24268 17116 24308 17156
rect 24474 17116 24514 17156
rect 844 17032 884 17072
rect 940 17023 980 17063
rect 1315 17032 1355 17072
rect 1996 17032 2036 17072
rect 2233 17032 2273 17072
rect 2380 17032 2420 17072
rect 2553 17032 2593 17072
rect 2764 17032 2804 17072
rect 2947 17032 2987 17072
rect 4195 17032 4235 17072
rect 4535 17032 4575 17072
rect 4780 17032 4820 17072
rect 5063 17032 5103 17072
rect 5251 17032 5291 17072
rect 6028 17032 6068 17072
rect 6988 17032 7028 17072
rect 8140 17032 8180 17072
rect 8443 17032 8483 17072
rect 8899 17032 8939 17072
rect 9004 17023 9044 17063
rect 9279 17032 9319 17072
rect 9460 17032 9500 17072
rect 10507 17032 10547 17072
rect 10732 17032 10772 17072
rect 11298 17007 11338 17047
rect 11491 17032 11531 17072
rect 11799 17032 11839 17072
rect 12460 17032 12500 17072
rect 12787 17032 12827 17072
rect 13027 17032 13067 17072
rect 13564 17032 13604 17072
rect 13900 17032 13940 17072
rect 14872 17032 14912 17072
rect 15235 17023 15275 17063
rect 16003 17032 16043 17072
rect 16300 17032 16340 17072
rect 16780 17032 16820 17072
rect 17356 17032 17396 17072
rect 17659 17032 17699 17072
rect 17827 17032 17867 17072
rect 17932 17023 17972 17063
rect 18206 17032 18246 17072
rect 18387 17032 18427 17072
rect 18628 17032 18668 17072
rect 18787 17032 18827 17072
rect 18904 17032 18944 17072
rect 19075 17032 19115 17072
rect 19197 17032 19237 17072
rect 19852 17032 19892 17072
rect 20087 17032 20127 17072
rect 20332 17032 20372 17072
rect 20620 17032 20660 17072
rect 20803 17032 20843 17072
rect 21388 17032 21428 17072
rect 21517 17032 21557 17072
rect 21772 17032 21812 17072
rect 22540 17032 22580 17072
rect 22819 17023 22859 17063
rect 23692 17032 23732 17072
rect 23875 17032 23915 17072
rect 23980 17032 24020 17072
rect 24174 17032 24214 17072
rect 25324 17032 25364 17072
rect 25942 17032 25982 17072
rect 28579 17032 28619 17072
rect 30028 17032 30068 17072
rect 1132 16948 1172 16988
rect 1708 16948 1748 16988
rect 2131 16939 2171 16979
rect 3811 16948 3851 16988
rect 4387 16948 4427 16988
rect 4675 16948 4715 16988
rect 10627 16948 10667 16988
rect 14707 16948 14747 16988
rect 15388 16948 15428 16988
rect 20227 16948 20267 16988
rect 22972 16948 23012 16988
rect 27043 16948 27083 16988
rect 28963 16948 29003 16988
rect 1612 16864 1652 16904
rect 3907 16864 3947 16904
rect 13123 16864 13163 16904
rect 16588 16864 16628 16904
rect 19459 16864 19499 16904
rect 20803 16864 20843 16904
rect 21100 16864 21140 16904
rect 30412 16864 30452 16904
rect 30604 16864 30644 16904
rect 643 16780 683 16820
rect 2380 16780 2420 16820
rect 2947 16780 2987 16820
rect 12652 16780 12692 16820
rect 13699 16780 13739 16820
rect 15820 16780 15860 16820
rect 17548 16780 17588 16820
rect 17827 16780 17867 16820
rect 22147 16780 22187 16820
rect 23980 16780 24020 16820
rect 24460 16780 24500 16820
rect 24931 16780 24971 16820
rect 26668 16780 26708 16820
rect 3112 16612 3480 16652
rect 10886 16612 11254 16652
rect 18660 16612 19028 16652
rect 26434 16612 26802 16652
rect 2659 16444 2699 16484
rect 4300 16444 4340 16484
rect 6691 16444 6731 16484
rect 7363 16444 7403 16484
rect 9964 16444 10004 16484
rect 12067 16444 12107 16484
rect 16099 16444 16139 16484
rect 16588 16444 16628 16484
rect 17827 16444 17867 16484
rect 24556 16444 24596 16484
rect 26092 16444 26132 16484
rect 28972 16444 29012 16484
rect 29356 16444 29396 16484
rect 9004 16360 9044 16400
rect 22828 16360 22868 16400
rect 28396 16360 28436 16400
rect 1420 16276 1460 16316
rect 1612 16276 1652 16316
rect 1843 16267 1883 16307
rect 6979 16276 7019 16316
rect 7180 16276 7220 16316
rect 1079 16192 1119 16232
rect 1219 16192 1259 16232
rect 1324 16192 1364 16232
rect 1708 16192 1748 16232
rect 1945 16192 1985 16232
rect 2188 16192 2228 16232
rect 2307 16192 2347 16232
rect 2425 16192 2465 16232
rect 2956 16192 2996 16232
rect 4003 16192 4043 16232
rect 4314 16192 4354 16232
rect 5587 16234 5627 16274
rect 10732 16276 10772 16316
rect 19315 16276 19355 16316
rect 21484 16276 21524 16316
rect 4481 16192 4521 16232
rect 4786 16192 4826 16232
rect 5395 16192 5435 16232
rect 5764 16192 5804 16232
rect 5937 16192 5977 16232
rect 6067 16192 6107 16232
rect 6179 16192 6219 16232
rect 6307 16192 6347 16232
rect 6508 16192 6548 16232
rect 6691 16192 6731 16232
rect 6839 16192 6879 16232
rect 7084 16192 7124 16232
rect 7355 16192 7395 16232
rect 7519 16192 7559 16232
rect 7647 16192 7687 16232
rect 7747 16192 7787 16232
rect 7924 16192 7964 16232
rect 8758 16192 8798 16232
rect 9187 16192 9227 16232
rect 9484 16192 9524 16232
rect 9667 16192 9707 16232
rect 10391 16192 10431 16232
rect 10531 16192 10571 16232
rect 10636 16192 10676 16232
rect 11926 16192 11966 16232
rect 12268 16192 12308 16232
rect 12364 16192 12404 16232
rect 13036 16192 13076 16232
rect 13155 16192 13195 16232
rect 13273 16192 13313 16232
rect 13750 16192 13790 16232
rect 14860 16192 14900 16232
rect 15244 16192 15284 16232
rect 15571 16192 15611 16232
rect 16097 16192 16137 16232
rect 16396 16192 16436 16232
rect 16588 16192 16628 16232
rect 16780 16192 16820 16232
rect 19507 16234 19547 16274
rect 23587 16276 23627 16316
rect 17644 16192 17684 16232
rect 17827 16192 17867 16232
rect 19660 16192 19700 16232
rect 19852 16192 19892 16232
rect 20515 16192 20555 16232
rect 21004 16192 21044 16232
rect 21580 16192 21620 16232
rect 21964 16192 22004 16232
rect 22082 16192 22122 16232
rect 22871 16192 22911 16232
rect 23011 16183 23051 16223
rect 23116 16192 23156 16232
rect 23447 16192 23487 16232
rect 23692 16192 23732 16232
rect 23932 16192 23972 16232
rect 24067 16192 24107 16232
rect 24172 16192 24212 16232
rect 24460 16192 24500 16232
rect 25795 16192 25835 16232
rect 26428 16192 26468 16232
rect 26620 16192 26660 16232
rect 26764 16234 26804 16274
rect 27820 16276 27860 16316
rect 31267 16276 31307 16316
rect 26956 16192 26996 16232
rect 27148 16192 27188 16232
rect 28012 16192 28052 16232
rect 28204 16192 28244 16232
rect 30883 16192 30923 16232
rect 2654 16108 2694 16148
rect 4579 16108 4619 16148
rect 9772 16108 9812 16148
rect 9975 16108 10015 16148
rect 12062 16108 12102 16148
rect 15436 16108 15476 16148
rect 19756 16108 19796 16148
rect 23779 16108 23819 16148
rect 26103 16108 26143 16148
rect 2092 16024 2132 16064
rect 2860 16024 2900 16064
rect 4099 16024 4139 16064
rect 4684 16024 4724 16064
rect 5827 16024 5867 16064
rect 8563 16024 8603 16064
rect 11731 16024 11771 16064
rect 12268 16024 12308 16064
rect 12940 16024 12980 16064
rect 13555 16024 13595 16064
rect 14668 16024 14708 16064
rect 16300 16024 16340 16064
rect 20332 16024 20372 16064
rect 24259 16024 24299 16064
rect 25891 16024 25931 16064
rect 26275 16024 26315 16064
rect 26860 16024 26900 16064
rect 28108 16024 28148 16064
rect 4352 15856 4720 15896
rect 12126 15856 12494 15896
rect 19900 15856 20268 15896
rect 27674 15856 28042 15896
rect 2956 15688 2996 15728
rect 4588 15688 4628 15728
rect 6316 15688 6356 15728
rect 8428 15688 8468 15728
rect 9283 15688 9323 15728
rect 11683 15688 11723 15728
rect 13420 15688 13460 15728
rect 15052 15688 15092 15728
rect 15619 15688 15659 15728
rect 16099 15688 16139 15728
rect 16771 15688 16811 15728
rect 17356 15688 17396 15728
rect 18139 15688 18179 15728
rect 18595 15688 18635 15728
rect 21100 15688 21140 15728
rect 23692 15688 23732 15728
rect 24700 15688 24740 15728
rect 24940 15688 24980 15728
rect 26860 15688 26900 15728
rect 27235 15688 27275 15728
rect 3379 15604 3419 15644
rect 8908 15604 8948 15644
rect 12748 15604 12788 15644
rect 14659 15604 14699 15644
rect 14846 15604 14886 15644
rect 16579 15595 16619 15635
rect 17153 15604 17193 15644
rect 27340 15604 27380 15644
rect 31267 15604 31307 15644
rect 1804 15520 1844 15560
rect 2092 15520 2132 15560
rect 2750 15520 2790 15560
rect 3052 15511 3092 15551
rect 3544 15520 3584 15560
rect 3820 15520 3860 15560
rect 4195 15520 4235 15560
rect 4302 15493 4342 15533
rect 5452 15520 5492 15560
rect 5709 15520 5749 15560
rect 6163 15520 6203 15560
rect 6412 15520 6452 15560
rect 3676 15436 3716 15476
rect 5596 15436 5636 15476
rect 5864 15478 5904 15518
rect 6531 15520 6571 15560
rect 6649 15520 6689 15560
rect 7324 15520 7364 15560
rect 7795 15520 7835 15560
rect 8140 15520 8180 15560
rect 6028 15436 6068 15476
rect 7468 15478 7508 15518
rect 8282 15488 8322 15528
rect 8812 15520 8852 15560
rect 9004 15520 9044 15560
rect 9263 15520 9303 15560
rect 9379 15520 9419 15560
rect 9523 15520 9563 15560
rect 9667 15520 9707 15560
rect 9772 15509 9812 15549
rect 10060 15520 10100 15560
rect 10252 15520 10292 15560
rect 11351 15520 11391 15560
rect 11596 15520 11636 15560
rect 12141 15520 12181 15560
rect 12303 15520 12343 15560
rect 12844 15520 12884 15560
rect 7660 15436 7700 15476
rect 11491 15436 11531 15476
rect 12595 15478 12635 15518
rect 13081 15520 13121 15560
rect 13219 15520 13259 15560
rect 13324 15520 13364 15560
rect 13527 15520 13567 15560
rect 14327 15520 14367 15560
rect 14572 15520 14612 15560
rect 15148 15511 15188 15551
rect 15287 15520 15327 15560
rect 15532 15520 15572 15560
rect 15767 15520 15807 15560
rect 16012 15520 16052 15560
rect 16291 15520 16331 15560
rect 16396 15511 16436 15551
rect 16670 15520 16710 15560
rect 16852 15520 16892 15560
rect 17452 15511 17492 15551
rect 17920 15511 17960 15551
rect 18019 15520 18059 15560
rect 18283 15520 18323 15560
rect 18508 15520 18548 15560
rect 19651 15520 19691 15560
rect 20899 15520 20939 15560
rect 23596 15520 23636 15560
rect 23788 15520 23828 15560
rect 24043 15520 24083 15560
rect 24268 15520 24308 15560
rect 24844 15520 24884 15560
rect 24988 15520 25028 15560
rect 25367 15520 25407 15560
rect 25507 15511 25547 15551
rect 25612 15520 25652 15560
rect 26044 15520 26084 15560
rect 26223 15520 26263 15560
rect 26501 15520 26541 15560
rect 26657 15520 26697 15560
rect 26956 15511 26996 15551
rect 27139 15520 27179 15560
rect 27447 15520 27487 15560
rect 28780 15520 28820 15560
rect 30883 15520 30923 15560
rect 12460 15436 12500 15476
rect 12979 15427 13019 15467
rect 14467 15436 14507 15476
rect 15427 15436 15467 15476
rect 15907 15436 15947 15476
rect 18403 15436 18443 15476
rect 24163 15436 24203 15476
rect 24364 15436 24404 15476
rect 26380 15436 26420 15476
rect 1804 15352 1844 15392
rect 5932 15352 5972 15392
rect 7564 15352 7604 15392
rect 10051 15352 10091 15392
rect 12364 15352 12404 15392
rect 26284 15352 26324 15392
rect 2755 15268 2795 15308
rect 14851 15268 14891 15308
rect 17155 15268 17195 15308
rect 17635 15268 17675 15308
rect 20044 15268 20084 15308
rect 21292 15268 21332 15308
rect 25324 15268 25364 15308
rect 26659 15268 26699 15308
rect 28108 15268 28148 15308
rect 28972 15268 29012 15308
rect 29356 15268 29396 15308
rect 3112 15100 3480 15140
rect 10886 15100 11254 15140
rect 18660 15100 19028 15140
rect 26434 15100 26802 15140
rect 4003 14932 4043 14972
rect 7171 14932 7211 14972
rect 7948 14932 7988 14972
rect 9859 14932 9899 14972
rect 11500 14932 11540 14972
rect 12988 14932 13028 14972
rect 18019 14932 18059 14972
rect 18499 14932 18539 14972
rect 24268 14932 24308 14972
rect 24940 14932 24980 14972
rect 28003 14932 28043 14972
rect 28387 14932 28427 14972
rect 4876 14848 4916 14888
rect 6691 14848 6731 14888
rect 6940 14839 6980 14879
rect 10348 14848 10388 14888
rect 20044 14848 20084 14888
rect 26668 14848 26708 14888
rect 27235 14848 27275 14888
rect 30700 14848 30740 14888
rect 31084 14848 31124 14888
rect 4515 14764 4555 14804
rect 10252 14764 10292 14804
rect 11059 14764 11099 14804
rect 14115 14764 14155 14804
rect 14787 14764 14827 14804
rect 16611 14764 16651 14804
rect 21484 14764 21524 14804
rect 24652 14764 24692 14804
rect 25324 14764 25364 14804
rect 25555 14755 25595 14795
rect 28402 14764 28442 14804
rect 1228 14680 1268 14720
rect 1372 14680 1412 14720
rect 2380 14680 2420 14720
rect 2755 14671 2795 14711
rect 3052 14680 3092 14720
rect 3715 14680 3755 14720
rect 3820 14680 3860 14720
rect 4405 14680 4445 14720
rect 4636 14680 4676 14720
rect 4775 14661 4815 14701
rect 4972 14680 5012 14720
rect 5764 14680 5804 14720
rect 5937 14680 5977 14720
rect 6067 14680 6107 14720
rect 6188 14691 6228 14731
rect 6307 14680 6347 14720
rect 6508 14680 6548 14720
rect 6691 14680 6731 14720
rect 6979 14680 7019 14720
rect 7388 14691 7428 14731
rect 7555 14680 7595 14720
rect 7672 14680 7712 14720
rect 7843 14680 7883 14720
rect 7965 14680 8005 14720
rect 8140 14680 8180 14720
rect 8332 14680 8372 14720
rect 9187 14680 9227 14720
rect 9484 14680 9524 14720
rect 9676 14680 9716 14720
rect 9859 14680 9899 14720
rect 10108 14680 10148 14720
rect 10423 14680 10463 14720
rect 10579 14680 10619 14720
rect 11224 14680 11264 14720
rect 11404 14680 11444 14720
rect 12844 14680 12884 14720
rect 13123 14680 13163 14720
rect 13241 14680 13281 14720
rect 13407 14680 13447 14720
rect 13507 14680 13547 14720
rect 13684 14680 13724 14720
rect 13996 14680 14036 14720
rect 14233 14680 14273 14720
rect 14668 14680 14708 14720
rect 14905 14680 14945 14720
rect 16216 14680 16256 14720
rect 16492 14680 16532 14720
rect 16709 14680 16749 14720
rect 16876 14680 16916 14720
rect 17068 14680 17108 14720
rect 17243 14680 17283 14720
rect 17369 14680 17409 14720
rect 17539 14671 17579 14711
rect 17643 14680 17683 14720
rect 17812 14680 17852 14720
rect 18322 14680 18362 14720
rect 18700 14680 18740 14720
rect 18802 14680 18842 14720
rect 19372 14680 19412 14720
rect 19627 14680 19667 14720
rect 19747 14680 19787 14720
rect 20995 14680 21035 14720
rect 21100 14680 21140 14720
rect 21580 14680 21620 14720
rect 22060 14680 22100 14720
rect 22548 14680 22588 14720
rect 23308 14680 23348 14720
rect 23980 14680 24020 14720
rect 24102 14680 24142 14720
rect 24212 14713 24252 14753
rect 24556 14680 24596 14720
rect 24777 14680 24817 14720
rect 24895 14680 24935 14720
rect 25420 14680 25460 14720
rect 25651 14680 25691 14720
rect 26711 14680 26751 14720
rect 26851 14671 26891 14711
rect 26956 14680 26996 14720
rect 27244 14680 27284 14720
rect 27436 14680 27476 14720
rect 27820 14680 27860 14720
rect 28003 14680 28043 14720
rect 28492 14680 28532 14720
rect 28972 14680 29012 14720
rect 30508 14680 30548 14720
rect 30700 14680 30740 14720
rect 30892 14680 30932 14720
rect 1027 14596 1067 14636
rect 2563 14596 2603 14636
rect 2860 14596 2900 14636
rect 4300 14596 4340 14636
rect 8236 14596 8276 14636
rect 9004 14596 9044 14636
rect 18017 14596 18057 14636
rect 18494 14596 18534 14636
rect 29644 14596 29684 14636
rect 1324 14512 1364 14552
rect 1708 14512 1748 14552
rect 2956 14512 2996 14552
rect 5827 14512 5867 14552
rect 13507 14512 13547 14552
rect 13900 14512 13940 14552
rect 14572 14512 14612 14552
rect 16051 14512 16091 14552
rect 16396 14512 16436 14552
rect 16972 14512 17012 14552
rect 17731 14512 17771 14552
rect 18220 14512 18260 14552
rect 22732 14512 22772 14552
rect 23452 14512 23492 14552
rect 29836 14512 29876 14552
rect 4352 14344 4720 14384
rect 12126 14344 12494 14384
rect 19900 14344 20268 14384
rect 27674 14344 28042 14384
rect 1795 14176 1835 14216
rect 1900 14176 1940 14216
rect 3715 14176 3755 14216
rect 4876 14176 4916 14216
rect 5635 14176 5675 14216
rect 9964 14176 10004 14216
rect 10636 14176 10676 14216
rect 14188 14176 14228 14216
rect 14755 14176 14795 14216
rect 15340 14176 15380 14216
rect 16483 14176 16523 14216
rect 19372 14176 19412 14216
rect 22243 14176 22283 14216
rect 24940 14176 24980 14216
rect 25612 14176 25652 14216
rect 26092 14176 26132 14216
rect 26956 14176 26996 14216
rect 27244 14176 27284 14216
rect 1123 14092 1163 14132
rect 2010 14092 2050 14132
rect 2659 14092 2699 14132
rect 14860 14092 14900 14132
rect 15447 14092 15487 14132
rect 16771 14083 16811 14123
rect 20140 14092 20180 14132
rect 21484 14092 21524 14132
rect 23884 14092 23924 14132
rect 24556 14092 24596 14132
rect 24663 14092 24703 14132
rect 1036 14008 1076 14048
rect 1208 14008 1248 14048
rect 1324 14008 1364 14048
rect 1699 14008 1739 14048
rect 2323 14008 2363 14048
rect 2518 14008 2558 14048
rect 3292 14008 3332 14048
rect 3530 14008 3570 14048
rect 3724 14008 3764 14048
rect 4972 14008 5012 14048
rect 5091 14008 5131 14048
rect 5209 14008 5249 14048
rect 5548 14008 5588 14048
rect 5932 14008 5972 14048
rect 6169 14008 6209 14048
rect 6316 14008 6356 14048
rect 6508 14008 6548 14048
rect 10060 14008 10100 14048
rect 10297 14008 10337 14048
rect 10732 14008 10772 14048
rect 10969 14008 11009 14048
rect 11203 14008 11243 14048
rect 12652 14008 12692 14048
rect 12844 14008 12884 14048
rect 14231 14008 14271 14048
rect 14371 13999 14411 14039
rect 14476 14008 14516 14048
rect 14657 14008 14697 14048
rect 14956 13999 14996 14039
rect 15139 14008 15179 14048
rect 15244 14008 15284 14048
rect 16483 14008 16523 14048
rect 16588 13999 16628 14039
rect 16867 14008 16907 14048
rect 17044 14008 17084 14048
rect 18892 14008 18932 14048
rect 19084 14008 19124 14048
rect 19276 14008 19316 14048
rect 19468 14008 19508 14048
rect 20249 14008 20289 14048
rect 20524 14008 20564 14048
rect 20812 14008 20852 14048
rect 20995 14008 21035 14048
rect 21148 14008 21188 14048
rect 21593 14008 21633 14048
rect 21868 14008 21908 14048
rect 22531 14008 22571 14048
rect 23277 14008 23317 14048
rect 23731 14008 23771 14048
rect 23980 14008 24020 14048
rect 5836 13924 5876 13964
rect 6051 13924 6091 13964
rect 10179 13924 10219 13964
rect 10851 13924 10891 13964
rect 11692 13924 11732 13964
rect 23432 13966 23472 14006
rect 24197 14008 24237 14048
rect 24355 14008 24395 14048
rect 24460 14008 24500 14048
rect 24940 14008 24980 14048
rect 25137 14008 25177 14048
rect 25276 14008 25316 14048
rect 25466 13984 25506 14024
rect 25804 14008 25844 14048
rect 26143 14008 26183 14048
rect 26668 14008 26708 14048
rect 27007 14008 27047 14048
rect 27405 13987 27445 14027
rect 27523 13999 27563 14039
rect 27632 14008 27672 14048
rect 28204 14008 28244 14048
rect 28588 14008 28628 14048
rect 30883 14008 30923 14048
rect 12940 13924 12980 13964
rect 22147 13924 22187 13964
rect 22723 13924 22763 13964
rect 23596 13924 23636 13964
rect 24099 13924 24139 13964
rect 26026 13924 26066 13964
rect 26890 13924 26930 13964
rect 29347 13924 29387 13964
rect 31267 13924 31307 13964
rect 844 13840 884 13880
rect 6316 13840 6356 13880
rect 11175 13840 11215 13880
rect 20995 13840 21035 13880
rect 23500 13840 23540 13880
rect 26764 13840 26804 13880
rect 28828 13840 28868 13880
rect 5356 13756 5396 13796
rect 11395 13756 11435 13796
rect 11932 13756 11972 13796
rect 18892 13756 18932 13796
rect 19852 13756 19892 13796
rect 25900 13756 25940 13796
rect 28972 13756 29012 13796
rect 3112 13588 3480 13628
rect 10886 13588 11254 13628
rect 18660 13588 19028 13628
rect 26434 13588 26802 13628
rect 2956 13420 2996 13460
rect 3820 13420 3860 13460
rect 14476 13420 14516 13460
rect 16483 13420 16523 13460
rect 17059 13420 17099 13460
rect 20716 13420 20756 13460
rect 21964 13420 22004 13460
rect 23683 13420 23723 13460
rect 24460 13420 24500 13460
rect 25804 13420 25844 13460
rect 26956 13420 26996 13460
rect 5548 13336 5588 13376
rect 6124 13336 6164 13376
rect 6796 13336 6836 13376
rect 8812 13336 8852 13376
rect 9283 13336 9323 13376
rect 10828 13336 10868 13376
rect 13132 13336 13172 13376
rect 13703 13336 13743 13376
rect 15532 13336 15572 13376
rect 19660 13336 19700 13376
rect 27244 13336 27284 13376
rect 29932 13336 29972 13376
rect 652 13252 692 13292
rect 2572 13252 2612 13292
rect 4771 13252 4811 13292
rect 4972 13252 5012 13292
rect 5644 13252 5684 13292
rect 6028 13252 6068 13292
rect 6892 13252 6932 13292
rect 8227 13252 8267 13292
rect 8716 13252 8756 13292
rect 10371 13252 10411 13292
rect 10732 13252 10772 13292
rect 12115 13252 12155 13292
rect 12675 13252 12715 13292
rect 13036 13252 13076 13292
rect 1027 13168 1067 13208
rect 3619 13168 3659 13208
rect 3724 13168 3764 13208
rect 4651 13168 4691 13208
rect 4876 13168 4916 13208
rect 5487 13168 5527 13208
rect 5347 13126 5387 13166
rect 5779 13168 5819 13208
rect 5884 13168 5924 13208
rect 6185 13168 6225 13208
rect 6556 13168 6596 13208
rect 6307 13126 6347 13166
rect 6721 13168 6761 13208
rect 7027 13168 7067 13208
rect 7439 13168 7479 13208
rect 7569 13168 7609 13208
rect 7672 13168 7712 13208
rect 7793 13179 7833 13219
rect 7945 13168 7985 13208
rect 8087 13168 8127 13208
rect 8332 13168 8372 13208
rect 8563 13126 8603 13166
rect 9043 13168 9083 13208
rect 9292 13168 9332 13208
rect 8880 13126 8920 13166
rect 9484 13168 9524 13208
rect 10252 13168 10292 13208
rect 10469 13168 10509 13208
rect 10588 13168 10628 13208
rect 10903 13168 10943 13208
rect 11043 13168 11083 13208
rect 11308 13168 11348 13208
rect 11596 13168 11636 13208
rect 12280 13168 12320 13208
rect 12556 13168 12596 13208
rect 12773 13168 12813 13208
rect 12892 13168 12932 13208
rect 13193 13168 13233 13208
rect 13468 13168 13508 13208
rect 13612 13210 13652 13250
rect 13806 13252 13846 13292
rect 14860 13252 14900 13292
rect 15628 13252 15668 13292
rect 22659 13252 22699 13292
rect 27109 13252 27149 13292
rect 27676 13252 27716 13292
rect 30796 13252 30836 13292
rect 10156 13084 10196 13124
rect 11404 13084 11444 13124
rect 13315 13126 13355 13166
rect 14380 13168 14420 13208
rect 13939 13126 13979 13166
rect 14572 13168 14612 13208
rect 14731 13168 14771 13208
rect 15031 13168 15071 13208
rect 15471 13168 15511 13208
rect 15139 13126 15179 13166
rect 15331 13126 15371 13166
rect 15749 13168 15789 13208
rect 16300 13168 16340 13208
rect 16483 13168 16523 13208
rect 16684 13168 16724 13208
rect 16876 13168 16916 13208
rect 17059 13168 17099 13208
rect 17177 13168 17217 13208
rect 17337 13168 17377 13208
rect 17443 13168 17483 13208
rect 17589 13168 17629 13208
rect 17827 13168 17867 13208
rect 17982 13168 18022 13208
rect 18085 13168 18125 13208
rect 18211 13168 18251 13208
rect 18345 13168 18385 13208
rect 18988 13168 19028 13208
rect 20044 13159 20084 13199
rect 20332 13168 20372 13208
rect 21004 13168 21044 13208
rect 21100 13159 21140 13199
rect 21388 13168 21428 13208
rect 21964 13168 22004 13208
rect 22252 13168 22292 13208
rect 22540 13168 22580 13208
rect 22757 13168 22797 13208
rect 23203 13168 23243 13208
rect 23678 13168 23718 13208
rect 23980 13168 24020 13208
rect 24172 13168 24212 13208
rect 24307 13168 24347 13208
rect 24421 13168 24461 13208
rect 25228 13168 25268 13208
rect 25411 13168 25451 13208
rect 25516 13168 25556 13208
rect 25708 13168 25748 13208
rect 25900 13168 25940 13208
rect 27017 13168 27057 13208
rect 27340 13168 27380 13208
rect 27571 13168 27611 13208
rect 28780 13168 28820 13208
rect 28972 13168 29012 13208
rect 30124 13168 30164 13208
rect 12460 13084 12500 13124
rect 16780 13084 16820 13124
rect 7459 13000 7499 13040
rect 8419 13000 8459 13040
rect 14947 13042 14987 13082
rect 18689 13084 18729 13124
rect 19948 13084 19988 13124
rect 22444 13084 22484 13124
rect 23404 13084 23444 13124
rect 23514 13084 23554 13124
rect 25315 13084 25355 13124
rect 28876 13084 28916 13124
rect 9484 13000 9524 13040
rect 18115 13000 18155 13040
rect 18787 13000 18827 13040
rect 18892 13000 18932 13040
rect 23299 13000 23339 13040
rect 23884 13000 23924 13040
rect 30556 13000 30596 13040
rect 4352 12832 4720 12872
rect 12126 12832 12494 12872
rect 19900 12832 20268 12872
rect 27674 12832 28042 12872
rect 3340 12664 3380 12704
rect 4204 12664 4244 12704
rect 4876 12664 4916 12704
rect 5740 12664 5780 12704
rect 6892 12664 6932 12704
rect 7468 12664 7508 12704
rect 9004 12664 9044 12704
rect 11404 12664 11444 12704
rect 13027 12664 13067 12704
rect 14563 12664 14603 12704
rect 14947 12664 14987 12704
rect 17068 12664 17108 12704
rect 19075 12664 19115 12704
rect 22051 12664 22091 12704
rect 23836 12664 23876 12704
rect 24259 12664 24299 12704
rect 25420 12664 25460 12704
rect 25804 12664 25844 12704
rect 26476 12664 26516 12704
rect 26620 12664 26660 12704
rect 26947 12664 26987 12704
rect 27724 12664 27764 12704
rect 28492 12664 28532 12704
rect 1324 12496 1364 12536
rect 1516 12496 1556 12536
rect 2860 12496 2900 12536
rect 3148 12496 3188 12536
rect 4300 12496 4340 12536
rect 4517 12496 4557 12536
rect 4673 12496 4713 12536
rect 4972 12487 5012 12527
rect 5836 12496 5876 12536
rect 6053 12496 6093 12536
rect 6988 12496 7028 12536
rect 4419 12412 4459 12452
rect 5971 12403 6011 12443
rect 7107 12412 7147 12452
rect 7228 12454 7268 12494
rect 7372 12496 7412 12536
rect 7563 12496 7603 12536
rect 7756 12496 7796 12536
rect 7953 12491 7993 12531
rect 8107 12496 8147 12536
rect 8393 12496 8433 12536
rect 8547 12496 8587 12536
rect 9100 12496 9140 12536
rect 9337 12496 9377 12536
rect 10492 12496 10532 12536
rect 10657 12496 10697 12536
rect 10963 12496 11003 12536
rect 11116 12496 11156 12536
rect 11257 12464 11297 12504
rect 12715 12496 12755 12536
rect 12940 12496 12980 12536
rect 13699 12496 13739 12536
rect 14380 12496 14420 12536
rect 14572 12496 14612 12536
rect 14764 12496 14804 12536
rect 14956 12496 14996 12536
rect 16588 12496 16628 12536
rect 16780 12496 16820 12536
rect 16972 12496 17012 12536
rect 17164 12496 17204 12536
rect 18480 12538 18520 12578
rect 23020 12580 23060 12620
rect 8236 12412 8276 12452
rect 9219 12412 9259 12452
rect 18172 12454 18212 12494
rect 18627 12496 18667 12536
rect 18763 12496 18803 12536
rect 18988 12496 19028 12536
rect 21100 12496 21140 12536
rect 21209 12496 21249 12536
rect 21484 12496 21524 12536
rect 21868 12496 21908 12536
rect 22060 12496 22100 12536
rect 23116 12496 23156 12536
rect 10828 12412 10868 12452
rect 12835 12412 12875 12452
rect 18316 12412 18356 12452
rect 18883 12412 18923 12452
rect 23235 12412 23275 12452
rect 23356 12454 23396 12494
rect 23500 12496 23540 12536
rect 23692 12496 23732 12536
rect 23980 12496 24020 12536
rect 24172 12496 24212 12536
rect 24460 12496 24500 12536
rect 25324 12496 25364 12536
rect 25516 12496 25556 12536
rect 25708 12496 25748 12536
rect 25900 12496 25940 12536
rect 26092 12496 26132 12536
rect 26214 12496 26254 12536
rect 26325 12496 26365 12536
rect 26431 12487 26471 12527
rect 26764 12496 26804 12536
rect 27100 12496 27140 12536
rect 27251 12496 27291 12536
rect 27767 12496 27807 12536
rect 27907 12487 27947 12527
rect 28012 12496 28052 12536
rect 28201 12496 28241 12536
rect 28326 12496 28366 12536
rect 28444 12478 28484 12518
rect 30595 12496 30635 12536
rect 29059 12412 29099 12452
rect 30979 12412 31019 12452
rect 1900 12328 1940 12368
rect 8332 12328 8372 12368
rect 10732 12328 10772 12368
rect 13744 12328 13784 12368
rect 18412 12328 18452 12368
rect 20812 12328 20852 12368
rect 27724 12328 27764 12368
rect 1324 12244 1364 12284
rect 4675 12244 4715 12284
rect 7852 12244 7892 12284
rect 13516 12244 13556 12284
rect 16588 12244 16628 12284
rect 23500 12244 23540 12284
rect 24172 12244 24212 12284
rect 28684 12244 28724 12284
rect 3112 12076 3480 12116
rect 10886 12076 11254 12116
rect 18660 12076 19028 12116
rect 26434 12076 26802 12116
rect 4483 11908 4523 11948
rect 9475 11908 9515 11948
rect 12172 11908 12212 11948
rect 3244 11824 3284 11864
rect 7564 11866 7604 11906
rect 13027 11908 13067 11948
rect 16771 11908 16811 11948
rect 18307 11908 18347 11948
rect 23308 11908 23348 11948
rect 25612 11908 25652 11948
rect 26188 11908 26228 11948
rect 26380 11908 26420 11948
rect 28012 11908 28052 11948
rect 29740 11908 29780 11948
rect 8140 11824 8180 11864
rect 10156 11824 10196 11864
rect 11404 11824 11444 11864
rect 13996 11824 14036 11864
rect 14764 11824 14804 11864
rect 16396 11824 16436 11864
rect 18076 11815 18116 11855
rect 2860 11740 2900 11780
rect 4498 11740 4538 11780
rect 5251 11740 5291 11780
rect 6979 11740 7019 11780
rect 7468 11740 7508 11780
rect 1315 11656 1355 11696
rect 4108 11656 4148 11696
rect 4588 11656 4628 11696
rect 5111 11656 5151 11696
rect 5356 11656 5396 11696
rect 5692 11667 5732 11707
rect 5827 11656 5867 11696
rect 5971 11656 6011 11696
rect 6076 11656 6116 11696
rect 6211 11656 6251 11696
rect 6407 11656 6447 11696
rect 6598 11656 6638 11696
rect 6844 11698 6884 11738
rect 8044 11740 8084 11780
rect 10924 11740 10964 11780
rect 11500 11740 11540 11780
rect 13900 11740 13940 11780
rect 15724 11740 15764 11780
rect 16485 11740 16525 11780
rect 20332 11740 20372 11780
rect 7084 11656 7124 11696
rect 7324 11656 7364 11696
rect 7625 11656 7665 11696
rect 7915 11656 7955 11696
rect 931 11572 971 11612
rect 7747 11614 7787 11654
rect 8371 11656 8411 11696
rect 9142 11656 9182 11696
rect 9484 11656 9524 11696
rect 8208 11614 8248 11654
rect 9591 11656 9631 11696
rect 10156 11656 10196 11696
rect 10483 11656 10523 11696
rect 11107 11656 11147 11696
rect 11780 11656 11820 11696
rect 12652 11656 12692 11696
rect 12835 11656 12875 11696
rect 13027 11656 13067 11696
rect 13183 11656 13223 11696
rect 13285 11656 13325 11696
rect 13406 11656 13446 11696
rect 13545 11656 13585 11696
rect 13756 11656 13796 11696
rect 14071 11656 14111 11696
rect 14227 11656 14267 11696
rect 14572 11656 14612 11696
rect 14947 11656 14987 11696
rect 15065 11656 15105 11696
rect 15197 11656 15237 11696
rect 15331 11656 15371 11696
rect 15465 11656 15505 11696
rect 15820 11656 15860 11696
rect 15955 11647 15995 11687
rect 16060 11656 16100 11696
rect 16163 11656 16203 11696
rect 16335 11656 16375 11696
rect 16613 11656 16653 11696
rect 16771 11656 16811 11696
rect 16915 11656 16955 11696
rect 17163 11656 17203 11696
rect 17332 11656 17372 11696
rect 18115 11656 18155 11696
rect 19363 11656 19403 11696
rect 19852 11656 19892 11696
rect 20428 11656 20468 11696
rect 20812 11656 20852 11696
rect 20930 11656 20970 11696
rect 21868 11656 21908 11696
rect 22051 11656 22091 11696
rect 22204 11656 22244 11696
rect 22376 11698 22416 11738
rect 22540 11740 22580 11780
rect 23116 11740 23156 11780
rect 28419 11740 28459 11780
rect 22661 11656 22701 11696
rect 22803 11656 22843 11696
rect 22915 11656 22955 11696
rect 23020 11656 23060 11696
rect 23308 11656 23348 11696
rect 23609 11656 23649 11696
rect 24460 11656 24500 11696
rect 25324 11656 25364 11696
rect 25446 11656 25486 11696
rect 25564 11656 25604 11696
rect 25996 11656 26036 11696
rect 26380 11656 26420 11696
rect 26577 11656 26617 11696
rect 26860 11656 26900 11696
rect 27715 11656 27755 11696
rect 27820 11656 27860 11696
rect 28300 11656 28340 11696
rect 28517 11656 28557 11696
rect 28876 11656 28916 11696
rect 29548 11656 29588 11696
rect 29740 11656 29780 11696
rect 29932 11656 29972 11696
rect 30124 11656 30164 11696
rect 30316 11656 30356 11696
rect 30691 11656 30731 11696
rect 6508 11572 6548 11612
rect 8947 11572 8987 11612
rect 11404 11572 11444 11612
rect 12748 11572 12788 11612
rect 17059 11605 17099 11645
rect 21964 11572 22004 11612
rect 3436 11488 3476 11528
rect 5443 11488 5483 11528
rect 5731 11488 5771 11528
rect 7171 11488 7211 11528
rect 13507 11488 13547 11528
rect 14467 11488 14507 11528
rect 15427 11488 15467 11528
rect 19180 11488 19220 11528
rect 22458 11530 22498 11570
rect 26476 11572 26516 11612
rect 28026 11572 28066 11612
rect 28204 11572 28244 11612
rect 30220 11572 30260 11612
rect 23788 11488 23828 11528
rect 25891 11488 25931 11528
rect 27532 11488 27572 11528
rect 30892 11488 30932 11528
rect 4352 11320 4720 11360
rect 12126 11320 12494 11360
rect 19900 11320 20268 11360
rect 27674 11320 28042 11360
rect 4195 11152 4235 11192
rect 4771 11152 4811 11192
rect 5164 11152 5204 11192
rect 6940 11152 6980 11192
rect 7276 11152 7316 11192
rect 8044 11152 8084 11192
rect 8908 11152 8948 11192
rect 10555 11152 10595 11192
rect 11395 11152 11435 11192
rect 11692 11152 11732 11192
rect 12604 11152 12644 11192
rect 13516 11152 13556 11192
rect 14371 11152 14411 11192
rect 15619 11152 15659 11192
rect 16684 11152 16724 11192
rect 17836 11152 17876 11192
rect 19180 11152 19220 11192
rect 19468 11152 19508 11192
rect 21868 11152 21908 11192
rect 26668 11152 26708 11192
rect 26995 11152 27035 11192
rect 27916 11152 27956 11192
rect 3907 11068 3947 11108
rect 14860 11068 14900 11108
rect 17260 11068 17300 11108
rect 22252 11068 22292 11108
rect 23404 11068 23444 11108
rect 31267 11068 31307 11108
rect 1132 10984 1172 11024
rect 1257 10984 1297 11024
rect 1420 10984 1460 11024
rect 2956 10984 2996 11024
rect 3448 10984 3488 11024
rect 4108 10984 4148 11024
rect 4420 10984 4460 11024
rect 4557 10984 4597 11024
rect 4696 10984 4736 11024
rect 4862 10984 4902 11024
rect 4963 10984 5003 11024
rect 5260 10984 5300 11024
rect 5497 10984 5537 11024
rect 6412 10984 6452 11024
rect 6595 10984 6635 11024
rect 7084 10984 7124 11024
rect 7372 10984 7412 11024
rect 7609 10984 7649 11024
rect 8140 10984 8180 11024
rect 8357 10984 8397 11024
rect 8620 10984 8660 11024
rect 8742 10984 8782 11024
rect 8869 10984 8909 11024
rect 9261 10975 9301 11015
rect 9379 10975 9419 11015
rect 9489 10984 9529 11024
rect 10336 10975 10376 11015
rect 10435 10984 10475 11024
rect 11063 10984 11103 11024
rect 11306 10984 11346 11024
rect 11596 10984 11636 11024
rect 11788 10984 11828 11024
rect 13132 10984 13172 11024
rect 13301 10984 13341 11024
rect 3283 10900 3323 10940
rect 5395 10891 5435 10931
rect 7507 10891 7547 10931
rect 8259 10900 8299 10940
rect 11203 10900 11243 10940
rect 12364 10900 12404 10940
rect 13612 10942 13652 10982
rect 13829 10984 13869 11024
rect 14270 10984 14310 11024
rect 14476 10984 14516 11024
rect 14572 10975 14612 11015
rect 14956 10984 14996 11024
rect 15193 10984 15233 11024
rect 15427 10984 15467 11024
rect 15772 10984 15812 11024
rect 16243 10984 16283 11024
rect 16780 10984 16820 11024
rect 16099 10942 16139 10982
rect 17017 10984 17057 11024
rect 17356 10984 17396 11024
rect 17593 10984 17633 11024
rect 17740 10984 17780 11024
rect 17932 10984 17972 11024
rect 18691 10984 18731 11024
rect 19084 10984 19124 11024
rect 19276 10984 19316 11024
rect 19651 10984 19691 11024
rect 20140 10975 20180 11015
rect 20620 10984 20660 11024
rect 21100 10984 21140 11024
rect 21218 10984 21258 11024
rect 21772 10984 21812 11024
rect 21955 10984 21995 11024
rect 22156 10984 22196 11024
rect 22348 10984 22388 11024
rect 22723 10984 22763 11024
rect 22828 10984 22868 11024
rect 23308 10984 23348 11024
rect 23491 10984 23531 11024
rect 23884 10984 23924 11024
rect 24067 10984 24107 11024
rect 24178 10972 24218 11012
rect 24739 10984 24779 11024
rect 27190 10984 27230 11024
rect 27523 10984 27563 11024
rect 27628 10984 27668 11024
rect 28108 10984 28148 11024
rect 30883 10984 30923 11024
rect 13731 10900 13771 10940
rect 15091 10891 15131 10931
rect 15916 10900 15956 10940
rect 16915 10891 16955 10931
rect 17491 10891 17531 10931
rect 18307 10900 18347 10940
rect 18883 10900 18923 10940
rect 20716 10900 20756 10940
rect 24364 10900 24404 10940
rect 26284 10900 26324 10940
rect 1132 10816 1172 10856
rect 9100 10816 9140 10856
rect 10051 10816 10091 10856
rect 15399 10816 15439 10856
rect 16012 10816 16052 10856
rect 18403 10816 18443 10856
rect 24172 10816 24212 10856
rect 2284 10732 2324 10772
rect 6595 10732 6635 10772
rect 13315 10732 13355 10772
rect 23011 10732 23051 10772
rect 28780 10732 28820 10772
rect 28972 10732 29012 10772
rect 29356 10732 29396 10772
rect 3112 10564 3480 10604
rect 10886 10564 11254 10604
rect 18660 10564 19028 10604
rect 26434 10564 26802 10604
rect 652 10396 692 10436
rect 4876 10396 4916 10436
rect 5731 10396 5771 10436
rect 9475 10396 9515 10436
rect 14947 10396 14987 10436
rect 21100 10396 21140 10436
rect 22444 10396 22484 10436
rect 24748 10396 24788 10436
rect 27148 10396 27188 10436
rect 29932 10396 29972 10436
rect 2371 10312 2411 10352
rect 7180 10312 7220 10352
rect 12268 10312 12308 10352
rect 18796 10312 18836 10352
rect 25036 10312 25076 10352
rect 25420 10312 25460 10352
rect 28387 10312 28427 10352
rect 3052 10228 3092 10268
rect 6220 10228 6260 10268
rect 6451 10219 6491 10259
rect 6915 10228 6955 10268
rect 7651 10228 7691 10268
rect 7852 10228 7892 10268
rect 8428 10228 8468 10268
rect 10755 10228 10795 10268
rect 844 10144 884 10184
rect 1420 10144 1460 10184
rect 1555 10144 1595 10184
rect 2083 10144 2123 10184
rect 2188 10144 2228 10184
rect 2711 10144 2751 10184
rect 2851 10144 2891 10184
rect 2956 10144 2996 10184
rect 3532 10144 3572 10184
rect 3916 10144 3956 10184
rect 4316 10155 4356 10195
rect 4507 10144 4547 10184
rect 4627 10144 4667 10184
rect 4766 10144 4806 10184
rect 4867 10144 4907 10184
rect 5443 10144 5483 10184
rect 5548 10144 5588 10184
rect 6316 10144 6356 10184
rect 6547 10144 6587 10184
rect 6796 10144 6836 10184
rect 7033 10144 7073 10184
rect 7180 10144 7220 10184
rect 7377 10144 7417 10184
rect 7531 10144 7571 10184
rect 7756 10144 7796 10184
rect 8044 10144 8084 10184
rect 8236 10144 8276 10184
rect 8524 10144 8564 10184
rect 8643 10144 8683 10184
rect 8761 10144 8801 10184
rect 9238 10144 9278 10184
rect 9868 10144 9908 10184
rect 10636 10144 10676 10184
rect 10867 10144 10907 10184
rect 10972 10186 11012 10226
rect 11093 10228 11133 10268
rect 11308 10228 11348 10268
rect 11884 10228 11924 10268
rect 12364 10228 12404 10268
rect 13315 10228 13355 10268
rect 13516 10228 13556 10268
rect 11205 10144 11245 10184
rect 11543 10144 11583 10184
rect 11683 10144 11723 10184
rect 11788 10144 11828 10184
rect 12045 10144 12085 10184
rect 12499 10186 12539 10226
rect 14419 10228 14459 10268
rect 15436 10228 15476 10268
rect 15667 10219 15707 10259
rect 16492 10228 16532 10268
rect 16723 10219 16763 10259
rect 17187 10228 17227 10268
rect 31036 10228 31076 10268
rect 12193 10144 12233 10184
rect 13203 10144 13243 10184
rect 13420 10144 13460 10184
rect 14614 10144 14654 10184
rect 14851 10135 14891 10175
rect 15148 10144 15188 10184
rect 15532 10144 15572 10184
rect 15769 10144 15809 10184
rect 16588 10144 16628 10184
rect 16825 10144 16865 10184
rect 17068 10144 17108 10184
rect 17305 10144 17345 10184
rect 17447 10144 17487 10184
rect 17635 10144 17675 10184
rect 18604 10144 18644 10184
rect 18719 10144 18759 10184
rect 18892 10144 18932 10184
rect 19084 10144 19124 10184
rect 19276 10144 19316 10184
rect 19948 10144 19988 10184
rect 20044 10144 20084 10184
rect 20320 10144 20360 10184
rect 21148 10144 21188 10184
rect 21292 10144 21332 10184
rect 21772 10144 21812 10184
rect 22636 10144 22676 10184
rect 23500 10144 23540 10184
rect 24556 10144 24596 10184
rect 24940 10144 24980 10184
rect 26668 10144 26708 10184
rect 26860 10144 26900 10184
rect 27052 10144 27092 10184
rect 28108 10144 28148 10184
rect 28396 10144 28436 10184
rect 28588 10144 28628 10184
rect 29068 10144 29108 10184
rect 29932 10144 29972 10184
rect 30047 10144 30087 10184
rect 30220 10144 30260 10184
rect 30355 10144 30395 10184
rect 30850 10144 30890 10184
rect 4156 10060 4196 10100
rect 9043 10060 9083 10100
rect 10540 10060 10580 10100
rect 16972 10060 17012 10100
rect 19180 10060 19220 10100
rect 19742 10060 19782 10100
rect 20476 10060 20516 10100
rect 26764 10060 26804 10100
rect 29740 10060 29780 10100
rect 30556 10060 30596 10100
rect 931 9976 971 10016
rect 1708 9976 1748 10016
rect 5836 9976 5876 10016
rect 6700 9976 6740 10016
rect 8227 9976 8267 10016
rect 17548 9976 17588 10016
rect 19843 9976 19883 10016
rect 23308 9976 23348 10016
rect 24172 9976 24212 10016
rect 24451 9976 24491 10016
rect 27436 9976 27476 10016
rect 4352 9808 4720 9848
rect 12126 9808 12494 9848
rect 19900 9808 20268 9848
rect 27674 9808 28042 9848
rect 1603 9640 1643 9680
rect 1900 9640 1940 9680
rect 2851 9640 2891 9680
rect 5836 9640 5876 9680
rect 6403 9640 6443 9680
rect 7459 9640 7499 9680
rect 8419 9640 8459 9680
rect 8524 9640 8564 9680
rect 8908 9640 8948 9680
rect 10483 9640 10523 9680
rect 11107 9640 11147 9680
rect 11779 9640 11819 9680
rect 13597 9640 13637 9680
rect 14428 9640 14468 9680
rect 15532 9640 15572 9680
rect 15964 9640 16004 9680
rect 18835 9640 18875 9680
rect 19372 9640 19412 9680
rect 20524 9640 20564 9680
rect 25612 9640 25652 9680
rect 27619 9640 27659 9680
rect 27724 9640 27764 9680
rect 28780 9640 28820 9680
rect 28972 9640 29012 9680
rect 2956 9556 2996 9596
rect 6618 9556 6658 9596
rect 6892 9556 6932 9596
rect 7852 9556 7892 9596
rect 8321 9556 8361 9596
rect 11212 9556 11252 9596
rect 11932 9556 11972 9596
rect 20131 9556 20171 9596
rect 24211 9556 24251 9596
rect 31267 9556 31307 9596
rect 1123 9472 1163 9512
rect 1420 9472 1460 9512
rect 1708 9472 1748 9512
rect 2059 9472 2099 9512
rect 2345 9472 2385 9512
rect 2515 9472 2555 9512
rect 2755 9472 2795 9512
rect 3063 9472 3103 9512
rect 5932 9472 5972 9512
rect 6149 9472 6189 9512
rect 6307 9472 6347 9512
rect 6412 9472 6452 9512
rect 6796 9472 6836 9512
rect 6979 9472 7019 9512
rect 7127 9472 7167 9512
rect 7372 9472 7412 9512
rect 7948 9472 7988 9512
rect 8182 9472 8222 9512
rect 8620 9463 8660 9503
rect 8812 9472 8852 9512
rect 9004 9472 9044 9512
rect 10648 9472 10688 9512
rect 11006 9472 11046 9512
rect 11308 9463 11348 9503
rect 11447 9472 11487 9512
rect 11692 9472 11732 9512
rect 12076 9472 12116 9512
rect 12844 9472 12884 9512
rect 13228 9472 13268 9512
rect 13699 9472 13739 9512
rect 13804 9463 13844 9503
rect 14275 9463 14315 9503
rect 14755 9463 14795 9503
rect 15436 9472 15476 9512
rect 15619 9472 15659 9512
rect 15811 9463 15851 9503
rect 16588 9472 16628 9512
rect 16703 9472 16743 9512
rect 16876 9472 16916 9512
rect 17591 9472 17631 9512
rect 17836 9472 17876 9512
rect 19030 9472 19070 9512
rect 19468 9472 19508 9512
rect 19819 9472 19859 9512
rect 20037 9472 20077 9512
rect 22435 9472 22475 9512
rect 23416 9472 23456 9512
rect 23596 9472 23636 9512
rect 2188 9388 2228 9428
rect 6051 9388 6091 9428
rect 7267 9388 7307 9428
rect 8083 9379 8123 9419
rect 11587 9388 11627 9428
rect 14908 9388 14948 9428
rect 17731 9388 17771 9428
rect 17932 9388 17972 9428
rect 19587 9388 19627 9428
rect 19708 9430 19748 9470
rect 23779 9472 23819 9512
rect 24376 9472 24416 9512
rect 24855 9445 24895 9485
rect 25804 9472 25844 9512
rect 26092 9472 26132 9512
rect 26214 9472 26254 9512
rect 26341 9472 26381 9512
rect 26572 9472 26612 9512
rect 26755 9472 26795 9512
rect 26860 9472 26900 9512
rect 27379 9472 27419 9512
rect 27523 9472 27563 9512
rect 27834 9472 27874 9512
rect 19925 9388 19965 9428
rect 20899 9388 20939 9428
rect 22819 9388 22859 9428
rect 23251 9388 23291 9428
rect 28481 9445 28521 9485
rect 28627 9472 28667 9512
rect 30883 9472 30923 9512
rect 24754 9388 24794 9428
rect 27187 9388 27227 9428
rect 29347 9388 29387 9428
rect 2284 9304 2324 9344
rect 16588 9304 16628 9344
rect 26380 9304 26420 9344
rect 1420 9220 1460 9260
rect 6604 9220 6644 9260
rect 13468 9220 13508 9260
rect 14092 9220 14132 9260
rect 23779 9220 23819 9260
rect 24652 9220 24692 9260
rect 26860 9220 26900 9260
rect 3112 9052 3480 9092
rect 10886 9052 11254 9092
rect 18660 9052 19028 9092
rect 26434 9052 26802 9092
rect 1219 8884 1259 8924
rect 3907 8884 3947 8924
rect 4876 8884 4916 8924
rect 5635 8884 5675 8924
rect 8323 8884 8363 8924
rect 12652 8884 12692 8924
rect 13900 8884 13940 8924
rect 14467 8884 14507 8924
rect 20035 8884 20075 8924
rect 23452 8884 23492 8924
rect 27100 8884 27140 8924
rect 28972 8884 29012 8924
rect 29932 8884 29972 8924
rect 11203 8800 11243 8840
rect 17788 8791 17828 8831
rect 19852 8800 19892 8840
rect 21772 8800 21812 8840
rect 26572 8800 26612 8840
rect 31084 8800 31124 8840
rect 2563 8716 2603 8756
rect 2764 8716 2804 8756
rect 4978 8716 5018 8756
rect 9196 8716 9236 8756
rect 11587 8716 11627 8756
rect 11788 8716 11828 8756
rect 15532 8716 15572 8756
rect 15747 8716 15787 8756
rect 17203 8707 17243 8747
rect 18220 8716 18260 8756
rect 18451 8707 18491 8747
rect 30034 8716 30074 8756
rect 1612 8632 1652 8672
rect 2092 8632 2132 8672
rect 2284 8632 2324 8672
rect 2423 8632 2463 8672
rect 2668 8632 2708 8672
rect 2947 8632 2987 8672
rect 3244 8632 3284 8672
rect 3619 8632 3659 8672
rect 3724 8632 3764 8672
rect 4195 8632 4235 8672
rect 4300 8632 4340 8672
rect 5068 8632 5108 8672
rect 6028 8632 6068 8672
rect 6883 8632 6923 8672
rect 6988 8632 7028 8672
rect 8035 8632 8075 8672
rect 8140 8632 8180 8672
rect 8707 8632 8747 8672
rect 8812 8632 8852 8672
rect 9292 8632 9332 8672
rect 9772 8632 9812 8672
rect 10291 8632 10331 8672
rect 10915 8632 10955 8672
rect 11020 8632 11060 8672
rect 11467 8632 11507 8672
rect 11692 8632 11732 8672
rect 12259 8632 12299 8672
rect 12368 8665 12408 8705
rect 13603 8632 13643 8672
rect 13708 8632 13748 8672
rect 14764 8632 14804 8672
rect 15040 8632 15080 8672
rect 15628 8632 15668 8672
rect 15865 8632 15905 8672
rect 16195 8632 16235 8672
rect 16300 8643 16340 8683
rect 16445 8632 16485 8672
rect 16575 8632 16615 8672
rect 16713 8632 16753 8672
rect 17068 8632 17108 8672
rect 17305 8632 17345 8672
rect 17827 8632 17867 8672
rect 18315 8632 18355 8672
rect 18553 8632 18593 8672
rect 19180 8632 19220 8672
rect 19459 8632 19499 8672
rect 20236 8632 20276 8672
rect 20338 8632 20378 8672
rect 23788 8632 23828 8672
rect 24076 8632 24116 8672
rect 24643 8674 24683 8714
rect 24455 8632 24495 8672
rect 24844 8632 24884 8672
rect 26956 8632 26996 8672
rect 28108 8632 28148 8672
rect 29644 8632 29684 8672
rect 30124 8632 30164 8672
rect 30547 8632 30587 8672
rect 4503 8548 4543 8588
rect 5731 8548 5771 8588
rect 13914 8548 13954 8588
rect 14465 8548 14505 8588
rect 18028 8548 18068 8588
rect 19564 8548 19604 8588
rect 20030 8548 20070 8588
rect 24556 8548 24596 8588
rect 2275 8464 2315 8504
rect 3148 8464 3188 8504
rect 4396 8464 4436 8504
rect 7276 8464 7316 8504
rect 10444 8464 10484 8504
rect 12163 8455 12203 8495
rect 14668 8464 14708 8504
rect 15196 8464 15236 8504
rect 16675 8464 16715 8504
rect 16972 8464 17012 8504
rect 28780 8464 28820 8504
rect 30748 8464 30788 8504
rect 4352 8296 4720 8336
rect 12126 8296 12494 8336
rect 19900 8296 20268 8336
rect 27674 8296 28042 8336
rect 2476 8128 2516 8168
rect 3235 8128 3275 8168
rect 4195 8128 4235 8168
rect 4492 8128 4532 8168
rect 5164 8128 5204 8168
rect 5395 8128 5435 8168
rect 6988 8128 7028 8168
rect 7459 8128 7499 8168
rect 11875 8128 11915 8168
rect 12259 8128 12299 8168
rect 13324 8128 13364 8168
rect 13900 8128 13940 8168
rect 16588 8128 16628 8168
rect 16876 8128 16916 8168
rect 18019 8128 18059 8168
rect 18124 8128 18164 8168
rect 18412 8128 18452 8168
rect 19363 8128 19403 8168
rect 19468 8128 19508 8168
rect 19747 8128 19787 8168
rect 22060 8128 22100 8168
rect 25420 8128 25460 8168
rect 27916 8128 27956 8168
rect 29164 8128 29204 8168
rect 30124 8128 30164 8168
rect 7756 8044 7796 8084
rect 12090 8044 12130 8084
rect 17356 8044 17396 8084
rect 17921 8044 17961 8084
rect 23107 8044 23147 8084
rect 25603 8044 25643 8084
rect 940 7960 980 8000
rect 1132 7960 1172 8000
rect 1507 7960 1547 8000
rect 1612 7960 1652 8000
rect 2380 7960 2420 8000
rect 2903 7960 2943 8000
rect 2563 7918 2603 7958
rect 3148 7960 3188 8000
rect 4300 7960 4340 8000
rect 4684 7960 4724 8000
rect 5068 7960 5108 8000
rect 5539 7960 5579 8000
rect 5644 7951 5684 7991
rect 6595 7960 6635 8000
rect 6700 7960 6740 8000
rect 7127 7960 7167 8000
rect 7372 7960 7412 8000
rect 7660 7960 7700 8000
rect 7852 7960 7892 8000
rect 9580 7960 9620 8000
rect 11779 7960 11819 8000
rect 11884 7960 11924 8000
rect 12445 7960 12485 8000
rect 12556 7960 12596 8000
rect 13036 7960 13076 8000
rect 13178 7928 13218 7968
rect 14092 7960 14132 8000
rect 14668 7960 14708 8000
rect 14860 7960 14900 8000
rect 16492 7960 16532 8000
rect 16675 7960 16715 8000
rect 16876 7960 16916 8000
rect 17068 7960 17108 8000
rect 17260 7960 17300 8000
rect 17452 7960 17492 8000
rect 18220 7951 18260 7991
rect 18508 7960 18548 8000
rect 3043 7876 3083 7916
rect 7267 7876 7307 7916
rect 18627 7876 18667 7916
rect 18748 7918 18788 7958
rect 19265 7960 19305 8000
rect 19564 7951 19604 7991
rect 20044 7960 20084 8000
rect 21676 7951 21716 7991
rect 21787 7951 21827 7991
rect 21907 7951 21947 7991
rect 22339 7960 22379 8000
rect 22732 7960 22772 8000
rect 23491 7960 23531 8000
rect 25987 7960 26027 8000
rect 28771 7960 28811 8000
rect 28876 7960 28916 8000
rect 29731 7960 29771 8000
rect 29838 7960 29878 8000
rect 30499 7960 30539 8000
rect 30604 7960 30644 8000
rect 19954 7876 19994 7916
rect 27532 7876 27572 7916
rect 1036 7792 1076 7832
rect 5932 7792 5972 7832
rect 31084 7792 31124 7832
rect 1795 7708 1835 7748
rect 9436 7708 9476 7748
rect 12076 7708 12116 7748
rect 14764 7708 14804 7748
rect 25036 7708 25076 7748
rect 30700 7708 30740 7748
rect 3112 7540 3480 7580
rect 10886 7540 11254 7580
rect 18660 7540 19028 7580
rect 26434 7540 26802 7580
rect 1507 7372 1547 7412
rect 3148 7372 3188 7412
rect 4972 7372 5012 7412
rect 6883 7372 6923 7412
rect 9964 7372 10004 7412
rect 11980 7372 12020 7412
rect 12739 7372 12779 7412
rect 14755 7372 14795 7412
rect 18220 7372 18260 7412
rect 20419 7372 20459 7412
rect 21292 7372 21332 7412
rect 22060 7372 22100 7412
rect 30508 7372 30548 7412
rect 8131 7288 8171 7328
rect 19459 7288 19499 7328
rect 19612 7288 19652 7328
rect 24652 7288 24692 7328
rect 28876 7288 28916 7328
rect 29644 7288 29684 7328
rect 1891 7204 1931 7244
rect 2092 7204 2132 7244
rect 4435 7195 4475 7235
rect 8908 7204 8948 7244
rect 9484 7204 9524 7244
rect 12499 7232 12539 7272
rect 18499 7204 18539 7244
rect 18700 7204 18740 7244
rect 1219 7120 1259 7160
rect 1324 7120 1364 7160
rect 1751 7120 1791 7160
rect 1996 7120 2036 7160
rect 2284 7120 2324 7160
rect 2476 7120 2516 7160
rect 2851 7120 2891 7160
rect 2956 7120 2996 7160
rect 4300 7120 4340 7160
rect 4534 7120 4574 7160
rect 4686 7153 4726 7193
rect 27571 7204 27611 7244
rect 29923 7204 29963 7244
rect 30124 7204 30164 7244
rect 4983 7120 5023 7160
rect 6700 7120 6740 7160
rect 6883 7120 6923 7160
rect 7843 7120 7883 7160
rect 7948 7120 7988 7160
rect 8375 7120 8415 7160
rect 8515 7120 8555 7160
rect 8620 7120 8660 7160
rect 9091 7120 9131 7160
rect 10045 7120 10085 7160
rect 10156 7153 10196 7193
rect 30610 7204 30650 7244
rect 10967 7120 11007 7160
rect 11107 7120 11147 7160
rect 11212 7120 11252 7160
rect 12172 7120 12212 7160
rect 12547 7120 12587 7160
rect 13228 7120 13268 7160
rect 13423 7120 13463 7160
rect 14467 7120 14507 7160
rect 14572 7120 14612 7160
rect 15196 7120 15236 7160
rect 15340 7120 15380 7160
rect 18013 7120 18053 7160
rect 18359 7120 18399 7160
rect 18604 7120 18644 7160
rect 19276 7120 19316 7160
rect 19459 7120 19499 7160
rect 19948 7120 19988 7160
rect 20236 7120 20276 7160
rect 20414 7120 20454 7160
rect 20716 7120 20756 7160
rect 21340 7120 21380 7160
rect 21484 7120 21524 7160
rect 22141 7120 22181 7160
rect 22252 7120 22292 7160
rect 23308 7120 23348 7160
rect 23500 7120 23540 7160
rect 23776 7120 23816 7160
rect 24268 7120 24308 7160
rect 25024 7120 25064 7160
rect 25180 7120 25220 7160
rect 27766 7120 27806 7160
rect 28588 7120 28628 7160
rect 28876 7120 28916 7160
rect 28991 7120 29031 7160
rect 29164 7120 29204 7160
rect 29356 7120 29396 7160
rect 29478 7120 29518 7160
rect 29596 7153 29636 7193
rect 29783 7120 29823 7160
rect 30028 7120 30068 7160
rect 30700 7120 30740 7160
rect 2380 7036 2420 7076
rect 3159 7036 3199 7076
rect 4204 7036 4244 7076
rect 9388 7036 9428 7076
rect 23203 7036 23243 7076
rect 28195 7036 28235 7076
rect 4771 6952 4811 6992
rect 8707 6952 8747 6992
rect 11299 6952 11339 6992
rect 12259 6952 12299 6992
rect 13411 6952 13451 6992
rect 15043 6952 15083 6992
rect 17923 6952 17963 6992
rect 20620 6952 20660 6992
rect 23500 6952 23540 6992
rect 23932 6952 23972 6992
rect 24364 6952 24404 6992
rect 4352 6784 4720 6824
rect 12126 6784 12494 6824
rect 19900 6784 20268 6824
rect 27674 6784 28042 6824
rect 1900 6616 1940 6656
rect 2668 6616 2708 6656
rect 3916 6616 3956 6656
rect 4684 6616 4724 6656
rect 6211 6616 6251 6656
rect 7468 6616 7508 6656
rect 8035 6616 8075 6656
rect 9292 6616 9332 6656
rect 10156 6616 10196 6656
rect 10828 6616 10868 6656
rect 12547 6616 12587 6656
rect 13516 6616 13556 6656
rect 16972 6616 17012 6656
rect 18211 6616 18251 6656
rect 21571 6616 21611 6656
rect 22492 6616 22532 6656
rect 23500 6616 23540 6656
rect 23683 6616 23723 6656
rect 26755 6616 26795 6656
rect 28780 6616 28820 6656
rect 29539 6616 29579 6656
rect 6604 6532 6644 6572
rect 6711 6532 6751 6572
rect 8140 6532 8180 6572
rect 14092 6532 14132 6572
rect 15043 6532 15083 6572
rect 29251 6532 29291 6572
rect 29751 6532 29791 6572
rect 1507 6448 1547 6488
rect 1612 6448 1652 6488
rect 2188 6448 2228 6488
rect 2476 6448 2516 6488
rect 2956 6448 2996 6488
rect 3148 6448 3188 6488
rect 3523 6448 3563 6488
rect 3628 6448 3668 6488
rect 4291 6448 4331 6488
rect 4396 6448 4436 6488
rect 4876 6448 4916 6488
rect 5068 6448 5108 6488
rect 3052 6364 3092 6404
rect 5884 6406 5924 6446
rect 6124 6448 6164 6488
rect 6403 6448 6443 6488
rect 6508 6448 6548 6488
rect 6988 6448 7028 6488
rect 7276 6448 7316 6488
rect 7934 6448 7974 6488
rect 8236 6439 8276 6479
rect 9196 6448 9236 6488
rect 9388 6448 9428 6488
rect 9676 6448 9716 6488
rect 9964 6448 10004 6488
rect 10540 6448 10580 6488
rect 10679 6448 10719 6488
rect 11875 6448 11915 6488
rect 11980 6448 12020 6488
rect 12748 6448 12788 6488
rect 13036 6448 13076 6488
rect 13612 6448 13652 6488
rect 13731 6448 13771 6488
rect 13849 6448 13889 6488
rect 13996 6448 14036 6488
rect 14179 6448 14219 6488
rect 14711 6448 14751 6488
rect 14956 6448 14996 6488
rect 15811 6448 15851 6488
rect 15916 6448 15956 6488
rect 16673 6448 16713 6488
rect 16819 6448 16859 6488
rect 17443 6448 17483 6488
rect 17740 6448 17780 6488
rect 17884 6406 17924 6446
rect 18125 6448 18165 6488
rect 19084 6448 19124 6488
rect 20323 6448 20363 6488
rect 21772 6448 21812 6488
rect 22060 6448 22100 6488
rect 22348 6448 22388 6488
rect 23107 6448 23147 6488
rect 23212 6448 23252 6488
rect 23980 6448 24020 6488
rect 25219 6448 25259 6488
rect 25948 6448 25988 6488
rect 26092 6448 26132 6488
rect 27052 6448 27092 6488
rect 27820 6448 27860 6488
rect 28060 6448 28100 6488
rect 28300 6448 28340 6488
rect 28444 6448 28484 6488
rect 28588 6448 28628 6488
rect 28919 6448 28959 6488
rect 29164 6448 29204 6488
rect 29443 6448 29483 6488
rect 30604 6448 30644 6488
rect 6019 6364 6059 6404
rect 14851 6364 14891 6404
rect 18019 6364 18059 6404
rect 23890 6364 23930 6404
rect 25036 6364 25076 6404
rect 25612 6364 25652 6404
rect 26962 6364 27002 6404
rect 27475 6364 27515 6404
rect 29059 6364 29099 6404
rect 30514 6364 30554 6404
rect 12163 6280 12203 6320
rect 25516 6280 25556 6320
rect 4972 6196 5012 6236
rect 16099 6196 16139 6236
rect 17740 6196 17780 6236
rect 18691 6196 18731 6236
rect 20716 6196 20756 6236
rect 25987 6196 26027 6236
rect 29740 6196 29780 6236
rect 30412 6196 30452 6236
rect 3112 6028 3480 6068
rect 10886 6028 11254 6068
rect 18660 6028 19028 6068
rect 26434 6028 26802 6068
rect 4348 5860 4388 5900
rect 16483 5860 16523 5900
rect 20908 5860 20948 5900
rect 21475 5860 21515 5900
rect 25411 5860 25451 5900
rect 27907 5860 27947 5900
rect 29260 5860 29300 5900
rect 30595 5860 30635 5900
rect 4684 5776 4724 5816
rect 6268 5767 6308 5807
rect 7276 5776 7316 5816
rect 9580 5776 9620 5816
rect 22051 5776 22091 5816
rect 2467 5692 2507 5732
rect 2668 5692 2708 5732
rect 4588 5692 4628 5732
rect 6787 5692 6827 5732
rect 6988 5692 7028 5732
rect 652 5608 692 5648
rect 1036 5608 1076 5648
rect 1603 5608 1643 5648
rect 1708 5608 1748 5648
rect 2327 5608 2367 5648
rect 2572 5608 2612 5648
rect 2860 5608 2900 5648
rect 3052 5608 3092 5648
rect 3436 5608 3476 5648
rect 3628 5608 3668 5648
rect 4771 5650 4811 5690
rect 4204 5608 4244 5648
rect 4899 5608 4939 5648
rect 4435 5566 4475 5606
rect 5452 5608 5492 5648
rect 5740 5608 5780 5648
rect 6307 5608 6347 5648
rect 6647 5608 6687 5648
rect 6892 5608 6932 5648
rect 7180 5608 7220 5648
rect 7852 5608 7892 5648
rect 8236 5608 8276 5648
rect 8764 5608 8804 5648
rect 8908 5608 8948 5648
rect 9340 5650 9380 5690
rect 9484 5692 9524 5732
rect 10867 5692 10907 5732
rect 13228 5692 13268 5732
rect 18691 5692 18731 5732
rect 18892 5692 18932 5732
rect 9811 5608 9851 5648
rect 11059 5608 11099 5648
rect 11203 5608 11243 5648
rect 12449 5608 12489 5648
rect 2956 5524 2996 5564
rect 6508 5524 6548 5564
rect 9648 5566 9688 5606
rect 12748 5608 12788 5648
rect 12892 5608 12932 5648
rect 13027 5608 13067 5648
rect 13132 5608 13172 5648
rect 13996 5608 14036 5648
rect 14284 5608 14324 5648
rect 14620 5608 14660 5648
rect 14764 5608 14804 5648
rect 15235 5608 15275 5648
rect 15340 5608 15380 5648
rect 16195 5608 16235 5648
rect 16300 5641 16340 5681
rect 21490 5692 21530 5732
rect 29731 5692 29771 5732
rect 29932 5692 29972 5732
rect 17548 5608 17588 5648
rect 17692 5641 17732 5681
rect 18124 5608 18164 5648
rect 18263 5608 18303 5648
rect 18551 5608 18591 5648
rect 18796 5608 18836 5648
rect 20140 5608 20180 5648
rect 20428 5608 20468 5648
rect 20611 5608 20651 5648
rect 20716 5608 20756 5648
rect 21580 5608 21620 5648
rect 22336 5641 22376 5681
rect 22435 5608 22475 5648
rect 24460 5608 24500 5648
rect 24748 5608 24788 5648
rect 25228 5608 25268 5648
rect 25411 5608 25451 5648
rect 25804 5608 25844 5648
rect 25911 5608 25951 5648
rect 27619 5608 27659 5648
rect 27724 5608 27764 5648
rect 28483 5608 28523 5648
rect 28972 5608 29012 5648
rect 29094 5608 29134 5648
rect 29221 5608 29261 5648
rect 29591 5608 29631 5648
rect 29837 5608 29877 5648
rect 30124 5608 30164 5648
rect 30263 5641 30303 5681
rect 30892 5608 30932 5648
rect 11511 5524 11551 5564
rect 12547 5524 12587 5564
rect 15436 5524 15476 5564
rect 15543 5524 15583 5564
rect 20919 5524 20959 5564
rect 28794 5524 28834 5564
rect 30590 5524 30630 5564
rect 1132 5440 1172 5480
rect 1996 5440 2036 5480
rect 3619 5440 3659 5480
rect 5932 5440 5972 5480
rect 8332 5440 8372 5480
rect 8611 5440 8651 5480
rect 11299 5440 11339 5480
rect 11404 5440 11444 5480
rect 12652 5440 12692 5480
rect 13795 5440 13835 5480
rect 14467 5440 14507 5480
rect 17836 5440 17876 5480
rect 18412 5440 18452 5480
rect 19939 5440 19979 5480
rect 20707 5440 20747 5480
rect 22555 5440 22595 5480
rect 24940 5440 24980 5480
rect 25603 5440 25643 5480
rect 28579 5440 28619 5480
rect 28684 5440 28724 5480
rect 30412 5440 30452 5480
rect 30796 5440 30836 5480
rect 4352 5272 4720 5312
rect 12126 5272 12494 5312
rect 19900 5272 20268 5312
rect 27674 5272 28042 5312
rect 3244 5104 3284 5144
rect 3916 5104 3956 5144
rect 5740 5104 5780 5144
rect 8044 5104 8084 5144
rect 9772 5104 9812 5144
rect 10540 5104 10580 5144
rect 11011 5104 11051 5144
rect 12268 5104 12308 5144
rect 12451 5104 12491 5144
rect 14467 5104 14507 5144
rect 14764 5104 14804 5144
rect 15724 5104 15764 5144
rect 16492 5104 16532 5144
rect 17356 5104 17396 5144
rect 18412 5104 18452 5144
rect 19276 5104 19316 5144
rect 20140 5104 20180 5144
rect 20419 5104 20459 5144
rect 20716 5104 20756 5144
rect 21571 5104 21611 5144
rect 21868 5104 21908 5144
rect 22915 5104 22955 5144
rect 24172 5104 24212 5144
rect 24355 5104 24395 5144
rect 25795 5104 25835 5144
rect 26659 5104 26699 5144
rect 28012 5104 28052 5144
rect 28387 5104 28427 5144
rect 30316 5104 30356 5144
rect 30499 5104 30539 5144
rect 1708 5020 1748 5060
rect 4483 5020 4523 5060
rect 7651 5020 7691 5060
rect 7838 5020 7878 5060
rect 16684 5020 16724 5060
rect 17251 5020 17291 5060
rect 19171 5020 19211 5060
rect 28492 5020 28532 5060
rect 1612 4936 1652 4976
rect 1804 4936 1844 4976
rect 2851 4936 2891 4976
rect 2956 4936 2996 4976
rect 3436 4936 3476 4976
rect 3724 4936 3764 4976
rect 4151 4936 4191 4976
rect 4396 4936 4436 4976
rect 5347 4936 5387 4976
rect 5452 4936 5492 4976
rect 7339 4936 7379 4976
rect 7564 4936 7604 4976
rect 8140 4927 8180 4967
rect 8812 4936 8852 4976
rect 9379 4936 9419 4976
rect 9484 4936 9524 4976
rect 10147 4936 10187 4976
rect 10252 4936 10292 4976
rect 10699 4936 10739 4976
rect 10924 4936 10964 4976
rect 11875 4936 11915 4976
rect 11986 4936 12026 4976
rect 12604 4936 12644 4976
rect 12748 4936 12788 4976
rect 13175 4936 13215 4976
rect 13420 4936 13460 4976
rect 14572 4936 14612 4976
rect 15331 4936 15371 4976
rect 15436 4936 15476 4976
rect 16099 4936 16139 4976
rect 16204 4936 16244 4976
rect 16780 4936 16820 4976
rect 17011 4936 17051 4976
rect 17153 4936 17193 4976
rect 17458 4936 17498 4976
rect 18019 4936 18059 4976
rect 18124 4936 18164 4976
rect 18700 4936 18740 4976
rect 18917 4936 18957 4976
rect 19073 4936 19113 4976
rect 19372 4927 19412 4967
rect 19660 4936 19700 4976
rect 20044 4936 20084 4976
rect 20524 4936 20564 4976
rect 21676 4936 21716 4976
rect 23116 4936 23156 4976
rect 23443 4936 23483 4976
rect 23779 4936 23819 4976
rect 23884 4936 23924 4976
rect 24541 4936 24581 4976
rect 24652 4936 24692 4976
rect 25981 4936 26021 4976
rect 26092 4936 26132 4976
rect 26860 4936 26900 4976
rect 27148 4936 27188 4976
rect 27811 4936 27851 4976
rect 28108 4936 28148 4976
rect 28289 4936 28329 4976
rect 28588 4927 28628 4967
rect 29080 4936 29120 4976
rect 29356 4936 29396 4976
rect 29539 4936 29579 4976
rect 29923 4936 29963 4976
rect 30028 4936 30068 4976
rect 30652 4936 30692 4976
rect 30796 4936 30836 4976
rect 4291 4852 4331 4892
rect 7459 4852 7499 4892
rect 10819 4852 10859 4892
rect 13315 4852 13355 4892
rect 13516 4852 13556 4892
rect 16915 4843 16955 4883
rect 18604 4852 18644 4892
rect 18819 4852 18859 4892
rect 28915 4852 28955 4892
rect 7843 4684 7883 4724
rect 8956 4684 8996 4724
rect 29539 4684 29579 4724
rect 3112 4516 3480 4556
rect 10886 4516 11254 4556
rect 18660 4516 19028 4556
rect 26434 4516 26802 4556
rect 3436 4348 3476 4388
rect 7372 4348 7412 4388
rect 9100 4348 9140 4388
rect 13132 4348 13172 4388
rect 16300 4348 16340 4388
rect 18412 4348 18452 4388
rect 21676 4348 21716 4388
rect 25891 4348 25931 4388
rect 26659 4348 26699 4388
rect 27331 4348 27371 4388
rect 5068 4264 5108 4304
rect 5347 4264 5387 4304
rect 10636 4264 10676 4304
rect 21283 4264 21323 4304
rect 28204 4264 28244 4304
rect 30220 4264 30260 4304
rect 5251 4180 5291 4220
rect 5500 4180 5540 4220
rect 7843 4180 7883 4220
rect 9202 4180 9242 4220
rect 10915 4180 10955 4220
rect 17635 4180 17675 4220
rect 19666 4180 19706 4220
rect 21778 4180 21818 4220
rect 29635 4180 29675 4220
rect 30700 4180 30740 4220
rect 748 4096 788 4136
rect 931 4096 971 4136
rect 1432 4096 1472 4136
rect 1655 4096 1695 4136
rect 1795 4096 1835 4136
rect 1900 4096 1940 4136
rect 2188 4096 2228 4136
rect 2380 4096 2420 4136
rect 3340 4096 3380 4136
rect 3532 4096 3572 4136
rect 4876 4096 4916 4136
rect 5635 4096 5675 4136
rect 6220 4096 6260 4136
rect 6604 4096 6644 4136
rect 7171 4096 7211 4136
rect 7276 4096 7316 4136
rect 7703 4096 7743 4136
rect 7948 4096 7988 4136
rect 8515 4096 8555 4136
rect 9292 4096 9332 4136
rect 9964 4096 10004 4136
rect 10339 4096 10379 4136
rect 10636 4096 10676 4136
rect 10775 4096 10815 4136
rect 11020 4096 11060 4136
rect 11452 4096 11492 4136
rect 11596 4096 11636 4136
rect 12364 4096 12404 4136
rect 12506 4096 12546 4136
rect 13036 4096 13076 4136
rect 13228 4096 13268 4136
rect 14092 4096 14132 4136
rect 14476 4096 14516 4136
rect 16003 4096 16043 4136
rect 16492 4096 16532 4136
rect 16684 4096 16724 4136
rect 17515 4096 17555 4136
rect 17740 4096 17780 4136
rect 18211 4096 18251 4136
rect 18316 4096 18356 4136
rect 19756 4096 19796 4136
rect 20995 4096 21035 4136
rect 21100 4096 21140 4136
rect 21868 4096 21908 4136
rect 23500 4096 23540 4136
rect 23692 4096 23732 4136
rect 24940 4096 24980 4136
rect 25324 4096 25364 4136
rect 25875 4107 25915 4147
rect 26019 4096 26059 4136
rect 26315 4096 26355 4136
rect 26452 4096 26492 4136
rect 26956 4096 26996 4136
rect 27160 4096 27200 4136
rect 27339 4096 27379 4136
rect 27684 4096 27724 4136
rect 27820 4096 27860 4136
rect 27998 4096 28038 4136
rect 28137 4096 28177 4136
rect 28300 4096 28340 4136
rect 29356 4096 29396 4136
rect 29500 4138 29540 4178
rect 29740 4096 29780 4136
rect 30359 4096 30399 4136
rect 30499 4096 30539 4136
rect 30604 4096 30644 4136
rect 30892 4096 30932 4136
rect 31084 4096 31124 4136
rect 844 4012 884 4052
rect 2284 4012 2324 4052
rect 8826 4012 8866 4052
rect 9763 4012 9803 4052
rect 16314 4012 16354 4052
rect 16588 4012 16628 4052
rect 17827 4012 17867 4052
rect 26179 4045 26219 4085
rect 26654 4012 26694 4052
rect 29827 4012 29867 4052
rect 30988 4012 31028 4052
rect 1267 3928 1307 3968
rect 1987 3928 2027 3968
rect 4771 3928 4811 3968
rect 6700 3928 6740 3968
rect 8035 3928 8075 3968
rect 8611 3928 8651 3968
rect 8716 3928 8756 3968
rect 10051 3928 10091 3968
rect 11107 3928 11147 3968
rect 11299 3928 11339 3968
rect 12652 3928 12692 3968
rect 14572 3928 14612 3968
rect 16099 3928 16139 3968
rect 19459 3928 19499 3968
rect 23596 3928 23636 3968
rect 24835 3928 24875 3968
rect 26860 3928 26900 3968
rect 27523 3928 27563 3968
rect 28684 3928 28724 3968
rect 4352 3760 4720 3800
rect 12126 3760 12494 3800
rect 19900 3760 20268 3800
rect 27674 3760 28042 3800
rect 4876 3592 4916 3632
rect 5644 3592 5684 3632
rect 5923 3592 5963 3632
rect 7747 3592 7787 3632
rect 9868 3592 9908 3632
rect 11020 3592 11060 3632
rect 11980 3592 12020 3632
rect 12652 3592 12692 3632
rect 13315 3592 13355 3632
rect 13996 3592 14036 3632
rect 14275 3592 14315 3632
rect 16588 3592 16628 3632
rect 17356 3592 17396 3632
rect 17971 3592 18011 3632
rect 19171 3592 19211 3632
rect 19747 3592 19787 3632
rect 20515 3592 20555 3632
rect 21475 3592 21515 3632
rect 22243 3592 22283 3632
rect 22915 3592 22955 3632
rect 23683 3592 23723 3632
rect 25420 3592 25460 3632
rect 25699 3592 25739 3632
rect 25996 3592 26036 3632
rect 27820 3592 27860 3632
rect 28972 3592 29012 3632
rect 31267 3508 31307 3548
rect 1132 3424 1172 3464
rect 1795 3424 1835 3464
rect 4396 3424 4436 3464
rect 4684 3424 4724 3464
rect 5164 3424 5204 3464
rect 5548 3424 5588 3464
rect 6028 3424 6068 3464
rect 7555 3424 7595 3464
rect 9475 3424 9515 3464
rect 9580 3424 9620 3464
rect 10627 3424 10667 3464
rect 10732 3424 10772 3464
rect 11587 3424 11627 3464
rect 11692 3424 11732 3464
rect 12172 3424 12212 3464
rect 12460 3424 12500 3464
rect 13003 3424 13043 3464
rect 13228 3424 13268 3464
rect 13793 3424 13833 3464
rect 14092 3415 14132 3455
rect 14461 3424 14501 3464
rect 15312 3466 15352 3506
rect 14572 3424 14612 3464
rect 15019 3424 15059 3464
rect 15475 3424 15515 3464
rect 16108 3424 16148 3464
rect 16492 3424 16532 3464
rect 16876 3424 16916 3464
rect 17164 3424 17204 3464
rect 18136 3424 18176 3464
rect 18307 3424 18347 3464
rect 18604 3424 18644 3464
rect 19276 3424 19316 3464
rect 19852 3424 19892 3464
rect 20236 3424 20276 3464
rect 20620 3424 20660 3464
rect 21004 3424 21044 3464
rect 21676 3424 21716 3464
rect 21964 3424 22004 3464
rect 22348 3424 22388 3464
rect 22732 3424 22772 3464
rect 23212 3424 23252 3464
rect 23980 3424 24020 3464
rect 24460 3424 24500 3464
rect 24652 3424 24692 3464
rect 24940 3424 24980 3464
rect 25324 3424 25364 3464
rect 25804 3424 25844 3464
rect 27427 3424 27467 3464
rect 27532 3424 27572 3464
rect 28396 3424 28436 3464
rect 28780 3424 28820 3464
rect 30883 3424 30923 3464
rect 1276 3340 1316 3380
rect 1420 3340 1460 3380
rect 13123 3340 13163 3380
rect 15148 3340 15188 3380
rect 23122 3340 23162 3380
rect 23890 3340 23930 3380
rect 7527 3256 7567 3296
rect 15244 3256 15284 3296
rect 3340 3172 3380 3212
rect 3724 3172 3764 3212
rect 6220 3172 6260 3212
rect 13795 3172 13835 3212
rect 14467 3172 14507 3212
rect 18604 3172 18644 3212
rect 19468 3172 19508 3212
rect 24556 3172 24596 3212
rect 28156 3172 28196 3212
rect 29356 3172 29396 3212
rect 3112 3004 3480 3044
rect 10886 3004 11254 3044
rect 18660 3004 19028 3044
rect 26434 3004 26802 3044
rect 1900 2836 1940 2876
rect 3916 2836 3956 2876
rect 7363 2836 7403 2876
rect 9475 2836 9515 2876
rect 13420 2836 13460 2876
rect 18508 2836 18548 2876
rect 20236 2836 20276 2876
rect 21187 2836 21227 2876
rect 23164 2836 23204 2876
rect 24844 2836 24884 2876
rect 28771 2836 28811 2876
rect 2476 2752 2516 2792
rect 6700 2752 6740 2792
rect 22828 2752 22868 2792
rect 25564 2752 25604 2792
rect 26860 2752 26900 2792
rect 30316 2752 30356 2792
rect 1132 2668 1172 2708
rect 1347 2668 1387 2708
rect 9859 2668 9899 2708
rect 12451 2668 12491 2708
rect 12652 2668 12692 2708
rect 1228 2584 1268 2624
rect 1465 2584 1505 2624
rect 1603 2584 1643 2624
rect 1708 2584 1748 2624
rect 3052 2584 3092 2624
rect 3244 2584 3284 2624
rect 3523 2584 3563 2624
rect 4588 2584 4628 2624
rect 4894 2584 4934 2624
rect 6028 2584 6068 2624
rect 6307 2584 6347 2624
rect 6424 2617 6464 2657
rect 14956 2668 14996 2708
rect 15916 2668 15956 2708
rect 7075 2584 7115 2624
rect 7180 2584 7220 2624
rect 7660 2584 7700 2624
rect 7799 2617 7839 2657
rect 8419 2584 8459 2624
rect 8524 2584 8564 2624
rect 9187 2584 9227 2624
rect 9292 2584 9332 2624
rect 9719 2584 9759 2624
rect 9964 2584 10004 2624
rect 10732 2584 10772 2624
rect 12311 2584 12351 2624
rect 12556 2584 12596 2624
rect 13123 2584 13163 2624
rect 13434 2584 13474 2624
rect 14615 2584 14655 2624
rect 14755 2584 14795 2624
rect 14860 2584 14900 2624
rect 16012 2584 16052 2624
rect 16131 2584 16171 2624
rect 16252 2626 16292 2666
rect 17746 2668 17786 2708
rect 18610 2668 18650 2708
rect 23587 2668 23627 2708
rect 23788 2668 23828 2708
rect 16435 2584 16475 2624
rect 16538 2584 16578 2624
rect 17164 2584 17204 2624
rect 17836 2584 17876 2624
rect 18700 2584 18740 2624
rect 19939 2584 19979 2624
rect 20247 2584 20287 2624
rect 21484 2584 21524 2624
rect 21676 2584 21716 2624
rect 22540 2584 22580 2624
rect 22662 2584 22702 2624
rect 22789 2584 22829 2624
rect 23308 2584 23348 2624
rect 23467 2584 23507 2624
rect 23692 2584 23732 2624
rect 23980 2584 24020 2624
rect 24163 2584 24203 2624
rect 24364 2584 24404 2624
rect 24508 2584 24548 2624
rect 24652 2584 24692 2624
rect 25324 2584 25364 2624
rect 25420 2584 25460 2624
rect 25756 2584 25796 2624
rect 28204 2584 28244 2624
rect 28396 2584 28436 2624
rect 28588 2584 28628 2624
rect 28771 2584 28811 2624
rect 28963 2584 29003 2624
rect 29260 2584 29300 2624
rect 29443 2584 29483 2624
rect 30124 2584 30164 2624
rect 1914 2500 1954 2540
rect 4684 2500 4724 2540
rect 13228 2500 13268 2540
rect 16865 2500 16905 2540
rect 20044 2500 20084 2540
rect 21182 2500 21222 2540
rect 24076 2500 24116 2540
rect 25121 2500 25161 2540
rect 3235 2416 3275 2456
rect 4780 2416 4820 2456
rect 5068 2416 5108 2456
rect 5356 2416 5396 2456
rect 6211 2407 6251 2447
rect 7948 2416 7988 2456
rect 8812 2416 8852 2456
rect 10051 2416 10091 2456
rect 10627 2416 10667 2456
rect 10924 2416 10964 2456
rect 16684 2416 16724 2456
rect 16963 2416 17003 2456
rect 17068 2416 17108 2456
rect 17539 2416 17579 2456
rect 21388 2416 21428 2456
rect 22348 2416 22388 2456
rect 22828 2416 22868 2456
rect 25219 2416 25259 2456
rect 28300 2416 28340 2456
rect 29164 2416 29204 2456
rect 4352 2248 4720 2288
rect 12126 2248 12494 2288
rect 19900 2248 20268 2288
rect 27674 2248 28042 2288
rect 4195 2080 4235 2120
rect 5260 2080 5300 2120
rect 6796 2080 6836 2120
rect 9004 2080 9044 2120
rect 10348 2080 10388 2120
rect 10723 2080 10763 2120
rect 12268 2080 12308 2120
rect 13132 2080 13172 2120
rect 13747 2080 13787 2120
rect 13996 2080 14036 2120
rect 14275 2080 14315 2120
rect 14899 2080 14939 2120
rect 16204 2080 16244 2120
rect 18019 2080 18059 2120
rect 18604 2080 18644 2120
rect 21484 2080 21524 2120
rect 24652 2080 24692 2120
rect 28108 2080 28148 2120
rect 28579 2080 28619 2120
rect 31084 2080 31124 2120
rect 1324 1996 1364 2036
rect 1603 1996 1643 2036
rect 18234 1996 18274 2036
rect 28684 1996 28724 2036
rect 1228 1912 1268 1952
rect 1411 1912 1451 1952
rect 1987 1912 2027 1952
rect 4300 1912 4340 1952
rect 4684 1912 4724 1952
rect 5452 1912 5492 1952
rect 6412 1912 6452 1952
rect 6979 1912 7019 1952
rect 9004 1912 9044 1952
rect 9196 1912 9236 1952
rect 9868 1912 9908 1952
rect 10252 1912 10292 1952
rect 10828 1912 10868 1952
rect 11212 1912 11252 1952
rect 11788 1912 11828 1952
rect 12172 1912 12212 1952
rect 12739 1912 12779 1952
rect 12844 1912 12884 1952
rect 13324 1912 13364 1952
rect 13516 1912 13556 1952
rect 13804 1912 13844 1952
rect 14380 1912 14420 1952
rect 14764 1912 14804 1952
rect 15043 1912 15083 1952
rect 15148 1903 15188 1943
rect 16300 1912 16340 1952
rect 17923 1912 17963 1952
rect 18028 1912 18068 1952
rect 18595 1912 18635 1952
rect 18700 1912 18740 1952
rect 19555 1912 19595 1952
rect 21811 1912 21851 1952
rect 22006 1912 22046 1952
rect 22723 1912 22763 1952
rect 22827 1914 22867 1954
rect 23308 1912 23348 1952
rect 23500 1912 23540 1952
rect 24163 1912 24203 1952
rect 24460 1912 24500 1952
rect 25324 1912 25364 1952
rect 26179 1912 26219 1952
rect 28478 1912 28518 1952
rect 28780 1903 28820 1943
rect 29836 1912 29876 1952
rect 30124 1912 30164 1952
rect 30988 1912 31028 1952
rect 31180 1912 31220 1952
rect 3532 1828 3572 1868
rect 19180 1828 19220 1868
rect 25804 1828 25844 1868
rect 27724 1828 27764 1868
rect 29155 1828 29195 1868
rect 3916 1744 3956 1784
rect 7024 1744 7064 1784
rect 7564 1744 7604 1784
rect 15436 1744 15476 1784
rect 16780 1744 16820 1784
rect 21100 1744 21140 1784
rect 23011 1744 23051 1784
rect 23788 1744 23828 1784
rect 24460 1744 24500 1784
rect 5059 1660 5099 1700
rect 5740 1660 5780 1700
rect 13420 1660 13460 1700
rect 18220 1660 18260 1700
rect 18892 1660 18932 1700
rect 23308 1660 23348 1700
rect 30796 1660 30836 1700
rect 3112 1492 3480 1532
rect 10886 1492 11254 1532
rect 18660 1492 19028 1532
rect 26434 1492 26802 1532
rect 8428 1324 8468 1364
rect 10348 1324 10388 1364
rect 11212 1324 11252 1364
rect 12844 1324 12884 1364
rect 17644 1324 17684 1364
rect 25228 1324 25268 1364
rect 28492 1324 28532 1364
rect 2668 1240 2708 1280
rect 4387 1240 4427 1280
rect 4828 1240 4868 1280
rect 10540 1240 10580 1280
rect 18988 1240 19028 1280
rect 20908 1240 20948 1280
rect 21676 1240 21716 1280
rect 25036 1240 25076 1280
rect 5059 1156 5099 1196
rect 6508 1156 6548 1196
rect 24652 1156 24692 1196
rect 26851 1156 26891 1196
rect 30787 1156 30827 1196
rect 4204 1072 4244 1112
rect 4387 1072 4427 1112
rect 4684 1072 4724 1112
rect 4919 1072 4959 1112
rect 5165 1072 5205 1112
rect 5443 1072 5483 1112
rect 5923 1105 5963 1145
rect 6883 1072 6923 1112
rect 9196 1072 9236 1112
rect 9868 1072 9908 1112
rect 10147 1072 10187 1112
rect 10915 1072 10955 1112
rect 11392 1072 11432 1112
rect 11548 1072 11588 1112
rect 12643 1072 12683 1112
rect 12748 1072 12788 1112
rect 13175 1072 13215 1112
rect 13315 1072 13355 1112
rect 13420 1072 13460 1112
rect 14284 1072 14324 1112
rect 14467 1072 14507 1112
rect 14812 1072 14852 1112
rect 14956 1072 14996 1112
rect 16099 1072 16139 1112
rect 18796 1072 18836 1112
rect 18911 1072 18951 1112
rect 19084 1072 19124 1112
rect 20044 1072 20084 1112
rect 20716 1072 20756 1112
rect 21475 1072 21515 1112
rect 23107 1072 23147 1112
rect 25852 1072 25892 1112
rect 26092 1072 26132 1112
rect 26284 1072 26324 1112
rect 27532 1072 27572 1112
rect 30403 1072 30443 1112
rect 5644 988 5684 1028
rect 5754 988 5794 1028
rect 11020 988 11060 1028
rect 11226 988 11266 1028
rect 13507 988 13547 1028
rect 15715 988 15755 1028
rect 22723 988 22763 1028
rect 26188 988 26228 1028
rect 5251 904 5291 944
rect 5539 904 5579 944
rect 6076 904 6116 944
rect 8812 904 8852 944
rect 13036 904 13076 944
rect 14380 904 14420 944
rect 14659 904 14699 944
rect 18028 904 18068 944
rect 21676 904 21716 944
rect 4352 736 4720 776
rect 12126 736 12494 776
rect 19900 736 20268 776
rect 27674 736 28042 776
<< metal2 >>
rect 16387 28624 16396 28664
rect 16436 28624 30068 28664
rect 30028 28580 30068 28624
rect 13891 28540 13900 28580
rect 13940 28540 23308 28580
rect 23348 28540 23357 28580
rect 30019 28540 30028 28580
rect 30068 28540 30077 28580
rect 12355 28372 12364 28412
rect 12404 28372 17644 28412
rect 17684 28372 17693 28412
rect 10051 28204 10060 28244
rect 10100 28204 20428 28244
rect 20468 28204 20477 28244
rect 14659 28120 14668 28160
rect 14708 28120 21388 28160
rect 21428 28120 21437 28160
rect 15427 28036 15436 28076
rect 15476 28036 20524 28076
rect 20564 28036 20573 28076
rect 4343 27952 4352 27992
rect 4720 27952 4729 27992
rect 12117 27952 12126 27992
rect 12494 27952 12503 27992
rect 19891 27952 19900 27992
rect 20268 27952 20277 27992
rect 27665 27952 27674 27992
rect 28042 27952 28051 27992
rect 9283 27868 9292 27908
rect 9332 27868 11788 27908
rect 11828 27868 11837 27908
rect 16195 27868 16204 27908
rect 16244 27868 21100 27908
rect 21140 27868 21149 27908
rect 11587 27784 11596 27824
rect 11636 27784 17836 27824
rect 17876 27784 17885 27824
rect 24172 27784 25940 27824
rect 29251 27784 29260 27824
rect 29300 27784 30932 27824
rect 3628 27700 8524 27740
rect 8564 27700 8660 27740
rect 11194 27700 11203 27740
rect 11243 27700 11692 27740
rect 11732 27700 11741 27740
rect 16396 27700 18164 27740
rect 22330 27700 22339 27740
rect 22379 27700 23980 27740
rect 24020 27700 24029 27740
rect 3628 27656 3668 27700
rect 6124 27656 6164 27700
rect 8620 27656 8660 27700
rect 16396 27656 16436 27700
rect 18124 27656 18164 27700
rect 24172 27656 24212 27784
rect 25114 27700 25123 27740
rect 25163 27700 25507 27740
rect 25547 27700 25556 27740
rect 25900 27656 25940 27784
rect 26947 27700 26956 27740
rect 26996 27700 28148 27740
rect 28483 27700 28492 27740
rect 28532 27700 29876 27740
rect 28108 27656 28148 27700
rect 29836 27656 29876 27700
rect 3610 27616 3619 27656
rect 3668 27616 3799 27656
rect 6106 27616 6115 27656
rect 6155 27616 6164 27656
rect 8602 27616 8611 27656
rect 8651 27616 8660 27656
rect 11578 27616 11587 27656
rect 11636 27616 11767 27656
rect 14179 27616 14188 27656
rect 14228 27616 15148 27656
rect 15188 27616 15197 27656
rect 16378 27616 16387 27656
rect 16427 27616 16436 27656
rect 16937 27616 17068 27656
rect 17108 27616 17117 27656
rect 18106 27616 18115 27656
rect 18155 27616 19084 27656
rect 19124 27616 20140 27656
rect 20180 27616 20189 27656
rect 22714 27616 22723 27656
rect 22772 27616 24212 27656
rect 25027 27616 25036 27656
rect 25076 27616 25085 27656
rect 25210 27616 25219 27656
rect 25259 27616 25268 27656
rect 25315 27616 25324 27656
rect 25364 27616 25612 27656
rect 25652 27616 25661 27656
rect 25882 27616 25891 27656
rect 25940 27616 26071 27656
rect 27916 27616 28012 27656
rect 28052 27616 28061 27656
rect 28108 27647 28916 27656
rect 28108 27616 28867 27647
rect 3235 27532 3244 27572
rect 3284 27532 3293 27572
rect 3523 27532 3532 27572
rect 3572 27532 3581 27572
rect 5609 27532 5740 27572
rect 5780 27532 5789 27572
rect 6691 27532 6700 27572
rect 6740 27532 6749 27572
rect 8105 27532 8236 27572
rect 8276 27532 8285 27572
rect 9283 27532 9292 27572
rect 9332 27532 9341 27572
rect 3017 27448 3052 27488
rect 3092 27448 3148 27488
rect 3188 27448 3197 27488
rect 3244 27404 3284 27532
rect 12844 27488 12884 27552
rect 15715 27532 15724 27572
rect 15764 27532 15773 27572
rect 16762 27532 16771 27572
rect 16820 27532 16951 27572
rect 17609 27532 17740 27572
rect 17780 27532 17789 27572
rect 19372 27488 19412 27552
rect 24000 27532 24460 27572
rect 24500 27532 24509 27572
rect 25036 27488 25076 27616
rect 12844 27448 13708 27488
rect 13748 27448 13757 27488
rect 19372 27448 20236 27488
rect 20276 27448 20285 27488
rect 20681 27448 20812 27488
rect 20852 27448 20861 27488
rect 24460 27448 25076 27488
rect 25228 27488 25268 27616
rect 27168 27532 27820 27572
rect 27860 27532 27869 27572
rect 27916 27488 27956 27616
rect 28858 27607 28867 27616
rect 28907 27607 28916 27647
rect 29225 27647 29356 27656
rect 29225 27616 29347 27647
rect 29396 27616 29405 27656
rect 29818 27647 29876 27656
rect 28858 27606 28916 27607
rect 29338 27607 29347 27616
rect 29387 27607 29396 27616
rect 29338 27606 29396 27607
rect 29818 27607 29827 27647
rect 29867 27607 29876 27647
rect 29818 27606 29876 27607
rect 30892 27572 30932 27784
rect 28963 27532 28972 27572
rect 29012 27532 29020 27572
rect 29060 27532 29143 27572
rect 29443 27532 29452 27572
rect 29492 27532 29500 27572
rect 29540 27532 29623 27572
rect 29923 27532 29932 27572
rect 29972 27532 29980 27572
rect 30020 27532 30103 27572
rect 30883 27532 30892 27572
rect 30932 27532 30941 27572
rect 25228 27448 25652 27488
rect 3244 27364 3724 27404
rect 3764 27364 3773 27404
rect 5539 27364 5548 27404
rect 5588 27364 7468 27404
rect 7508 27364 7517 27404
rect 8035 27364 8044 27404
rect 8084 27364 9676 27404
rect 9716 27364 9725 27404
rect 10409 27364 10540 27404
rect 10580 27364 10589 27404
rect 13315 27364 13324 27404
rect 13364 27364 13516 27404
rect 13556 27364 13565 27404
rect 13795 27364 13804 27404
rect 13844 27364 14044 27404
rect 14084 27364 14093 27404
rect 14345 27364 14476 27404
rect 14516 27364 14525 27404
rect 14659 27364 14668 27404
rect 14708 27364 16924 27404
rect 16964 27364 16973 27404
rect 19651 27364 19660 27404
rect 19700 27364 20044 27404
rect 20084 27364 20093 27404
rect 24460 27320 24500 27448
rect 25612 27404 25652 27448
rect 27820 27448 27956 27488
rect 30185 27448 30316 27488
rect 30356 27448 30365 27488
rect 30953 27448 31084 27488
rect 31124 27448 31133 27488
rect 27820 27404 27860 27448
rect 24643 27364 24652 27404
rect 24692 27364 25516 27404
rect 25556 27364 25565 27404
rect 25612 27364 26132 27404
rect 27139 27364 27148 27404
rect 27188 27364 27820 27404
rect 27860 27364 27869 27404
rect 28553 27364 28684 27404
rect 28724 27364 28733 27404
rect 30403 27364 30412 27404
rect 30452 27364 30652 27404
rect 30692 27364 30701 27404
rect 20899 27280 20908 27320
rect 20948 27280 24500 27320
rect 3103 27196 3112 27236
rect 3480 27196 3489 27236
rect 10877 27196 10886 27236
rect 11254 27196 11263 27236
rect 18651 27196 18660 27236
rect 19028 27196 19037 27236
rect 8707 27112 8716 27152
rect 8756 27112 18068 27152
rect 18115 27112 18124 27152
rect 18164 27112 24940 27152
rect 24980 27112 24989 27152
rect 18028 27068 18068 27112
rect 26092 27068 26132 27364
rect 26425 27196 26434 27236
rect 26802 27196 26811 27236
rect 3148 27028 3916 27068
rect 3956 27028 3965 27068
rect 11561 27028 11692 27068
rect 11732 27028 11741 27068
rect 14074 27028 14083 27068
rect 14123 27028 14132 27068
rect 16771 27028 16780 27068
rect 16820 27028 17068 27068
rect 17108 27028 17117 27068
rect 17731 27028 17740 27068
rect 17780 27028 17932 27068
rect 17972 27028 17981 27068
rect 18028 27028 20716 27068
rect 20756 27028 20765 27068
rect 26092 27028 26851 27068
rect 26891 27028 26900 27068
rect 26947 27028 26956 27068
rect 26996 27028 30796 27068
rect 30836 27028 30845 27068
rect 3148 26984 3188 27028
rect 14092 26984 14132 27028
rect 2755 26944 2764 26984
rect 2804 26944 2813 26984
rect 3139 26944 3148 26984
rect 3188 26944 3197 26984
rect 3401 26944 3532 26984
rect 3572 26944 3581 26984
rect 3715 26944 3724 26984
rect 3764 26944 3895 26984
rect 5417 26944 5452 26984
rect 5492 26944 5548 26984
rect 5588 26944 5597 26984
rect 6569 26944 6700 26984
rect 6740 26944 6749 26984
rect 9161 26944 9292 26984
rect 9332 26944 9341 26984
rect 10348 26944 11884 26984
rect 11924 26944 11933 26984
rect 12556 26944 13324 26984
rect 13364 26944 13373 26984
rect 13577 26944 13708 26984
rect 13748 26944 13757 26984
rect 14092 26944 14516 26984
rect 15593 26944 15724 26984
rect 15764 26944 15773 26984
rect 17731 26944 17740 26984
rect 17780 26944 17789 26984
rect 24329 26944 24460 26984
rect 24500 26944 24509 26984
rect 26179 26944 26188 26984
rect 26228 26944 27284 26984
rect 27689 26944 27820 26984
rect 27860 26944 27869 26984
rect 2764 26040 2804 26944
rect 10348 26900 10388 26944
rect 8393 26860 8476 26900
rect 8516 26860 8524 26900
rect 8564 26860 8573 26900
rect 10252 26860 10388 26900
rect 10697 26860 10828 26900
rect 10868 26860 12460 26900
rect 12500 26860 12509 26900
rect 10252 26816 10292 26860
rect 10828 26816 10868 26860
rect 12556 26816 12596 26944
rect 14380 26816 14420 26825
rect 14476 26816 14516 26944
rect 15235 26860 15244 26900
rect 15284 26860 16780 26900
rect 16820 26860 16829 26900
rect 17740 26816 17780 26944
rect 19468 26860 19660 26900
rect 19700 26860 19709 26900
rect 20803 26860 20812 26900
rect 20852 26860 20861 26900
rect 23107 26860 23116 26900
rect 23156 26860 23308 26900
rect 23348 26860 23357 26900
rect 23788 26860 24835 26900
rect 24875 26860 24884 26900
rect 24940 26860 27188 26900
rect 19468 26816 19508 26860
rect 23788 26816 23828 26860
rect 24940 26816 24980 26860
rect 25900 26816 25940 26860
rect 27148 26816 27188 26860
rect 3715 26776 3724 26816
rect 3764 26776 3773 26816
rect 3907 26776 3916 26816
rect 3956 26776 4876 26816
rect 4916 26776 4925 26816
rect 6185 26776 6316 26816
rect 6356 26776 6365 26816
rect 7337 26776 7468 26816
rect 7508 26776 7517 26816
rect 8311 26776 8320 26816
rect 8360 26776 10100 26816
rect 10243 26776 10252 26816
rect 10292 26776 10301 26816
rect 10387 26776 10396 26816
rect 10436 26776 10732 26816
rect 10772 26776 10781 26816
rect 11011 26776 11020 26816
rect 11060 26776 11069 26816
rect 12547 26776 12556 26816
rect 12596 26776 12605 26816
rect 12739 26776 12748 26816
rect 12788 26776 12919 26816
rect 14249 26776 14380 26816
rect 14420 26776 14429 26816
rect 14476 26776 14572 26816
rect 14612 26776 14621 26816
rect 16073 26776 16108 26816
rect 16148 26776 16204 26816
rect 16244 26776 16253 26816
rect 16937 26776 17068 26816
rect 17108 26776 17117 26816
rect 17338 26776 17347 26816
rect 17387 26776 17396 26816
rect 17740 26776 18604 26816
rect 18644 26776 18653 26816
rect 19459 26776 19468 26816
rect 19508 26776 19517 26816
rect 19564 26776 19892 26816
rect 20122 26776 20131 26816
rect 20180 26776 20311 26816
rect 23788 26776 23800 26816
rect 23840 26776 23849 26816
rect 23959 26776 23968 26816
rect 24008 26776 24020 26816
rect 24163 26776 24172 26816
rect 24212 26776 24980 26816
rect 25385 26776 25516 26816
rect 25556 26776 25565 26816
rect 25891 26776 25900 26816
rect 25940 26776 25949 26816
rect 25996 26776 26021 26816
rect 26061 26776 26083 26816
rect 26275 26776 26284 26816
rect 26363 26776 26455 26816
rect 26921 26776 27052 26816
rect 27092 26776 27101 26816
rect 27244 26816 27284 26944
rect 27427 26860 27436 26900
rect 27476 26860 28780 26900
rect 28820 26860 28963 26900
rect 29003 26860 29012 26900
rect 31075 26860 31084 26900
rect 31124 26860 31133 26900
rect 27244 26776 27283 26816
rect 27323 26776 27332 26816
rect 27619 26776 27628 26816
rect 27668 26776 28387 26816
rect 28427 26776 28436 26816
rect 28483 26776 28492 26816
rect 28532 26776 28663 26816
rect 30761 26776 30883 26816
rect 30932 26776 30941 26816
rect 3724 26564 3764 26776
rect 4300 26692 4780 26732
rect 4820 26692 4829 26732
rect 4972 26692 5452 26732
rect 5492 26692 5501 26732
rect 5548 26692 6220 26732
rect 6260 26692 6269 26732
rect 8131 26692 8140 26732
rect 8180 26692 9196 26732
rect 9236 26692 9245 26732
rect 4300 26648 4340 26692
rect 4972 26648 5012 26692
rect 5548 26648 5588 26692
rect 4291 26608 4300 26648
rect 4340 26608 4349 26648
rect 4675 26608 4684 26648
rect 4724 26608 5012 26648
rect 5059 26608 5068 26648
rect 5108 26608 5588 26648
rect 5635 26608 5644 26648
rect 5684 26608 5693 26648
rect 7267 26608 7276 26648
rect 7316 26608 7756 26648
rect 7796 26608 7805 26648
rect 8611 26608 8620 26648
rect 8660 26608 8812 26648
rect 8852 26608 8861 26648
rect 3724 26524 4780 26564
rect 4820 26524 4829 26564
rect 4343 26440 4352 26480
rect 4720 26440 4729 26480
rect 4714 26272 4723 26312
rect 4763 26272 5108 26312
rect 3715 26188 3724 26228
rect 3764 26188 3956 26228
rect 3916 26144 3956 26188
rect 5068 26144 5108 26272
rect 5644 26228 5684 26608
rect 10060 26396 10100 26776
rect 10828 26767 10868 26776
rect 10243 26692 10252 26732
rect 10292 26692 10526 26732
rect 10566 26692 10575 26732
rect 11020 26648 11060 26776
rect 14380 26767 14420 26776
rect 10618 26608 10627 26648
rect 10667 26608 11060 26648
rect 11116 26692 14078 26732
rect 14118 26692 14127 26732
rect 11116 26564 11156 26692
rect 12835 26608 12844 26648
rect 12884 26608 13420 26648
rect 13460 26608 13469 26648
rect 14275 26608 14284 26648
rect 14324 26608 14668 26648
rect 14708 26608 14717 26648
rect 17356 26564 17396 26776
rect 17443 26692 17452 26732
rect 17492 26692 18787 26732
rect 18827 26692 18836 26732
rect 10435 26524 10444 26564
rect 10484 26524 11156 26564
rect 11395 26524 11404 26564
rect 11444 26524 17396 26564
rect 19564 26480 19604 26776
rect 19852 26732 19892 26776
rect 23980 26732 24020 26776
rect 25996 26732 26036 26776
rect 27148 26732 27188 26776
rect 19738 26692 19747 26732
rect 19787 26692 19796 26732
rect 19852 26692 23788 26732
rect 23828 26692 23837 26732
rect 23884 26692 24020 26732
rect 25577 26692 25699 26732
rect 25748 26692 25757 26732
rect 25987 26692 25996 26732
rect 26036 26692 26045 26732
rect 26284 26692 26846 26732
rect 26886 26692 26895 26732
rect 27148 26692 27532 26732
rect 27572 26692 27581 26732
rect 31258 26692 31267 26732
rect 31307 26692 31316 26732
rect 12117 26440 12126 26480
rect 12494 26440 12503 26480
rect 12931 26440 12940 26480
rect 12980 26440 13804 26480
rect 13844 26440 13853 26480
rect 16099 26440 16108 26480
rect 16148 26440 19604 26480
rect 10060 26356 11980 26396
rect 12020 26356 16972 26396
rect 17012 26356 17021 26396
rect 17155 26356 17164 26396
rect 17204 26356 18892 26396
rect 18932 26356 19276 26396
rect 19316 26356 19325 26396
rect 19756 26312 19796 26692
rect 23884 26648 23924 26692
rect 22051 26608 22060 26648
rect 22100 26608 22109 26648
rect 23059 26608 23068 26648
rect 23108 26608 23116 26648
rect 23156 26608 23239 26648
rect 23587 26608 23596 26648
rect 23675 26608 23924 26648
rect 24067 26608 24076 26648
rect 24116 26608 24124 26648
rect 24164 26608 24247 26648
rect 25993 26608 26002 26648
rect 26042 26608 26051 26648
rect 19891 26440 19900 26480
rect 20268 26440 20277 26480
rect 22060 26312 22100 26608
rect 25996 26564 26036 26608
rect 26284 26564 26324 26692
rect 26515 26608 26524 26648
rect 26564 26608 26573 26648
rect 27331 26608 27340 26648
rect 27380 26608 27484 26648
rect 27524 26608 27533 26648
rect 28771 26608 28780 26648
rect 28820 26608 28829 26648
rect 25603 26524 25612 26564
rect 25652 26524 26324 26564
rect 26524 26480 26564 26608
rect 23395 26440 23404 26480
rect 23444 26440 26564 26480
rect 27665 26440 27674 26480
rect 28042 26440 28051 26480
rect 7939 26272 7948 26312
rect 7988 26272 7997 26312
rect 8227 26272 8236 26312
rect 8276 26272 8284 26312
rect 8324 26272 8407 26312
rect 8585 26272 8716 26312
rect 8756 26272 8765 26312
rect 9545 26272 9667 26312
rect 9716 26272 9725 26312
rect 9955 26272 9964 26312
rect 10004 26272 10013 26312
rect 10147 26272 10156 26312
rect 10196 26272 10484 26312
rect 11273 26272 11395 26312
rect 11444 26272 11453 26312
rect 11587 26272 11596 26312
rect 11636 26272 11923 26312
rect 11963 26272 13172 26312
rect 15017 26272 15148 26312
rect 15188 26272 16916 26312
rect 17321 26272 17443 26312
rect 17492 26272 17501 26312
rect 17993 26272 18115 26312
rect 18164 26272 18173 26312
rect 18787 26272 18796 26312
rect 18836 26272 19564 26312
rect 19604 26272 19613 26312
rect 19747 26272 19756 26312
rect 19796 26272 19805 26312
rect 19939 26272 19948 26312
rect 19988 26272 22100 26312
rect 23849 26272 23971 26312
rect 24020 26272 24029 26312
rect 26083 26272 26092 26312
rect 26132 26272 26188 26312
rect 26228 26272 26263 26312
rect 7948 26228 7988 26272
rect 9964 26228 10004 26272
rect 10444 26228 10484 26272
rect 5155 26188 5164 26228
rect 5204 26188 5396 26228
rect 5626 26188 5635 26228
rect 5675 26188 5684 26228
rect 5827 26188 5836 26228
rect 5876 26188 6356 26228
rect 7948 26188 8756 26228
rect 5356 26144 5396 26188
rect 6316 26144 6356 26188
rect 8716 26144 8756 26188
rect 9057 26188 9100 26228
rect 9140 26188 9149 26228
rect 9964 26188 10314 26228
rect 9057 26144 9097 26188
rect 10274 26146 10314 26188
rect 10426 26219 10484 26228
rect 10426 26179 10435 26219
rect 10475 26179 10484 26219
rect 10426 26178 10484 26179
rect 10540 26188 11884 26228
rect 11924 26188 11933 26228
rect 12268 26188 12556 26228
rect 12596 26188 12605 26228
rect 12713 26188 12835 26228
rect 12884 26188 12893 26228
rect 3497 26104 3619 26144
rect 3668 26104 3677 26144
rect 3916 26135 4520 26144
rect 3916 26104 4480 26135
rect 4570 26104 4579 26144
rect 4619 26104 4628 26144
rect 4937 26104 5068 26144
rect 5108 26104 5117 26144
rect 5164 26104 5260 26144
rect 5300 26104 5309 26144
rect 5356 26104 5740 26144
rect 5780 26104 5789 26144
rect 6010 26104 6019 26144
rect 6059 26104 6220 26144
rect 6260 26104 6269 26144
rect 6316 26104 8140 26144
rect 8180 26104 8189 26144
rect 8294 26104 8332 26144
rect 8372 26104 8425 26144
rect 8465 26104 8474 26144
rect 8542 26137 8551 26144
rect 8524 26104 8551 26137
rect 8591 26104 8600 26144
rect 8668 26104 8677 26144
rect 8717 26104 8756 26144
rect 8899 26104 8908 26144
rect 8948 26104 8957 26144
rect 9039 26104 9048 26144
rect 9088 26104 9097 26144
rect 9148 26104 9157 26144
rect 9236 26104 9337 26144
rect 9763 26104 9772 26144
rect 9812 26104 9964 26144
rect 10004 26104 10013 26144
rect 10138 26104 10147 26144
rect 10187 26104 10196 26144
rect 4480 26086 4520 26095
rect 4588 26060 4628 26104
rect 5164 26060 5204 26104
rect 8524 26097 8599 26104
rect 8686 26097 8756 26104
rect 8524 26060 8564 26097
rect 8908 26060 8948 26104
rect 10156 26060 10196 26104
rect 10252 26135 10314 26146
rect 10540 26144 10580 26188
rect 12268 26144 12308 26188
rect 13132 26144 13172 26272
rect 15523 26188 15532 26228
rect 15572 26188 16820 26228
rect 16780 26144 16820 26188
rect 16876 26144 16916 26272
rect 17347 26188 17356 26228
rect 17396 26188 18590 26228
rect 18630 26188 18639 26228
rect 18682 26188 18691 26228
rect 18731 26188 20468 26228
rect 20428 26144 20468 26188
rect 22060 26144 22100 26272
rect 28780 26228 28820 26608
rect 31276 26312 31316 26692
rect 30499 26272 30508 26312
rect 30548 26272 31316 26312
rect 23945 26188 24076 26228
rect 24116 26188 24748 26228
rect 24788 26188 25996 26228
rect 26036 26188 26284 26228
rect 26324 26188 27052 26228
rect 27092 26188 27293 26228
rect 26845 26144 26885 26188
rect 27253 26144 27293 26188
rect 10292 26106 10314 26135
rect 10522 26104 10531 26144
rect 10571 26104 10580 26144
rect 10627 26104 10636 26144
rect 10705 26104 10807 26144
rect 11177 26104 11308 26144
rect 11348 26104 11357 26144
rect 11971 26104 11980 26144
rect 12020 26104 12088 26144
rect 12128 26104 12151 26144
rect 12228 26104 12237 26144
rect 12277 26104 12308 26144
rect 12390 26104 12399 26144
rect 12439 26104 12460 26144
rect 12500 26104 12570 26144
rect 12643 26104 12652 26144
rect 12731 26104 12940 26144
rect 12980 26104 12989 26144
rect 13132 26104 13219 26144
rect 13259 26104 13268 26144
rect 14467 26104 14476 26144
rect 14516 26104 15436 26144
rect 15476 26104 15485 26144
rect 15619 26104 15628 26144
rect 15668 26104 15820 26144
rect 15860 26104 15869 26144
rect 15994 26104 16003 26144
rect 16043 26104 16052 26144
rect 16099 26104 16108 26144
rect 16148 26104 16279 26144
rect 16457 26104 16555 26144
rect 16628 26104 16637 26144
rect 16771 26104 16780 26144
rect 16820 26104 16829 26144
rect 16876 26104 17548 26144
rect 17588 26104 17597 26144
rect 17897 26104 17932 26144
rect 17972 26104 18028 26144
rect 18068 26104 18077 26144
rect 18211 26104 18220 26144
rect 18260 26104 18269 26144
rect 18761 26104 18892 26144
rect 18932 26104 18941 26144
rect 18988 26104 19070 26144
rect 19110 26104 19119 26144
rect 19267 26104 19276 26144
rect 19316 26104 19325 26144
rect 19372 26135 19468 26144
rect 10252 26086 10292 26095
rect 3994 26020 4003 26060
rect 4043 26020 4244 26060
rect 4588 26020 5164 26060
rect 5204 26020 5213 26060
rect 5539 26020 5548 26060
rect 5588 26020 5856 26060
rect 8476 26020 8564 26060
rect 8870 26020 8908 26060
rect 8948 26020 8957 26060
rect 9283 26020 9292 26060
rect 9332 26020 10196 26060
rect 4204 25976 4244 26020
rect 1699 25936 1708 25976
rect 1748 25936 2324 25976
rect 4186 25936 4195 25976
rect 4235 25936 4244 25976
rect 8476 25976 8516 26020
rect 10156 25976 10196 26020
rect 11020 26062 11068 26102
rect 11108 26062 11117 26102
rect 11020 25976 11060 26062
rect 15436 26060 15476 26104
rect 16012 26060 16052 26104
rect 17548 26060 17588 26104
rect 18220 26060 18260 26104
rect 18892 26086 18932 26095
rect 11194 26020 11203 26060
rect 11243 26020 11500 26060
rect 11540 26020 11549 26060
rect 12550 26020 12559 26060
rect 12599 26020 12844 26060
rect 12884 26020 12893 26060
rect 13699 26020 13708 26060
rect 13748 26020 13757 26060
rect 15436 26020 16204 26060
rect 16244 26020 16253 26060
rect 16666 26020 16675 26060
rect 16715 26020 16724 26060
rect 16867 26020 16876 26060
rect 16916 26020 16925 26060
rect 17548 26020 18260 26060
rect 16684 25976 16724 26020
rect 8476 25936 9004 25976
rect 9044 25936 9053 25976
rect 9187 25936 9196 25976
rect 9236 25936 10060 25976
rect 10100 25936 10109 25976
rect 10156 25936 10828 25976
rect 10868 25936 10877 25976
rect 11020 25936 11444 25976
rect 12451 25936 12460 25976
rect 12500 25936 12748 25976
rect 12788 25936 12797 25976
rect 15052 25936 15284 25976
rect 16282 25936 16291 25976
rect 16331 25936 16492 25976
rect 16532 25936 16724 25976
rect 16876 25976 16916 26020
rect 18988 25976 19028 26104
rect 16876 25936 17548 25976
rect 17588 25936 17597 25976
rect 18019 25936 18028 25976
rect 18068 25936 18412 25976
rect 18452 25936 19028 25976
rect 19276 25976 19316 26104
rect 19412 26104 19468 26135
rect 19508 26104 19948 26144
rect 19988 26104 19997 26144
rect 20419 26104 20428 26144
rect 20468 26104 20477 26144
rect 20585 26104 20716 26144
rect 20756 26104 20765 26144
rect 20944 26104 20953 26144
rect 20993 26104 21004 26144
rect 21044 26104 21133 26144
rect 21763 26104 21772 26144
rect 21812 26104 22100 26144
rect 23753 26104 23873 26144
rect 23924 26104 23933 26144
rect 24041 26104 24172 26144
rect 24212 26104 24221 26144
rect 24643 26104 24652 26144
rect 24692 26135 24823 26144
rect 24692 26104 24739 26135
rect 19372 26086 19412 26095
rect 24172 26086 24212 26095
rect 24730 26095 24739 26104
rect 24779 26104 24823 26135
rect 25411 26104 25420 26144
rect 25460 26135 25591 26144
rect 25460 26104 25507 26135
rect 24779 26095 24788 26104
rect 24730 26094 24788 26095
rect 25498 26095 25507 26104
rect 25547 26104 25591 26135
rect 25900 26104 25996 26144
rect 26036 26104 26045 26144
rect 26170 26104 26179 26144
rect 26219 26104 26228 26144
rect 26845 26104 26872 26144
rect 26912 26104 26921 26144
rect 27048 26104 27057 26144
rect 27097 26111 27106 26144
rect 27097 26104 27158 26111
rect 27235 26104 27244 26144
rect 27284 26104 27293 26144
rect 27375 26188 27859 26228
rect 27899 26188 27908 26228
rect 28108 26188 28684 26228
rect 28724 26188 28733 26228
rect 28780 26188 30452 26228
rect 25547 26095 25556 26104
rect 25498 26094 25556 26095
rect 20489 26020 20620 26060
rect 20660 26020 20669 26060
rect 20803 26020 20812 26060
rect 20875 26020 20983 26060
rect 24835 26020 24844 26060
rect 24884 26020 24892 26060
rect 24932 26020 25015 26060
rect 25651 26020 25660 26060
rect 25700 26020 25708 26060
rect 25748 26020 25831 26060
rect 25900 25976 25940 26104
rect 26188 26060 26228 26104
rect 27052 26071 27158 26104
rect 27375 26102 27415 26188
rect 28108 26144 28148 26188
rect 30412 26144 30452 26188
rect 27484 26104 27493 26144
rect 27533 26104 27628 26144
rect 27668 26104 27677 26144
rect 28045 26104 28054 26144
rect 28094 26104 28148 26144
rect 28195 26104 28204 26144
rect 28244 26104 28253 26144
rect 28299 26104 28387 26144
rect 28427 26104 28436 26144
rect 28483 26104 28492 26144
rect 28532 26104 28819 26144
rect 28859 26104 28868 26144
rect 29005 26104 29014 26144
rect 29054 26104 29155 26144
rect 29195 26104 29204 26144
rect 29260 26104 29836 26144
rect 29876 26104 29885 26144
rect 30403 26104 30412 26144
rect 30452 26104 30461 26144
rect 30595 26104 30604 26144
rect 30644 26104 31180 26144
rect 31220 26104 31229 26144
rect 27118 26060 27158 26071
rect 27357 26062 27366 26102
rect 27406 26062 27415 26102
rect 26083 26020 26092 26060
rect 26132 26020 26228 26060
rect 26659 26020 26668 26060
rect 26708 26020 26956 26060
rect 26996 26020 27005 26060
rect 27118 26020 27148 26060
rect 27188 26020 27197 26060
rect 27375 25976 27415 26062
rect 28204 26060 28244 26104
rect 28003 26020 28012 26060
rect 28052 26020 28244 26060
rect 28299 25976 28339 26104
rect 29260 25976 29300 26104
rect 30857 26020 30988 26060
rect 31028 26020 31037 26060
rect 19276 25936 19852 25976
rect 19892 25936 19901 25976
rect 22121 25936 22252 25976
rect 22292 25936 22301 25976
rect 24931 25936 24940 25976
rect 24980 25936 25940 25976
rect 25987 25936 25996 25976
rect 26036 25936 26428 25976
rect 26468 25936 26477 25976
rect 27235 25936 27244 25976
rect 27284 25936 27415 25976
rect 27523 25936 27532 25976
rect 27572 25936 27820 25976
rect 27860 25936 28339 25976
rect 28771 25936 28780 25976
rect 28820 25936 29300 25976
rect 29897 25936 30028 25976
rect 30068 25936 30077 25976
rect 30739 25936 30748 25976
rect 30788 25936 31084 25976
rect 31124 25936 31133 25976
rect 2284 25892 2324 25936
rect 11404 25892 11444 25936
rect 15052 25892 15092 25936
rect 2284 25852 8140 25892
rect 8180 25852 8189 25892
rect 10138 25852 10147 25892
rect 10187 25852 10444 25892
rect 10484 25852 10493 25892
rect 11395 25852 11404 25892
rect 11444 25852 11453 25892
rect 11971 25852 11980 25892
rect 12020 25852 15092 25892
rect 15244 25892 15284 25936
rect 15244 25852 18068 25892
rect 19066 25852 19075 25892
rect 19115 25852 19372 25892
rect 19412 25852 19421 25892
rect 20131 25852 20140 25892
rect 20180 25852 21100 25892
rect 21140 25852 21149 25892
rect 21196 25852 26036 25892
rect 26729 25852 26860 25892
rect 26900 25852 26909 25892
rect 28265 25852 28387 25892
rect 28436 25852 28445 25892
rect 18028 25808 18068 25852
rect 21196 25808 21236 25852
rect 4195 25768 4204 25808
rect 4244 25768 10100 25808
rect 11683 25768 11692 25808
rect 11732 25768 17972 25808
rect 18028 25768 19124 25808
rect 19171 25768 19180 25808
rect 19220 25768 21236 25808
rect 25996 25808 26036 25852
rect 25996 25768 27340 25808
rect 27380 25768 27389 25808
rect 10060 25724 10100 25768
rect 3103 25684 3112 25724
rect 3480 25684 3489 25724
rect 8323 25684 8332 25724
rect 8372 25684 9868 25724
rect 9908 25684 9917 25724
rect 10060 25684 10444 25724
rect 10484 25684 10493 25724
rect 10877 25684 10886 25724
rect 11254 25684 11263 25724
rect 15139 25684 15148 25724
rect 15188 25684 17068 25724
rect 17108 25684 17117 25724
rect 17932 25640 17972 25768
rect 19084 25724 19124 25768
rect 18651 25684 18660 25724
rect 19028 25684 19037 25724
rect 19084 25684 26036 25724
rect 26425 25684 26434 25724
rect 26802 25684 26811 25724
rect 26947 25684 26956 25724
rect 26996 25684 29932 25724
rect 29972 25684 29981 25724
rect 25996 25640 26036 25684
rect 9292 25600 17356 25640
rect 17396 25600 17405 25640
rect 17932 25600 25804 25640
rect 25844 25600 25853 25640
rect 25996 25600 28972 25640
rect 29012 25600 29021 25640
rect 9292 25556 9332 25600
rect 5530 25516 5539 25556
rect 5579 25516 6316 25556
rect 6356 25516 6365 25556
rect 9274 25516 9283 25556
rect 9323 25516 9332 25556
rect 10147 25516 10156 25556
rect 10196 25516 10772 25556
rect 10819 25516 10828 25556
rect 10868 25516 11308 25556
rect 11348 25516 11357 25556
rect 12643 25516 12652 25556
rect 12692 25516 12844 25556
rect 12884 25516 12893 25556
rect 12940 25516 16156 25556
rect 16196 25516 16205 25556
rect 19555 25516 19564 25556
rect 19604 25516 19756 25556
rect 19796 25516 19900 25556
rect 19940 25516 19949 25556
rect 20323 25516 20332 25556
rect 20372 25516 23060 25556
rect 23779 25516 23788 25556
rect 23828 25516 25420 25556
rect 25460 25516 25612 25556
rect 25652 25516 26476 25556
rect 26516 25516 27244 25556
rect 27284 25516 27293 25556
rect 10732 25472 10772 25516
rect 12940 25472 12980 25516
rect 23020 25472 23060 25516
rect 4684 25432 5068 25472
rect 5108 25432 5155 25472
rect 5195 25432 5204 25472
rect 6761 25432 6892 25472
rect 6932 25432 6941 25472
rect 10601 25432 10732 25472
rect 10772 25432 11348 25472
rect 11491 25432 11500 25472
rect 11540 25432 12980 25472
rect 13027 25432 13036 25472
rect 13076 25432 13207 25472
rect 14537 25432 14668 25472
rect 14708 25432 14717 25472
rect 19843 25432 19852 25472
rect 19892 25432 21196 25472
rect 21236 25432 21245 25472
rect 23020 25432 23596 25472
rect 23636 25432 24308 25472
rect 3043 25348 3052 25388
rect 3092 25348 3101 25388
rect 4684 25304 4724 25432
rect 5164 25348 5644 25388
rect 5684 25348 5693 25388
rect 8899 25348 8908 25388
rect 8948 25348 9964 25388
rect 10004 25348 10100 25388
rect 10531 25348 10540 25388
rect 10580 25348 10676 25388
rect 11033 25348 11116 25388
rect 11195 25348 11213 25388
rect 2563 25264 2572 25304
rect 2612 25264 3139 25304
rect 3179 25264 3188 25304
rect 4472 25264 4481 25304
rect 4521 25264 4724 25304
rect 4771 25289 4780 25329
rect 4820 25289 4842 25329
rect 5164 25304 5204 25348
rect 9542 25304 9582 25348
rect 10060 25304 10100 25348
rect 10636 25304 10676 25348
rect 11308 25346 11348 25432
rect 11500 25348 21332 25388
rect 22243 25348 22252 25388
rect 22292 25348 22301 25388
rect 23753 25348 23884 25388
rect 23924 25348 23933 25388
rect 11308 25306 11347 25346
rect 11387 25306 11396 25346
rect 11500 25304 11540 25348
rect 4780 25220 4820 25289
rect 4963 25264 4972 25304
rect 5012 25264 5021 25304
rect 5146 25264 5155 25304
rect 5195 25264 5204 25304
rect 5251 25264 5260 25304
rect 5300 25264 5356 25304
rect 5396 25264 5431 25304
rect 5530 25264 5539 25304
rect 5588 25264 5740 25304
rect 5780 25264 5789 25304
rect 6499 25264 6508 25304
rect 6548 25264 6557 25304
rect 8227 25264 8236 25304
rect 8276 25264 9004 25304
rect 9044 25264 9053 25304
rect 9161 25264 9283 25304
rect 9332 25264 9341 25304
rect 9402 25264 9411 25304
rect 9451 25264 9460 25304
rect 9524 25264 9533 25304
rect 9573 25264 9582 25304
rect 9658 25264 9667 25304
rect 9707 25264 9716 25304
rect 9835 25264 9844 25304
rect 9884 25264 10004 25304
rect 10060 25264 10540 25304
rect 10580 25264 10589 25304
rect 10636 25264 10662 25304
rect 10702 25264 10711 25304
rect 10780 25264 10789 25304
rect 10868 25264 10969 25304
rect 11479 25264 11488 25304
rect 11528 25264 11540 25304
rect 11587 25264 11596 25304
rect 11636 25264 11980 25304
rect 12020 25264 12029 25304
rect 12346 25264 12355 25304
rect 12395 25264 12404 25304
rect 12643 25264 12652 25304
rect 12703 25264 12823 25304
rect 13315 25264 13324 25304
rect 13364 25264 14284 25304
rect 14324 25264 14333 25304
rect 14467 25264 14476 25304
rect 14516 25264 14647 25304
rect 15209 25264 15340 25304
rect 15380 25264 15389 25304
rect 16361 25264 16492 25304
rect 16532 25264 16541 25304
rect 16771 25264 16780 25304
rect 16820 25264 16829 25304
rect 17225 25264 17347 25304
rect 17396 25264 17405 25304
rect 17453 25264 17462 25304
rect 17502 25264 17548 25304
rect 17588 25264 17633 25304
rect 18077 25264 18109 25304
rect 18149 25264 18164 25304
rect 18211 25264 18220 25304
rect 18260 25264 18269 25304
rect 18569 25264 18700 25304
rect 18740 25264 18749 25304
rect 18883 25264 18892 25304
rect 18932 25264 19063 25304
rect 19337 25264 19372 25304
rect 19412 25264 19468 25304
rect 19508 25264 19517 25304
rect 19651 25264 19660 25304
rect 19700 25264 19852 25304
rect 19892 25264 19901 25304
rect 20009 25264 20044 25304
rect 20084 25264 20140 25304
rect 20180 25264 20189 25304
rect 20323 25264 20332 25304
rect 20372 25264 20381 25304
rect 20489 25264 20611 25304
rect 20660 25264 20669 25304
rect 4972 25220 5012 25264
rect 5260 25220 5300 25264
rect 6508 25220 6548 25264
rect 3514 25180 3523 25220
rect 3563 25180 3572 25220
rect 4771 25180 4780 25220
rect 4820 25180 4829 25220
rect 4972 25180 5300 25220
rect 5548 25180 6548 25220
rect 3532 25136 3572 25180
rect 4972 25136 5012 25180
rect 1219 25096 1228 25136
rect 1268 25096 1277 25136
rect 3532 25096 4579 25136
rect 4619 25096 4628 25136
rect 4675 25096 4684 25136
rect 4724 25096 5012 25136
rect 1228 24800 1268 25096
rect 4343 24928 4352 24968
rect 4720 24928 4729 24968
rect 4771 24844 4780 24884
rect 4820 24844 5452 24884
rect 5492 24844 5501 24884
rect 4972 24800 5012 24844
rect 5548 24800 5588 25180
rect 5705 25096 5836 25136
rect 5876 25096 5885 25136
rect 6979 25096 6988 25136
rect 7028 25096 7276 25136
rect 7316 25096 7325 25136
rect 8009 25096 8131 25136
rect 8180 25096 8189 25136
rect 8419 25096 8428 25136
rect 8468 25096 8524 25136
rect 8564 25096 8599 25136
rect 9410 24968 9450 25264
rect 9676 25052 9716 25264
rect 9964 25136 10004 25264
rect 11500 25220 11540 25264
rect 12364 25220 12404 25264
rect 16780 25220 16820 25264
rect 18124 25220 18164 25264
rect 18220 25220 18260 25264
rect 20332 25220 20372 25264
rect 21292 25220 21332 25348
rect 24268 25346 24308 25432
rect 24211 25306 24220 25346
rect 24260 25306 24308 25346
rect 24395 25337 24435 25516
rect 24652 25432 24844 25472
rect 24884 25432 24893 25472
rect 25507 25432 25516 25472
rect 25556 25432 26956 25472
rect 26996 25432 27005 25472
rect 28090 25432 28099 25472
rect 28139 25432 28628 25472
rect 24547 25348 24556 25388
rect 24596 25348 24605 25388
rect 21562 25264 21571 25304
rect 21611 25264 22732 25304
rect 22772 25264 22781 25304
rect 23971 25264 23980 25304
rect 24020 25264 24029 25304
rect 24076 25264 24099 25304
rect 24139 25264 24148 25304
rect 24556 25304 24596 25348
rect 24652 25304 24692 25432
rect 28588 25388 28628 25432
rect 24739 25348 24748 25388
rect 24788 25348 24797 25388
rect 24931 25348 24940 25388
rect 24980 25348 25018 25388
rect 24748 25304 24788 25348
rect 24978 25304 25018 25348
rect 25546 25379 26092 25388
rect 25546 25339 25555 25379
rect 25595 25348 26092 25379
rect 26132 25348 26141 25388
rect 26275 25348 26284 25388
rect 26324 25348 26668 25388
rect 26708 25348 26717 25388
rect 26947 25348 26956 25388
rect 26996 25348 27031 25388
rect 27773 25348 27820 25388
rect 27860 25348 27869 25388
rect 27927 25348 28012 25388
rect 28052 25348 28061 25388
rect 28570 25348 28579 25388
rect 28619 25348 28628 25388
rect 30307 25348 30316 25388
rect 30356 25348 30365 25388
rect 25595 25339 25604 25348
rect 25128 25304 25137 25339
rect 24395 25288 24435 25297
rect 24509 25295 24596 25304
rect 24509 25264 24547 25295
rect 23980 25220 24020 25264
rect 24076 25220 24116 25264
rect 24538 25255 24547 25264
rect 24587 25255 24596 25295
rect 24643 25264 24652 25304
rect 24692 25264 24701 25304
rect 24748 25264 24844 25304
rect 24884 25264 24893 25304
rect 24960 25264 24969 25304
rect 25009 25264 25018 25304
rect 25109 25264 25118 25304
rect 25177 25299 25268 25339
rect 25546 25338 25604 25339
rect 26284 25304 26324 25348
rect 26991 25304 27031 25348
rect 27820 25304 27860 25348
rect 27927 25304 27967 25348
rect 25158 25264 25268 25299
rect 25315 25264 25324 25304
rect 25364 25264 25373 25304
rect 25654 25264 25663 25304
rect 25703 25264 25844 25304
rect 25891 25264 25900 25304
rect 25940 25264 26071 25304
rect 26284 25264 26371 25304
rect 26411 25264 26420 25304
rect 26467 25264 26476 25304
rect 26516 25264 26572 25304
rect 26612 25264 26647 25304
rect 26729 25264 26860 25304
rect 26900 25264 26909 25304
rect 26973 25264 26982 25304
rect 27022 25264 27043 25304
rect 27100 25264 27109 25304
rect 27149 25264 27158 25304
rect 27802 25264 27811 25304
rect 27851 25264 27860 25304
rect 27909 25264 27918 25304
rect 27958 25264 27967 25304
rect 28195 25264 28204 25304
rect 28244 25264 28439 25304
rect 28479 25264 28488 25304
rect 28675 25264 28684 25304
rect 28724 25264 28855 25304
rect 29338 25264 29347 25304
rect 29387 25264 30892 25304
rect 30932 25264 30941 25304
rect 24538 25254 24596 25255
rect 25324 25220 25364 25264
rect 10540 25180 11540 25220
rect 11635 25180 11644 25220
rect 11684 25180 11924 25220
rect 11971 25180 11980 25220
rect 12020 25180 12404 25220
rect 14371 25180 14380 25220
rect 14420 25180 16588 25220
rect 16628 25180 16820 25220
rect 17260 25180 17932 25220
rect 17972 25180 17981 25220
rect 18115 25180 18124 25220
rect 18164 25180 18173 25220
rect 18220 25180 19220 25220
rect 19267 25180 19276 25220
rect 19316 25180 20372 25220
rect 20707 25180 20716 25220
rect 20756 25180 20765 25220
rect 21178 25180 21187 25220
rect 21227 25180 21236 25220
rect 21292 25180 23980 25220
rect 24020 25180 24029 25220
rect 24076 25180 24500 25220
rect 24931 25180 24940 25220
rect 24980 25180 25612 25220
rect 25652 25180 25661 25220
rect 10540 25136 10580 25180
rect 11884 25136 11924 25180
rect 9964 25096 10156 25136
rect 10196 25096 10580 25136
rect 10636 25096 11692 25136
rect 11732 25096 11741 25136
rect 11875 25096 11884 25136
rect 11924 25096 12451 25136
rect 12491 25096 12500 25136
rect 15881 25096 16012 25136
rect 16052 25096 16061 25136
rect 10636 25052 10676 25096
rect 17260 25052 17300 25180
rect 19180 25136 19220 25180
rect 17609 25096 17644 25136
rect 17684 25096 17740 25136
rect 17780 25096 17789 25136
rect 17914 25096 17923 25136
rect 17963 25096 17972 25136
rect 18761 25096 18883 25136
rect 18932 25096 18941 25136
rect 19162 25096 19171 25136
rect 19211 25096 19220 25136
rect 17932 25052 17972 25096
rect 19276 25052 19316 25180
rect 9545 25012 9676 25052
rect 9716 25012 10676 25052
rect 10915 25012 10924 25052
rect 10964 25012 11308 25052
rect 11348 25012 17300 25052
rect 17347 25012 17356 25052
rect 17396 25012 17972 25052
rect 18211 25012 18220 25052
rect 18260 25012 19316 25052
rect 9292 24928 9450 24968
rect 9859 24928 9868 24968
rect 9908 24928 11500 24968
rect 11540 24928 11549 24968
rect 12117 24928 12126 24968
rect 12494 24928 12503 24968
rect 14467 24928 14476 24968
rect 14516 24928 18356 24968
rect 19891 24928 19900 24968
rect 20268 24928 20277 24968
rect 9292 24800 9332 24928
rect 18316 24884 18356 24928
rect 1228 24760 4099 24800
rect 4139 24760 4148 24800
rect 4963 24760 4972 24800
rect 5012 24760 5021 24800
rect 5539 24760 5548 24800
rect 5588 24760 5597 24800
rect 8131 24760 8140 24800
rect 8180 24760 8899 24800
rect 8939 24760 8948 24800
rect 9187 24760 9196 24800
rect 9236 24760 9332 24800
rect 9484 24844 12980 24884
rect 4867 24676 4876 24716
rect 4916 24676 5492 24716
rect 8323 24676 8332 24716
rect 8372 24676 8397 24716
rect 8449 24676 8908 24716
rect 8948 24676 8957 24716
rect 5452 24632 5492 24676
rect 8332 24632 8372 24676
rect 8449 24632 8489 24676
rect 2057 24592 2188 24632
rect 2228 24592 2237 24632
rect 4073 24592 4204 24632
rect 4244 24592 4253 24632
rect 4387 24592 4396 24632
rect 4436 24592 4588 24632
rect 4628 24592 4637 24632
rect 4771 24592 4780 24632
rect 4820 24592 4972 24632
rect 5012 24592 5021 24632
rect 5146 24592 5155 24632
rect 5204 24592 5335 24632
rect 5443 24592 5452 24632
rect 5492 24592 5501 24632
rect 5626 24592 5635 24632
rect 5684 24592 5815 24632
rect 6202 24592 6211 24632
rect 6260 24592 6391 24632
rect 8292 24592 8301 24632
rect 8341 24592 8372 24632
rect 8428 24592 8449 24632
rect 8489 24592 8498 24632
rect 8707 24592 8716 24632
rect 8781 24592 8887 24632
rect 8995 24592 9004 24632
rect 9044 24592 9175 24632
rect 8428 24548 8468 24592
rect 9484 24548 9524 24844
rect 10435 24760 10444 24800
rect 10484 24760 10627 24800
rect 10667 24760 10676 24800
rect 12940 24716 12980 24844
rect 17452 24844 18260 24884
rect 18316 24844 20332 24884
rect 20372 24844 20381 24884
rect 17452 24800 17492 24844
rect 18220 24800 18260 24844
rect 14746 24760 14755 24800
rect 14795 24760 15340 24800
rect 15380 24760 15389 24800
rect 16810 24760 16819 24800
rect 16859 24760 17492 24800
rect 17539 24760 17548 24800
rect 17588 24760 17827 24800
rect 17867 24760 17876 24800
rect 17923 24760 17932 24800
rect 17972 24760 18124 24800
rect 18164 24760 18173 24800
rect 18220 24760 18740 24800
rect 18883 24760 18892 24800
rect 18932 24760 20236 24800
rect 20276 24760 20285 24800
rect 18700 24716 18740 24760
rect 19564 24716 19604 24760
rect 9929 24676 9964 24716
rect 10004 24707 10100 24716
rect 10004 24676 10051 24707
rect 10042 24667 10051 24676
rect 10091 24667 10100 24707
rect 10147 24676 10156 24716
rect 10196 24676 10205 24716
rect 11587 24676 11596 24716
rect 11636 24676 12404 24716
rect 12940 24676 14612 24716
rect 10042 24666 10100 24667
rect 10156 24632 10196 24676
rect 12364 24632 12404 24676
rect 14572 24632 14612 24676
rect 14668 24676 16052 24716
rect 17908 24676 18028 24716
rect 18079 24676 18088 24716
rect 18211 24676 18220 24716
rect 18260 24676 18297 24716
rect 18700 24676 18988 24716
rect 19028 24676 19037 24716
rect 19546 24707 19604 24716
rect 14668 24632 14708 24676
rect 9571 24592 9580 24632
rect 9620 24592 9763 24632
rect 9803 24592 9812 24632
rect 9868 24623 9908 24632
rect 10146 24592 10155 24632
rect 10195 24592 10243 24632
rect 10315 24592 10324 24632
rect 10364 24592 10772 24632
rect 10906 24592 10915 24632
rect 10964 24592 11095 24632
rect 11395 24592 11404 24632
rect 11444 24592 11447 24632
rect 11487 24592 11575 24632
rect 11683 24592 11692 24632
rect 11732 24592 11863 24632
rect 12346 24592 12355 24632
rect 12395 24592 12404 24632
rect 14292 24592 14380 24632
rect 14420 24592 14423 24632
rect 14463 24592 14472 24632
rect 14554 24592 14563 24632
rect 14603 24592 14612 24632
rect 14659 24592 14668 24632
rect 14708 24592 14717 24632
rect 14851 24592 14860 24632
rect 14900 24623 15031 24632
rect 14900 24592 14947 24623
rect 9868 24548 9908 24583
rect 5827 24508 5836 24548
rect 5876 24508 5885 24548
rect 6883 24508 6892 24548
rect 6932 24508 6941 24548
rect 8227 24508 8236 24548
rect 8276 24508 8468 24548
rect 8515 24508 8524 24548
rect 8564 24508 8620 24548
rect 8660 24508 8695 24548
rect 8812 24508 9524 24548
rect 9763 24508 9772 24548
rect 9812 24508 9908 24548
rect 10060 24508 10252 24548
rect 10292 24508 10301 24548
rect 10409 24508 10531 24548
rect 10580 24508 10589 24548
rect 5836 24464 5876 24508
rect 8812 24464 8852 24508
rect 10060 24464 10100 24508
rect 1769 24424 1900 24464
rect 1940 24424 1949 24464
rect 2921 24424 3052 24464
rect 3092 24424 3101 24464
rect 4387 24424 4396 24464
rect 4436 24424 5068 24464
rect 5108 24424 5117 24464
rect 5191 24424 5200 24464
rect 5240 24424 5644 24464
rect 5684 24424 5693 24464
rect 5789 24424 5836 24464
rect 5876 24424 5885 24464
rect 8515 24424 8524 24464
rect 8564 24424 8852 24464
rect 9772 24424 10100 24464
rect 10732 24464 10772 24592
rect 14938 24583 14947 24592
rect 14987 24592 15031 24623
rect 14987 24583 14996 24592
rect 14938 24582 14996 24583
rect 16012 24548 16052 24676
rect 16099 24592 16108 24632
rect 16148 24592 16279 24632
rect 16963 24592 16972 24632
rect 17024 24592 17143 24632
rect 17443 24592 17452 24632
rect 17492 24592 17731 24632
rect 17771 24592 17780 24632
rect 18220 24627 18260 24676
rect 18700 24632 18740 24676
rect 19546 24667 19555 24707
rect 19595 24667 19604 24707
rect 19546 24666 19604 24667
rect 19660 24676 20516 24716
rect 19660 24632 19700 24676
rect 20476 24632 20516 24676
rect 18206 24587 18215 24627
rect 18255 24587 18264 24627
rect 18403 24592 18412 24632
rect 18452 24592 18583 24632
rect 18691 24592 18700 24632
rect 18740 24592 18749 24632
rect 18979 24592 18988 24632
rect 19028 24592 19037 24632
rect 19123 24592 19132 24632
rect 19172 24592 19267 24632
rect 19307 24592 19316 24632
rect 19372 24623 19412 24632
rect 18988 24548 19028 24592
rect 19642 24592 19651 24632
rect 19691 24592 19700 24632
rect 19747 24592 19756 24632
rect 19825 24592 19996 24632
rect 20036 24592 20045 24632
rect 20166 24592 20236 24632
rect 20276 24592 20297 24632
rect 20337 24592 20346 24632
rect 20458 24592 20467 24632
rect 20507 24592 20660 24632
rect 19372 24548 19412 24583
rect 10985 24508 11107 24548
rect 11156 24508 11165 24548
rect 11578 24508 11587 24548
rect 11627 24508 11636 24548
rect 11779 24508 11788 24548
rect 11828 24508 11980 24548
rect 12020 24508 12029 24548
rect 13027 24508 13036 24548
rect 13076 24508 13085 24548
rect 15091 24508 15100 24548
rect 15140 24508 15148 24548
rect 15188 24508 15271 24548
rect 16012 24508 18164 24548
rect 18307 24508 18316 24548
rect 18356 24508 18365 24548
rect 18988 24508 19084 24548
rect 19124 24508 19133 24548
rect 19296 24508 19372 24548
rect 19412 24508 20140 24548
rect 20180 24508 20189 24548
rect 11596 24464 11636 24508
rect 18124 24464 18164 24508
rect 18316 24464 18356 24508
rect 20620 24464 20660 24592
rect 20716 24548 20756 25180
rect 21043 25096 21052 25136
rect 21092 25096 21140 25136
rect 21100 24632 21140 25096
rect 21196 24800 21236 25180
rect 24460 25136 24500 25180
rect 22819 25096 22828 25136
rect 22868 25096 23500 25136
rect 23540 25096 23549 25136
rect 24233 25096 24364 25136
rect 24404 25096 24413 25136
rect 24460 25096 25132 25136
rect 25172 25096 25181 25136
rect 25411 25096 25420 25136
rect 25460 25096 25591 25136
rect 25804 25052 25844 25264
rect 27118 25220 27158 25264
rect 26275 25180 26284 25220
rect 26324 25180 26659 25220
rect 26699 25180 26708 25220
rect 26947 25180 26956 25220
rect 26996 25180 27158 25220
rect 28762 25180 28771 25220
rect 28811 25180 28963 25220
rect 29003 25180 29012 25220
rect 26345 25096 26380 25136
rect 26420 25096 26476 25136
rect 26516 25096 26525 25136
rect 31267 25096 31276 25136
rect 31316 25096 31325 25136
rect 25804 25012 26380 25052
rect 26420 25012 26429 25052
rect 27665 24928 27674 24968
rect 28042 24928 28051 24968
rect 26092 24844 26860 24884
rect 26900 24844 26909 24884
rect 27967 24844 28916 24884
rect 21187 24760 21196 24800
rect 21236 24760 21245 24800
rect 23491 24760 23500 24800
rect 23540 24760 25036 24800
rect 25076 24760 25085 24800
rect 25315 24760 25324 24800
rect 25364 24760 25652 24800
rect 25612 24716 25652 24760
rect 21187 24676 21196 24716
rect 21236 24676 24940 24716
rect 24980 24676 24989 24716
rect 25210 24676 25219 24716
rect 25259 24676 25268 24716
rect 25411 24676 25420 24716
rect 25460 24676 25556 24716
rect 25612 24676 25804 24716
rect 25844 24676 25991 24716
rect 23596 24632 23636 24676
rect 21100 24592 21868 24632
rect 21908 24592 21917 24632
rect 22697 24592 22828 24632
rect 22868 24592 22877 24632
rect 23587 24592 23596 24632
rect 23636 24592 23645 24632
rect 24233 24592 24333 24632
rect 24404 24592 24413 24632
rect 24486 24592 24495 24632
rect 24535 24592 24556 24632
rect 24596 24592 24666 24632
rect 24739 24592 24748 24632
rect 24813 24592 24919 24632
rect 24987 24592 25036 24632
rect 25076 24592 25118 24632
rect 25158 24592 25167 24632
rect 25228 24548 25268 24676
rect 25516 24629 25556 24676
rect 25951 24632 25991 24676
rect 26092 24632 26132 24844
rect 26249 24760 26380 24800
rect 26420 24760 26429 24800
rect 26563 24760 26572 24800
rect 26612 24760 27052 24800
rect 27092 24760 27101 24800
rect 27967 24716 28007 24844
rect 28876 24800 28916 24844
rect 28090 24760 28099 24800
rect 28139 24760 28684 24800
rect 28724 24760 28733 24800
rect 28867 24760 28876 24800
rect 28916 24760 28925 24800
rect 31276 24716 31316 25096
rect 26179 24676 26188 24716
rect 26228 24676 26237 24716
rect 26332 24676 26764 24716
rect 26804 24676 26813 24716
rect 27148 24676 27436 24716
rect 27476 24676 27485 24716
rect 27967 24676 28148 24716
rect 26188 24632 26228 24676
rect 26332 24632 26372 24676
rect 27148 24632 27188 24676
rect 28108 24632 28148 24676
rect 28308 24676 28396 24716
rect 28436 24676 28445 24716
rect 30220 24676 31316 24716
rect 28308 24659 28348 24676
rect 25417 24589 25426 24629
rect 25466 24589 25556 24629
rect 25603 24592 25612 24632
rect 25652 24623 25889 24632
rect 25652 24592 25849 24623
rect 20716 24508 22147 24548
rect 22187 24508 22196 24548
rect 22252 24508 23500 24548
rect 23540 24508 23549 24548
rect 24643 24508 24652 24548
rect 24692 24508 25268 24548
rect 25942 24592 25951 24632
rect 25991 24592 26000 24632
rect 26074 24623 26132 24632
rect 22252 24464 22292 24508
rect 25849 24464 25889 24583
rect 26074 24583 26083 24623
rect 26123 24583 26132 24623
rect 26179 24592 26188 24632
rect 26228 24592 26275 24632
rect 26332 24592 26369 24632
rect 26409 24592 26418 24632
rect 26568 24592 26577 24632
rect 26617 24592 26708 24632
rect 26825 24592 26956 24632
rect 26996 24592 27005 24632
rect 27130 24592 27139 24632
rect 27179 24592 27188 24632
rect 27331 24592 27340 24632
rect 27380 24592 27436 24632
rect 27476 24592 27511 24632
rect 27619 24592 27628 24632
rect 27668 24592 27724 24632
rect 27764 24592 27799 24632
rect 27907 24592 27916 24632
rect 27956 24592 27965 24632
rect 28099 24592 28108 24632
rect 28148 24592 28157 24632
rect 28289 24619 28298 24659
rect 28338 24619 28348 24659
rect 30220 24632 30260 24676
rect 28483 24592 28492 24632
rect 28532 24592 28541 24632
rect 29417 24592 29548 24632
rect 29588 24592 30260 24632
rect 30787 24592 30796 24632
rect 30836 24592 30845 24632
rect 26074 24582 26132 24583
rect 26668 24548 26708 24592
rect 26659 24508 26668 24548
rect 26708 24508 26717 24548
rect 26845 24464 26885 24592
rect 27916 24548 27956 24592
rect 28492 24548 28532 24592
rect 30796 24548 30836 24592
rect 27715 24508 27724 24548
rect 27764 24508 28108 24548
rect 28148 24508 28157 24548
rect 28265 24508 28396 24548
rect 28436 24508 28445 24548
rect 28492 24508 31276 24548
rect 31316 24508 31325 24548
rect 28492 24464 28532 24508
rect 10732 24424 11500 24464
rect 11540 24424 11549 24464
rect 11596 24424 11884 24464
rect 11924 24424 11933 24464
rect 14124 24424 14188 24464
rect 14228 24424 14284 24464
rect 14324 24424 15572 24464
rect 17033 24424 17164 24464
rect 17204 24424 17213 24464
rect 18124 24424 18356 24464
rect 19171 24424 19180 24464
rect 19220 24424 20236 24464
rect 20276 24424 20285 24464
rect 20620 24424 22292 24464
rect 22889 24424 22924 24464
rect 22964 24424 23020 24464
rect 23060 24424 23124 24464
rect 23203 24424 23212 24464
rect 23252 24424 23444 24464
rect 24425 24424 24556 24464
rect 24596 24424 24605 24464
rect 25849 24424 26885 24464
rect 27523 24424 27532 24464
rect 27572 24424 28532 24464
rect 29801 24424 29932 24464
rect 29972 24424 29981 24464
rect 30595 24424 30604 24464
rect 30644 24424 30988 24464
rect 31028 24424 31037 24464
rect 9772 24380 9812 24424
rect 11596 24380 11636 24424
rect 15532 24380 15572 24424
rect 23404 24380 23444 24424
rect 2851 24340 2860 24380
rect 2900 24340 3532 24380
rect 3572 24340 3581 24380
rect 4579 24340 4588 24380
rect 4628 24340 5356 24380
rect 5396 24340 5405 24380
rect 9754 24340 9763 24380
rect 9803 24340 9812 24380
rect 10435 24340 10444 24380
rect 10484 24340 11636 24380
rect 13769 24340 13900 24380
rect 13940 24340 13949 24380
rect 15235 24340 15244 24380
rect 15284 24340 15436 24380
rect 15476 24340 15485 24380
rect 15532 24340 19084 24380
rect 19124 24340 19133 24380
rect 19258 24340 19267 24380
rect 19307 24340 21580 24380
rect 21620 24340 21629 24380
rect 22252 24340 23348 24380
rect 23404 24340 24596 24380
rect 24643 24340 24652 24380
rect 24692 24340 25804 24380
rect 25844 24340 25900 24380
rect 25940 24340 25949 24380
rect 27017 24340 27139 24380
rect 27188 24340 27197 24380
rect 28771 24340 28780 24380
rect 28820 24340 30124 24380
rect 30164 24340 30173 24380
rect 22252 24296 22292 24340
rect 23308 24296 23348 24340
rect 24556 24296 24596 24340
rect 3619 24256 3628 24296
rect 3668 24256 16916 24296
rect 16963 24256 16972 24296
rect 17012 24256 22292 24296
rect 22339 24256 22348 24296
rect 22388 24256 23212 24296
rect 23252 24256 23261 24296
rect 23308 24256 24460 24296
rect 24500 24256 24509 24296
rect 24556 24256 29452 24296
rect 29492 24256 29501 24296
rect 3103 24172 3112 24212
rect 3480 24172 3489 24212
rect 3724 24172 8084 24212
rect 8611 24172 8620 24212
rect 8660 24172 10444 24212
rect 10484 24172 10493 24212
rect 10877 24172 10886 24212
rect 11254 24172 11263 24212
rect 2956 23920 3148 23960
rect 3188 23920 3197 23960
rect 2956 23876 2996 23920
rect 1891 23836 1900 23876
rect 1940 23836 1949 23876
rect 2938 23836 2947 23876
rect 2987 23836 2996 23876
rect 2441 23752 2563 23792
rect 2612 23752 2621 23792
rect 3401 23752 3532 23792
rect 3572 23752 3581 23792
rect 3532 23734 3572 23743
rect 634 23668 643 23708
rect 683 23668 2188 23708
rect 2228 23668 2237 23708
rect 3427 23668 3436 23708
rect 3476 23668 3485 23708
rect 3436 23624 3476 23668
rect 3436 23584 3628 23624
rect 3668 23584 3677 23624
rect 3724 23372 3764 24172
rect 8044 24128 8084 24172
rect 16876 24128 16916 24256
rect 18651 24172 18660 24212
rect 19028 24172 19037 24212
rect 19084 24172 24844 24212
rect 24884 24172 24893 24212
rect 26425 24172 26434 24212
rect 26802 24172 26811 24212
rect 19084 24128 19124 24172
rect 5155 24088 5164 24128
rect 5204 24088 7988 24128
rect 8044 24088 13420 24128
rect 13460 24088 13469 24128
rect 16876 24088 19124 24128
rect 20803 24088 20812 24128
rect 20852 24088 27340 24128
rect 27380 24088 27444 24128
rect 7948 24044 7988 24088
rect 5129 24004 5251 24044
rect 5300 24004 5309 24044
rect 7930 24004 7939 24044
rect 7979 24004 7988 24044
rect 8140 24004 9292 24044
rect 9332 24004 9341 24044
rect 9667 24004 9676 24044
rect 9716 24004 10540 24044
rect 10580 24004 10589 24044
rect 11683 24004 11692 24044
rect 11732 24004 12268 24044
rect 12308 24004 12317 24044
rect 15532 24004 16012 24044
rect 16052 24004 16061 24044
rect 18403 24004 18412 24044
rect 18452 24004 18604 24044
rect 18644 24004 18653 24044
rect 19267 24004 19276 24044
rect 19316 24004 19459 24044
rect 19499 24004 19508 24044
rect 22723 24004 22732 24044
rect 22772 24004 26956 24044
rect 26996 24004 27005 24044
rect 4780 23920 5108 23960
rect 3820 23836 4243 23876
rect 4283 23836 4396 23876
rect 4436 23836 4445 23876
rect 3820 23792 3860 23836
rect 4780 23792 4820 23920
rect 5068 23876 5108 23920
rect 5002 23867 5108 23876
rect 5002 23827 5011 23867
rect 5051 23836 5108 23867
rect 5303 23920 6220 23960
rect 6260 23920 6269 23960
rect 6953 23920 7084 23960
rect 7124 23920 7133 23960
rect 5051 23827 5060 23836
rect 5002 23826 5060 23827
rect 5303 23792 5343 23920
rect 5548 23792 5588 23801
rect 8140 23792 8180 24004
rect 8969 23920 9100 23960
rect 9140 23920 9149 23960
rect 9283 23920 9292 23960
rect 9332 23920 10828 23960
rect 10868 23920 11636 23960
rect 11962 23920 11971 23960
rect 12011 23920 14324 23960
rect 11596 23876 11636 23920
rect 3811 23752 3820 23792
rect 3860 23752 3869 23792
rect 4195 23752 4204 23792
rect 4244 23752 4438 23792
rect 4478 23752 4820 23792
rect 4866 23752 4875 23792
rect 4915 23752 4924 23792
rect 5104 23752 5113 23792
rect 5153 23752 5343 23792
rect 5417 23752 5548 23792
rect 5588 23752 5597 23792
rect 6883 23752 6892 23792
rect 6932 23752 7468 23792
rect 7508 23752 7517 23792
rect 7928 23752 7937 23792
rect 7977 23752 8180 23792
rect 8236 23836 9004 23876
rect 9044 23836 9716 23876
rect 8236 23792 8276 23836
rect 9676 23792 9716 23836
rect 9868 23836 10060 23876
rect 10100 23836 10109 23876
rect 11596 23836 11828 23876
rect 11875 23836 11884 23876
rect 11924 23836 12116 23876
rect 12425 23836 12547 23876
rect 12596 23836 12605 23876
rect 9868 23792 9908 23836
rect 11788 23792 11828 23836
rect 12076 23792 12116 23836
rect 14284 23792 14324 23920
rect 15532 23876 15572 24004
rect 18761 23951 18892 23960
rect 18761 23920 18860 23951
rect 18932 23920 18941 23960
rect 19075 23920 19084 23960
rect 19124 23920 19468 23960
rect 19508 23920 19517 23960
rect 24268 23920 24556 23960
rect 24596 23920 24605 23960
rect 25132 23920 25516 23960
rect 25556 23920 25565 23960
rect 26563 23920 26572 23960
rect 26612 23920 27148 23960
rect 27188 23920 27197 23960
rect 18860 23902 18900 23911
rect 14371 23836 14380 23876
rect 14420 23836 14515 23876
rect 14555 23836 14564 23876
rect 15139 23836 15148 23876
rect 15188 23836 15197 23876
rect 15427 23836 15436 23876
rect 15476 23836 15572 23876
rect 17088 23836 17164 23876
rect 17204 23836 17213 23876
rect 19795 23836 19804 23876
rect 19844 23836 20812 23876
rect 20852 23836 20861 23876
rect 22915 23836 22924 23876
rect 22964 23836 22973 23876
rect 23098 23836 23107 23876
rect 23147 23836 24212 23876
rect 15148 23792 15188 23836
rect 8515 23752 8524 23792
rect 8564 23752 8573 23792
rect 8707 23752 8716 23792
rect 8756 23752 8765 23792
rect 9161 23752 9292 23792
rect 9332 23752 9341 23792
rect 9475 23752 9484 23792
rect 9524 23752 9533 23792
rect 9667 23752 9676 23792
rect 9716 23752 9725 23792
rect 9859 23752 9868 23792
rect 9908 23752 9917 23792
rect 10435 23752 10444 23792
rect 10484 23752 10684 23792
rect 10724 23752 10733 23792
rect 10793 23752 10924 23792
rect 10964 23752 10973 23792
rect 11779 23752 11788 23792
rect 11828 23752 11837 23792
rect 11962 23752 11971 23792
rect 12011 23752 12020 23792
rect 12076 23752 12155 23792
rect 12195 23752 12204 23792
rect 12355 23752 12364 23792
rect 12404 23752 12413 23792
rect 13219 23752 13228 23792
rect 13268 23752 13900 23792
rect 13940 23752 13949 23792
rect 14057 23752 14188 23792
rect 14228 23752 14237 23792
rect 14284 23752 14680 23792
rect 14720 23752 14860 23792
rect 14900 23752 14909 23792
rect 15038 23752 15047 23792
rect 15087 23752 15188 23792
rect 15235 23752 15244 23792
rect 15284 23752 15415 23792
rect 15802 23752 15811 23792
rect 15851 23752 15860 23792
rect 17801 23752 17932 23792
rect 17972 23752 17981 23792
rect 18403 23752 18412 23792
rect 18452 23752 18883 23792
rect 18923 23752 18932 23792
rect 18979 23752 18988 23792
rect 19028 23752 19276 23792
rect 19316 23752 19325 23792
rect 19450 23752 19459 23792
rect 19499 23752 19508 23792
rect 19639 23752 19648 23792
rect 19700 23752 19828 23792
rect 22601 23752 22723 23792
rect 22772 23752 22781 23792
rect 23404 23752 23452 23792
rect 23492 23752 23501 23792
rect 23587 23752 23596 23792
rect 23636 23752 24076 23792
rect 24116 23752 24125 23792
rect 4649 23668 4780 23708
rect 4820 23668 4829 23708
rect 4343 23416 4352 23456
rect 4720 23416 4729 23456
rect 2179 23332 2188 23372
rect 2228 23332 3764 23372
rect 3148 23120 3188 23332
rect 4876 23288 4916 23752
rect 5107 23708 5147 23752
rect 5548 23743 5588 23752
rect 8236 23743 8276 23752
rect 8524 23708 8564 23752
rect 8716 23708 8756 23752
rect 9484 23708 9524 23752
rect 4963 23668 4972 23708
rect 5012 23668 5147 23708
rect 5240 23668 5249 23708
rect 5289 23668 5356 23708
rect 5396 23668 5420 23708
rect 8524 23668 8620 23708
rect 8660 23668 8669 23708
rect 8716 23668 9428 23708
rect 9484 23668 10051 23708
rect 10091 23668 10100 23708
rect 9388 23624 9428 23668
rect 11980 23624 12020 23752
rect 12364 23708 12404 23752
rect 15820 23708 15860 23752
rect 12364 23668 13507 23708
rect 13547 23668 13556 23708
rect 13603 23668 13612 23708
rect 13652 23668 15860 23708
rect 19468 23708 19508 23752
rect 19468 23668 20332 23708
rect 20372 23668 20381 23708
rect 5251 23584 5260 23624
rect 5300 23584 5452 23624
rect 5492 23584 5501 23624
rect 7980 23584 8044 23624
rect 8084 23584 8140 23624
rect 8180 23584 8332 23624
rect 8372 23584 8381 23624
rect 8585 23584 8707 23624
rect 8756 23584 8765 23624
rect 9388 23584 10540 23624
rect 10580 23584 10589 23624
rect 11203 23584 11212 23624
rect 11252 23584 11596 23624
rect 11636 23584 11645 23624
rect 11980 23584 12844 23624
rect 12884 23584 12893 23624
rect 15226 23584 15235 23624
rect 15275 23584 15284 23624
rect 5251 23416 5260 23456
rect 5300 23416 11692 23456
rect 11732 23416 11741 23456
rect 12117 23416 12126 23456
rect 12494 23416 12503 23456
rect 12556 23372 12596 23584
rect 15244 23372 15284 23584
rect 5644 23332 10484 23372
rect 4745 23248 4867 23288
rect 4907 23248 5012 23288
rect 5059 23248 5068 23288
rect 5108 23248 5588 23288
rect 4829 23164 4876 23204
rect 4916 23164 4925 23204
rect 4876 23120 4916 23164
rect 4972 23120 5012 23248
rect 5548 23204 5588 23248
rect 5530 23164 5539 23204
rect 5579 23164 5588 23204
rect 5644 23120 5684 23332
rect 7843 23248 7852 23288
rect 7892 23248 10252 23288
rect 10292 23248 10301 23288
rect 8410 23164 8419 23204
rect 8459 23164 8908 23204
rect 8948 23164 8957 23204
rect 10444 23120 10484 23332
rect 12316 23332 12596 23372
rect 12844 23332 15284 23372
rect 10915 23248 10924 23288
rect 10964 23248 11356 23288
rect 11396 23248 11405 23288
rect 10531 23164 10540 23204
rect 10580 23164 11059 23204
rect 11099 23164 11108 23204
rect 11203 23164 11212 23204
rect 11252 23164 11261 23204
rect 11212 23120 11252 23164
rect 12316 23122 12356 23332
rect 12547 23248 12556 23288
rect 12596 23248 12788 23288
rect 12268 23120 12356 23122
rect 835 23080 844 23120
rect 884 23080 2284 23120
rect 2324 23080 2333 23120
rect 3139 23080 3148 23120
rect 3188 23080 3197 23120
rect 3497 23080 3532 23120
rect 3572 23080 3628 23120
rect 3668 23080 3677 23120
rect 4588 23080 4684 23120
rect 4724 23080 4733 23120
rect 4867 23080 4876 23120
rect 4916 23080 4925 23120
rect 4972 23080 5164 23120
rect 5204 23080 5213 23120
rect 5392 23080 5401 23120
rect 5441 23080 5684 23120
rect 5914 23080 5923 23120
rect 5972 23080 6220 23120
rect 6260 23080 6269 23120
rect 7363 23080 7372 23120
rect 7412 23080 8044 23120
rect 8084 23080 8093 23120
rect 8794 23080 8803 23120
rect 8852 23080 8983 23120
rect 10444 23080 11116 23120
rect 11156 23080 11165 23120
rect 11212 23080 11224 23120
rect 11264 23080 11299 23120
rect 11491 23080 11500 23120
rect 11540 23080 11774 23120
rect 11814 23080 11823 23120
rect 11877 23080 11886 23120
rect 11926 23080 11935 23120
rect 11980 23080 12076 23120
rect 12116 23080 12125 23120
rect 12259 23080 12268 23120
rect 12308 23082 12356 23120
rect 12399 23164 12460 23204
rect 12500 23164 12509 23204
rect 12399 23099 12439 23164
rect 12748 23120 12788 23248
rect 12844 23120 12884 23332
rect 15724 23288 15764 23668
rect 17731 23584 17740 23624
rect 17780 23584 17932 23624
rect 17972 23584 17981 23624
rect 18953 23584 19075 23624
rect 19124 23584 19133 23624
rect 20803 23584 20812 23624
rect 20852 23584 22252 23624
rect 22292 23584 23060 23624
rect 23177 23584 23299 23624
rect 23348 23584 23357 23624
rect 23020 23540 23060 23584
rect 23404 23540 23444 23752
rect 24172 23708 24212 23836
rect 24268 23792 24308 23920
rect 24691 23836 24700 23876
rect 24740 23836 24940 23876
rect 24980 23836 24989 23876
rect 24364 23792 24404 23801
rect 25132 23792 25172 23920
rect 27244 23792 27284 24088
rect 28195 24004 28204 24044
rect 28244 24004 28492 24044
rect 28532 24004 28541 24044
rect 31145 24004 31276 24044
rect 31316 24004 31325 24044
rect 27523 23920 27532 23960
rect 27572 23920 29012 23960
rect 28972 23876 29012 23920
rect 27532 23836 28492 23876
rect 28532 23836 28541 23876
rect 28963 23836 28972 23876
rect 29012 23836 29021 23876
rect 30019 23836 30028 23876
rect 30068 23836 30077 23876
rect 27532 23792 27572 23836
rect 24259 23752 24268 23792
rect 24308 23752 24317 23792
rect 24451 23752 24460 23792
rect 24539 23752 24631 23792
rect 24835 23752 24844 23792
rect 24884 23752 24983 23792
rect 25023 23752 25032 23792
rect 25114 23752 25123 23792
rect 25163 23752 25172 23792
rect 25217 23752 25226 23792
rect 25266 23752 25275 23792
rect 25420 23752 25516 23792
rect 25556 23752 25565 23792
rect 25649 23752 25658 23792
rect 25698 23752 25804 23792
rect 25844 23752 25853 23792
rect 25900 23752 26188 23792
rect 26228 23752 26237 23792
rect 26371 23752 26380 23792
rect 26420 23752 26551 23792
rect 26659 23752 26668 23792
rect 26708 23752 26860 23792
rect 26900 23752 26909 23792
rect 27235 23752 27244 23792
rect 27284 23752 27293 23792
rect 27418 23752 27427 23792
rect 27467 23752 27476 23792
rect 27523 23752 27532 23792
rect 27572 23752 27581 23792
rect 27737 23752 27820 23792
rect 27860 23752 27868 23792
rect 27908 23752 27917 23792
rect 28002 23752 28011 23792
rect 28051 23752 28300 23792
rect 28340 23752 28387 23792
rect 28427 23752 28471 23792
rect 28649 23752 28698 23792
rect 28738 23752 28780 23792
rect 28820 23752 28829 23792
rect 29338 23752 29347 23792
rect 29396 23752 29527 23792
rect 23587 23668 23596 23708
rect 23636 23668 24062 23708
rect 24102 23668 24111 23708
rect 24154 23668 24163 23708
rect 24203 23668 24212 23708
rect 23683 23584 23692 23624
rect 23732 23584 24268 23624
rect 24308 23584 24317 23624
rect 15811 23500 15820 23540
rect 15860 23500 22348 23540
rect 22388 23500 22397 23540
rect 23020 23500 23444 23540
rect 24364 23540 24404 23752
rect 25228 23708 25268 23752
rect 24547 23668 24556 23708
rect 24596 23668 25268 23708
rect 25420 23624 25460 23752
rect 25900 23708 25940 23752
rect 25891 23668 25900 23708
rect 25940 23668 25949 23708
rect 24643 23584 24652 23624
rect 24692 23584 25315 23624
rect 25355 23584 25460 23624
rect 25795 23584 25804 23624
rect 25844 23584 25853 23624
rect 26057 23584 26188 23624
rect 26228 23584 26237 23624
rect 26441 23584 26563 23624
rect 26612 23584 26621 23624
rect 26729 23584 26860 23624
rect 26900 23584 26909 23624
rect 25804 23540 25844 23584
rect 26572 23540 26612 23584
rect 24364 23500 25844 23540
rect 26092 23500 26612 23540
rect 27436 23540 27476 23752
rect 28030 23668 28588 23708
rect 28628 23668 28637 23708
rect 27523 23584 27532 23624
rect 27572 23584 27916 23624
rect 27956 23584 27965 23624
rect 28030 23540 28070 23668
rect 28474 23584 28483 23624
rect 28523 23584 28684 23624
rect 28724 23584 28733 23624
rect 27436 23500 28070 23540
rect 26092 23456 26132 23500
rect 19891 23416 19900 23456
rect 20268 23416 20277 23456
rect 20419 23416 20428 23456
rect 20468 23416 25516 23456
rect 25556 23416 25565 23456
rect 26083 23416 26092 23456
rect 26132 23416 26141 23456
rect 27665 23416 27674 23456
rect 28042 23416 28051 23456
rect 24067 23332 24076 23372
rect 24116 23332 24460 23372
rect 24500 23332 24940 23372
rect 24980 23332 24989 23372
rect 15523 23248 15532 23288
rect 15572 23248 15581 23288
rect 15724 23248 16531 23288
rect 16571 23248 16588 23288
rect 16628 23248 16740 23288
rect 17923 23248 17932 23288
rect 17972 23248 20180 23288
rect 20297 23248 20332 23288
rect 20372 23248 20419 23288
rect 20459 23248 20477 23288
rect 23465 23248 23596 23288
rect 23636 23248 23645 23288
rect 23692 23248 25940 23288
rect 26947 23248 26956 23288
rect 26996 23248 27763 23288
rect 27803 23248 29356 23288
rect 29396 23248 29405 23288
rect 30979 23248 30988 23288
rect 31028 23248 31276 23288
rect 31316 23248 31325 23288
rect 15532 23204 15572 23248
rect 20140 23204 20180 23248
rect 23692 23204 23732 23248
rect 12931 23164 12940 23204
rect 12980 23164 13028 23204
rect 15532 23164 16108 23204
rect 16148 23164 18892 23204
rect 18932 23164 19276 23204
rect 19316 23164 19325 23204
rect 20140 23164 20612 23204
rect 12988 23120 13028 23164
rect 18316 23120 18356 23164
rect 20572 23120 20612 23164
rect 20716 23164 23732 23204
rect 24172 23164 24364 23204
rect 24404 23164 24413 23204
rect 25315 23164 25324 23204
rect 25364 23164 25844 23204
rect 20716 23120 20756 23164
rect 21538 23120 21578 23164
rect 21868 23120 21908 23164
rect 24172 23120 24212 23164
rect 25804 23120 25844 23164
rect 25900 23120 25940 23248
rect 25987 23164 25996 23204
rect 26036 23164 26324 23204
rect 26284 23120 26324 23164
rect 26554 23195 27148 23204
rect 26554 23155 26563 23195
rect 26603 23164 27148 23195
rect 27188 23164 27197 23204
rect 27427 23164 27436 23204
rect 27476 23164 30508 23204
rect 30548 23164 30557 23204
rect 26603 23155 26612 23164
rect 26554 23154 26612 23155
rect 27916 23120 27956 23164
rect 12308 23080 12317 23082
rect 4588 23036 4628 23080
rect 4291 22996 4300 23036
rect 4340 22996 5283 23036
rect 5323 22996 5548 23036
rect 5588 22996 5597 23036
rect 7075 22996 7084 23036
rect 7124 22996 7133 23036
rect 7337 22996 7468 23036
rect 7508 22996 7517 23036
rect 9091 22996 9100 23036
rect 9140 22996 9149 23036
rect 10313 22996 10348 23036
rect 10388 22996 10444 23036
rect 10484 22996 10493 23036
rect 11587 22996 11596 23036
rect 11636 22996 11732 23036
rect 11692 22952 11732 22996
rect 1961 22912 2092 22952
rect 2132 22912 2141 22952
rect 7721 22912 7852 22952
rect 7892 22912 7901 22952
rect 10723 22912 10732 22952
rect 10772 22912 11020 22952
rect 11060 22912 11069 22952
rect 11683 22912 11692 22952
rect 11732 22912 11741 22952
rect 11884 22868 11924 23080
rect 11980 23036 12020 23080
rect 12399 23059 12412 23099
rect 12452 23059 12461 23099
rect 12508 23080 12517 23120
rect 12596 23080 12697 23120
rect 12739 23080 12748 23120
rect 12788 23080 12797 23120
rect 12844 23080 12871 23120
rect 12911 23080 12920 23120
rect 12979 23080 12988 23120
rect 13028 23080 13037 23120
rect 13594 23080 13603 23120
rect 13652 23080 13783 23120
rect 16003 23080 16012 23120
rect 16052 23080 16726 23120
rect 16766 23080 16972 23120
rect 17012 23080 17021 23120
rect 17225 23080 17356 23120
rect 17396 23080 17405 23120
rect 17513 23111 17644 23120
rect 17513 23080 17635 23111
rect 17684 23080 17693 23120
rect 17779 23080 17788 23120
rect 17828 23080 17932 23120
rect 17972 23080 17981 23120
rect 18298 23080 18307 23120
rect 18347 23080 18356 23120
rect 18403 23080 18412 23120
rect 18452 23080 18583 23120
rect 18876 23080 18988 23120
rect 19028 23080 19036 23120
rect 19076 23080 19085 23120
rect 19171 23080 19180 23120
rect 19220 23080 19351 23120
rect 19776 23080 19843 23120
rect 19883 23080 19892 23120
rect 19939 23080 19948 23120
rect 19988 23080 20332 23120
rect 20372 23080 20381 23120
rect 20563 23080 20572 23120
rect 20612 23080 20621 23120
rect 20707 23080 20716 23120
rect 20756 23080 20765 23120
rect 20899 23080 20908 23120
rect 20948 23080 21292 23120
rect 21332 23080 21341 23120
rect 21520 23080 21529 23120
rect 21569 23080 21578 23120
rect 21662 23080 21671 23120
rect 21711 23080 21812 23120
rect 21859 23080 21868 23120
rect 21908 23080 21917 23120
rect 22121 23080 22252 23120
rect 22292 23080 22301 23120
rect 22915 23080 22924 23120
rect 22964 23080 23500 23120
rect 23540 23080 23549 23120
rect 23674 23080 23683 23120
rect 23732 23080 23863 23120
rect 24163 23080 24172 23120
rect 24212 23080 24221 23120
rect 24329 23080 24460 23120
rect 24500 23080 24509 23120
rect 24634 23080 24643 23120
rect 24692 23080 24823 23120
rect 24931 23080 24940 23120
rect 24980 23080 25219 23120
rect 25259 23080 25268 23120
rect 25385 23080 25507 23120
rect 25556 23080 25565 23120
rect 25795 23080 25804 23120
rect 25844 23080 25853 23120
rect 25900 23080 25996 23120
rect 26036 23080 26083 23120
rect 26277 23080 26286 23120
rect 26326 23080 26335 23120
rect 26380 23111 26420 23120
rect 17626 23071 17635 23080
rect 17675 23071 17684 23080
rect 17626 23070 17684 23071
rect 11971 22996 11980 23036
rect 12020 22996 12029 23036
rect 13219 22996 13228 23036
rect 13268 22996 13277 23036
rect 14659 22996 14668 23036
rect 14708 22996 14717 23036
rect 13228 22952 13268 22996
rect 18988 22952 19028 23080
rect 19852 23036 19892 23080
rect 19363 22996 19372 23036
rect 19412 22996 19892 23036
rect 11971 22912 11980 22952
rect 12020 22912 12460 22952
rect 12500 22912 12509 22952
rect 13027 22912 13036 22952
rect 13076 22912 13268 22952
rect 18586 22912 18595 22952
rect 18635 22912 19028 22952
rect 20572 22952 20612 23080
rect 21772 23036 21812 23080
rect 25996 23036 26036 23080
rect 26650 23080 26659 23120
rect 26699 23080 26755 23120
rect 26827 23080 26836 23120
rect 26900 23080 27016 23120
rect 27139 23080 27148 23120
rect 27188 23080 27197 23120
rect 27331 23080 27340 23120
rect 27380 23080 27860 23120
rect 27916 23080 27928 23120
rect 27968 23080 27977 23120
rect 28099 23080 28108 23120
rect 28148 23080 28724 23120
rect 28771 23080 28780 23120
rect 28820 23080 28972 23120
rect 29012 23080 29021 23120
rect 29338 23080 29347 23120
rect 29396 23080 29527 23120
rect 26380 23036 26420 23071
rect 26668 23036 26708 23080
rect 27148 23036 27188 23080
rect 21091 22996 21100 23036
rect 21140 22996 21196 23036
rect 21236 22996 21271 23036
rect 21402 22996 21411 23036
rect 21451 22996 21812 23036
rect 24307 22996 24316 23036
rect 24356 22996 24556 23036
rect 24596 22996 24605 23036
rect 25027 22996 25036 23036
rect 25076 22996 25268 23036
rect 21411 22952 21451 22996
rect 20572 22912 21451 22952
rect 24617 22912 24643 22952
rect 24683 22912 24748 22952
rect 24788 22912 24797 22952
rect 25228 22868 25268 22996
rect 25420 22996 25612 23036
rect 25652 22996 25661 23036
rect 25987 22996 25996 23036
rect 26036 22996 26045 23036
rect 26333 22996 26380 23036
rect 26420 22996 26429 23036
rect 26659 22996 26668 23036
rect 26708 22996 26717 23036
rect 27148 22996 27340 23036
rect 27380 22996 27389 23036
rect 2947 22828 2956 22868
rect 2996 22828 3628 22868
rect 3668 22828 3677 22868
rect 3763 22828 3772 22868
rect 3812 22828 8132 22868
rect 8179 22828 8188 22868
rect 8228 22828 8332 22868
rect 8372 22828 8381 22868
rect 10636 22828 11924 22868
rect 16771 22828 16780 22868
rect 16820 22828 16963 22868
rect 17003 22828 17012 22868
rect 19066 22828 19075 22868
rect 19115 22828 19564 22868
rect 19604 22828 19613 22868
rect 20122 22828 20131 22868
rect 20171 22828 20332 22868
rect 20372 22828 20381 22868
rect 21641 22828 21772 22868
rect 21812 22828 21821 22868
rect 25219 22828 25228 22868
rect 25268 22828 25277 22868
rect 8092 22784 8132 22828
rect 10636 22784 10676 22828
rect 8092 22744 10636 22784
rect 10676 22744 10685 22784
rect 25420 22700 25460 22996
rect 25673 22828 25804 22868
rect 25844 22828 25853 22868
rect 26266 22828 26275 22868
rect 26315 22828 26324 22868
rect 27113 22828 27244 22868
rect 27284 22828 27293 22868
rect 26284 22700 26324 22828
rect 27820 22784 27860 23080
rect 28684 22868 28724 23080
rect 29923 22996 29932 23036
rect 29972 22996 29981 23036
rect 28684 22828 30836 22868
rect 30883 22828 30892 22868
rect 30932 22828 30941 22868
rect 30796 22784 30836 22828
rect 27820 22744 28972 22784
rect 29012 22744 29021 22784
rect 30787 22744 30796 22784
rect 30836 22744 30845 22784
rect 30892 22700 30932 22828
rect 3103 22660 3112 22700
rect 3480 22660 3489 22700
rect 10877 22660 10886 22700
rect 11254 22660 11263 22700
rect 18651 22660 18660 22700
rect 19028 22660 19037 22700
rect 25420 22660 26324 22700
rect 26425 22660 26434 22700
rect 26802 22660 26811 22700
rect 30115 22660 30124 22700
rect 30164 22660 30932 22700
rect 12067 22576 12076 22616
rect 12116 22576 14476 22616
rect 14516 22576 14525 22616
rect 18604 22576 20180 22616
rect 18604 22532 18644 22576
rect 20140 22532 20180 22576
rect 25132 22576 27628 22616
rect 27668 22576 28204 22616
rect 28244 22576 30220 22616
rect 30260 22576 30269 22616
rect 25132 22532 25172 22576
rect 713 22492 844 22532
rect 884 22492 893 22532
rect 1420 22492 7660 22532
rect 7700 22492 7709 22532
rect 12739 22492 12748 22532
rect 12788 22492 14851 22532
rect 14891 22492 14900 22532
rect 18595 22492 18604 22532
rect 18644 22492 18653 22532
rect 19241 22492 19372 22532
rect 19412 22492 19421 22532
rect 20140 22492 24596 22532
rect 24643 22492 24652 22532
rect 24692 22492 25172 22532
rect 25219 22492 25228 22532
rect 25268 22492 25603 22532
rect 25643 22492 25652 22532
rect 0 22364 400 22384
rect 1420 22364 1460 22492
rect 24556 22448 24596 22492
rect 4003 22408 4012 22448
rect 4052 22408 6028 22448
rect 6068 22408 6077 22448
rect 6377 22408 6508 22448
rect 6548 22408 6557 22448
rect 8140 22408 9676 22448
rect 9716 22408 9725 22448
rect 10627 22408 10636 22448
rect 10676 22408 11356 22448
rect 11396 22408 11404 22448
rect 11444 22408 11556 22448
rect 12809 22408 12844 22448
rect 12884 22408 12940 22448
rect 12980 22408 12989 22448
rect 18700 22408 19276 22448
rect 19316 22408 19325 22448
rect 19747 22408 19756 22448
rect 19796 22408 22388 22448
rect 24556 22439 25028 22448
rect 24556 22408 24988 22439
rect 0 22324 1460 22364
rect 2083 22324 2092 22364
rect 2132 22324 2141 22364
rect 4253 22324 4300 22364
rect 4340 22324 4349 22364
rect 4396 22324 7516 22364
rect 7556 22324 7565 22364
rect 0 22304 400 22324
rect 4300 22280 4340 22324
rect 4396 22280 4436 22324
rect 8140 22280 8180 22408
rect 8506 22324 8515 22364
rect 8555 22324 8620 22364
rect 8660 22324 8695 22364
rect 10444 22324 12076 22364
rect 12116 22324 12125 22364
rect 12451 22324 12460 22364
rect 12500 22324 12966 22364
rect 10444 22280 10484 22324
rect 10924 22280 10964 22324
rect 12926 22280 12966 22324
rect 18700 22280 18740 22408
rect 22348 22364 22388 22408
rect 25193 22408 25219 22448
rect 25259 22408 25324 22448
rect 25364 22408 25373 22448
rect 25746 22408 26708 22448
rect 26921 22408 27052 22448
rect 27092 22408 27101 22448
rect 28474 22408 28483 22448
rect 28523 22408 30740 22448
rect 24988 22364 25028 22399
rect 25746 22364 25786 22408
rect 26668 22364 26708 22408
rect 30700 22364 30740 22408
rect 19075 22324 19084 22364
rect 19124 22324 19171 22364
rect 21292 22324 21772 22364
rect 21812 22324 21821 22364
rect 21868 22324 22292 22364
rect 22348 22324 22930 22364
rect 22970 22324 23540 22364
rect 19084 22280 19124 22324
rect 21292 22280 21332 22324
rect 21868 22280 21908 22324
rect 22252 22280 22292 22324
rect 23500 22280 23540 22324
rect 24460 22324 24844 22364
rect 24884 22324 24893 22364
rect 24988 22324 25786 22364
rect 25900 22324 26188 22364
rect 26228 22324 26237 22364
rect 26668 22324 27532 22364
rect 27572 22324 27581 22364
rect 28204 22324 28396 22364
rect 28436 22324 28445 22364
rect 30211 22324 30220 22364
rect 30260 22324 30548 22364
rect 30682 22324 30691 22364
rect 30731 22324 30740 22364
rect 30787 22324 30796 22364
rect 30836 22324 30892 22364
rect 30932 22324 30967 22364
rect 24460 22280 24500 22324
rect 25900 22322 25940 22324
rect 25882 22313 25940 22322
rect 2563 22240 2572 22280
rect 2612 22240 2755 22280
rect 2795 22240 2804 22280
rect 3497 22240 3619 22280
rect 3668 22240 3677 22280
rect 4282 22240 4291 22280
rect 4331 22240 4340 22280
rect 4387 22240 4396 22280
rect 4436 22240 4445 22280
rect 4841 22240 4972 22280
rect 5012 22240 5021 22280
rect 5539 22240 5548 22280
rect 5588 22240 5836 22280
rect 5876 22240 5885 22280
rect 6019 22240 6028 22280
rect 6068 22240 6199 22280
rect 7651 22240 7660 22280
rect 7700 22240 8044 22280
rect 8084 22240 8180 22280
rect 8244 22240 8332 22280
rect 8372 22240 8375 22280
rect 8415 22240 8424 22280
rect 8611 22240 8620 22280
rect 8660 22240 8716 22280
rect 8756 22240 8791 22280
rect 10147 22240 10156 22280
rect 10196 22240 10205 22280
rect 10435 22240 10444 22280
rect 10484 22240 10493 22280
rect 10804 22240 10813 22280
rect 10853 22240 10868 22280
rect 10915 22240 10924 22280
rect 10964 22240 10973 22280
rect 11299 22240 11308 22280
rect 11348 22240 11500 22280
rect 11540 22240 11549 22280
rect 11779 22240 11788 22280
rect 11828 22240 12172 22280
rect 12212 22240 12221 22280
rect 12307 22240 12316 22280
rect 12356 22240 12364 22280
rect 12404 22240 12487 22280
rect 12748 22240 12760 22280
rect 12800 22240 12809 22280
rect 12917 22240 12926 22280
rect 12966 22240 12975 22280
rect 13027 22240 13036 22280
rect 13076 22240 13085 22280
rect 13229 22240 13238 22280
rect 13278 22240 13324 22280
rect 13364 22240 13409 22280
rect 15113 22240 15244 22280
rect 15284 22240 15293 22280
rect 15977 22240 16099 22280
rect 16148 22240 16157 22280
rect 18691 22240 18700 22280
rect 18740 22240 18749 22280
rect 19066 22240 19075 22280
rect 19115 22240 19124 22280
rect 19171 22240 19180 22280
rect 19220 22240 19351 22280
rect 20969 22240 21100 22280
rect 21140 22240 21149 22280
rect 21283 22240 21292 22280
rect 21332 22240 21341 22280
rect 21388 22240 21431 22280
rect 21471 22240 21480 22280
rect 21562 22240 21571 22280
rect 21611 22240 21620 22280
rect 21667 22240 21676 22280
rect 21716 22240 21908 22280
rect 21955 22240 21964 22280
rect 22004 22240 22147 22280
rect 22187 22240 22196 22280
rect 22243 22240 22252 22280
rect 22292 22240 22423 22280
rect 23011 22240 23020 22280
rect 23060 22240 23069 22280
rect 23491 22240 23500 22280
rect 23540 22240 23549 22280
rect 23683 22240 23692 22280
rect 23732 22240 23863 22280
rect 24329 22240 24460 22280
rect 24500 22240 24509 22280
rect 24754 22240 24763 22280
rect 24803 22240 24812 22280
rect 25001 22240 25027 22280
rect 25067 22240 25132 22280
rect 25172 22240 25181 22280
rect 25882 22273 25891 22313
rect 25931 22273 25940 22313
rect 26668 22280 26708 22324
rect 28204 22280 28244 22324
rect 30508 22280 30548 22324
rect 25882 22272 25940 22273
rect 25987 22240 25996 22280
rect 26036 22240 26092 22280
rect 26132 22240 26176 22280
rect 26554 22240 26563 22280
rect 26603 22240 26612 22280
rect 26668 22240 26755 22280
rect 26795 22240 26804 22280
rect 27178 22240 27187 22280
rect 27227 22240 27293 22280
rect 27374 22240 27383 22280
rect 27423 22240 27432 22280
rect 27496 22240 27505 22280
rect 27545 22240 27572 22280
rect 27619 22240 27628 22280
rect 27668 22240 27724 22280
rect 27764 22240 27799 22280
rect 28073 22240 28108 22280
rect 28148 22240 28195 22280
rect 28235 22240 28244 22280
rect 28291 22240 28300 22280
rect 28340 22240 28349 22280
rect 29321 22240 29452 22280
rect 29492 22240 29501 22280
rect 30115 22240 30124 22280
rect 30164 22240 30412 22280
rect 30452 22240 30461 22280
rect 30508 22240 30551 22280
rect 30591 22240 30600 22280
rect 30787 22240 30796 22280
rect 30836 22240 30845 22280
rect 30953 22240 31084 22280
rect 31124 22240 31133 22280
rect 31267 22240 31276 22280
rect 31316 22240 31325 22280
rect 3130 22156 3139 22196
rect 3179 22156 4492 22196
rect 4532 22156 4541 22196
rect 4593 22156 4602 22196
rect 4642 22156 5932 22196
rect 5972 22156 5981 22196
rect 6028 22112 6068 22240
rect 10156 22196 10196 22240
rect 10828 22196 10868 22240
rect 8698 22156 8707 22196
rect 8747 22156 8908 22196
rect 8948 22156 8957 22196
rect 10156 22156 10868 22196
rect 5513 22072 5644 22112
rect 5684 22072 5693 22112
rect 6028 22072 9292 22112
rect 9332 22072 9341 22112
rect 9833 22072 9955 22112
rect 10004 22072 10013 22112
rect 10147 22072 10156 22112
rect 10196 22072 10627 22112
rect 10667 22072 10676 22112
rect 10828 22028 10868 22156
rect 12172 22112 12212 22240
rect 12748 22196 12788 22240
rect 13036 22196 13076 22240
rect 21388 22196 21428 22240
rect 21580 22196 21620 22240
rect 23020 22196 23060 22240
rect 23692 22196 23732 22240
rect 24763 22196 24803 22240
rect 26572 22196 26612 22240
rect 12521 22156 12595 22196
rect 12635 22156 12652 22196
rect 12692 22156 12701 22196
rect 12748 22156 12844 22196
rect 12884 22156 12893 22196
rect 12989 22156 13036 22196
rect 13076 22156 13085 22196
rect 16483 22156 16492 22196
rect 16532 22156 17644 22196
rect 17684 22156 17693 22196
rect 18892 22156 19386 22196
rect 19426 22156 20908 22196
rect 20948 22156 20957 22196
rect 21388 22156 21484 22196
rect 21524 22156 21533 22196
rect 21580 22156 22060 22196
rect 22100 22156 22109 22196
rect 23020 22156 23732 22196
rect 23971 22156 23980 22196
rect 24020 22156 24803 22196
rect 25891 22156 25900 22196
rect 25940 22156 26188 22196
rect 26228 22156 26612 22196
rect 18892 22112 18932 22156
rect 21580 22112 21620 22156
rect 27253 22112 27293 22240
rect 27375 22196 27415 22240
rect 27375 22156 27436 22196
rect 27476 22156 27485 22196
rect 12172 22072 16244 22112
rect 18473 22072 18595 22112
rect 18644 22072 18653 22112
rect 18883 22072 18892 22112
rect 18932 22072 18941 22112
rect 19756 22072 20620 22112
rect 20660 22072 20669 22112
rect 21274 22072 21283 22112
rect 21323 22072 21620 22112
rect 21754 22072 21763 22112
rect 21803 22072 21812 22112
rect 22409 22072 22540 22112
rect 22580 22072 22589 22112
rect 22714 22072 22723 22112
rect 22763 22072 22924 22112
rect 22964 22072 22973 22112
rect 23561 22072 23683 22112
rect 23732 22072 23741 22112
rect 25795 22072 25804 22112
rect 25844 22072 26107 22112
rect 26147 22072 26156 22112
rect 27253 22072 27340 22112
rect 27380 22072 27389 22112
rect 2860 21988 6412 22028
rect 6452 21988 6461 22028
rect 10828 21988 13228 22028
rect 13268 21988 13277 22028
rect 0 21944 400 21964
rect 2860 21944 2900 21988
rect 16204 21944 16244 22072
rect 19756 21944 19796 22072
rect 21772 22028 21812 22072
rect 27532 22028 27572 22240
rect 28300 22196 28340 22240
rect 30796 22196 30836 22240
rect 28300 22156 29731 22196
rect 29771 22156 29780 22196
rect 30796 22156 31180 22196
rect 31220 22156 31229 22196
rect 31276 22112 31316 22240
rect 28649 22072 28780 22112
rect 28820 22072 28829 22112
rect 31180 22072 31316 22112
rect 21772 21988 23500 22028
rect 23540 21988 23549 22028
rect 27331 21988 27340 22028
rect 27380 21988 31084 22028
rect 31124 21988 31133 22028
rect 31180 21944 31220 22072
rect 0 21904 2900 21944
rect 4343 21904 4352 21944
rect 4720 21904 4729 21944
rect 12117 21904 12126 21944
rect 12494 21904 12503 21944
rect 16204 21904 19796 21944
rect 19891 21904 19900 21944
rect 20268 21904 20277 21944
rect 20332 21904 25612 21944
rect 25652 21904 25661 21944
rect 26380 21904 27183 21944
rect 27665 21904 27674 21944
rect 28042 21904 28051 21944
rect 28387 21904 28396 21944
rect 28436 21904 31220 21944
rect 0 21884 400 21904
rect 20332 21860 20372 21904
rect 26380 21860 26420 21904
rect 2860 21820 17876 21860
rect 2860 21776 2900 21820
rect 17836 21776 17876 21820
rect 20044 21820 20372 21860
rect 20572 21820 26420 21860
rect 27143 21860 27183 21904
rect 27143 21820 30412 21860
rect 30452 21820 30461 21860
rect 20044 21776 20084 21820
rect 20572 21776 20612 21820
rect 355 21736 364 21776
rect 404 21736 2900 21776
rect 5260 21736 7756 21776
rect 7796 21736 7805 21776
rect 11683 21736 11692 21776
rect 11732 21736 12748 21776
rect 12788 21736 12797 21776
rect 13123 21736 13132 21776
rect 13172 21736 16579 21776
rect 16619 21736 16628 21776
rect 17338 21736 17347 21776
rect 17387 21736 17740 21776
rect 17780 21736 17789 21776
rect 17836 21736 18172 21776
rect 18212 21736 18221 21776
rect 20026 21736 20035 21776
rect 20075 21736 20084 21776
rect 4186 21652 4195 21692
rect 4235 21652 4972 21692
rect 5012 21652 5021 21692
rect 5260 21608 5300 21736
rect 5434 21652 5443 21692
rect 5483 21652 5644 21692
rect 5684 21652 5693 21692
rect 9100 21652 9908 21692
rect 643 21568 652 21608
rect 692 21568 1708 21608
rect 1748 21568 2860 21608
rect 2900 21568 2909 21608
rect 3977 21568 4108 21608
rect 4148 21568 4157 21608
rect 4282 21568 4291 21608
rect 4331 21568 4340 21608
rect 0 21524 400 21544
rect 0 21484 4012 21524
rect 4052 21484 4061 21524
rect 0 21464 400 21484
rect 4300 21440 4340 21568
rect 4393 21536 4402 21576
rect 4442 21536 4457 21576
rect 4570 21568 4579 21608
rect 4619 21568 4684 21608
rect 4724 21568 4759 21608
rect 4860 21568 4869 21608
rect 4909 21568 5012 21608
rect 5059 21568 5068 21608
rect 5108 21568 5117 21608
rect 5251 21568 5260 21608
rect 5300 21568 5309 21608
rect 5818 21568 5827 21608
rect 5867 21568 8812 21608
rect 8852 21568 8861 21608
rect 4417 21524 4457 21536
rect 4972 21524 5012 21568
rect 5068 21524 5108 21568
rect 9100 21524 9140 21652
rect 9868 21608 9908 21652
rect 17740 21608 17780 21736
rect 20044 21692 20084 21736
rect 20140 21736 20275 21776
rect 20315 21736 20612 21776
rect 21833 21736 21964 21776
rect 22004 21736 22013 21776
rect 22243 21736 22252 21776
rect 22292 21736 22780 21776
rect 22820 21736 22829 21776
rect 24931 21736 24940 21776
rect 24980 21736 25228 21776
rect 25268 21736 25277 21776
rect 25498 21736 25507 21776
rect 25547 21736 26092 21776
rect 26132 21736 26228 21776
rect 20140 21692 20180 21736
rect 26188 21692 26228 21736
rect 26956 21736 27340 21776
rect 27380 21736 27389 21776
rect 28841 21736 28972 21776
rect 29012 21736 29021 21776
rect 29443 21736 29452 21776
rect 29492 21736 29923 21776
rect 29963 21736 29972 21776
rect 30211 21736 30220 21776
rect 30260 21736 30460 21776
rect 30500 21736 30892 21776
rect 30932 21736 30941 21776
rect 19843 21652 19852 21692
rect 19892 21652 20084 21692
rect 20131 21652 20140 21692
rect 20180 21652 20189 21692
rect 21379 21652 21388 21692
rect 21428 21652 23980 21692
rect 24020 21652 24820 21692
rect 20044 21608 20084 21652
rect 9187 21568 9196 21608
rect 9236 21568 9245 21608
rect 9379 21568 9388 21608
rect 9428 21568 9772 21608
rect 9812 21568 9821 21608
rect 9868 21568 11212 21608
rect 11252 21568 11261 21608
rect 11491 21568 11500 21608
rect 11540 21599 11692 21608
rect 11540 21568 11587 21599
rect 4417 21484 4916 21524
rect 4963 21484 4972 21524
rect 5012 21484 5021 21524
rect 5068 21484 5356 21524
rect 5396 21484 5405 21524
rect 6499 21484 6508 21524
rect 6548 21484 6557 21524
rect 7180 21484 9140 21524
rect 9196 21524 9236 21568
rect 11578 21559 11587 21568
rect 11627 21568 11692 21599
rect 11732 21568 11796 21608
rect 11875 21568 11884 21608
rect 11924 21568 13036 21608
rect 13076 21568 13085 21608
rect 13193 21568 13324 21608
rect 13364 21568 13373 21608
rect 13481 21568 13612 21608
rect 13652 21568 13661 21608
rect 14092 21568 16108 21608
rect 16148 21568 16867 21608
rect 16907 21568 16916 21608
rect 17513 21568 17635 21608
rect 17684 21568 17693 21608
rect 17740 21599 18068 21608
rect 17740 21568 18019 21599
rect 11627 21559 11636 21568
rect 11578 21558 11636 21559
rect 14092 21524 14132 21568
rect 18010 21559 18019 21568
rect 18059 21559 18068 21599
rect 18979 21568 18988 21608
rect 19028 21568 19276 21608
rect 19316 21568 19372 21608
rect 19412 21568 19421 21608
rect 19817 21568 19948 21608
rect 19988 21568 19997 21608
rect 20044 21568 20332 21608
rect 20372 21568 20381 21608
rect 20524 21568 20995 21608
rect 21035 21568 21044 21608
rect 21571 21568 21580 21608
rect 21620 21568 21868 21608
rect 21908 21568 21917 21608
rect 22042 21568 22051 21608
rect 22100 21568 22231 21608
rect 22793 21568 22924 21608
rect 22964 21568 22973 21608
rect 24521 21568 24652 21608
rect 24692 21568 24701 21608
rect 24780 21605 24820 21652
rect 26188 21652 26380 21692
rect 26420 21652 26429 21692
rect 26524 21652 26860 21692
rect 26900 21652 26909 21692
rect 26188 21608 26228 21652
rect 26524 21608 26564 21652
rect 26956 21608 26996 21736
rect 28972 21692 29012 21736
rect 27340 21652 28108 21692
rect 28148 21652 28157 21692
rect 28483 21652 28492 21692
rect 28532 21652 28916 21692
rect 28972 21652 29822 21692
rect 29862 21652 29871 21692
rect 30019 21652 30028 21692
rect 30068 21652 30931 21692
rect 30971 21652 30980 21692
rect 27340 21608 27380 21652
rect 18010 21558 18068 21559
rect 9196 21484 9682 21524
rect 9722 21484 9964 21524
rect 10004 21484 10013 21524
rect 10723 21484 10732 21524
rect 10772 21484 11308 21524
rect 11348 21484 11357 21524
rect 11770 21484 11779 21524
rect 11819 21484 12364 21524
rect 12404 21484 14132 21524
rect 14188 21484 16060 21524
rect 16100 21484 16109 21524
rect 16291 21484 16300 21524
rect 16340 21484 16349 21524
rect 16474 21484 16483 21524
rect 16532 21484 16868 21524
rect 16937 21484 17059 21524
rect 17108 21484 17117 21524
rect 17242 21484 17251 21524
rect 17291 21484 17548 21524
rect 17588 21484 17597 21524
rect 17705 21484 17827 21524
rect 17876 21484 17885 21524
rect 4876 21440 4916 21484
rect 2537 21400 2572 21440
rect 2612 21400 2668 21440
rect 2708 21400 2717 21440
rect 4300 21400 4532 21440
rect 4867 21400 4876 21440
rect 4916 21400 4925 21440
rect 5155 21400 5164 21440
rect 5204 21400 5213 21440
rect 4492 21356 4532 21400
rect 5164 21356 5204 21400
rect 7180 21356 7220 21484
rect 14188 21440 14228 21484
rect 16300 21440 16340 21484
rect 16828 21440 16868 21484
rect 17260 21440 17300 21484
rect 20524 21440 20564 21568
rect 21004 21524 21044 21568
rect 24771 21565 24780 21605
rect 24820 21565 24829 21605
rect 25481 21568 25516 21608
rect 25556 21568 25612 21608
rect 25652 21568 25661 21608
rect 25900 21568 25996 21608
rect 26036 21568 26045 21608
rect 26179 21568 26188 21608
rect 26228 21568 26237 21608
rect 26284 21568 26385 21608
rect 26425 21568 26434 21608
rect 26506 21568 26515 21608
rect 26555 21568 26564 21608
rect 26611 21568 26620 21608
rect 26660 21568 26669 21608
rect 26719 21599 26996 21608
rect 21004 21484 22348 21524
rect 22388 21484 22397 21524
rect 25123 21484 25132 21524
rect 25172 21484 25181 21524
rect 7948 21400 8948 21440
rect 8995 21400 9004 21440
rect 9044 21400 9812 21440
rect 10435 21400 10444 21440
rect 10484 21400 11404 21440
rect 11444 21400 11453 21440
rect 11971 21400 11980 21440
rect 12020 21400 12305 21440
rect 12355 21400 12364 21440
rect 12404 21400 14228 21440
rect 14345 21400 14476 21440
rect 14516 21400 14525 21440
rect 16300 21400 16579 21440
rect 16619 21400 16628 21440
rect 16828 21400 17300 21440
rect 17356 21400 19756 21440
rect 19796 21400 19805 21440
rect 20515 21400 20524 21440
rect 20564 21400 20573 21440
rect 22313 21400 22444 21440
rect 22484 21400 22493 21440
rect 7948 21356 7988 21400
rect 8908 21356 8948 21400
rect 9772 21356 9812 21400
rect 12265 21356 12305 21400
rect 17356 21356 17396 21400
rect 2371 21316 2380 21356
rect 2420 21316 2764 21356
rect 2804 21316 2813 21356
rect 4492 21316 5068 21356
rect 5108 21316 5117 21356
rect 5164 21316 7220 21356
rect 7267 21316 7276 21356
rect 7316 21316 7372 21356
rect 7412 21316 7447 21356
rect 7747 21316 7756 21356
rect 7796 21316 7948 21356
rect 7988 21316 7997 21356
rect 8323 21316 8332 21356
rect 8372 21316 8803 21356
rect 8843 21316 8852 21356
rect 8908 21316 9388 21356
rect 9428 21316 9437 21356
rect 9545 21316 9667 21356
rect 9716 21316 9725 21356
rect 9772 21316 12124 21356
rect 12164 21316 12173 21356
rect 12265 21316 12988 21356
rect 13028 21316 13037 21356
rect 16387 21316 16396 21356
rect 16436 21316 17396 21356
rect 19049 21316 19180 21356
rect 19220 21316 19229 21356
rect 20995 21316 21004 21356
rect 21044 21316 21196 21356
rect 21236 21316 21245 21356
rect 1987 21232 1996 21272
rect 2036 21232 24748 21272
rect 24788 21232 24797 21272
rect 3103 21148 3112 21188
rect 3480 21148 3489 21188
rect 4675 21148 4684 21188
rect 4724 21148 9004 21188
rect 9044 21148 9053 21188
rect 10877 21148 10886 21188
rect 11254 21148 11263 21188
rect 11395 21148 11404 21188
rect 11444 21148 16396 21188
rect 16436 21148 16445 21188
rect 18651 21148 18660 21188
rect 19028 21148 19037 21188
rect 0 21104 400 21124
rect 0 21064 4052 21104
rect 4099 21064 4108 21104
rect 4148 21064 12364 21104
rect 12404 21064 12413 21104
rect 12940 21064 24652 21104
rect 24692 21064 24701 21104
rect 0 21044 400 21064
rect 521 20980 652 21020
rect 692 20980 701 21020
rect 4012 20936 4052 21064
rect 12940 21020 12980 21064
rect 25132 21020 25172 21484
rect 25363 21400 25372 21440
rect 25412 21400 25804 21440
rect 25844 21400 25853 21440
rect 25673 21316 25708 21356
rect 25748 21316 25804 21356
rect 25844 21316 25853 21356
rect 25900 21020 25940 21568
rect 26284 21524 26324 21568
rect 26620 21524 26660 21568
rect 26759 21568 26996 21599
rect 27139 21568 27148 21608
rect 27188 21568 27197 21608
rect 27322 21568 27331 21608
rect 27371 21568 27380 21608
rect 27427 21568 27436 21608
rect 27476 21568 27523 21608
rect 27563 21568 27628 21608
rect 27668 21568 27677 21608
rect 27811 21568 27820 21608
rect 27860 21568 27869 21608
rect 28099 21568 28108 21608
rect 28148 21568 28244 21608
rect 28290 21568 28299 21608
rect 28339 21568 28348 21608
rect 28474 21568 28483 21608
rect 28523 21568 28532 21608
rect 28579 21568 28588 21608
rect 28628 21568 28759 21608
rect 26719 21550 26759 21559
rect 26275 21484 26284 21524
rect 26324 21484 26333 21524
rect 26563 21484 26572 21524
rect 26612 21484 26660 21524
rect 27148 21524 27188 21568
rect 27820 21524 27860 21568
rect 27148 21484 27340 21524
rect 27380 21484 27389 21524
rect 27820 21484 28148 21524
rect 27139 21400 27148 21440
rect 27188 21400 27820 21440
rect 27860 21400 27869 21440
rect 25987 21316 25996 21356
rect 26036 21316 26167 21356
rect 26659 21316 26668 21356
rect 26708 21316 26717 21356
rect 27322 21316 27331 21356
rect 27371 21316 28012 21356
rect 28052 21316 28061 21356
rect 26668 21272 26708 21316
rect 28108 21272 28148 21484
rect 28204 21440 28244 21568
rect 28300 21524 28340 21568
rect 28492 21524 28532 21568
rect 28876 21524 28916 21652
rect 29513 21568 29644 21608
rect 29684 21568 29693 21608
rect 30124 21599 30164 21608
rect 30124 21524 30164 21559
rect 30298 21599 30508 21608
rect 30298 21559 30307 21599
rect 30347 21568 30508 21599
rect 30548 21568 30557 21608
rect 30974 21568 30988 21608
rect 31028 21568 31096 21608
rect 31136 21568 31154 21608
rect 30347 21559 30356 21568
rect 30298 21558 30356 21559
rect 28291 21484 28300 21524
rect 28340 21484 28386 21524
rect 28492 21484 28780 21524
rect 28820 21484 28829 21524
rect 28876 21484 30164 21524
rect 28204 21400 30220 21440
rect 30260 21400 30269 21440
rect 28579 21316 28588 21356
rect 28628 21316 28780 21356
rect 28820 21316 28829 21356
rect 26668 21232 27436 21272
rect 27476 21232 27485 21272
rect 28108 21232 30124 21272
rect 30164 21232 30173 21272
rect 26425 21148 26434 21188
rect 26802 21148 26811 21188
rect 4963 20980 4972 21020
rect 5012 20980 6220 21020
rect 6260 20980 6269 21020
rect 8044 20980 11212 21020
rect 11252 20980 11261 21020
rect 11491 20980 11500 21020
rect 11540 20980 12980 21020
rect 13603 20980 13612 21020
rect 13652 20980 15052 21020
rect 15092 20980 15724 21020
rect 15764 20980 15773 21020
rect 16099 20980 16108 21020
rect 16148 20980 23404 21020
rect 23444 20980 23453 21020
rect 23683 20980 23692 21020
rect 23732 20980 25172 21020
rect 25891 20980 25900 21020
rect 25940 20980 25949 21020
rect 25996 20980 26572 21020
rect 26612 20980 26621 21020
rect 26755 20980 26764 21020
rect 26804 20980 26860 21020
rect 26900 20980 26935 21020
rect 27427 20980 27436 21020
rect 27476 20980 27572 21020
rect 28073 20980 28204 21020
rect 28244 20980 28588 21020
rect 28628 20980 28637 21020
rect 29635 20980 29644 21020
rect 29684 20980 31276 21020
rect 31316 20980 31325 21020
rect 8044 20936 8084 20980
rect 3763 20896 3772 20936
rect 3812 20896 3956 20936
rect 4012 20896 8084 20936
rect 8140 20896 9244 20936
rect 9284 20896 9293 20936
rect 10828 20896 11404 20936
rect 11444 20896 11540 20936
rect 11674 20896 11683 20936
rect 11723 20896 11980 20936
rect 12020 20896 12029 20936
rect 13219 20896 13228 20936
rect 13268 20896 13460 20936
rect 3916 20852 3956 20896
rect 8140 20852 8180 20896
rect 10828 20852 10868 20896
rect 11500 20852 11540 20896
rect 13420 20852 13460 20896
rect 15820 20896 16588 20936
rect 16628 20896 21524 20936
rect 2659 20812 2668 20852
rect 2708 20812 2717 20852
rect 3916 20812 4340 20852
rect 4474 20812 4483 20852
rect 4523 20812 5443 20852
rect 5483 20812 5740 20852
rect 5780 20812 5789 20852
rect 6892 20812 7180 20852
rect 7220 20812 7229 20852
rect 7843 20812 7852 20852
rect 7892 20812 8131 20852
rect 8171 20812 8180 20852
rect 8873 20812 9004 20852
rect 9044 20812 9053 20852
rect 10339 20812 10348 20852
rect 10388 20812 10819 20852
rect 10859 20812 10868 20852
rect 11386 20812 11395 20852
rect 11435 20812 11444 20852
rect 11500 20812 11587 20852
rect 11627 20812 11636 20852
rect 11683 20812 11692 20852
rect 11732 20812 12163 20852
rect 12203 20812 12212 20852
rect 13411 20812 13420 20852
rect 13460 20812 13469 20852
rect 14467 20812 14476 20852
rect 14516 20812 14525 20852
rect 15139 20812 15148 20852
rect 15188 20812 15340 20852
rect 15380 20812 15389 20852
rect 4300 20768 4340 20812
rect 6892 20768 6932 20812
rect 11404 20768 11444 20812
rect 15820 20768 15860 20896
rect 16291 20812 16300 20852
rect 16340 20812 16492 20852
rect 16532 20812 16541 20852
rect 17129 20812 17260 20852
rect 17300 20812 17309 20852
rect 17539 20812 17548 20852
rect 17588 20812 17836 20852
rect 17876 20812 17885 20852
rect 19267 20812 19276 20852
rect 19355 20812 19447 20852
rect 19660 20812 20140 20852
rect 20180 20812 20189 20852
rect 20515 20812 20524 20852
rect 20564 20812 20643 20852
rect 20683 20812 20695 20852
rect 20873 20812 20995 20852
rect 21044 20812 21053 20852
rect 19660 20768 19700 20812
rect 2441 20728 2563 20768
rect 2612 20728 2621 20768
rect 2851 20728 2860 20768
rect 2900 20728 3148 20768
rect 3188 20728 3197 20768
rect 3427 20728 3436 20768
rect 3476 20728 3532 20768
rect 3572 20728 4204 20768
rect 4244 20728 4253 20768
rect 4300 20728 4436 20768
rect 4553 20728 4684 20768
rect 4724 20728 4733 20768
rect 5172 20728 5260 20768
rect 5300 20728 5303 20768
rect 5343 20728 5396 20768
rect 5443 20728 5452 20768
rect 5492 20728 5548 20768
rect 5588 20728 6740 20768
rect 6883 20728 6892 20768
rect 6932 20728 6941 20768
rect 7267 20728 7276 20768
rect 7316 20728 8011 20768
rect 8084 20728 8093 20768
rect 8227 20728 8236 20768
rect 8276 20728 10444 20768
rect 10484 20728 10493 20768
rect 10540 20728 10563 20768
rect 10603 20728 10612 20768
rect 10672 20728 10681 20768
rect 10721 20728 10732 20768
rect 10772 20728 10861 20768
rect 11194 20728 11203 20768
rect 11243 20728 11252 20768
rect 11404 20728 11596 20768
rect 11636 20728 11645 20768
rect 11962 20728 11971 20768
rect 12011 20728 12020 20768
rect 12547 20728 12556 20768
rect 12596 20728 12605 20768
rect 12826 20728 12835 20768
rect 12875 20728 13556 20768
rect 13786 20728 13795 20768
rect 13835 20728 15860 20768
rect 15950 20728 15959 20768
rect 15999 20728 16008 20768
rect 16090 20728 16099 20768
rect 16139 20728 16148 20768
rect 16195 20728 16204 20768
rect 16244 20728 16396 20768
rect 16436 20728 16445 20768
rect 17434 20728 17443 20768
rect 17483 20728 17492 20768
rect 17722 20728 17731 20768
rect 17771 20728 17932 20768
rect 18011 20728 18132 20768
rect 19501 20728 19510 20768
rect 19550 20728 19604 20768
rect 19651 20728 19660 20768
rect 19700 20728 19709 20768
rect 19843 20728 19852 20768
rect 19892 20728 20023 20768
rect 20393 20728 20428 20768
rect 20468 20728 20524 20768
rect 20564 20728 20573 20768
rect 20620 20728 20741 20768
rect 20781 20728 20790 20768
rect 20861 20728 20875 20768
rect 20915 20728 20948 20768
rect 0 20684 400 20704
rect 4396 20684 4436 20728
rect 5356 20684 5396 20728
rect 6700 20684 6740 20728
rect 8236 20684 8276 20728
rect 10540 20684 10580 20728
rect 11212 20684 11252 20728
rect 11980 20684 12020 20728
rect 0 20644 1228 20684
rect 1268 20644 1277 20684
rect 2938 20644 2947 20684
rect 2996 20644 3127 20684
rect 4169 20644 4291 20684
rect 4340 20644 4349 20684
rect 4396 20644 5164 20684
rect 5204 20644 5213 20684
rect 5356 20644 6316 20684
rect 6356 20644 6365 20684
rect 6700 20644 8276 20684
rect 9235 20644 9244 20684
rect 9284 20644 11020 20684
rect 11060 20644 11069 20684
rect 11212 20644 12020 20684
rect 12556 20684 12596 20728
rect 13516 20684 13556 20728
rect 15959 20684 15999 20728
rect 12556 20644 12748 20684
rect 12788 20644 12797 20684
rect 12931 20644 12940 20684
rect 12980 20644 13111 20684
rect 13516 20644 14380 20684
rect 14420 20644 14429 20684
rect 15907 20644 15916 20684
rect 15956 20644 15999 20684
rect 16108 20684 16148 20728
rect 17452 20684 17492 20728
rect 19564 20684 19604 20728
rect 20620 20684 20660 20728
rect 20908 20684 20948 20728
rect 21004 20728 21100 20768
rect 21140 20728 21149 20768
rect 21484 20749 21524 20896
rect 22435 20812 22444 20852
rect 22484 20812 22493 20852
rect 23884 20768 23924 20980
rect 25996 20936 26036 20980
rect 24931 20896 24940 20936
rect 24980 20896 25036 20936
rect 25076 20896 25111 20936
rect 25612 20896 26036 20936
rect 26083 20896 26092 20936
rect 26132 20896 26324 20936
rect 25612 20852 25652 20896
rect 24163 20812 24172 20852
rect 24212 20812 25612 20852
rect 25652 20812 25661 20852
rect 25738 20843 25804 20852
rect 25738 20803 25747 20843
rect 25787 20812 25804 20843
rect 25844 20812 26132 20852
rect 25787 20803 25796 20812
rect 25738 20802 25796 20803
rect 26092 20768 26132 20812
rect 26284 20768 26324 20896
rect 26369 20810 26409 20980
rect 26467 20896 26476 20936
rect 26516 20896 26612 20936
rect 26659 20896 26668 20936
rect 26708 20896 27476 20936
rect 26572 20852 26612 20896
rect 27436 20852 27476 20896
rect 26572 20812 27188 20852
rect 27235 20812 27244 20852
rect 27284 20812 27327 20852
rect 27418 20812 27427 20852
rect 27467 20812 27476 20852
rect 26369 20801 26412 20810
rect 26369 20770 26372 20801
rect 21676 20749 21763 20768
rect 21484 20728 21763 20749
rect 21803 20728 21812 20768
rect 23875 20728 23884 20768
rect 23924 20728 23933 20768
rect 24547 20728 24556 20768
rect 24596 20728 24835 20768
rect 24875 20728 24884 20768
rect 25507 20728 25516 20768
rect 25556 20728 25687 20768
rect 25846 20728 25855 20768
rect 25895 20728 25900 20768
rect 25940 20728 26035 20768
rect 26083 20728 26092 20768
rect 26132 20728 26141 20768
rect 26245 20728 26254 20768
rect 26294 20728 26324 20768
rect 27148 20768 27188 20812
rect 27287 20768 27327 20812
rect 27532 20768 27572 20980
rect 28003 20812 28012 20852
rect 28052 20812 28148 20852
rect 28291 20812 28300 20852
rect 28340 20812 28588 20852
rect 28628 20812 28637 20852
rect 28771 20812 28780 20852
rect 28820 20812 28972 20852
rect 29012 20812 29021 20852
rect 30595 20812 30604 20852
rect 30644 20812 30653 20852
rect 28108 20768 28148 20812
rect 26372 20752 26412 20761
rect 26465 20728 26474 20768
rect 26516 20728 26647 20768
rect 26860 20728 26903 20768
rect 26943 20728 26952 20768
rect 27034 20759 27092 20768
rect 16108 20644 17644 20684
rect 17684 20644 18988 20684
rect 19028 20644 19037 20684
rect 19564 20644 19756 20684
rect 19796 20644 19805 20684
rect 19939 20644 19948 20684
rect 19988 20644 20428 20684
rect 20468 20644 20477 20684
rect 20611 20644 20620 20684
rect 20660 20644 20669 20684
rect 20899 20644 20908 20684
rect 20948 20644 20957 20684
rect 0 20624 400 20644
rect 5539 20560 5548 20600
rect 5588 20560 5635 20600
rect 5675 20560 5719 20600
rect 8131 20560 8140 20600
rect 8180 20560 8323 20600
rect 8363 20560 8372 20600
rect 10793 20560 10915 20600
rect 10964 20560 10973 20600
rect 11212 20516 11252 20644
rect 21004 20600 21044 20728
rect 21484 20709 21716 20728
rect 21178 20644 21187 20684
rect 21227 20644 21379 20684
rect 21419 20644 21428 20684
rect 24547 20644 24556 20684
rect 24596 20644 25172 20684
rect 25132 20600 25172 20644
rect 26860 20600 26900 20728
rect 27034 20719 27043 20759
rect 27083 20719 27092 20759
rect 27139 20728 27148 20768
rect 27188 20728 27197 20768
rect 27278 20728 27287 20768
rect 27327 20728 27336 20768
rect 27523 20728 27532 20768
rect 27572 20728 27581 20768
rect 27689 20728 27820 20768
rect 27860 20728 27869 20768
rect 28012 20728 28021 20768
rect 28061 20728 28148 20768
rect 28195 20728 28204 20768
rect 28244 20728 28253 20768
rect 28361 20728 28492 20768
rect 28532 20728 28541 20768
rect 29338 20728 29347 20768
rect 29387 20728 30220 20768
rect 30260 20728 30269 20768
rect 27034 20718 27092 20719
rect 27052 20600 27092 20718
rect 28204 20684 28244 20728
rect 27427 20644 27436 20684
rect 27476 20644 28244 20684
rect 14083 20560 14092 20600
rect 14132 20560 18172 20600
rect 18212 20560 18221 20600
rect 21004 20560 22636 20600
rect 22676 20560 25036 20600
rect 25076 20560 25085 20600
rect 25132 20560 25612 20600
rect 25652 20560 25661 20600
rect 25795 20560 25804 20600
rect 25844 20560 26900 20600
rect 27043 20560 27052 20600
rect 27092 20560 27101 20600
rect 27331 20560 27340 20600
rect 27380 20560 27619 20600
rect 27659 20560 27668 20600
rect 27811 20560 27820 20600
rect 27860 20560 28300 20600
rect 28340 20560 28349 20600
rect 10060 20476 11252 20516
rect 11875 20476 11884 20516
rect 11924 20476 23444 20516
rect 10060 20432 10100 20476
rect 451 20392 460 20432
rect 500 20392 4244 20432
rect 4343 20392 4352 20432
rect 4720 20392 4729 20432
rect 8995 20392 9004 20432
rect 9044 20392 10100 20432
rect 12117 20392 12126 20432
rect 12494 20392 12503 20432
rect 19891 20392 19900 20432
rect 20268 20392 20277 20432
rect 4204 20348 4244 20392
rect 23404 20348 23444 20476
rect 24652 20392 25172 20432
rect 27665 20392 27674 20432
rect 28042 20392 28051 20432
rect 1315 20308 1324 20348
rect 1364 20308 4108 20348
rect 4148 20308 4157 20348
rect 4204 20308 11980 20348
rect 12020 20308 12029 20348
rect 19171 20308 19180 20348
rect 19220 20308 23060 20348
rect 23404 20308 24556 20348
rect 24596 20308 24605 20348
rect 0 20264 400 20284
rect 23020 20264 23060 20308
rect 24652 20264 24692 20392
rect 24739 20308 24748 20348
rect 24788 20308 25076 20348
rect 25036 20264 25076 20308
rect 0 20224 1420 20264
rect 1460 20224 1469 20264
rect 1516 20224 10924 20264
rect 10964 20224 10973 20264
rect 12730 20224 12739 20264
rect 12779 20224 12788 20264
rect 13289 20224 13411 20264
rect 13460 20224 13469 20264
rect 14467 20224 14476 20264
rect 14516 20224 15715 20264
rect 15755 20224 15764 20264
rect 16771 20224 16780 20264
rect 16820 20224 17068 20264
rect 17108 20224 17117 20264
rect 17251 20224 17260 20264
rect 17300 20224 17539 20264
rect 17579 20224 17588 20264
rect 17705 20224 17740 20264
rect 17780 20224 17836 20264
rect 17876 20224 17885 20264
rect 20371 20224 20380 20264
rect 20420 20224 20908 20264
rect 20948 20224 20957 20264
rect 23020 20224 24692 20264
rect 25018 20224 25027 20264
rect 25067 20224 25076 20264
rect 25132 20264 25172 20392
rect 25219 20308 25228 20348
rect 25268 20308 26764 20348
rect 26804 20308 26813 20348
rect 26860 20308 27052 20348
rect 27092 20308 27101 20348
rect 26860 20264 26900 20308
rect 25132 20224 26668 20264
rect 26708 20224 26717 20264
rect 26851 20224 26860 20264
rect 26900 20224 26909 20264
rect 27017 20224 27139 20264
rect 27188 20224 27197 20264
rect 27427 20224 27436 20264
rect 27476 20224 31180 20264
rect 31220 20224 31284 20264
rect 0 20204 400 20224
rect 1516 20180 1556 20224
rect 12748 20180 12788 20224
rect 931 20140 940 20180
rect 980 20140 1556 20180
rect 2188 20140 2668 20180
rect 2708 20140 3436 20180
rect 3476 20140 3820 20180
rect 3860 20140 3869 20180
rect 6691 20140 6700 20180
rect 6740 20140 6871 20180
rect 8515 20140 8524 20180
rect 8564 20140 8707 20180
rect 8747 20140 8756 20180
rect 10051 20140 10060 20180
rect 10100 20140 13516 20180
rect 13556 20140 13844 20180
rect 14249 20140 14371 20180
rect 14420 20140 14429 20180
rect 16483 20140 16492 20180
rect 16532 20140 17972 20180
rect 18979 20140 18988 20180
rect 19028 20140 19037 20180
rect 19468 20140 23116 20180
rect 23156 20140 23165 20180
rect 24652 20140 25364 20180
rect 2188 20096 2228 20140
rect 13804 20096 13844 20140
rect 17932 20096 17972 20140
rect 1673 20056 1804 20096
rect 1844 20056 1853 20096
rect 2032 20056 2041 20096
rect 2081 20056 2228 20096
rect 2275 20056 2284 20096
rect 2324 20056 2455 20096
rect 2537 20056 2563 20096
rect 2603 20056 2668 20096
rect 2708 20056 2717 20096
rect 2851 20056 2860 20096
rect 2900 20056 3379 20096
rect 3419 20056 3428 20096
rect 3497 20056 3574 20096
rect 3614 20056 3628 20096
rect 3668 20056 3677 20096
rect 3785 20056 3820 20096
rect 3860 20056 3916 20096
rect 3956 20056 3965 20096
rect 4048 20056 4057 20096
rect 4097 20056 4300 20096
rect 4340 20056 4349 20096
rect 4483 20056 4492 20096
rect 4532 20056 4663 20096
rect 5033 20056 5155 20096
rect 5204 20056 5923 20096
rect 5963 20056 5972 20096
rect 6316 20056 6494 20096
rect 6534 20056 6543 20096
rect 6796 20087 6836 20096
rect 6316 20012 6356 20056
rect 6979 20056 6988 20096
rect 7028 20056 7084 20096
rect 7124 20056 7159 20096
rect 7267 20056 7276 20096
rect 7316 20056 7447 20096
rect 7625 20056 7747 20096
rect 7796 20056 8995 20096
rect 9044 20056 9053 20096
rect 9370 20087 9428 20096
rect 6796 20012 6836 20047
rect 9370 20047 9379 20087
rect 9419 20047 9428 20087
rect 9370 20046 9428 20047
rect 1577 19972 1708 20012
rect 1748 19972 1757 20012
rect 1930 20003 3340 20012
rect 1930 19963 1939 20003
rect 1979 19972 3340 20003
rect 3380 19972 3389 20012
rect 3593 19972 3724 20012
rect 3764 19972 3773 20012
rect 3946 20003 4204 20012
rect 1979 19963 1988 19972
rect 1930 19962 1988 19963
rect 3946 19963 3955 20003
rect 3995 19972 4204 20003
rect 4244 19972 4253 20012
rect 4579 19972 4588 20012
rect 4628 19972 4637 20012
rect 4841 19972 4972 20012
rect 5012 19972 5021 20012
rect 5417 19972 5548 20012
rect 5588 19972 5597 20012
rect 5731 19972 5740 20012
rect 5780 19972 5789 20012
rect 6307 19972 6316 20012
rect 6356 19972 6365 20012
rect 6787 19972 6796 20012
rect 6836 19972 6883 20012
rect 7555 19972 7564 20012
rect 7604 19972 7735 20012
rect 8009 19972 8140 20012
rect 8180 19972 8611 20012
rect 8651 19972 8660 20012
rect 8707 19972 8716 20012
rect 8756 19972 9187 20012
rect 9227 19972 9236 20012
rect 3995 19963 4004 19972
rect 3946 19962 4004 19963
rect 4588 19928 4628 19972
rect 1219 19888 1228 19928
rect 1268 19888 1844 19928
rect 2947 19888 2956 19928
rect 2996 19888 3127 19928
rect 4588 19888 4876 19928
rect 4916 19888 4925 19928
rect 5443 19888 5452 19928
rect 5492 19888 5501 19928
rect 0 19844 400 19864
rect 1804 19844 1844 19888
rect 0 19804 1324 19844
rect 1364 19804 1373 19844
rect 1804 19804 2380 19844
rect 2420 19804 2429 19844
rect 0 19784 400 19804
rect 5452 19760 5492 19888
rect 5548 19844 5588 19972
rect 5740 19928 5780 19972
rect 5740 19888 5836 19928
rect 5876 19888 5885 19928
rect 6089 19888 6124 19928
rect 6164 19888 6220 19928
rect 6260 19888 6269 19928
rect 6316 19844 6356 19972
rect 9388 19928 9428 20046
rect 10060 20056 10444 20096
rect 10484 20056 10493 20096
rect 10601 20056 10636 20096
rect 10676 20056 10732 20096
rect 10772 20056 10781 20096
rect 10889 20056 11011 20096
rect 11060 20056 11069 20096
rect 11203 20056 11212 20096
rect 11252 20056 11299 20096
rect 11339 20056 11383 20096
rect 13097 20056 13219 20096
rect 13268 20056 13277 20096
rect 13786 20056 13795 20096
rect 13835 20056 13844 20096
rect 14921 20056 15052 20096
rect 15092 20056 15101 20096
rect 15811 20056 15820 20096
rect 15860 20056 15991 20096
rect 16265 20056 16396 20096
rect 16436 20056 16445 20096
rect 16570 20056 16579 20096
rect 16628 20056 16759 20096
rect 16866 20056 16875 20096
rect 16915 20056 16924 20096
rect 16976 20056 17107 20096
rect 17147 20056 17156 20096
rect 17203 20056 17212 20096
rect 17252 20056 17261 20096
rect 17443 20056 17452 20096
rect 17492 20056 17836 20096
rect 17876 20056 17885 20096
rect 17932 20056 17955 20096
rect 17995 20056 18004 20096
rect 18064 20056 18073 20096
rect 18113 20056 18124 20096
rect 18164 20056 18253 20096
rect 18377 20087 18508 20096
rect 18377 20056 18499 20087
rect 18548 20056 18557 20096
rect 10060 20012 10100 20056
rect 15562 20014 15571 20054
rect 15611 20014 15668 20054
rect 15628 20012 15668 20014
rect 7066 19888 7075 19928
rect 7115 19888 7180 19928
rect 7220 19888 7255 19928
rect 7913 19888 8044 19928
rect 8084 19888 8093 19928
rect 8419 19888 8428 19928
rect 8468 19888 9428 19928
rect 9484 19972 9532 20012
rect 9572 19972 10100 20012
rect 10819 19972 10828 20012
rect 10868 19972 10877 20012
rect 11273 19972 11404 20012
rect 11444 19972 11453 20012
rect 13027 19972 13036 20012
rect 13076 19972 13085 20012
rect 13577 19972 13708 20012
rect 13748 19972 13757 20012
rect 15370 19972 15379 20012
rect 15419 19972 15428 20012
rect 15628 19972 16052 20012
rect 9484 19844 9524 19972
rect 10828 19928 10868 19972
rect 10723 19888 10732 19928
rect 10772 19888 10868 19928
rect 13036 19928 13076 19972
rect 13036 19888 13804 19928
rect 13844 19888 13853 19928
rect 15388 19844 15428 19972
rect 16012 19928 16052 19972
rect 16003 19888 16012 19928
rect 16052 19888 16061 19928
rect 5548 19804 6356 19844
rect 6403 19804 6412 19844
rect 6452 19804 6499 19844
rect 6539 19804 6583 19844
rect 6979 19804 6988 19844
rect 7028 19804 9524 19844
rect 10435 19804 10444 19844
rect 10484 19804 11500 19844
rect 11540 19804 11549 19844
rect 13027 19804 13036 19844
rect 13076 19804 15428 19844
rect 739 19720 748 19760
rect 788 19720 2860 19760
rect 2900 19720 2909 19760
rect 4579 19720 4588 19760
rect 4628 19720 5492 19760
rect 7852 19720 10100 19760
rect 3103 19636 3112 19676
rect 3480 19636 3489 19676
rect 7852 19592 7892 19720
rect 835 19552 844 19592
rect 884 19552 7892 19592
rect 10060 19592 10100 19720
rect 15388 19676 15428 19804
rect 16876 19760 16916 20056
rect 16986 19972 16995 20012
rect 17035 19972 17044 20012
rect 16995 19844 17035 19972
rect 17212 19928 17252 20056
rect 17338 19972 17347 20012
rect 17396 19972 17527 20012
rect 18124 19928 18164 20056
rect 18490 20047 18499 20056
rect 18539 20047 18548 20056
rect 18490 20046 18548 20047
rect 18988 20012 19028 20140
rect 19468 20096 19508 20140
rect 20236 20096 20276 20140
rect 24652 20096 24692 20140
rect 25324 20096 25364 20140
rect 25516 20140 25996 20180
rect 26036 20140 26045 20180
rect 26572 20140 27340 20180
rect 27380 20140 27389 20180
rect 27436 20140 27628 20180
rect 27668 20140 28052 20180
rect 28157 20140 28204 20180
rect 28244 20140 28253 20180
rect 28300 20140 29635 20180
rect 29675 20140 29684 20180
rect 25516 20096 25556 20140
rect 26572 20096 26612 20140
rect 27436 20096 27476 20140
rect 19145 20056 19276 20096
rect 19316 20056 19325 20096
rect 19459 20056 19468 20096
rect 19508 20056 19703 20096
rect 19743 20056 19752 20096
rect 19843 20056 19852 20096
rect 19892 20056 19948 20096
rect 19988 20056 20023 20096
rect 20227 20056 20236 20096
rect 20276 20056 20285 20096
rect 20419 20056 20428 20096
rect 20468 20056 20707 20096
rect 20747 20056 20852 20096
rect 20986 20056 20995 20096
rect 21035 20087 21332 20096
rect 21035 20056 21283 20087
rect 18643 19972 18652 20012
rect 18692 19972 18701 20012
rect 18988 19972 19843 20012
rect 19883 19972 19892 20012
rect 20035 19972 20044 20012
rect 20084 19972 20236 20012
rect 20276 19972 20285 20012
rect 18652 19928 18692 19972
rect 19852 19928 19892 19972
rect 20428 19928 20468 20056
rect 20812 20012 20852 20056
rect 21274 20047 21283 20056
rect 21323 20047 21332 20087
rect 24451 20056 24460 20096
rect 24500 20056 24509 20096
rect 24634 20056 24643 20096
rect 24683 20056 24692 20096
rect 24739 20056 24748 20096
rect 24788 20056 24797 20096
rect 24905 20056 25027 20096
rect 25076 20056 25085 20096
rect 25193 20056 25315 20096
rect 25364 20056 25373 20096
rect 25498 20056 25507 20096
rect 25547 20056 25556 20096
rect 25690 20056 25699 20096
rect 25748 20056 25879 20096
rect 26563 20056 26572 20096
rect 26612 20056 26621 20096
rect 27043 20056 27052 20096
rect 27092 20056 27101 20096
rect 27298 20056 27307 20096
rect 27347 20056 27476 20096
rect 27523 20056 27532 20096
rect 27572 20056 27703 20096
rect 21274 20046 21332 20047
rect 24460 20012 24500 20056
rect 24748 20012 24788 20056
rect 27052 20012 27092 20056
rect 28012 20012 28052 20140
rect 28204 20096 28244 20140
rect 28300 20096 28340 20140
rect 31084 20096 31124 20224
rect 28186 20056 28195 20096
rect 28235 20056 28244 20096
rect 28291 20056 28300 20096
rect 28340 20056 28349 20096
rect 29321 20056 29452 20096
rect 29492 20056 29501 20096
rect 30185 20056 30316 20096
rect 30356 20056 30365 20096
rect 30490 20087 30508 20096
rect 30490 20047 30499 20087
rect 30548 20056 30679 20096
rect 30979 20056 30988 20096
rect 31028 20056 31037 20096
rect 31084 20056 31180 20096
rect 31220 20056 31229 20096
rect 30539 20047 30548 20056
rect 30490 20046 30548 20047
rect 20515 19972 20524 20012
rect 20564 19972 20695 20012
rect 20812 19972 20908 20012
rect 20948 19972 20957 20012
rect 21091 19972 21100 20012
rect 21140 19972 21149 20012
rect 21388 19972 21436 20012
rect 21476 19972 21485 20012
rect 24460 19972 24596 20012
rect 24748 19972 26428 20012
rect 26468 19972 26477 20012
rect 26563 19972 26572 20012
rect 26612 19972 27052 20012
rect 27092 19972 27101 20012
rect 27418 19972 27427 20012
rect 27467 19972 27476 20012
rect 27619 19972 27628 20012
rect 27668 19972 27677 20012
rect 28012 19972 28876 20012
rect 28916 19972 28925 20012
rect 30643 19972 30652 20012
rect 30692 19972 30892 20012
rect 30932 19972 30941 20012
rect 17212 19888 17260 19928
rect 17300 19888 17309 19928
rect 18124 19888 19660 19928
rect 19700 19888 19709 19928
rect 19852 19888 20468 19928
rect 20707 19888 20716 19928
rect 20756 19888 21004 19928
rect 21044 19888 21053 19928
rect 21100 19844 21140 19972
rect 16995 19804 17644 19844
rect 17684 19804 17693 19844
rect 19267 19804 19276 19844
rect 19316 19804 19468 19844
rect 19508 19804 19517 19844
rect 20227 19804 20236 19844
rect 20276 19804 21100 19844
rect 21140 19804 21149 19844
rect 16876 19720 17452 19760
rect 17492 19720 17501 19760
rect 10877 19636 10886 19676
rect 11254 19636 11263 19676
rect 11587 19636 11596 19676
rect 11636 19636 11980 19676
rect 12020 19636 12029 19676
rect 15388 19636 16972 19676
rect 17012 19636 17021 19676
rect 18651 19636 18660 19676
rect 19028 19636 19037 19676
rect 21388 19592 21428 19972
rect 24556 19928 24596 19972
rect 24556 19888 25036 19928
rect 25076 19888 25085 19928
rect 26153 19888 26284 19928
rect 26324 19888 26333 19928
rect 24617 19804 24748 19844
rect 24788 19804 24797 19844
rect 26425 19636 26434 19676
rect 26802 19636 26811 19676
rect 10060 19552 21428 19592
rect 27436 19508 27476 19972
rect 2947 19468 2956 19508
rect 2996 19468 4156 19508
rect 4196 19468 4204 19508
rect 4244 19468 5164 19508
rect 5204 19468 5213 19508
rect 7267 19468 7276 19508
rect 7316 19468 7325 19508
rect 7377 19468 7756 19508
rect 7796 19468 7805 19508
rect 9763 19468 9772 19508
rect 9812 19468 11884 19508
rect 11924 19468 11933 19508
rect 16186 19468 16195 19508
rect 16235 19468 16396 19508
rect 16436 19468 16445 19508
rect 16666 19468 16675 19508
rect 16715 19468 17356 19508
rect 17396 19468 17405 19508
rect 17513 19468 17635 19508
rect 17684 19468 17693 19508
rect 19459 19468 19468 19508
rect 19508 19468 20468 19508
rect 26170 19468 26179 19508
rect 26219 19468 27476 19508
rect 0 19424 400 19444
rect 7276 19424 7316 19468
rect 0 19384 1324 19424
rect 1364 19384 1373 19424
rect 1795 19384 1804 19424
rect 1844 19384 3572 19424
rect 3619 19384 3628 19424
rect 3668 19384 4436 19424
rect 4483 19384 4492 19424
rect 4532 19384 6988 19424
rect 7028 19384 7037 19424
rect 7084 19384 7316 19424
rect 0 19364 400 19384
rect 1001 19300 1132 19340
rect 1172 19300 1181 19340
rect 1577 19300 1708 19340
rect 1748 19300 1757 19340
rect 1306 19216 1315 19256
rect 1355 19216 1364 19256
rect 1885 19249 1894 19289
rect 1934 19249 1943 19289
rect 2764 19256 2804 19265
rect 3004 19256 3044 19384
rect 3532 19340 3572 19384
rect 4396 19340 4436 19384
rect 3139 19300 3148 19340
rect 3211 19300 3319 19340
rect 3532 19300 3916 19340
rect 3956 19300 3965 19340
rect 4387 19300 4396 19340
rect 4436 19300 4780 19340
rect 4820 19300 4829 19340
rect 5705 19300 5836 19340
rect 5876 19300 5885 19340
rect 6124 19256 6164 19384
rect 7084 19340 7124 19384
rect 7377 19340 7417 19468
rect 11884 19424 11924 19468
rect 7651 19384 7660 19424
rect 7700 19384 8140 19424
rect 8180 19384 8189 19424
rect 10540 19384 10924 19424
rect 10964 19384 10973 19424
rect 11789 19384 11924 19424
rect 11971 19384 11980 19424
rect 12020 19384 12151 19424
rect 14921 19384 14956 19424
rect 14996 19384 15052 19424
rect 15092 19384 15101 19424
rect 19651 19384 19660 19424
rect 19700 19384 20276 19424
rect 10540 19340 10580 19384
rect 6307 19300 6316 19340
rect 6356 19300 6395 19340
rect 6676 19300 7124 19340
rect 7244 19300 7253 19340
rect 7293 19300 7417 19340
rect 7459 19300 7468 19340
rect 7508 19300 7660 19340
rect 7700 19300 7709 19340
rect 8131 19300 8140 19340
rect 8180 19300 8236 19340
rect 8276 19300 8311 19340
rect 8800 19300 8908 19340
rect 8971 19300 8980 19340
rect 9737 19300 9772 19340
rect 9812 19300 9859 19340
rect 9899 19300 9917 19340
rect 10522 19300 10531 19340
rect 10571 19300 10580 19340
rect 10723 19300 10732 19340
rect 10772 19300 10924 19340
rect 10964 19300 10973 19340
rect 11146 19331 11308 19340
rect 6316 19256 6356 19300
rect 6676 19256 6716 19300
rect 7084 19298 7124 19300
rect 7084 19258 7132 19298
rect 7172 19258 7181 19298
rect 11146 19291 11155 19331
rect 11195 19300 11308 19331
rect 11348 19300 11357 19340
rect 11491 19300 11500 19340
rect 11540 19300 11636 19340
rect 11195 19291 11204 19300
rect 11146 19290 11204 19291
rect 9964 19256 10100 19259
rect 11596 19256 11636 19300
rect 11789 19256 11829 19384
rect 13219 19300 13228 19340
rect 13268 19300 13277 19340
rect 13411 19300 13420 19340
rect 13460 19300 14860 19340
rect 14900 19300 15092 19340
rect 13228 19256 13268 19300
rect 15052 19256 15092 19300
rect 15916 19300 16244 19340
rect 17129 19300 17260 19340
rect 17300 19300 18508 19340
rect 18548 19300 18557 19340
rect 1324 19088 1364 19216
rect 1900 19172 1940 19249
rect 2083 19216 2092 19256
rect 2132 19216 2199 19256
rect 2239 19216 2462 19256
rect 2502 19216 2511 19256
rect 2633 19216 2764 19256
rect 2804 19216 2813 19256
rect 3004 19216 3052 19256
rect 3092 19216 3101 19256
rect 3148 19216 3269 19256
rect 3309 19216 3318 19256
rect 3427 19216 3436 19256
rect 3476 19216 3485 19256
rect 3610 19216 3619 19256
rect 3659 19216 4492 19256
rect 4532 19216 4541 19256
rect 5501 19216 5515 19256
rect 5555 19216 5564 19256
rect 5626 19216 5635 19256
rect 5675 19216 5684 19256
rect 5731 19216 5740 19256
rect 5780 19216 5911 19256
rect 6115 19216 6124 19256
rect 6164 19216 6173 19256
rect 6299 19216 6308 19256
rect 6348 19216 6357 19256
rect 6516 19216 6604 19256
rect 6644 19216 6667 19256
rect 6707 19216 6716 19256
rect 6778 19216 6787 19256
rect 6827 19216 6836 19256
rect 6883 19216 6892 19256
rect 6932 19216 6941 19256
rect 7363 19216 7372 19256
rect 7412 19216 7421 19256
rect 7721 19216 7843 19256
rect 7892 19216 7901 19256
rect 7948 19216 8812 19256
rect 8852 19216 8861 19256
rect 9040 19216 9049 19256
rect 9089 19216 9280 19256
rect 9332 19216 9341 19256
rect 9710 19216 9719 19256
rect 9759 19216 9768 19256
rect 9833 19216 9964 19256
rect 10004 19219 10391 19256
rect 10004 19216 10013 19219
rect 10060 19216 10391 19219
rect 10431 19216 10440 19256
rect 10627 19216 10636 19256
rect 10676 19216 11020 19256
rect 11060 19216 11069 19256
rect 11248 19216 11257 19256
rect 11297 19216 11404 19256
rect 11444 19216 11500 19256
rect 11540 19216 11549 19256
rect 11596 19216 11619 19256
rect 11659 19216 11668 19256
rect 11728 19216 11737 19256
rect 11777 19216 11829 19256
rect 11875 19216 11884 19256
rect 11924 19216 11933 19256
rect 12067 19216 12076 19256
rect 12116 19216 12125 19256
rect 12259 19216 12268 19256
rect 12308 19216 12317 19256
rect 12451 19216 12460 19256
rect 12500 19216 12631 19256
rect 13123 19216 13132 19256
rect 13172 19216 13268 19256
rect 13315 19216 13324 19256
rect 13364 19216 13516 19256
rect 13556 19216 13565 19256
rect 13673 19216 13804 19256
rect 13844 19216 13853 19256
rect 14345 19216 14419 19256
rect 14459 19216 14476 19256
rect 14516 19216 14525 19256
rect 14605 19216 14614 19256
rect 14654 19216 14697 19256
rect 2764 19207 2804 19216
rect 3148 19172 3188 19216
rect 3436 19172 3476 19216
rect 5524 19172 5564 19216
rect 1481 19132 1516 19172
rect 1556 19132 1612 19172
rect 1652 19132 1661 19172
rect 1889 19132 1900 19172
rect 1940 19132 1949 19172
rect 1996 19132 2188 19172
rect 2228 19132 2237 19172
rect 2371 19132 2380 19172
rect 2420 19132 2563 19172
rect 2603 19132 2612 19172
rect 2851 19132 2860 19172
rect 2900 19132 2909 19172
rect 3043 19132 3052 19172
rect 3092 19132 3340 19172
rect 3380 19132 3389 19172
rect 3436 19132 3820 19172
rect 3860 19132 3869 19172
rect 5524 19132 5548 19172
rect 5588 19132 5597 19172
rect 1996 19088 2036 19132
rect 2860 19088 2900 19132
rect 5644 19088 5684 19216
rect 5897 19132 6019 19172
rect 6068 19132 6077 19172
rect 1027 19048 1036 19088
rect 1076 19048 1987 19088
rect 2027 19048 2036 19088
rect 2083 19048 2092 19088
rect 2132 19048 2141 19088
rect 2659 19048 2668 19088
rect 2708 19048 2900 19088
rect 2947 19048 2956 19088
rect 2996 19048 3005 19088
rect 3523 19048 3532 19088
rect 3572 19048 3581 19088
rect 5644 19048 6700 19088
rect 6740 19048 6749 19088
rect 2092 19004 2132 19048
rect 2956 19004 2996 19048
rect 1795 18964 1804 19004
rect 1844 18964 2132 19004
rect 2860 18964 2996 19004
rect 2860 18920 2900 18964
rect 3532 18920 3572 19048
rect 6796 19004 6836 19216
rect 6892 19172 6932 19216
rect 7372 19172 7412 19216
rect 7948 19172 7988 19216
rect 8812 19172 8852 19216
rect 9719 19172 9759 19216
rect 11020 19172 11060 19216
rect 11884 19172 11924 19216
rect 12076 19172 12116 19216
rect 6892 19132 7988 19172
rect 8585 19132 8716 19172
rect 8756 19132 8765 19172
rect 8812 19132 9004 19172
rect 9044 19132 9053 19172
rect 9317 19132 9759 19172
rect 9868 19132 10868 19172
rect 11020 19132 11404 19172
rect 11444 19132 11924 19172
rect 11971 19132 11980 19172
rect 12020 19132 12116 19172
rect 12268 19172 12308 19216
rect 12268 19132 12556 19172
rect 12596 19132 12605 19172
rect 13123 19132 13132 19172
rect 13172 19132 13603 19172
rect 13643 19132 13652 19172
rect 9317 19088 9357 19132
rect 9868 19088 9908 19132
rect 6970 19048 6979 19088
rect 7019 19048 7564 19088
rect 7604 19048 7613 19088
rect 8803 19048 8812 19088
rect 8852 19048 9357 19088
rect 9427 19048 9436 19088
rect 9476 19048 9908 19088
rect 10042 19048 10051 19088
rect 10091 19048 10100 19088
rect 10714 19048 10723 19088
rect 10763 19048 10772 19088
rect 9436 19004 9476 19048
rect 6796 18964 6892 19004
rect 6932 18964 6941 19004
rect 7267 18964 7276 19004
rect 7316 18964 9476 19004
rect 10060 18920 10100 19048
rect 1603 18880 1612 18920
rect 1652 18880 2900 18920
rect 2956 18880 3572 18920
rect 4343 18880 4352 18920
rect 4720 18880 4729 18920
rect 8995 18880 9004 18920
rect 9044 18880 10100 18920
rect 10732 18920 10772 19048
rect 10828 19004 10868 19132
rect 14657 19088 14697 19216
rect 14746 19247 14996 19256
rect 14746 19207 14755 19247
rect 14795 19216 14996 19247
rect 15043 19216 15052 19256
rect 15092 19216 15436 19256
rect 15476 19216 15820 19256
rect 15860 19216 15869 19256
rect 14795 19207 14804 19216
rect 14746 19206 14804 19207
rect 14956 19172 14996 19216
rect 14956 19132 15052 19172
rect 15092 19132 15380 19172
rect 15340 19088 15380 19132
rect 10915 19048 10924 19088
rect 10964 19048 12364 19088
rect 12404 19048 12413 19088
rect 13882 19048 13891 19088
rect 13931 19048 14476 19088
rect 14516 19048 14525 19088
rect 14657 19048 15148 19088
rect 15188 19048 15197 19088
rect 15322 19048 15331 19088
rect 15371 19048 15436 19088
rect 15476 19048 15540 19088
rect 15610 19048 15619 19088
rect 15659 19048 15724 19088
rect 15764 19048 15799 19088
rect 15916 19004 15956 19300
rect 16204 19256 16244 19300
rect 16003 19216 16012 19256
rect 16052 19216 16061 19256
rect 16186 19216 16195 19256
rect 16235 19216 16244 19256
rect 16972 19256 17012 19265
rect 17260 19256 17300 19300
rect 19660 19256 19700 19384
rect 19747 19300 19756 19340
rect 19796 19300 19939 19340
rect 19979 19300 19988 19340
rect 20236 19256 20276 19384
rect 20428 19340 20468 19468
rect 20515 19384 20524 19424
rect 20564 19384 20660 19424
rect 21187 19384 21196 19424
rect 21236 19384 21292 19424
rect 21332 19384 21868 19424
rect 21908 19384 21917 19424
rect 23002 19384 23011 19424
rect 23051 19384 23060 19424
rect 23386 19384 23395 19424
rect 23435 19384 24212 19424
rect 24547 19384 24556 19424
rect 24596 19384 24844 19424
rect 24884 19384 24893 19424
rect 20620 19340 20660 19384
rect 23020 19340 23060 19384
rect 24172 19340 24212 19384
rect 20410 19300 20419 19340
rect 20459 19300 20468 19340
rect 20611 19300 20620 19340
rect 20660 19300 20669 19340
rect 20803 19300 20812 19340
rect 20852 19300 20983 19340
rect 21091 19300 21100 19340
rect 21140 19300 21388 19340
rect 21428 19300 21437 19340
rect 22732 19300 22828 19340
rect 22868 19300 22877 19340
rect 23020 19300 23299 19340
rect 23339 19300 23348 19340
rect 23491 19300 23500 19340
rect 23540 19300 23548 19340
rect 23588 19300 23671 19340
rect 24172 19300 24308 19340
rect 24643 19300 24652 19340
rect 24692 19300 25036 19340
rect 25076 19300 25085 19340
rect 25900 19300 27476 19340
rect 22732 19256 22772 19300
rect 24268 19298 24308 19300
rect 24268 19289 24312 19298
rect 24268 19258 24272 19289
rect 17251 19216 17260 19256
rect 17300 19216 17309 19256
rect 17356 19216 17379 19256
rect 17419 19216 17428 19256
rect 17488 19216 17497 19256
rect 17537 19216 17548 19256
rect 17588 19216 17780 19256
rect 17929 19216 17938 19256
rect 17978 19216 18220 19256
rect 18260 19216 18269 19256
rect 19049 19216 19171 19256
rect 19220 19216 19229 19256
rect 19348 19216 19468 19256
rect 19519 19216 19528 19256
rect 19660 19216 19799 19256
rect 19839 19216 19848 19256
rect 20035 19216 20044 19256
rect 20084 19216 20160 19256
rect 20236 19216 20279 19256
rect 20319 19216 20328 19256
rect 20515 19216 20524 19256
rect 20564 19216 20573 19256
rect 20899 19216 20908 19256
rect 20948 19216 20995 19256
rect 21035 19216 21079 19256
rect 21379 19216 21388 19256
rect 21428 19216 21523 19256
rect 21563 19216 21572 19256
rect 22714 19216 22723 19256
rect 22763 19216 22772 19256
rect 22819 19216 22828 19256
rect 22868 19216 23588 19256
rect 23681 19216 23690 19256
rect 23732 19216 23863 19256
rect 24041 19216 24163 19256
rect 24212 19216 24221 19256
rect 25900 19256 25940 19300
rect 24272 19240 24312 19249
rect 25193 19216 25219 19256
rect 25259 19216 25324 19256
rect 25364 19216 25373 19256
rect 25882 19216 25891 19256
rect 25931 19216 25940 19256
rect 25987 19216 25996 19256
rect 26036 19216 26045 19256
rect 26467 19216 26476 19256
rect 26516 19216 26525 19256
rect 16012 19088 16052 19216
rect 16972 19172 17012 19216
rect 17356 19172 17396 19216
rect 17740 19172 17780 19216
rect 20044 19172 20084 19216
rect 20524 19172 20564 19216
rect 16099 19132 16108 19172
rect 16148 19132 16670 19172
rect 16710 19132 16876 19172
rect 16916 19132 16925 19172
rect 16972 19132 17164 19172
rect 17204 19132 17213 19172
rect 17332 19132 17356 19172
rect 17396 19132 17630 19172
rect 17670 19132 17679 19172
rect 17740 19132 18988 19172
rect 19028 19132 19037 19172
rect 19363 19132 19372 19172
rect 19412 19132 20564 19172
rect 23548 19172 23588 19216
rect 24172 19172 24212 19216
rect 25996 19172 26036 19216
rect 26476 19172 26516 19216
rect 27436 19172 27476 19300
rect 27628 19256 27668 19972
rect 30988 19928 31028 20056
rect 28474 19888 28483 19928
rect 28523 19888 31028 19928
rect 28649 19804 28780 19844
rect 28820 19804 28829 19844
rect 30979 19804 30988 19844
rect 31028 19804 31037 19844
rect 30988 19508 31028 19804
rect 28963 19468 28972 19508
rect 29012 19468 30316 19508
rect 30356 19468 30365 19508
rect 30988 19468 31220 19508
rect 31180 19340 31220 19468
rect 28099 19300 28108 19340
rect 28148 19300 28340 19340
rect 29827 19300 29836 19340
rect 29876 19300 29885 19340
rect 31180 19300 31267 19340
rect 31307 19300 31316 19340
rect 28300 19256 28340 19300
rect 27628 19216 28108 19256
rect 28148 19216 28157 19256
rect 28282 19216 28291 19256
rect 28331 19216 28340 19256
rect 30761 19216 30883 19256
rect 30932 19216 30941 19256
rect 23548 19132 24212 19172
rect 25027 19132 25036 19172
rect 25076 19132 26036 19172
rect 26083 19132 26092 19172
rect 26132 19132 26516 19172
rect 27139 19132 27148 19172
rect 27188 19132 27340 19172
rect 27380 19132 27389 19172
rect 27436 19132 28300 19172
rect 28340 19132 28349 19172
rect 28468 19132 28492 19172
rect 28532 19132 28599 19172
rect 28639 19132 28648 19172
rect 16012 19048 16108 19088
rect 16148 19048 16157 19088
rect 16675 19048 16684 19088
rect 16724 19048 16876 19088
rect 16916 19048 16925 19088
rect 17155 19048 17164 19088
rect 17204 19048 17452 19088
rect 17492 19048 17501 19088
rect 17635 19048 17644 19088
rect 17684 19048 17836 19088
rect 17876 19048 17885 19088
rect 19145 19048 19267 19088
rect 19316 19048 19325 19088
rect 20122 19048 20131 19088
rect 20171 19048 20908 19088
rect 20948 19048 20957 19088
rect 21715 19048 21724 19088
rect 21764 19048 21773 19088
rect 23020 19048 23116 19088
rect 23156 19048 23165 19088
rect 23273 19048 23395 19088
rect 23444 19048 23453 19088
rect 23945 19079 24076 19088
rect 23945 19048 24067 19079
rect 24116 19048 24125 19088
rect 24617 19048 24739 19088
rect 24788 19048 24797 19088
rect 27305 19048 27436 19088
rect 27476 19048 27485 19088
rect 28378 19048 28387 19088
rect 28427 19048 28436 19088
rect 28483 19048 28492 19088
rect 28532 19048 28588 19088
rect 28628 19048 28663 19088
rect 28963 19048 28972 19088
rect 29012 19048 29021 19088
rect 19276 19004 19316 19048
rect 10819 18964 10828 19004
rect 10868 18964 11404 19004
rect 11444 18964 11453 19004
rect 14563 18964 14572 19004
rect 14612 18964 19316 19004
rect 10732 18880 11692 18920
rect 11732 18880 11741 18920
rect 12117 18880 12126 18920
rect 12494 18880 12503 18920
rect 19891 18880 19900 18920
rect 20268 18880 20277 18920
rect 2956 18836 2996 18880
rect 21724 18836 21764 19048
rect 67 18796 76 18836
rect 116 18796 2092 18836
rect 2132 18796 2141 18836
rect 2558 18796 2996 18836
rect 3139 18796 3148 18836
rect 3188 18796 21764 18836
rect 1123 18712 1132 18752
rect 1172 18712 1411 18752
rect 1451 18712 1460 18752
rect 1769 18712 1891 18752
rect 1940 18712 1949 18752
rect 2558 18668 2598 18796
rect 23020 18752 23060 19048
rect 24058 19039 24067 19048
rect 24107 19039 24116 19048
rect 24058 19038 24116 19039
rect 28396 19004 28436 19048
rect 28972 19004 29012 19048
rect 27043 18964 27052 19004
rect 27092 18964 29012 19004
rect 27665 18880 27674 18920
rect 28042 18880 28051 18920
rect 2755 18712 2764 18752
rect 2804 18712 3052 18752
rect 3092 18712 3101 18752
rect 4073 18712 4204 18752
rect 4244 18712 4253 18752
rect 4963 18712 4972 18752
rect 5012 18712 5251 18752
rect 5291 18712 5300 18752
rect 5356 18712 5740 18752
rect 5780 18712 6412 18752
rect 6452 18712 6461 18752
rect 6883 18712 6892 18752
rect 6932 18712 7276 18752
rect 7316 18712 7325 18752
rect 7564 18712 7988 18752
rect 8131 18712 8140 18752
rect 8180 18712 8660 18752
rect 8777 18712 8899 18752
rect 8948 18712 8957 18752
rect 9235 18712 9244 18752
rect 9284 18712 9292 18752
rect 9332 18712 9415 18752
rect 11011 18712 11020 18752
rect 11060 18712 11069 18752
rect 11177 18712 11308 18752
rect 11348 18712 11357 18752
rect 13411 18712 13420 18752
rect 13460 18712 13891 18752
rect 13931 18712 14476 18752
rect 14516 18712 14525 18752
rect 16553 18712 16684 18752
rect 16724 18712 16733 18752
rect 17801 18712 17923 18752
rect 17972 18712 17981 18752
rect 18211 18712 18220 18752
rect 18260 18712 18403 18752
rect 18443 18712 18452 18752
rect 19241 18712 19363 18752
rect 19412 18712 20236 18752
rect 20276 18712 20285 18752
rect 22915 18712 22924 18752
rect 22964 18712 23060 18752
rect 27139 18712 27148 18752
rect 27188 18712 27763 18752
rect 27803 18712 28492 18752
rect 28532 18712 28541 18752
rect 28963 18712 28972 18752
rect 29012 18712 29452 18752
rect 29492 18712 29501 18752
rect 5356 18668 5396 18712
rect 7564 18668 7604 18712
rect 7948 18668 7988 18712
rect 8620 18668 8660 18712
rect 11020 18668 11060 18712
rect 1324 18628 2092 18668
rect 2132 18628 2141 18668
rect 2284 18628 2558 18668
rect 2598 18628 2607 18668
rect 2650 18628 2659 18668
rect 2699 18628 3307 18668
rect 3715 18628 3724 18668
rect 3764 18628 3998 18668
rect 4038 18628 4047 18668
rect 4108 18628 4780 18668
rect 4820 18628 5012 18668
rect 1324 18584 1364 18628
rect 1804 18584 1844 18628
rect 940 18544 1079 18584
rect 1119 18544 1128 18584
rect 1315 18544 1324 18584
rect 1364 18544 1373 18584
rect 1795 18544 1804 18584
rect 1844 18544 1853 18584
rect 2057 18544 2092 18584
rect 2132 18544 2188 18584
rect 2228 18544 2237 18584
rect 940 18416 980 18544
rect 1555 18502 1564 18542
rect 1604 18502 1613 18542
rect 1097 18460 1219 18500
rect 1268 18460 1277 18500
rect 1564 18416 1604 18502
rect 2284 18500 2324 18628
rect 3267 18584 3307 18628
rect 4108 18584 4148 18628
rect 4972 18584 5012 18628
rect 5164 18628 5396 18668
rect 5635 18628 5644 18668
rect 5684 18628 5693 18668
rect 5923 18628 5932 18668
rect 5972 18628 7604 18668
rect 7651 18628 7660 18668
rect 7700 18628 7831 18668
rect 7948 18628 8179 18668
rect 8219 18628 8564 18668
rect 8620 18628 8798 18668
rect 8852 18628 8861 18668
rect 8995 18628 9004 18668
rect 9044 18628 9175 18668
rect 10732 18628 10828 18668
rect 10868 18628 10877 18668
rect 11020 18628 11980 18668
rect 12020 18628 12029 18668
rect 13594 18628 13603 18668
rect 13643 18628 13652 18668
rect 16841 18628 16876 18668
rect 16916 18628 16972 18668
rect 17012 18628 17021 18668
rect 18028 18628 18508 18668
rect 18548 18628 18557 18668
rect 19180 18628 19468 18668
rect 19508 18628 19517 18668
rect 19747 18628 19756 18668
rect 19796 18628 20180 18668
rect 20314 18628 20323 18668
rect 20363 18628 20812 18668
rect 20852 18628 20861 18668
rect 21257 18628 21388 18668
rect 21428 18628 21437 18668
rect 22924 18628 23692 18668
rect 23732 18628 23741 18668
rect 24329 18628 24451 18668
rect 24500 18628 24509 18668
rect 27305 18628 27331 18668
rect 27371 18628 27436 18668
rect 27476 18628 27485 18668
rect 27967 18628 28780 18668
rect 28820 18628 28829 18668
rect 5164 18584 5204 18628
rect 5644 18584 5684 18628
rect 8524 18584 8564 18628
rect 10732 18584 10772 18628
rect 13612 18584 13652 18628
rect 2416 18544 2425 18584
rect 2465 18544 2567 18584
rect 2633 18544 2668 18584
rect 2708 18544 2764 18584
rect 2804 18544 2813 18584
rect 2860 18575 2956 18584
rect 2527 18500 2567 18544
rect 2900 18544 2956 18575
rect 2996 18544 3031 18584
rect 3139 18544 3148 18584
rect 3188 18544 3197 18584
rect 3258 18544 3267 18584
rect 3307 18544 3316 18584
rect 3436 18544 4148 18584
rect 4291 18544 4300 18584
rect 4340 18544 4471 18584
rect 4930 18544 4939 18584
rect 4979 18544 5012 18584
rect 5155 18544 5164 18584
rect 5204 18544 5548 18584
rect 5588 18544 5597 18584
rect 5644 18544 5765 18584
rect 5805 18544 5814 18584
rect 5912 18544 5921 18584
rect 5961 18544 6068 18584
rect 6115 18544 6124 18584
rect 6164 18544 6173 18584
rect 6220 18575 6260 18584
rect 2860 18526 2900 18535
rect 1690 18460 1699 18500
rect 1748 18460 1879 18500
rect 2083 18460 2092 18500
rect 2132 18460 2141 18500
rect 2275 18460 2284 18500
rect 2347 18460 2455 18500
rect 2527 18460 2764 18500
rect 2804 18460 2813 18500
rect 2092 18416 2132 18460
rect 3148 18416 3188 18544
rect 3436 18542 3476 18544
rect 3379 18502 3388 18542
rect 3428 18502 3476 18542
rect 4300 18526 4340 18535
rect 940 18376 1662 18416
rect 2092 18376 3188 18416
rect 1622 18248 1662 18376
rect 3436 18332 3476 18502
rect 4780 18502 4819 18542
rect 4859 18502 4868 18542
rect 3811 18460 3820 18500
rect 3860 18460 3869 18500
rect 4553 18460 4627 18500
rect 4667 18460 4684 18500
rect 4724 18460 4733 18500
rect 3820 18416 3860 18460
rect 4780 18416 4820 18502
rect 6028 18500 6068 18544
rect 5050 18460 5059 18500
rect 5108 18460 5239 18500
rect 5443 18460 5452 18500
rect 5492 18460 5588 18500
rect 3820 18376 4820 18416
rect 2083 18292 2092 18332
rect 2132 18292 3580 18332
rect 3620 18292 3629 18332
rect 3881 18292 4003 18332
rect 4052 18292 4061 18332
rect 1622 18208 2188 18248
rect 2228 18208 2237 18248
rect 2860 18208 3956 18248
rect 2860 18080 2900 18208
rect 3103 18124 3112 18164
rect 3480 18124 3489 18164
rect 2284 18040 2900 18080
rect 3916 18080 3956 18208
rect 4780 18164 4820 18376
rect 5548 18248 5588 18460
rect 5674 18491 5972 18500
rect 5674 18451 5683 18491
rect 5723 18460 5972 18491
rect 6019 18460 6028 18500
rect 6068 18460 6077 18500
rect 5723 18451 5732 18460
rect 5674 18450 5732 18451
rect 5932 18332 5972 18460
rect 6124 18416 6164 18544
rect 6473 18544 6508 18584
rect 6548 18544 6604 18584
rect 6644 18544 6653 18584
rect 6736 18544 6745 18584
rect 6785 18544 6892 18584
rect 6932 18544 6941 18584
rect 7049 18544 7180 18584
rect 7220 18544 7229 18584
rect 7325 18544 7371 18584
rect 7411 18544 7420 18584
rect 7546 18544 7555 18584
rect 7604 18544 7735 18584
rect 7854 18544 7863 18584
rect 7903 18544 8140 18584
rect 8180 18544 8189 18584
rect 8365 18544 8374 18584
rect 8414 18544 8468 18584
rect 8515 18544 8524 18584
rect 8564 18544 8573 18584
rect 9100 18575 9140 18584
rect 6220 18500 6260 18535
rect 6211 18460 6220 18500
rect 6260 18460 6307 18500
rect 6496 18460 6508 18500
rect 6548 18460 6627 18500
rect 6667 18460 6676 18500
rect 7180 18416 7220 18544
rect 7372 18500 7412 18544
rect 7863 18500 7903 18544
rect 7363 18460 7372 18500
rect 7412 18460 7421 18500
rect 7660 18460 7903 18500
rect 8428 18500 8468 18544
rect 10723 18544 10732 18584
rect 10772 18544 10781 18584
rect 10865 18544 10874 18584
rect 10914 18544 11018 18584
rect 11081 18544 11212 18584
rect 11252 18544 11261 18584
rect 11386 18544 11395 18584
rect 11435 18544 11788 18584
rect 11828 18544 11837 18584
rect 12685 18544 12694 18584
rect 12734 18544 13132 18584
rect 13172 18544 13181 18584
rect 13315 18544 13324 18584
rect 13364 18544 13652 18584
rect 13699 18544 13708 18584
rect 13748 18544 13804 18584
rect 13844 18544 13879 18584
rect 14467 18544 14476 18584
rect 14516 18544 14668 18584
rect 14708 18544 14717 18584
rect 14851 18544 14860 18584
rect 14900 18544 15031 18584
rect 16195 18544 16204 18584
rect 16244 18544 16253 18584
rect 16364 18544 16373 18584
rect 16413 18544 16436 18584
rect 16483 18544 16492 18584
rect 16532 18544 16684 18584
rect 16724 18544 16733 18584
rect 16858 18544 16867 18584
rect 16907 18544 16916 18584
rect 9100 18500 9140 18535
rect 10978 18500 11018 18544
rect 8428 18460 8812 18500
rect 8852 18460 8861 18500
rect 9091 18460 9100 18500
rect 9140 18460 9187 18500
rect 9475 18460 9484 18500
rect 9524 18460 9533 18500
rect 10978 18460 11404 18500
rect 11444 18460 11453 18500
rect 11683 18460 11692 18500
rect 11732 18460 12499 18500
rect 12539 18460 16108 18500
rect 16148 18460 16157 18500
rect 7660 18416 7700 18460
rect 9484 18416 9524 18460
rect 6124 18376 6189 18416
rect 7180 18376 7700 18416
rect 7747 18376 7756 18416
rect 7796 18376 7805 18416
rect 9484 18376 15916 18416
rect 15956 18376 15965 18416
rect 5914 18292 5923 18332
rect 5963 18292 5972 18332
rect 6149 18332 6189 18376
rect 7756 18332 7796 18376
rect 6149 18292 6316 18332
rect 6356 18292 7660 18332
rect 7700 18292 7709 18332
rect 7756 18292 7852 18332
rect 7892 18292 7901 18332
rect 5548 18208 6796 18248
rect 6836 18208 6845 18248
rect 9484 18164 9524 18376
rect 11011 18292 11020 18332
rect 11060 18292 11540 18332
rect 13123 18292 13132 18332
rect 13172 18292 13612 18332
rect 13652 18292 13661 18332
rect 14633 18292 14764 18332
rect 14804 18292 14813 18332
rect 11500 18248 11540 18292
rect 11500 18208 13516 18248
rect 13556 18208 13565 18248
rect 4780 18124 9524 18164
rect 10877 18124 10886 18164
rect 11254 18124 11263 18164
rect 3916 18040 4972 18080
rect 5012 18040 5021 18080
rect 5155 18040 5164 18080
rect 5204 18040 12844 18080
rect 12884 18040 12893 18080
rect 1289 17956 1411 17996
rect 1460 17956 1469 17996
rect 1699 17956 1708 17996
rect 1748 17956 2179 17996
rect 2219 17956 2228 17996
rect 2284 17912 2324 18040
rect 16204 17996 16244 18544
rect 16396 18416 16436 18544
rect 16876 18500 16916 18544
rect 17068 18544 17175 18584
rect 17215 18544 17224 18584
rect 17290 18544 17299 18584
rect 17339 18544 17396 18584
rect 17705 18544 17827 18584
rect 17876 18544 17885 18584
rect 17068 18500 17108 18544
rect 17356 18500 17396 18544
rect 18028 18500 18068 18628
rect 18115 18544 18124 18584
rect 18175 18544 18302 18584
rect 18342 18544 18351 18584
rect 18604 18575 18644 18584
rect 16483 18460 16492 18500
rect 16532 18460 16916 18500
rect 17059 18460 17068 18500
rect 17108 18460 17117 18500
rect 17347 18460 17356 18500
rect 17396 18460 17405 18500
rect 17491 18460 17500 18500
rect 17540 18460 17548 18500
rect 17588 18460 18028 18500
rect 18068 18460 18077 18500
rect 17068 18416 17108 18460
rect 18124 18416 18164 18544
rect 18900 18544 18988 18584
rect 19028 18544 19031 18584
rect 19071 18544 19080 18584
rect 18604 18500 18644 18535
rect 19180 18500 19220 18628
rect 20140 18584 20180 18628
rect 22924 18584 22964 18628
rect 27967 18584 28007 18628
rect 28588 18584 28628 18628
rect 19265 18544 19274 18584
rect 19314 18544 19323 18584
rect 19546 18544 19555 18584
rect 19595 18544 19604 18584
rect 19651 18544 19660 18584
rect 19700 18544 19709 18584
rect 19854 18562 19863 18584
rect 19852 18544 19863 18562
rect 19903 18544 19912 18584
rect 19987 18544 19996 18584
rect 20036 18544 20045 18584
rect 20122 18544 20131 18584
rect 20171 18544 20180 18584
rect 20227 18544 20236 18584
rect 20276 18544 20407 18584
rect 20995 18544 21004 18584
rect 21044 18544 21091 18584
rect 21131 18544 21175 18584
rect 22906 18544 22915 18584
rect 22955 18544 22964 18584
rect 23011 18544 23020 18584
rect 23060 18544 23500 18584
rect 23540 18544 23549 18584
rect 24355 18544 24364 18584
rect 24404 18544 24413 18584
rect 24547 18544 24556 18584
rect 24596 18544 24748 18584
rect 24788 18544 24797 18584
rect 26825 18544 26947 18584
rect 26996 18544 27005 18584
rect 27946 18544 27955 18584
rect 27995 18544 28007 18584
rect 28066 18544 28075 18584
rect 28148 18544 28255 18584
rect 28522 18544 28531 18584
rect 28571 18544 28628 18584
rect 28745 18544 28780 18584
rect 28820 18544 28876 18584
rect 28916 18544 28925 18584
rect 30761 18544 30883 18584
rect 30932 18544 30941 18584
rect 19276 18500 19316 18544
rect 18307 18460 18316 18500
rect 18356 18460 18644 18500
rect 19162 18460 19171 18500
rect 19211 18460 19220 18500
rect 19267 18460 19276 18500
rect 19316 18460 19361 18500
rect 19564 18416 19604 18544
rect 16396 18376 16972 18416
rect 17012 18376 17021 18416
rect 17068 18376 18164 18416
rect 18211 18376 18220 18416
rect 18260 18376 19604 18416
rect 19660 18332 19700 18544
rect 19852 18522 19903 18544
rect 19852 18416 19892 18522
rect 19996 18500 20036 18544
rect 24364 18500 24404 18544
rect 28359 18502 28368 18542
rect 28408 18502 28436 18542
rect 28396 18500 28436 18502
rect 19939 18460 19948 18500
rect 19988 18460 20036 18500
rect 20777 18460 20908 18500
rect 20948 18460 20957 18500
rect 21091 18460 21100 18500
rect 21140 18460 21484 18500
rect 21524 18460 21533 18500
rect 21737 18460 21868 18500
rect 21908 18460 21917 18500
rect 24364 18460 25324 18500
rect 25364 18460 25373 18500
rect 26275 18460 26284 18500
rect 26324 18460 26333 18500
rect 28073 18460 28204 18500
rect 28244 18460 28253 18500
rect 28396 18460 28636 18500
rect 28676 18460 28685 18500
rect 30979 18460 30988 18500
rect 31028 18460 31037 18500
rect 31258 18460 31267 18500
rect 31307 18460 31316 18500
rect 19843 18376 19852 18416
rect 19892 18376 19901 18416
rect 20131 18376 20140 18416
rect 20180 18376 21812 18416
rect 22723 18376 22732 18416
rect 22772 18376 23212 18416
rect 23252 18376 23261 18416
rect 25027 18376 25036 18416
rect 25076 18376 25420 18416
rect 25460 18376 25469 18416
rect 28291 18376 28300 18416
rect 28340 18376 28349 18416
rect 21772 18332 21812 18376
rect 17129 18292 17164 18332
rect 17204 18292 17260 18332
rect 17300 18292 17309 18332
rect 18115 18292 18124 18332
rect 18164 18292 18173 18332
rect 19363 18292 19372 18332
rect 19412 18292 19700 18332
rect 19948 18292 21628 18332
rect 21668 18292 21677 18332
rect 21772 18292 23060 18332
rect 25027 18292 25036 18332
rect 25076 18292 26092 18332
rect 26132 18292 26141 18332
rect 3331 17956 3340 17996
rect 3380 17956 3724 17996
rect 3764 17956 3773 17996
rect 3820 17956 4684 17996
rect 4724 17956 4733 17996
rect 5059 17956 5068 17996
rect 5108 17956 5740 17996
rect 5780 17956 5789 17996
rect 6787 17956 6796 17996
rect 6836 17956 7555 17996
rect 7595 17956 7604 17996
rect 8851 17956 8860 17996
rect 8900 17956 9004 17996
rect 9044 17956 9053 17996
rect 9100 17956 11500 17996
rect 11540 17956 11549 17996
rect 16204 17956 16300 17996
rect 16340 17956 16349 17996
rect 1315 17872 1324 17912
rect 1364 17872 2324 17912
rect 3820 17828 3860 17956
rect 3907 17872 3916 17912
rect 3956 17872 8812 17912
rect 8852 17872 8861 17912
rect 9100 17828 9140 17956
rect 10732 17872 11780 17912
rect 2563 17788 2572 17828
rect 2612 17788 2995 17828
rect 3035 17788 3044 17828
rect 3772 17788 3860 17828
rect 4099 17788 4108 17828
rect 4148 17788 4300 17828
rect 4340 17788 4349 17828
rect 4522 17819 5164 17828
rect 1708 17744 1748 17753
rect 2476 17744 2516 17753
rect 3628 17744 3668 17753
rect 3772 17744 3812 17788
rect 4522 17779 4531 17819
rect 4571 17788 5164 17819
rect 5204 17788 5213 17828
rect 6787 17788 6796 17828
rect 6836 17788 6845 17828
rect 7276 17788 9140 17828
rect 9292 17788 9772 17828
rect 9812 17788 9821 17828
rect 4571 17779 4580 17788
rect 4522 17778 4580 17779
rect 6796 17744 6836 17788
rect 7276 17744 7316 17788
rect 9292 17744 9332 17788
rect 10732 17744 10772 17872
rect 11740 17828 11780 17872
rect 18124 17828 18164 18292
rect 18651 18124 18660 18164
rect 19028 18124 19037 18164
rect 18211 17956 18220 17996
rect 18260 17956 18391 17996
rect 19625 17956 19756 17996
rect 19796 17956 19805 17996
rect 10819 17788 10828 17828
rect 10868 17788 11212 17828
rect 11252 17788 11261 17828
rect 11722 17788 11731 17828
rect 11771 17788 11780 17828
rect 12988 17788 13036 17828
rect 13076 17788 13085 17828
rect 13132 17788 13708 17828
rect 13748 17788 13757 17828
rect 13891 17788 13900 17828
rect 13940 17788 15668 17828
rect 18124 17788 18836 17828
rect 12988 17744 13028 17788
rect 13132 17744 13172 17788
rect 15148 17744 15188 17788
rect 15628 17744 15668 17788
rect 18796 17744 18836 17788
rect 1577 17704 1708 17744
rect 1748 17704 1757 17744
rect 2153 17704 2177 17744
rect 2217 17704 2284 17744
rect 2324 17704 2333 17744
rect 3181 17704 3190 17744
rect 3230 17704 3532 17744
rect 3572 17704 3581 17744
rect 3763 17704 3772 17744
rect 3812 17704 3821 17744
rect 3898 17704 3907 17744
rect 3947 17704 3956 17744
rect 4003 17704 4012 17744
rect 4052 17704 4396 17744
rect 4436 17704 4445 17744
rect 4624 17704 4633 17744
rect 4673 17704 4780 17744
rect 4820 17704 4876 17744
rect 4916 17704 4925 17744
rect 4972 17704 4995 17744
rect 5035 17704 5044 17744
rect 5104 17704 5113 17744
rect 5153 17704 5260 17744
rect 5300 17704 5309 17744
rect 5609 17704 5740 17744
rect 5780 17704 5789 17744
rect 5868 17704 5932 17744
rect 5972 17704 6028 17744
rect 6068 17704 6508 17744
rect 6548 17704 6604 17744
rect 6644 17704 6653 17744
rect 6749 17704 6795 17744
rect 6835 17704 6844 17744
rect 6979 17704 6988 17744
rect 7028 17704 7037 17744
rect 7162 17704 7171 17744
rect 7211 17704 7316 17744
rect 7363 17704 7372 17744
rect 7412 17704 7488 17744
rect 7546 17704 7555 17744
rect 7595 17704 7604 17744
rect 7651 17704 7660 17744
rect 7700 17704 8083 17744
rect 8123 17704 8132 17744
rect 8269 17704 8278 17744
rect 8318 17704 8428 17744
rect 8468 17704 8477 17744
rect 8995 17704 9004 17744
rect 9044 17704 9053 17744
rect 9283 17704 9292 17744
rect 9332 17704 9341 17744
rect 9402 17704 9411 17744
rect 9451 17704 9460 17744
rect 9520 17704 9529 17744
rect 9569 17704 9676 17744
rect 9716 17704 9738 17744
rect 9859 17704 9868 17744
rect 9908 17704 10060 17744
rect 10100 17704 10109 17744
rect 10217 17704 10348 17744
rect 10388 17704 10397 17744
rect 10531 17704 10540 17744
rect 10580 17704 10732 17744
rect 10772 17704 10781 17744
rect 10915 17704 10924 17744
rect 10964 17704 10973 17744
rect 11054 17704 11063 17744
rect 11103 17704 11112 17744
rect 11194 17704 11203 17744
rect 11243 17704 11252 17744
rect 11299 17704 11308 17744
rect 11348 17704 11479 17744
rect 11917 17704 11926 17744
rect 11966 17704 13028 17744
rect 13114 17704 13123 17744
rect 13163 17704 13172 17744
rect 13289 17704 13420 17744
rect 13460 17704 13469 17744
rect 14797 17704 14806 17744
rect 14846 17704 15092 17744
rect 15139 17704 15148 17744
rect 15188 17704 15197 17744
rect 15305 17704 15436 17744
rect 15476 17704 15485 17744
rect 15619 17704 15628 17744
rect 15668 17704 15799 17744
rect 15994 17704 16003 17744
rect 16043 17704 16204 17744
rect 16244 17704 16492 17744
rect 16532 17704 16541 17744
rect 16675 17704 16684 17744
rect 16724 17704 16855 17744
rect 17417 17704 17548 17744
rect 17588 17704 17597 17744
rect 17708 17704 17717 17744
rect 17757 17704 17766 17744
rect 17914 17704 17923 17744
rect 17963 17704 18164 17744
rect 18211 17704 18220 17744
rect 18271 17704 18391 17744
rect 18796 17704 19459 17744
rect 19499 17704 19508 17744
rect 19721 17704 19770 17744
rect 19810 17704 19852 17744
rect 19892 17704 19901 17744
rect 1708 17695 1748 17704
rect 2476 17660 2516 17704
rect 3628 17660 3668 17704
rect 3916 17660 3956 17704
rect 4396 17660 4436 17704
rect 4972 17660 5012 17704
rect 6988 17660 7028 17704
rect 7448 17660 7488 17704
rect 1400 17620 1409 17660
rect 1449 17620 1612 17660
rect 1652 17620 1661 17660
rect 2476 17620 2572 17660
rect 2612 17620 2621 17660
rect 3209 17620 3329 17660
rect 3380 17620 3389 17660
rect 3628 17620 3860 17660
rect 3916 17620 4012 17660
rect 4052 17620 4061 17660
rect 4108 17620 4300 17660
rect 4340 17620 4349 17660
rect 4396 17620 4820 17660
rect 4867 17620 4876 17660
rect 4916 17620 5068 17660
rect 5108 17620 5172 17660
rect 6569 17620 6700 17660
rect 6740 17620 6749 17660
rect 6988 17620 7276 17660
rect 7316 17620 7488 17660
rect 7564 17660 7604 17704
rect 9004 17660 9044 17704
rect 9411 17660 9451 17704
rect 7564 17620 8716 17660
rect 8756 17620 8765 17660
rect 9004 17620 9196 17660
rect 9236 17620 9245 17660
rect 9411 17620 9484 17660
rect 9524 17620 9533 17660
rect 1603 17536 1612 17576
rect 1652 17536 1661 17576
rect 2345 17536 2380 17576
rect 2420 17536 2476 17576
rect 2516 17536 2525 17576
rect 2947 17536 2956 17576
rect 2996 17536 3427 17576
rect 3467 17536 3476 17576
rect 3523 17536 3532 17576
rect 3572 17536 3628 17576
rect 3668 17536 3703 17576
rect 1612 17492 1652 17536
rect 3532 17492 3572 17536
rect 1027 17452 1036 17492
rect 1076 17452 1324 17492
rect 1364 17452 3572 17492
rect 3820 17492 3860 17620
rect 4108 17492 4148 17620
rect 4780 17576 4820 17620
rect 7448 17576 7488 17620
rect 9580 17576 9620 17704
rect 10540 17660 10580 17704
rect 10924 17660 10964 17704
rect 11063 17660 11103 17704
rect 10060 17620 10580 17660
rect 10627 17620 10636 17660
rect 10676 17620 10964 17660
rect 11011 17620 11020 17660
rect 11060 17620 11103 17660
rect 10060 17576 10100 17620
rect 11212 17576 11252 17704
rect 15052 17660 15092 17704
rect 17717 17660 17757 17704
rect 18124 17660 18164 17704
rect 19948 17660 19988 18292
rect 23020 18248 23060 18292
rect 23020 18208 26188 18248
rect 26228 18208 26237 18248
rect 26425 18124 26434 18164
rect 26802 18124 26811 18164
rect 22505 17956 22636 17996
rect 22676 17956 26860 17996
rect 26900 17956 26909 17996
rect 27523 17956 27532 17996
rect 27572 17956 27724 17996
rect 27764 17956 27773 17996
rect 23404 17872 25324 17912
rect 25364 17872 25373 17912
rect 22636 17788 23156 17828
rect 22636 17744 22676 17788
rect 23116 17744 23156 17788
rect 23404 17744 23444 17872
rect 24172 17788 24884 17828
rect 24172 17744 24212 17788
rect 24844 17744 24884 17788
rect 25900 17788 27148 17828
rect 27188 17788 27197 17828
rect 25900 17744 25940 17788
rect 28300 17744 28340 18376
rect 31276 17996 31316 18460
rect 30691 17956 30700 17996
rect 30740 17956 31316 17996
rect 29705 17872 29836 17912
rect 29876 17872 29885 17912
rect 30857 17872 30892 17912
rect 30932 17872 30988 17912
rect 31028 17872 31037 17912
rect 28387 17788 28396 17828
rect 28436 17788 29300 17828
rect 29260 17744 29300 17788
rect 22339 17704 22348 17744
rect 22388 17704 22636 17744
rect 22676 17704 22685 17744
rect 22808 17704 22924 17744
rect 22979 17704 22988 17744
rect 23098 17735 23156 17744
rect 23098 17695 23107 17735
rect 23147 17695 23156 17735
rect 23395 17704 23404 17744
rect 23444 17704 23453 17744
rect 24163 17704 24172 17744
rect 24212 17704 24221 17744
rect 24329 17704 24460 17744
rect 24500 17704 24509 17744
rect 24713 17704 24844 17744
rect 24884 17704 24893 17744
rect 24979 17704 24988 17744
rect 25028 17704 25036 17744
rect 25076 17704 25159 17744
rect 25891 17704 25900 17744
rect 25940 17704 25949 17744
rect 26083 17704 26092 17744
rect 26132 17704 26263 17744
rect 27331 17704 27340 17744
rect 27380 17704 27628 17744
rect 27668 17704 27677 17744
rect 27811 17704 27820 17744
rect 27860 17704 27869 17744
rect 28300 17704 28396 17744
rect 28436 17704 28445 17744
rect 28570 17704 28579 17744
rect 28628 17704 28759 17744
rect 29251 17704 29260 17744
rect 29300 17704 29309 17744
rect 30019 17704 30028 17744
rect 30068 17704 30077 17744
rect 23098 17694 23156 17695
rect 11386 17620 11395 17660
rect 11444 17620 11575 17660
rect 12931 17620 12940 17660
rect 12980 17620 13900 17660
rect 13940 17620 13949 17660
rect 15052 17620 15532 17660
rect 15572 17620 15581 17660
rect 16305 17620 16314 17660
rect 16354 17620 16588 17660
rect 16628 17620 16637 17660
rect 17251 17620 17260 17660
rect 17300 17620 17836 17660
rect 17876 17620 17917 17660
rect 18115 17620 18124 17660
rect 18164 17620 18173 17660
rect 19372 17620 19988 17660
rect 23203 17620 23212 17660
rect 23252 17620 24364 17660
rect 24404 17620 24413 17660
rect 24521 17620 24643 17660
rect 24692 17620 24701 17660
rect 4649 17536 4780 17576
rect 4820 17536 4829 17576
rect 7075 17536 7084 17576
rect 7124 17536 7133 17576
rect 7448 17536 8948 17576
rect 9283 17536 9292 17576
rect 9332 17536 9620 17576
rect 9672 17536 10100 17576
rect 10435 17536 10444 17576
rect 10484 17536 10493 17576
rect 10723 17536 10732 17576
rect 10772 17536 11252 17576
rect 14467 17536 14476 17576
rect 14516 17536 14611 17576
rect 14651 17536 14660 17576
rect 14825 17536 14860 17576
rect 14900 17536 14956 17576
rect 14996 17536 15005 17576
rect 15226 17536 15235 17576
rect 15275 17536 15436 17576
rect 15476 17536 15485 17576
rect 16090 17536 16099 17576
rect 16139 17536 16148 17576
rect 17635 17536 17644 17576
rect 17684 17536 17693 17576
rect 17897 17536 18019 17576
rect 18068 17536 18077 17576
rect 7084 17492 7124 17536
rect 8908 17492 8948 17536
rect 9672 17492 9712 17536
rect 10444 17492 10484 17536
rect 16108 17492 16148 17536
rect 3820 17452 4148 17492
rect 4780 17452 7124 17492
rect 8899 17452 8908 17492
rect 8948 17452 9712 17492
rect 9955 17452 9964 17492
rect 10004 17452 10013 17492
rect 10444 17452 12556 17492
rect 12596 17452 12605 17492
rect 13507 17452 13516 17492
rect 13556 17452 16148 17492
rect 17644 17492 17684 17536
rect 17644 17452 19276 17492
rect 19316 17452 19325 17492
rect 4343 17368 4352 17408
rect 4720 17368 4729 17408
rect 4780 17240 4820 17452
rect 9964 17408 10004 17452
rect 19372 17408 19412 17620
rect 25900 17576 25940 17704
rect 27820 17660 27860 17704
rect 30028 17660 30068 17704
rect 27820 17620 28108 17660
rect 28148 17620 28300 17660
rect 28340 17620 28349 17660
rect 28483 17620 28492 17660
rect 28532 17620 30068 17660
rect 19546 17536 19555 17576
rect 19595 17536 19604 17576
rect 23587 17536 23596 17576
rect 23636 17536 23971 17576
rect 24011 17536 24020 17576
rect 24259 17536 24268 17576
rect 24308 17536 24460 17576
rect 24500 17536 24940 17576
rect 24980 17536 25940 17576
rect 25987 17536 25996 17576
rect 26036 17536 26045 17576
rect 29146 17536 29155 17576
rect 29195 17536 29204 17576
rect 29443 17536 29452 17576
rect 29492 17536 31276 17576
rect 31316 17536 31325 17576
rect 8419 17368 8428 17408
rect 8468 17368 10004 17408
rect 12117 17368 12126 17408
rect 12494 17368 12503 17408
rect 12556 17368 19412 17408
rect 12556 17324 12596 17368
rect 19564 17324 19604 17536
rect 19891 17368 19900 17408
rect 20268 17368 20277 17408
rect 25996 17324 26036 17536
rect 27665 17368 27674 17408
rect 28042 17368 28051 17408
rect 4963 17284 4972 17324
rect 5012 17284 12596 17324
rect 12931 17284 12940 17324
rect 12980 17284 13228 17324
rect 13268 17284 13277 17324
rect 17356 17284 19124 17324
rect 19564 17284 20564 17324
rect 13420 17240 13460 17249
rect 844 17200 1612 17240
rect 1652 17200 1661 17240
rect 2275 17200 2284 17240
rect 2324 17200 2708 17240
rect 844 17156 884 17200
rect 632 17116 641 17156
rect 681 17116 884 17156
rect 940 17116 1900 17156
rect 1940 17116 1949 17156
rect 2179 17116 2188 17156
rect 2228 17116 2282 17156
rect 835 17032 844 17072
rect 884 17032 893 17072
rect 940 17063 980 17116
rect 2242 17072 2282 17116
rect 844 16904 884 17032
rect 940 17014 980 17023
rect 1036 17032 1315 17072
rect 1364 17032 1373 17072
rect 1987 17032 1996 17072
rect 2036 17032 2092 17072
rect 2132 17032 2167 17072
rect 2224 17032 2233 17072
rect 2273 17032 2282 17072
rect 2345 17116 2476 17156
rect 2516 17116 2525 17156
rect 2345 17072 2385 17116
rect 2668 17072 2708 17200
rect 3532 17200 4820 17240
rect 5033 17200 5164 17240
rect 5204 17200 5213 17240
rect 6089 17200 6172 17240
rect 6212 17200 6220 17240
rect 6260 17200 6269 17240
rect 8969 17200 9100 17240
rect 9140 17200 9149 17240
rect 11011 17200 11020 17240
rect 11060 17200 11107 17240
rect 11147 17200 11191 17240
rect 11395 17200 11404 17240
rect 11444 17200 11587 17240
rect 11627 17200 11636 17240
rect 12460 17200 13420 17240
rect 13460 17200 13708 17240
rect 13748 17200 13757 17240
rect 16745 17200 16867 17240
rect 16916 17200 16925 17240
rect 3532 17072 3572 17200
rect 4396 17116 4867 17156
rect 4907 17116 4916 17156
rect 4963 17116 4972 17156
rect 5012 17116 6595 17156
rect 6635 17116 7124 17156
rect 8201 17116 8236 17156
rect 8276 17116 8332 17156
rect 8372 17116 8381 17156
rect 9065 17147 9196 17156
rect 9065 17116 9187 17147
rect 9236 17116 9245 17156
rect 10627 17116 10636 17156
rect 10676 17116 10685 17156
rect 10810 17116 10819 17156
rect 10859 17116 11006 17156
rect 11046 17116 11055 17156
rect 11175 17116 11212 17156
rect 11252 17116 11261 17156
rect 11683 17116 11692 17156
rect 11732 17116 11884 17156
rect 11924 17116 11933 17156
rect 2345 17032 2380 17072
rect 2420 17032 2429 17072
rect 2544 17032 2553 17072
rect 2593 17032 2602 17072
rect 2668 17032 2764 17072
rect 2804 17032 2813 17072
rect 2938 17032 2947 17072
rect 2987 17032 3572 17072
rect 3619 17032 3628 17072
rect 3668 17032 4195 17072
rect 4235 17032 4244 17072
rect 1036 16904 1076 17032
rect 2558 16988 2598 17032
rect 4396 16988 4436 17116
rect 7084 17072 7124 17116
rect 9178 17107 9187 17116
rect 9227 17107 9236 17116
rect 9178 17106 9236 17107
rect 10636 17072 10676 17116
rect 11175 17114 11215 17116
rect 11116 17074 11215 17114
rect 11116 17072 11156 17074
rect 12460 17072 12500 17200
rect 13420 17191 13460 17200
rect 13603 17116 13612 17156
rect 13652 17116 15284 17156
rect 15244 17072 15284 17116
rect 17356 17072 17396 17284
rect 19084 17240 19124 17284
rect 17923 17200 17932 17240
rect 17972 17200 18884 17240
rect 18970 17200 18979 17240
rect 19019 17200 19028 17240
rect 19084 17200 20428 17240
rect 20468 17200 20477 17240
rect 18844 17156 18884 17200
rect 18988 17156 19028 17200
rect 20524 17156 20564 17284
rect 23020 17284 26036 17324
rect 23020 17156 23060 17284
rect 29164 17240 29204 17536
rect 17827 17116 17836 17156
rect 17876 17116 17923 17156
rect 17993 17116 18028 17156
rect 18068 17147 18164 17156
rect 18068 17116 18115 17147
rect 17836 17072 17876 17116
rect 18106 17107 18115 17116
rect 18155 17107 18164 17147
rect 18211 17116 18220 17156
rect 18260 17116 18394 17156
rect 18844 17116 18944 17156
rect 18988 17116 20276 17156
rect 20410 17116 20419 17156
rect 20459 17116 20564 17156
rect 20611 17116 20620 17156
rect 20660 17116 20852 17156
rect 18106 17106 18164 17107
rect 18354 17072 18394 17116
rect 18904 17072 18944 17116
rect 20236 17072 20276 17116
rect 20812 17072 20852 17116
rect 21772 17116 23060 17156
rect 23692 17200 24556 17240
rect 24596 17200 25747 17240
rect 25787 17200 25796 17240
rect 29164 17200 29356 17240
rect 29396 17200 29405 17240
rect 21772 17072 21812 17116
rect 23692 17072 23732 17200
rect 23884 17116 23980 17156
rect 24020 17116 24029 17156
rect 24137 17116 24268 17156
rect 24308 17116 24317 17156
rect 24465 17116 24474 17156
rect 24514 17116 25036 17156
rect 25076 17116 25085 17156
rect 28588 17116 30892 17156
rect 30932 17116 30941 17156
rect 23884 17072 23924 17116
rect 28588 17072 28628 17116
rect 4483 17032 4492 17072
rect 4532 17032 4535 17072
rect 4575 17032 4663 17072
rect 4771 17032 4780 17072
rect 4820 17032 4829 17072
rect 5021 17032 5063 17072
rect 5103 17032 5112 17072
rect 5242 17032 5251 17072
rect 5291 17032 5300 17072
rect 5539 17032 5548 17072
rect 5588 17032 6028 17072
rect 6068 17032 6077 17072
rect 6979 17032 6988 17072
rect 7028 17032 7037 17072
rect 7084 17032 8140 17072
rect 8180 17032 8189 17072
rect 8236 17032 8443 17072
rect 8483 17032 8492 17072
rect 8777 17032 8899 17072
rect 8948 17032 8957 17072
rect 9004 17063 9044 17072
rect 4780 16988 4820 17032
rect 5068 16988 5108 17032
rect 5260 16988 5300 17032
rect 1123 16948 1132 16988
rect 1172 16948 1181 16988
rect 1603 16948 1612 16988
rect 1652 16948 1708 16988
rect 1748 16948 1783 16988
rect 2122 16979 2180 16988
rect 844 16864 1076 16904
rect 521 16780 643 16820
rect 692 16780 701 16820
rect 1132 16316 1172 16948
rect 2122 16939 2131 16979
rect 2171 16939 2180 16979
rect 2558 16948 2860 16988
rect 2900 16948 2909 16988
rect 3715 16948 3724 16988
rect 3764 16948 3811 16988
rect 3851 16948 3895 16988
rect 4378 16948 4387 16988
rect 4427 16948 4436 16988
rect 4666 16948 4675 16988
rect 4715 16948 4724 16988
rect 4771 16948 4780 16988
rect 4820 16948 4867 16988
rect 5059 16948 5068 16988
rect 5108 16948 5117 16988
rect 5260 16948 6700 16988
rect 6740 16948 6749 16988
rect 2122 16938 2180 16939
rect 2140 16904 2180 16938
rect 1603 16864 1612 16904
rect 1652 16864 1996 16904
rect 2036 16864 2045 16904
rect 2140 16864 2284 16904
rect 2324 16864 2333 16904
rect 3785 16864 3907 16904
rect 3956 16864 3965 16904
rect 2249 16780 2380 16820
rect 2420 16780 2429 16820
rect 2860 16780 2947 16820
rect 2987 16780 2996 16820
rect 2860 16736 2900 16780
rect 1219 16696 1228 16736
rect 1268 16696 2900 16736
rect 3103 16612 3112 16652
rect 3480 16612 3489 16652
rect 4684 16484 4724 16948
rect 6988 16904 7028 17032
rect 8236 16988 8276 17032
rect 9270 17032 9279 17072
rect 9319 17032 9332 17072
rect 9451 17032 9460 17072
rect 9524 17032 9640 17072
rect 10498 17032 10507 17072
rect 10547 17032 10676 17072
rect 10723 17032 10732 17072
rect 10772 17032 10828 17072
rect 10868 17032 10903 17072
rect 11011 17032 11020 17072
rect 11060 17032 11156 17072
rect 9004 16988 9044 17023
rect 9292 16988 9332 17032
rect 11266 17030 11298 17047
rect 11233 17007 11298 17030
rect 11338 17007 11347 17047
rect 11482 17032 11491 17072
rect 11531 17032 11540 17072
rect 11683 17032 11692 17072
rect 11732 17032 11799 17072
rect 11839 17032 11863 17072
rect 12451 17032 12460 17072
rect 12500 17032 12509 17072
rect 12778 17032 12787 17072
rect 12827 17032 13027 17072
rect 13067 17032 13420 17072
rect 13460 17032 13564 17072
rect 13604 17032 13613 17072
rect 13795 17032 13804 17072
rect 13844 17032 13900 17072
rect 13940 17032 13975 17072
rect 14755 17032 14764 17072
rect 14804 17032 14872 17072
rect 14912 17032 14935 17072
rect 15226 17063 15628 17072
rect 11233 16990 11306 17007
rect 11233 16988 11273 16990
rect 8227 16948 8236 16988
rect 8276 16948 8285 16988
rect 8995 16948 9004 16988
rect 9044 16948 9091 16988
rect 9283 16948 9292 16988
rect 9332 16948 9375 16988
rect 10505 16948 10627 16988
rect 10676 16948 10685 16988
rect 11203 16948 11212 16988
rect 11252 16948 11273 16988
rect 10636 16904 10676 16948
rect 11500 16904 11540 17032
rect 15226 17023 15235 17063
rect 15275 17032 15628 17063
rect 15668 17032 15677 17072
rect 15994 17032 16003 17072
rect 16043 17032 16052 17072
rect 16291 17032 16300 17072
rect 16340 17032 16780 17072
rect 16820 17032 17356 17072
rect 17396 17032 17405 17072
rect 17644 17032 17659 17072
rect 17699 17032 17708 17072
rect 17818 17032 17827 17072
rect 17867 17032 17876 17072
rect 17932 17063 17972 17072
rect 15275 17023 15284 17032
rect 15226 17022 15284 17023
rect 16012 16988 16052 17032
rect 17644 16988 17684 17032
rect 18197 17032 18206 17072
rect 18246 17032 18260 17072
rect 18354 17032 18387 17072
rect 18427 17032 18628 17072
rect 18668 17032 18677 17072
rect 18778 17047 18787 17072
rect 18719 17032 18787 17047
rect 18827 17032 18836 17072
rect 18895 17032 18904 17072
rect 18944 17032 18953 17072
rect 19036 17032 19075 17072
rect 19115 17032 19124 17072
rect 19188 17032 19197 17072
rect 19237 17032 19276 17072
rect 19316 17032 19377 17072
rect 19721 17032 19756 17072
rect 19796 17032 19852 17072
rect 19892 17032 19901 17072
rect 19948 17032 20087 17072
rect 20127 17032 20136 17072
rect 20236 17032 20332 17072
rect 20372 17032 20381 17072
rect 20611 17032 20620 17072
rect 20660 17032 20669 17072
rect 20794 17032 20803 17072
rect 20843 17032 21044 17072
rect 21257 17032 21388 17072
rect 21428 17032 21437 17072
rect 21508 17032 21517 17072
rect 21557 17032 21580 17072
rect 21620 17032 21697 17072
rect 21763 17032 21772 17072
rect 21812 17032 21821 17072
rect 22409 17032 22540 17072
rect 22580 17063 22868 17072
rect 22580 17032 22819 17063
rect 12451 16948 12460 16988
rect 12500 16948 14572 16988
rect 14612 16948 14707 16988
rect 14747 16948 14756 16988
rect 15379 16948 15388 16988
rect 15428 16948 16108 16988
rect 16148 16948 16876 16988
rect 16916 16948 17740 16988
rect 17780 16948 17789 16988
rect 17932 16904 17972 17023
rect 18220 16988 18260 17032
rect 18719 17007 18836 17032
rect 18719 16988 18759 17007
rect 18172 16948 18759 16988
rect 6988 16864 8908 16904
rect 8948 16864 8957 16904
rect 10636 16864 11540 16904
rect 13114 16864 13123 16904
rect 13163 16864 14284 16904
rect 14324 16864 14333 16904
rect 14755 16864 14764 16904
rect 14804 16864 16396 16904
rect 16436 16864 16588 16904
rect 16628 16864 16684 16904
rect 16724 16864 16788 16904
rect 17347 16864 17356 16904
rect 17396 16864 17932 16904
rect 17972 16864 17981 16904
rect 12521 16780 12652 16820
rect 12692 16780 12701 16820
rect 13315 16780 13324 16820
rect 13364 16780 13699 16820
rect 13739 16780 13748 16820
rect 13795 16780 13804 16820
rect 13844 16780 15244 16820
rect 15284 16780 15820 16820
rect 15860 16780 15869 16820
rect 17417 16780 17548 16820
rect 17588 16780 17597 16820
rect 17818 16780 17827 16820
rect 17867 16780 18028 16820
rect 18068 16780 18077 16820
rect 18172 16736 18212 16948
rect 8803 16696 8812 16736
rect 8852 16696 12556 16736
rect 12596 16696 12605 16736
rect 15139 16696 15148 16736
rect 15188 16696 18212 16736
rect 19036 16736 19076 17032
rect 19948 16988 19988 17032
rect 20620 16988 20660 17032
rect 19555 16948 19564 16988
rect 19604 16948 19988 16988
rect 20218 16948 20227 16988
rect 20267 16948 20524 16988
rect 20564 16948 20573 16988
rect 20620 16948 20948 16988
rect 19267 16864 19276 16904
rect 19316 16864 19459 16904
rect 19499 16864 19508 16904
rect 19747 16864 19756 16904
rect 19796 16864 20803 16904
rect 20843 16864 20852 16904
rect 20908 16820 20948 16948
rect 21004 16904 21044 17032
rect 22810 17023 22819 17032
rect 22859 17023 22868 17063
rect 23683 17032 23692 17072
rect 23732 17032 23741 17072
rect 23866 17032 23875 17072
rect 23915 17032 23924 17072
rect 23971 17032 23980 17072
rect 24020 17032 24029 17072
rect 24165 17032 24174 17072
rect 24214 17032 24844 17072
rect 24884 17032 24893 17072
rect 25315 17032 25324 17072
rect 25364 17032 25942 17072
rect 25982 17032 27148 17072
rect 27188 17032 27197 17072
rect 28570 17032 28579 17072
rect 28619 17032 28628 17072
rect 29356 17032 30028 17072
rect 30068 17032 30077 17072
rect 22810 17022 22868 17023
rect 23982 16988 24022 17032
rect 22963 16948 22972 16988
rect 23012 16948 23020 16988
rect 23060 16948 23143 16988
rect 23982 16948 24652 16988
rect 24692 16948 24701 16988
rect 24748 16948 27043 16988
rect 27083 16948 27092 16988
rect 28387 16948 28396 16988
rect 28436 16948 28445 16988
rect 28954 16948 28963 16988
rect 29003 16948 29012 16988
rect 24748 16904 24788 16948
rect 21004 16864 21100 16904
rect 21140 16864 21149 16904
rect 23299 16864 23308 16904
rect 23348 16864 24788 16904
rect 26284 16864 27183 16904
rect 20131 16780 20140 16820
rect 20180 16780 20948 16820
rect 22025 16780 22147 16820
rect 22196 16780 22205 16820
rect 23971 16780 23980 16820
rect 24020 16780 24268 16820
rect 24308 16780 24317 16820
rect 24451 16780 24460 16820
rect 24500 16780 24631 16820
rect 24835 16780 24844 16820
rect 24884 16780 24931 16820
rect 24971 16780 25015 16820
rect 19036 16696 19316 16736
rect 19276 16652 19316 16696
rect 10877 16612 10886 16652
rect 11254 16612 11263 16652
rect 11308 16612 12844 16652
rect 12884 16612 12893 16652
rect 18651 16612 18660 16652
rect 19028 16612 19037 16652
rect 19267 16612 19276 16652
rect 19316 16612 19325 16652
rect 19939 16612 19948 16652
rect 19988 16612 21868 16652
rect 21908 16612 21917 16652
rect 11308 16568 11348 16612
rect 8227 16528 8236 16568
rect 8276 16528 9484 16568
rect 9524 16528 9533 16568
rect 9763 16528 9772 16568
rect 9812 16528 11348 16568
rect 11404 16528 12212 16568
rect 11404 16484 11444 16528
rect 12172 16484 12212 16528
rect 19372 16528 24844 16568
rect 24884 16528 24893 16568
rect 2275 16444 2284 16484
rect 2324 16444 2659 16484
rect 2699 16444 2708 16484
rect 4291 16444 4300 16484
rect 4340 16444 4724 16484
rect 6569 16444 6691 16484
rect 6740 16444 6749 16484
rect 7241 16444 7363 16484
rect 7412 16444 7421 16484
rect 8995 16444 9004 16484
rect 9044 16444 9964 16484
rect 10004 16444 10013 16484
rect 10435 16444 10444 16484
rect 10484 16444 11444 16484
rect 11779 16444 11788 16484
rect 11828 16444 12067 16484
rect 12107 16444 12116 16484
rect 12172 16444 14188 16484
rect 14228 16444 14237 16484
rect 14371 16444 14380 16484
rect 14420 16444 16099 16484
rect 16139 16444 16148 16484
rect 16457 16444 16588 16484
rect 16628 16444 16637 16484
rect 17731 16444 17740 16484
rect 17780 16444 17827 16484
rect 17867 16444 17911 16484
rect 18019 16444 18028 16484
rect 18068 16444 18796 16484
rect 18836 16444 18845 16484
rect 19372 16400 19412 16528
rect 26284 16484 26324 16864
rect 27143 16820 27183 16864
rect 28972 16820 29012 16948
rect 26659 16780 26668 16820
rect 26708 16780 27052 16820
rect 27092 16780 27101 16820
rect 27143 16780 29012 16820
rect 26425 16612 26434 16652
rect 26802 16612 26811 16652
rect 29356 16568 29396 17032
rect 30281 16864 30412 16904
rect 30452 16864 30461 16904
rect 30595 16864 30604 16904
rect 30644 16864 30775 16904
rect 4684 16360 5068 16400
rect 5108 16360 5117 16400
rect 6508 16360 7276 16400
rect 7316 16360 7325 16400
rect 8995 16360 9004 16400
rect 9044 16360 9196 16400
rect 9236 16360 9245 16400
rect 9955 16360 9964 16400
rect 10004 16360 12117 16400
rect 12835 16360 12844 16400
rect 12884 16360 19412 16400
rect 19516 16444 19756 16484
rect 19796 16444 19805 16484
rect 21571 16444 21580 16484
rect 21620 16444 23060 16484
rect 23491 16444 23500 16484
rect 23540 16444 24556 16484
rect 24596 16444 24605 16484
rect 26083 16444 26092 16484
rect 26132 16444 26324 16484
rect 26956 16528 29396 16568
rect 1132 16276 1420 16316
rect 1460 16276 1469 16316
rect 1577 16276 1612 16316
rect 1652 16276 1708 16316
rect 1748 16276 1757 16316
rect 1834 16307 2764 16316
rect 1834 16267 1843 16307
rect 1883 16276 2764 16307
rect 2804 16276 2813 16316
rect 1883 16267 1892 16276
rect 1834 16266 1892 16267
rect 2956 16232 2996 16241
rect 4684 16232 4724 16360
rect 5644 16276 5972 16316
rect 5644 16274 5684 16276
rect 5578 16234 5587 16274
rect 5627 16234 5684 16274
rect 5932 16232 5972 16276
rect 6508 16232 6548 16360
rect 6857 16276 6892 16316
rect 6932 16276 6979 16316
rect 7019 16276 7037 16316
rect 7171 16276 7180 16316
rect 7220 16276 7679 16316
rect 7639 16232 7679 16276
rect 7756 16276 9004 16316
rect 9044 16276 9053 16316
rect 10601 16276 10732 16316
rect 10772 16276 10781 16316
rect 7756 16232 7796 16276
rect 10828 16232 10868 16360
rect 12077 16316 12117 16360
rect 12077 16276 12268 16316
rect 12308 16276 12317 16316
rect 18499 16276 18508 16316
rect 18548 16276 19276 16316
rect 19355 16276 19364 16316
rect 19516 16274 19556 16444
rect 23020 16400 23060 16444
rect 26956 16400 26996 16528
rect 29356 16484 29396 16528
rect 27139 16444 27148 16484
rect 27188 16444 28972 16484
rect 29012 16444 29021 16484
rect 29347 16444 29356 16484
rect 29396 16444 29405 16484
rect 20131 16360 20140 16400
rect 20180 16360 22828 16400
rect 22868 16360 22877 16400
rect 23020 16360 26996 16400
rect 28265 16360 28396 16400
rect 28436 16360 28445 16400
rect 19651 16276 19660 16316
rect 19700 16276 19709 16316
rect 21353 16276 21484 16316
rect 21524 16276 21533 16316
rect 21859 16276 21868 16316
rect 21908 16276 23396 16316
rect 23578 16276 23587 16316
rect 23636 16276 23767 16316
rect 23932 16276 24268 16316
rect 24308 16276 24317 16316
rect 26083 16276 26092 16316
rect 26132 16276 26660 16316
rect 12364 16232 12404 16241
rect 16396 16232 16436 16241
rect 19498 16234 19507 16274
rect 19547 16234 19556 16274
rect 19660 16232 19700 16276
rect 21004 16232 21044 16241
rect 23356 16232 23396 16276
rect 23932 16232 23972 16276
rect 26620 16232 26660 16276
rect 26845 16276 26860 16316
rect 26900 16276 26909 16316
rect 27043 16276 27052 16316
rect 27092 16276 27188 16316
rect 27811 16276 27820 16316
rect 27860 16276 28244 16316
rect 30595 16276 30604 16316
rect 30644 16276 30653 16316
rect 31258 16276 31267 16316
rect 31316 16276 31447 16316
rect 26845 16274 26885 16276
rect 26755 16234 26764 16274
rect 26804 16234 26885 16274
rect 27148 16232 27188 16276
rect 28204 16232 28244 16276
rect 948 16192 1036 16232
rect 1076 16192 1079 16232
rect 1119 16192 1128 16232
rect 1210 16192 1219 16232
rect 1259 16192 1268 16232
rect 1315 16192 1324 16232
rect 1364 16192 1708 16232
rect 1748 16192 1757 16232
rect 1936 16192 1945 16232
rect 1985 16192 2188 16232
rect 2228 16192 2237 16232
rect 2284 16192 2307 16232
rect 2347 16192 2356 16232
rect 2416 16192 2425 16232
rect 2465 16192 2668 16232
rect 2708 16192 2717 16232
rect 2996 16192 3628 16232
rect 3668 16192 3677 16232
rect 3881 16192 4003 16232
rect 4052 16192 4061 16232
rect 4305 16192 4314 16232
rect 4354 16192 4481 16232
rect 4521 16192 4724 16232
rect 4777 16192 4786 16232
rect 4826 16192 4876 16232
rect 4916 16192 4966 16232
rect 5321 16192 5395 16232
rect 5435 16192 5452 16232
rect 5492 16192 5501 16232
rect 5755 16192 5764 16232
rect 5804 16192 5876 16232
rect 5928 16192 5937 16232
rect 5977 16192 5986 16232
rect 6058 16192 6067 16232
rect 6107 16192 6116 16232
rect 6170 16192 6179 16232
rect 6219 16192 6239 16232
rect 6298 16192 6307 16232
rect 6347 16192 6508 16232
rect 6548 16192 6557 16232
rect 6682 16192 6691 16232
rect 6731 16192 6740 16232
rect 6787 16192 6796 16232
rect 6836 16192 6839 16232
rect 6879 16192 6967 16232
rect 7075 16192 7084 16232
rect 7124 16192 7180 16232
rect 7220 16192 7255 16232
rect 7346 16192 7355 16232
rect 7395 16192 7404 16232
rect 7510 16192 7519 16232
rect 7559 16192 7580 16232
rect 7638 16192 7647 16232
rect 7687 16192 7696 16232
rect 7738 16192 7747 16232
rect 7787 16192 7796 16232
rect 7915 16192 7924 16232
rect 7988 16192 8104 16232
rect 8681 16192 8758 16232
rect 8798 16192 8812 16232
rect 8852 16192 8861 16232
rect 8908 16192 9187 16232
rect 9227 16192 9428 16232
rect 9475 16192 9484 16232
rect 9524 16192 9667 16232
rect 9716 16192 9725 16232
rect 9955 16192 9964 16232
rect 10004 16192 10391 16232
rect 10431 16192 10440 16232
rect 10522 16192 10531 16232
rect 10571 16192 10580 16232
rect 10627 16192 10636 16232
rect 10676 16192 11212 16232
rect 11252 16192 11261 16232
rect 11917 16192 11926 16232
rect 11966 16192 12268 16232
rect 12308 16192 12317 16232
rect 12451 16192 12460 16232
rect 12500 16192 13036 16232
rect 13076 16192 13085 16232
rect 13146 16192 13155 16232
rect 13195 16192 13204 16232
rect 13264 16192 13273 16232
rect 13313 16192 13324 16232
rect 13364 16192 13453 16232
rect 13673 16192 13750 16232
rect 13790 16192 13804 16232
rect 13844 16192 13853 16232
rect 14825 16192 14860 16232
rect 14900 16192 14956 16232
rect 14996 16192 15005 16232
rect 15235 16192 15244 16232
rect 15284 16192 15293 16232
rect 15562 16192 15571 16232
rect 15611 16192 15820 16232
rect 15860 16192 15869 16232
rect 15977 16192 16097 16232
rect 16148 16192 16157 16232
rect 16436 16192 16439 16232
rect 16483 16192 16492 16232
rect 16532 16192 16588 16232
rect 16628 16192 16663 16232
rect 16771 16192 16780 16232
rect 16820 16192 16876 16232
rect 16916 16192 16951 16232
rect 17539 16192 17548 16232
rect 17588 16192 17644 16232
rect 17684 16192 17719 16232
rect 17818 16192 17827 16232
rect 17867 16192 18124 16232
rect 18164 16192 18173 16232
rect 19651 16192 19660 16232
rect 19700 16192 19747 16232
rect 19843 16192 19852 16232
rect 19892 16192 20180 16232
rect 20506 16192 20515 16232
rect 20555 16192 20908 16232
rect 20948 16192 20957 16232
rect 21091 16192 21100 16232
rect 21140 16192 21580 16232
rect 21620 16192 21629 16232
rect 21955 16192 21964 16232
rect 22004 16192 22013 16232
rect 22073 16192 22082 16232
rect 22122 16192 22444 16232
rect 22484 16192 22493 16232
rect 22862 16192 22871 16232
rect 22911 16192 22920 16232
rect 23002 16223 23060 16232
rect 1228 16148 1268 16192
rect 1219 16108 1228 16148
rect 1268 16108 1315 16148
rect 1708 16064 1748 16192
rect 2284 16148 2324 16192
rect 2956 16183 2996 16192
rect 5836 16148 5876 16192
rect 1795 16108 1804 16148
rect 1844 16108 2380 16148
rect 2420 16108 2654 16148
rect 2694 16108 2703 16148
rect 4291 16108 4300 16148
rect 4340 16108 4579 16148
rect 4619 16108 4628 16148
rect 5827 16108 5836 16148
rect 5876 16108 5885 16148
rect 1708 16024 2092 16064
rect 2132 16024 2141 16064
rect 2467 16024 2476 16064
rect 2516 16024 2860 16064
rect 2900 16024 4099 16064
rect 4139 16024 4684 16064
rect 4724 16024 4733 16064
rect 5705 16024 5740 16064
rect 5780 16024 5827 16064
rect 5867 16024 5885 16064
rect 5932 15896 5972 16192
rect 6067 16064 6107 16192
rect 6199 16148 6239 16192
rect 6700 16148 6740 16192
rect 7348 16148 7388 16192
rect 6199 16108 6508 16148
rect 6548 16108 6557 16148
rect 6653 16108 6700 16148
rect 6740 16108 6749 16148
rect 7267 16108 7276 16148
rect 7316 16108 7388 16148
rect 7540 16148 7580 16192
rect 7540 16108 7564 16148
rect 7604 16108 7613 16148
rect 7756 16064 7796 16192
rect 8908 16064 8948 16192
rect 6067 16024 7796 16064
rect 8515 16024 8524 16064
rect 8603 16024 8695 16064
rect 8803 16024 8812 16064
rect 8852 16024 8948 16064
rect 9388 15980 9428 16192
rect 10540 16148 10580 16192
rect 12364 16148 12404 16192
rect 13155 16148 13195 16192
rect 15244 16148 15284 16192
rect 16396 16183 16439 16192
rect 16399 16148 16439 16183
rect 20140 16148 20180 16192
rect 21004 16148 21044 16192
rect 21964 16148 22004 16192
rect 9641 16108 9772 16148
rect 9812 16108 9821 16148
rect 9868 16108 9975 16148
rect 10015 16108 10024 16148
rect 10540 16108 10636 16148
rect 10676 16108 10685 16148
rect 11683 16108 11692 16148
rect 11732 16108 12062 16148
rect 12102 16108 12111 16148
rect 12172 16108 12404 16148
rect 12460 16108 12556 16148
rect 12596 16108 13076 16148
rect 13155 16108 14380 16148
rect 14420 16108 14429 16148
rect 14563 16108 14572 16148
rect 14612 16108 15284 16148
rect 15427 16108 15436 16148
rect 15476 16108 15485 16148
rect 16399 16108 19756 16148
rect 19796 16108 19805 16148
rect 20140 16108 21196 16148
rect 21236 16108 21245 16148
rect 21571 16108 21580 16148
rect 21620 16108 22004 16148
rect 9868 16064 9908 16108
rect 12172 16064 12212 16108
rect 12460 16064 12500 16108
rect 13036 16064 13076 16108
rect 9475 16024 9484 16064
rect 9524 16024 10060 16064
rect 10100 16024 10109 16064
rect 11395 16024 11404 16064
rect 11444 16024 11731 16064
rect 11771 16024 11780 16064
rect 11971 16024 11980 16064
rect 12020 16024 12212 16064
rect 12259 16024 12268 16064
rect 12308 16024 12500 16064
rect 12931 16024 12940 16064
rect 12980 16024 12989 16064
rect 13036 16024 13324 16064
rect 13364 16024 13373 16064
rect 13507 16024 13516 16064
rect 13595 16024 14092 16064
rect 14132 16024 14141 16064
rect 14467 16024 14476 16064
rect 14516 16024 14668 16064
rect 14708 16024 14717 16064
rect 9388 15940 12844 15980
rect 12884 15940 12893 15980
rect 4343 15856 4352 15896
rect 4720 15856 4729 15896
rect 5932 15856 9964 15896
rect 10004 15856 11404 15896
rect 11444 15856 11453 15896
rect 12117 15856 12126 15896
rect 12494 15856 12503 15896
rect 12940 15812 12980 16024
rect 15436 15980 15476 16108
rect 22871 16064 22911 16192
rect 23002 16183 23011 16223
rect 23051 16183 23060 16223
rect 23107 16192 23116 16232
rect 23156 16192 23287 16232
rect 23340 16192 23447 16232
rect 23487 16192 23500 16232
rect 23540 16192 23549 16232
rect 23683 16192 23692 16232
rect 23732 16192 23863 16232
rect 23923 16192 23932 16232
rect 23972 16192 23981 16232
rect 24058 16212 24067 16232
rect 24023 16192 24067 16212
rect 24107 16192 24116 16232
rect 24163 16192 24172 16232
rect 24212 16192 24343 16232
rect 24425 16192 24460 16232
rect 24500 16192 24556 16232
rect 24596 16192 24605 16232
rect 25786 16192 25795 16232
rect 25835 16192 26324 16232
rect 26371 16192 26380 16232
rect 26420 16192 26428 16232
rect 26468 16192 26551 16232
rect 26611 16192 26620 16232
rect 26660 16192 26669 16232
rect 26947 16192 26956 16232
rect 26996 16192 27005 16232
rect 27139 16192 27148 16232
rect 27188 16192 27197 16232
rect 27331 16192 27340 16232
rect 27380 16192 28012 16232
rect 28052 16192 28061 16232
rect 28195 16192 28204 16232
rect 28244 16192 28253 16232
rect 30761 16192 30883 16232
rect 30932 16192 30941 16232
rect 23002 16182 23060 16183
rect 23020 16148 23060 16182
rect 24023 16172 24116 16192
rect 24023 16148 24063 16172
rect 23020 16108 23212 16148
rect 23252 16108 23261 16148
rect 23770 16108 23779 16148
rect 23819 16108 24063 16148
rect 26092 16108 26103 16148
rect 26143 16108 26152 16148
rect 16099 16024 16108 16064
rect 16148 16024 16300 16064
rect 16340 16024 16780 16064
rect 16820 16024 16829 16064
rect 20297 16024 20332 16064
rect 20372 16024 20428 16064
rect 20468 16024 21388 16064
rect 21428 16024 21437 16064
rect 22871 16024 23444 16064
rect 24250 16024 24259 16064
rect 24299 16024 24308 16064
rect 25882 16024 25891 16064
rect 25931 16024 26036 16064
rect 23404 15980 23444 16024
rect 24268 15980 24308 16024
rect 2860 15772 3724 15812
rect 3764 15772 3773 15812
rect 3916 15772 12980 15812
rect 13034 15940 15476 15980
rect 15532 15940 23308 15980
rect 23348 15940 23357 15980
rect 23404 15940 24308 15980
rect 2860 15728 2900 15772
rect 1324 15688 2900 15728
rect 2947 15688 2956 15728
rect 2996 15688 3820 15728
rect 3860 15688 3869 15728
rect 0 15644 400 15664
rect 1324 15644 1364 15688
rect 0 15604 1364 15644
rect 1411 15604 1420 15644
rect 1460 15604 3379 15644
rect 3419 15604 3428 15644
rect 0 15584 400 15604
rect 3916 15560 3956 15772
rect 13034 15728 13074 15940
rect 15532 15896 15572 15940
rect 25996 15896 26036 16024
rect 26092 15980 26132 16108
rect 26284 16064 26324 16192
rect 26620 16148 26660 16192
rect 26956 16148 26996 16192
rect 26620 16108 26996 16148
rect 26266 16024 26275 16064
rect 26315 16024 26324 16064
rect 26467 16024 26476 16064
rect 26516 16024 26860 16064
rect 26900 16024 26909 16064
rect 28099 16024 28108 16064
rect 28148 16024 28157 16064
rect 28108 15980 28148 16024
rect 26092 15940 28148 15980
rect 14179 15856 14188 15896
rect 14228 15856 15572 15896
rect 17740 15856 18740 15896
rect 18787 15856 18796 15896
rect 18836 15856 19276 15896
rect 19316 15856 19325 15896
rect 19891 15856 19900 15896
rect 20268 15856 20277 15896
rect 24748 15856 25748 15896
rect 25996 15856 26284 15896
rect 26324 15856 27340 15896
rect 27380 15856 27389 15896
rect 27665 15856 27674 15896
rect 28042 15856 28051 15896
rect 17740 15812 17780 15856
rect 18700 15812 18740 15856
rect 24748 15812 24788 15856
rect 25708 15812 25748 15856
rect 13123 15772 13132 15812
rect 13172 15772 17780 15812
rect 17836 15772 18644 15812
rect 18700 15772 19660 15812
rect 19700 15772 19709 15812
rect 23020 15772 24788 15812
rect 4579 15688 4588 15728
rect 4628 15688 4637 15728
rect 5827 15688 5836 15728
rect 5876 15688 6316 15728
rect 6356 15688 6365 15728
rect 7171 15688 7180 15728
rect 7220 15688 8428 15728
rect 8468 15688 8477 15728
rect 9161 15688 9283 15728
rect 9332 15688 9341 15728
rect 9388 15688 11116 15728
rect 11156 15688 11165 15728
rect 11561 15688 11683 15728
rect 11732 15688 11741 15728
rect 12193 15688 13074 15728
rect 13219 15688 13228 15728
rect 13268 15688 13420 15728
rect 13460 15688 13469 15728
rect 14755 15688 14764 15728
rect 14804 15688 15052 15728
rect 15092 15688 15101 15728
rect 15610 15688 15619 15728
rect 15659 15688 15668 15728
rect 16090 15688 16099 15728
rect 16139 15688 16492 15728
rect 16532 15688 16541 15728
rect 16745 15688 16771 15728
rect 16811 15688 16876 15728
rect 16916 15688 16925 15728
rect 17225 15688 17356 15728
rect 17396 15688 17405 15728
rect 4588 15644 4628 15688
rect 9388 15644 9428 15688
rect 4588 15604 6548 15644
rect 6508 15560 6548 15604
rect 7084 15604 7700 15644
rect 1673 15520 1804 15560
rect 1844 15520 1853 15560
rect 2083 15520 2092 15560
rect 2132 15520 2141 15560
rect 2371 15520 2380 15560
rect 2420 15520 2750 15560
rect 2790 15520 2799 15560
rect 3052 15551 3092 15560
rect 1219 15352 1228 15392
rect 1268 15352 1804 15392
rect 1844 15352 1853 15392
rect 0 15224 400 15244
rect 2092 15224 2132 15520
rect 3523 15520 3532 15560
rect 3584 15520 3703 15560
rect 3811 15520 3820 15560
rect 3860 15520 3956 15560
rect 4186 15557 4195 15560
rect 4156 15520 4195 15557
rect 4235 15520 4244 15560
rect 4483 15533 4492 15560
rect 3052 15476 3092 15511
rect 4156 15517 4244 15520
rect 4156 15476 4196 15517
rect 4293 15493 4302 15533
rect 4342 15520 4492 15533
rect 4532 15520 4541 15560
rect 5321 15520 5452 15560
rect 5492 15520 5501 15560
rect 5609 15520 5709 15560
rect 5780 15520 5789 15560
rect 6089 15520 6163 15560
rect 6203 15520 6220 15560
rect 6260 15520 6269 15560
rect 6403 15520 6412 15560
rect 6452 15520 6461 15560
rect 6508 15520 6531 15560
rect 6571 15520 6580 15560
rect 6640 15520 6649 15560
rect 6689 15520 6796 15560
rect 6836 15520 6845 15560
rect 4342 15493 4532 15520
rect 5836 15478 5864 15518
rect 5904 15478 5913 15518
rect 5836 15476 5876 15478
rect 3052 15436 3676 15476
rect 3716 15436 3725 15476
rect 4099 15436 4108 15476
rect 4148 15436 4196 15476
rect 5587 15436 5596 15476
rect 5636 15436 5876 15476
rect 6019 15436 6028 15476
rect 6068 15436 6199 15476
rect 6412 15392 6452 15520
rect 7084 15476 7124 15604
rect 7193 15520 7276 15560
rect 7316 15520 7324 15560
rect 7364 15520 7373 15560
rect 7459 15478 7468 15518
rect 7508 15478 7517 15518
rect 5923 15352 5932 15392
rect 5972 15352 6452 15392
rect 6604 15436 7124 15476
rect 2633 15268 2755 15308
rect 2804 15268 2813 15308
rect 6604 15224 6644 15436
rect 7468 15392 7508 15478
rect 7660 15476 7700 15604
rect 7804 15604 8908 15644
rect 8948 15604 8957 15644
rect 9004 15604 9100 15644
rect 9140 15604 9149 15644
rect 9288 15604 9428 15644
rect 9475 15604 9484 15644
rect 9524 15604 9908 15644
rect 9955 15604 9964 15644
rect 10004 15604 10100 15644
rect 11491 15604 11500 15644
rect 11540 15604 11732 15644
rect 7804 15560 7844 15604
rect 9004 15560 9044 15604
rect 9288 15560 9328 15604
rect 9676 15560 9716 15604
rect 7786 15520 7795 15560
rect 7835 15520 7844 15560
rect 8044 15520 8140 15560
rect 8180 15520 8189 15560
rect 8044 15476 8084 15520
rect 8273 15488 8282 15528
rect 8322 15488 8331 15528
rect 8803 15520 8812 15560
rect 8852 15520 8861 15560
rect 8995 15520 9004 15560
rect 9044 15520 9053 15560
rect 9100 15520 9263 15560
rect 9303 15520 9328 15560
rect 9370 15520 9379 15560
rect 9419 15520 9428 15560
rect 9514 15520 9523 15560
rect 9563 15520 9578 15560
rect 9658 15520 9667 15560
rect 9707 15520 9716 15560
rect 7651 15436 7660 15476
rect 7700 15436 7709 15476
rect 7939 15436 7948 15476
rect 7988 15436 8084 15476
rect 8291 15392 8331 15488
rect 6787 15352 6796 15392
rect 6836 15352 7180 15392
rect 7220 15352 7229 15392
rect 7276 15352 7508 15392
rect 7555 15352 7564 15392
rect 7604 15352 7735 15392
rect 8035 15352 8044 15392
rect 8084 15352 8331 15392
rect 8812 15392 8852 15520
rect 9100 15476 9140 15520
rect 9388 15476 9428 15520
rect 8899 15436 8908 15476
rect 8948 15436 9140 15476
rect 9187 15436 9196 15476
rect 9236 15436 9428 15476
rect 8812 15352 9388 15392
rect 9428 15352 9437 15392
rect 7276 15308 7316 15352
rect 7075 15268 7084 15308
rect 7124 15268 7316 15308
rect 7363 15268 7372 15308
rect 7412 15268 8236 15308
rect 8276 15268 8285 15308
rect 0 15184 1460 15224
rect 2092 15184 5452 15224
rect 5492 15184 5501 15224
rect 5731 15184 5740 15224
rect 5780 15184 6644 15224
rect 0 15164 400 15184
rect 1420 14972 1460 15184
rect 9538 15140 9578 15520
rect 9763 15509 9772 15549
rect 9812 15509 9821 15549
rect 3103 15100 3112 15140
rect 3480 15100 3489 15140
rect 3724 15100 5356 15140
rect 5396 15100 5405 15140
rect 9538 15100 9580 15140
rect 9620 15100 9629 15140
rect 3724 15056 3764 15100
rect 1699 15016 1708 15056
rect 1748 15016 3764 15056
rect 3820 15016 6124 15056
rect 6164 15016 6173 15056
rect 6220 15016 7756 15056
rect 7796 15016 7805 15056
rect 3820 14972 3860 15016
rect 1420 14932 3860 14972
rect 3977 14932 4003 14972
rect 4043 14932 4108 14972
rect 4148 14932 4157 14972
rect 4291 14932 4300 14972
rect 4340 14932 5740 14972
rect 5780 14932 5789 14972
rect 6220 14888 6260 15016
rect 9772 14972 9812 15509
rect 9868 15476 9908 15604
rect 10060 15560 10100 15604
rect 10051 15520 10060 15560
rect 10100 15520 10109 15560
rect 10243 15520 10252 15560
rect 10292 15520 10540 15560
rect 10580 15520 10589 15560
rect 10723 15520 10732 15560
rect 10772 15520 11351 15560
rect 11391 15520 11400 15560
rect 11587 15520 11596 15560
rect 11636 15520 11645 15560
rect 9868 15436 10156 15476
rect 10196 15436 10205 15476
rect 11369 15436 11491 15476
rect 11540 15436 11549 15476
rect 11596 15392 11636 15520
rect 9955 15352 9964 15392
rect 10004 15352 10051 15392
rect 10091 15352 10164 15392
rect 11203 15352 11212 15392
rect 11252 15352 11636 15392
rect 11692 15392 11732 15604
rect 12193 15560 12233 15688
rect 15628 15644 15668 15688
rect 12500 15604 12748 15644
rect 12788 15604 12797 15644
rect 13090 15604 13804 15644
rect 13844 15604 14188 15644
rect 14228 15604 14237 15644
rect 14650 15604 14659 15644
rect 14699 15604 14846 15644
rect 14886 15604 14895 15644
rect 15049 15604 15428 15644
rect 15628 15604 16292 15644
rect 16457 15635 16588 15644
rect 16457 15604 16579 15635
rect 16628 15604 16637 15644
rect 17144 15604 17153 15644
rect 17204 15604 17324 15644
rect 12500 15560 12540 15604
rect 13090 15560 13130 15604
rect 15049 15560 15089 15604
rect 15388 15560 15428 15604
rect 16252 15561 16292 15604
rect 16570 15595 16579 15604
rect 16619 15595 16628 15604
rect 16570 15594 16628 15595
rect 16252 15560 16340 15561
rect 17836 15560 17876 15772
rect 18604 15728 18644 15772
rect 18017 15688 18028 15728
rect 18068 15688 18139 15728
rect 18179 15688 18197 15728
rect 18586 15688 18595 15728
rect 18635 15688 18644 15728
rect 20899 15688 20908 15728
rect 20948 15688 21100 15728
rect 21140 15688 21149 15728
rect 23020 15644 23060 15772
rect 24748 15728 24788 15772
rect 23561 15688 23692 15728
rect 23732 15688 23741 15728
rect 24691 15688 24700 15728
rect 24740 15688 24788 15728
rect 24844 15772 25652 15812
rect 25708 15772 28684 15812
rect 28724 15772 28733 15812
rect 18211 15604 18220 15644
rect 18260 15604 18332 15644
rect 19843 15604 19852 15644
rect 19892 15604 23060 15644
rect 23788 15604 24212 15644
rect 18292 15560 18332 15604
rect 23788 15560 23828 15604
rect 24172 15560 24212 15604
rect 24844 15560 24884 15772
rect 24931 15688 24940 15728
rect 24980 15688 25228 15728
rect 25268 15688 25277 15728
rect 25036 15604 25556 15644
rect 25036 15560 25076 15604
rect 25516 15560 25556 15604
rect 25612 15560 25652 15772
rect 25987 15688 25996 15728
rect 26036 15688 26860 15728
rect 26900 15688 27235 15728
rect 27275 15688 27284 15728
rect 26249 15604 26380 15644
rect 26420 15604 27340 15644
rect 27380 15604 27389 15644
rect 28108 15604 31267 15644
rect 31307 15604 31316 15644
rect 26284 15560 26324 15604
rect 11779 15520 11788 15560
rect 11828 15520 12141 15560
rect 12181 15520 12233 15560
rect 12294 15520 12303 15560
rect 12343 15520 12540 15560
rect 12835 15520 12844 15560
rect 12884 15520 13015 15560
rect 13072 15520 13081 15560
rect 13121 15520 13130 15560
rect 13181 15520 13219 15560
rect 13259 15520 13268 15560
rect 13315 15520 13324 15560
rect 13364 15520 13373 15560
rect 13507 15520 13516 15560
rect 13567 15520 13687 15560
rect 14083 15520 14092 15560
rect 14132 15520 14327 15560
rect 14367 15520 14376 15560
rect 14563 15520 14572 15560
rect 14612 15520 15089 15560
rect 15148 15551 15188 15560
rect 12586 15478 12595 15518
rect 12635 15478 12692 15518
rect 12329 15436 12460 15476
rect 12500 15436 12509 15476
rect 12652 15392 12692 15478
rect 13228 15476 13268 15520
rect 13324 15476 13364 15520
rect 15278 15520 15287 15560
rect 15327 15520 15336 15560
rect 15388 15520 15532 15560
rect 15572 15520 15767 15560
rect 15807 15520 15816 15560
rect 15907 15520 15916 15560
rect 15956 15520 16012 15560
rect 16052 15520 16087 15560
rect 16252 15521 16291 15560
rect 16282 15520 16291 15521
rect 16331 15520 16340 15560
rect 16396 15551 16436 15560
rect 15148 15476 15188 15511
rect 15287 15476 15327 15520
rect 16661 15520 16670 15560
rect 16710 15520 16724 15560
rect 16843 15520 16852 15560
rect 16892 15520 17356 15560
rect 17396 15520 17405 15560
rect 17452 15551 17740 15560
rect 16396 15476 16436 15511
rect 12940 15467 13036 15476
rect 12940 15427 12979 15467
rect 13019 15436 13036 15467
rect 13076 15436 13159 15476
rect 13219 15436 13228 15476
rect 13268 15436 13277 15476
rect 13324 15436 13612 15476
rect 13652 15436 13661 15476
rect 14371 15436 14380 15476
rect 14420 15436 14467 15476
rect 14507 15436 15188 15476
rect 15235 15436 15244 15476
rect 15284 15436 15327 15476
rect 15418 15436 15427 15476
rect 15467 15436 15907 15476
rect 15947 15436 15956 15476
rect 16349 15436 16396 15476
rect 16436 15436 16445 15476
rect 13019 15427 13028 15436
rect 12940 15426 13028 15427
rect 12940 15392 12980 15426
rect 15916 15392 15956 15436
rect 11692 15352 12364 15392
rect 12404 15352 12413 15392
rect 12652 15352 12980 15392
rect 14659 15352 14668 15392
rect 14708 15352 15820 15392
rect 15860 15352 15869 15392
rect 15916 15352 16588 15392
rect 16628 15352 16637 15392
rect 16684 15308 16724 15520
rect 17492 15520 17740 15551
rect 17780 15520 17789 15560
rect 17836 15551 17960 15560
rect 17836 15520 17920 15551
rect 17452 15502 17492 15511
rect 18010 15520 18019 15560
rect 18068 15520 18199 15560
rect 18274 15520 18283 15560
rect 18323 15520 18332 15560
rect 18499 15520 18508 15560
rect 18548 15520 18557 15560
rect 19075 15520 19084 15560
rect 19124 15520 19651 15560
rect 19691 15520 20620 15560
rect 20660 15520 20669 15560
rect 20890 15520 20899 15560
rect 20939 15520 20948 15560
rect 21475 15520 21484 15560
rect 21524 15520 23596 15560
rect 23636 15520 23645 15560
rect 23779 15520 23788 15560
rect 23828 15520 23837 15560
rect 23982 15520 24043 15560
rect 24083 15520 24092 15560
rect 24137 15520 24172 15560
rect 24212 15520 24268 15560
rect 24308 15520 24317 15560
rect 24364 15520 24844 15560
rect 24884 15520 24893 15560
rect 24979 15520 24988 15560
rect 25028 15520 25036 15560
rect 25076 15520 25159 15560
rect 25219 15520 25228 15560
rect 25268 15520 25367 15560
rect 25407 15520 25416 15560
rect 25498 15551 25556 15560
rect 17920 15502 17960 15511
rect 18281 15436 18316 15476
rect 18356 15436 18403 15476
rect 18443 15436 18461 15476
rect 18508 15392 18548 15520
rect 20908 15476 20948 15520
rect 23982 15476 24022 15520
rect 24364 15476 24404 15520
rect 25498 15511 25507 15551
rect 25547 15511 25556 15551
rect 25603 15520 25612 15560
rect 25652 15520 25661 15560
rect 25891 15520 25900 15560
rect 25940 15520 26044 15560
rect 26084 15520 26093 15560
rect 26214 15520 26223 15560
rect 26263 15520 26324 15560
rect 26370 15520 26476 15560
rect 26541 15520 26550 15560
rect 26648 15520 26657 15560
rect 26697 15520 26860 15560
rect 26900 15520 26909 15560
rect 26956 15551 26996 15560
rect 25498 15510 25556 15511
rect 27043 15520 27052 15560
rect 27092 15520 27139 15560
rect 27179 15520 27223 15560
rect 27427 15520 27436 15560
rect 27487 15520 27607 15560
rect 26956 15476 26996 15511
rect 19651 15436 19660 15476
rect 19700 15436 20948 15476
rect 23683 15436 23692 15476
rect 23732 15436 24022 15476
rect 24154 15436 24163 15476
rect 24203 15436 24212 15476
rect 24355 15436 24364 15476
rect 24404 15436 24413 15476
rect 26371 15436 26380 15476
rect 26420 15436 26708 15476
rect 26909 15436 26956 15476
rect 26996 15436 27005 15476
rect 17164 15352 18548 15392
rect 18691 15352 18700 15392
rect 18740 15352 20428 15392
rect 20468 15352 20477 15392
rect 17164 15308 17204 15352
rect 14842 15268 14851 15308
rect 14891 15268 14956 15308
rect 14996 15268 15031 15308
rect 16675 15268 16684 15308
rect 16724 15268 16733 15308
rect 17146 15268 17155 15308
rect 17195 15268 17204 15308
rect 17513 15268 17635 15308
rect 17684 15268 17693 15308
rect 20035 15268 20044 15308
rect 20084 15268 20812 15308
rect 20852 15268 20861 15308
rect 21161 15268 21292 15308
rect 21332 15268 21341 15308
rect 19555 15184 19564 15224
rect 19604 15184 21580 15224
rect 21620 15184 21629 15224
rect 10877 15100 10886 15140
rect 11254 15100 11263 15140
rect 15811 15100 15820 15140
rect 15860 15100 16300 15140
rect 16340 15100 16349 15140
rect 18651 15100 18660 15140
rect 19028 15100 19037 15140
rect 19084 15100 22156 15140
rect 22196 15100 22205 15140
rect 19084 15056 19124 15100
rect 9964 15016 11788 15056
rect 11828 15016 11837 15056
rect 17347 15016 17356 15056
rect 17396 15016 18548 15056
rect 7075 14932 7084 14972
rect 7124 14932 7171 14972
rect 7211 14932 7255 14972
rect 7817 14932 7948 14972
rect 7988 14932 7997 14972
rect 9772 14932 9859 14972
rect 9899 14932 9908 14972
rect 9964 14888 10004 15016
rect 1219 14848 1228 14888
rect 1268 14848 1708 14888
rect 1748 14848 1757 14888
rect 3724 14848 4876 14888
rect 4916 14848 4925 14888
rect 5980 14848 6260 14888
rect 6682 14848 6691 14888
rect 6731 14879 6980 14888
rect 6731 14848 6940 14879
rect 0 14804 400 14824
rect 0 14764 2956 14804
rect 2996 14764 3005 14804
rect 0 14744 400 14764
rect 3724 14720 3764 14848
rect 5980 14804 6020 14848
rect 6940 14830 6980 14839
rect 7660 14848 8236 14888
rect 8276 14848 8285 14888
rect 9091 14848 9100 14888
rect 9140 14848 10004 14888
rect 10060 14932 10156 14972
rect 10196 14932 10205 14972
rect 4099 14764 4108 14804
rect 4148 14764 4515 14804
rect 4555 14764 4564 14804
rect 4972 14764 6020 14804
rect 6199 14764 6548 14804
rect 4972 14720 5012 14764
rect 5937 14720 5977 14764
rect 6199 14731 6239 14764
rect 1097 14680 1228 14720
rect 1268 14680 1277 14720
rect 1363 14680 1372 14720
rect 1412 14680 1804 14720
rect 1844 14680 1853 14720
rect 2249 14680 2380 14720
rect 2420 14680 2429 14720
rect 2746 14711 2804 14720
rect 2746 14671 2755 14711
rect 2795 14671 2804 14711
rect 2851 14680 2860 14720
rect 2900 14680 3052 14720
rect 3092 14680 3101 14720
rect 3523 14680 3532 14720
rect 3572 14680 3715 14720
rect 3755 14680 3764 14720
rect 3811 14680 3820 14720
rect 3860 14680 3869 14720
rect 4204 14680 4405 14720
rect 4445 14680 4454 14720
rect 4627 14680 4636 14720
rect 4676 14680 4685 14720
rect 2746 14670 2804 14671
rect 905 14596 1027 14636
rect 1076 14596 1085 14636
rect 1315 14596 1324 14636
rect 1364 14596 2563 14636
rect 2603 14596 2612 14636
rect 2764 14552 2804 14670
rect 3820 14636 3860 14680
rect 2851 14596 2860 14636
rect 2900 14596 3436 14636
rect 3476 14596 3485 14636
rect 3715 14596 3724 14636
rect 3764 14596 3860 14636
rect 1132 14512 1324 14552
rect 1364 14512 1373 14552
rect 1420 14512 1708 14552
rect 1748 14512 1757 14552
rect 1891 14512 1900 14552
rect 1940 14512 2804 14552
rect 2860 14512 2956 14552
rect 2996 14512 3005 14552
rect 0 14384 400 14404
rect 1132 14384 1172 14512
rect 1420 14468 1460 14512
rect 1219 14428 1228 14468
rect 1268 14428 1460 14468
rect 2860 14468 2900 14512
rect 2860 14428 4108 14468
rect 4148 14428 4157 14468
rect 0 14344 940 14384
rect 980 14344 989 14384
rect 1132 14344 2188 14384
rect 2228 14344 2764 14384
rect 2804 14344 2813 14384
rect 0 14324 400 14344
rect 2860 14300 2900 14428
rect 1673 14260 1804 14300
rect 1844 14260 2900 14300
rect 1804 14216 1844 14260
rect 4204 14216 4244 14680
rect 4636 14636 4676 14680
rect 4766 14661 4775 14701
rect 4815 14661 4824 14701
rect 4963 14680 4972 14720
rect 5012 14680 5021 14720
rect 5642 14680 5740 14720
rect 5804 14680 5822 14720
rect 5928 14680 5937 14720
rect 5977 14680 5986 14720
rect 6058 14680 6067 14720
rect 6107 14680 6116 14720
rect 6179 14691 6188 14731
rect 6228 14691 6239 14731
rect 6508 14720 6548 14764
rect 7379 14720 7388 14731
rect 6298 14680 6307 14720
rect 6347 14680 6356 14720
rect 6499 14680 6508 14720
rect 6548 14680 6557 14720
rect 6682 14680 6691 14720
rect 6731 14680 6796 14720
rect 6836 14680 6871 14720
rect 6953 14680 6979 14720
rect 7019 14680 7084 14720
rect 7124 14680 7133 14720
rect 7377 14691 7388 14720
rect 7428 14691 7437 14731
rect 7660 14720 7700 14848
rect 7747 14764 7756 14804
rect 7796 14764 7892 14804
rect 8131 14764 8140 14804
rect 8180 14764 8189 14804
rect 8515 14764 8524 14804
rect 8564 14764 9716 14804
rect 7852 14720 7892 14764
rect 8140 14720 8180 14764
rect 9676 14720 9716 14764
rect 10060 14720 10100 14932
rect 10217 14848 10348 14888
rect 10388 14848 10397 14888
rect 10243 14764 10252 14804
rect 10292 14764 10423 14804
rect 10588 14720 10628 15016
rect 18508 14972 18548 15016
rect 18700 15016 19124 15056
rect 19564 15016 21484 15056
rect 21524 15016 21533 15056
rect 18700 14972 18740 15016
rect 11465 14932 11500 14972
rect 11540 14932 11596 14972
rect 11636 14932 11884 14972
rect 11924 14932 11933 14972
rect 12979 14932 12988 14972
rect 13028 14932 13228 14972
rect 13268 14932 13277 14972
rect 17827 14932 17836 14972
rect 17876 14932 18019 14972
rect 18059 14932 18068 14972
rect 18490 14932 18499 14972
rect 18539 14932 18548 14972
rect 18691 14932 18700 14972
rect 18740 14932 18749 14972
rect 12844 14848 14155 14888
rect 11050 14764 11059 14804
rect 11099 14764 11444 14804
rect 11404 14720 11444 14764
rect 12844 14720 12884 14848
rect 12931 14764 12940 14804
rect 12980 14764 13268 14804
rect 13228 14720 13268 14764
rect 13406 14720 13446 14848
rect 14115 14804 14155 14848
rect 14106 14764 14115 14804
rect 14155 14764 14164 14804
rect 14656 14764 14764 14804
rect 14827 14764 14836 14804
rect 16480 14764 16492 14804
rect 16532 14764 16611 14804
rect 16651 14764 16660 14804
rect 16780 14764 17164 14804
rect 17204 14764 17268 14804
rect 17378 14764 17452 14804
rect 17492 14764 17501 14804
rect 17635 14764 17644 14804
rect 17684 14764 17693 14804
rect 18480 14764 18604 14804
rect 18644 14764 18653 14804
rect 16780 14720 16820 14764
rect 17068 14720 17108 14764
rect 17378 14720 17418 14764
rect 17644 14720 17684 14764
rect 18480 14720 18520 14764
rect 19564 14720 19604 15016
rect 24172 14972 24212 15436
rect 26153 15352 26284 15392
rect 26324 15352 26333 15392
rect 26668 15308 26708 15436
rect 28108 15392 28148 15604
rect 28771 15520 28780 15560
rect 28820 15520 28829 15560
rect 30761 15520 30883 15560
rect 30932 15520 30941 15560
rect 25193 15268 25324 15308
rect 25364 15268 25373 15308
rect 26650 15268 26659 15308
rect 26699 15268 26708 15308
rect 28012 15352 28148 15392
rect 26425 15100 26434 15140
rect 26802 15100 26811 15140
rect 24940 15016 25036 15056
rect 25076 15016 25085 15056
rect 24940 14972 24980 15016
rect 28012 14972 28052 15352
rect 28099 15268 28108 15308
rect 28148 15268 28157 15308
rect 24172 14932 24268 14972
rect 24308 14932 24317 14972
rect 24931 14932 24940 14972
rect 24980 14932 24989 14972
rect 26179 14932 26188 14972
rect 26228 14932 27284 14972
rect 27994 14932 28003 14972
rect 28043 14932 28052 14972
rect 27244 14888 27284 14932
rect 19747 14848 19756 14888
rect 19796 14848 20044 14888
rect 20084 14848 20093 14888
rect 21187 14848 21196 14888
rect 21236 14848 24596 14888
rect 26659 14848 26668 14888
rect 26708 14848 26717 14888
rect 27226 14848 27235 14888
rect 27275 14848 27284 14888
rect 19756 14764 20908 14804
rect 20948 14764 21100 14804
rect 21140 14764 21149 14804
rect 21353 14764 21484 14804
rect 21524 14764 21533 14804
rect 23308 14764 24237 14804
rect 19756 14720 19796 14764
rect 22060 14720 22100 14729
rect 23308 14720 23348 14764
rect 24197 14762 24237 14764
rect 24197 14753 24252 14762
rect 7377 14680 7428 14691
rect 7546 14680 7555 14720
rect 7595 14680 7604 14720
rect 7660 14680 7672 14720
rect 7712 14680 7721 14720
rect 7834 14680 7843 14720
rect 7883 14680 7892 14720
rect 7956 14680 7965 14720
rect 8005 14680 8084 14720
rect 8131 14680 8140 14720
rect 8180 14680 8227 14720
rect 8323 14680 8332 14720
rect 8372 14680 8503 14720
rect 9065 14680 9187 14720
rect 9236 14680 9245 14720
rect 9353 14680 9484 14720
rect 9524 14680 9533 14720
rect 9667 14680 9676 14720
rect 9716 14680 9725 14720
rect 9833 14680 9859 14720
rect 9899 14680 9964 14720
rect 10004 14680 10013 14720
rect 10060 14680 10108 14720
rect 10148 14680 10157 14720
rect 10313 14680 10423 14720
rect 10484 14680 10493 14720
rect 10570 14680 10579 14720
rect 10619 14680 10628 14720
rect 10723 14680 10732 14720
rect 10772 14680 11212 14720
rect 11264 14680 11273 14720
rect 11395 14680 11404 14720
rect 11444 14680 11575 14720
rect 12547 14680 12556 14720
rect 12596 14680 12844 14720
rect 12884 14680 12893 14720
rect 13001 14680 13123 14720
rect 13172 14680 13181 14720
rect 13228 14680 13241 14720
rect 13281 14680 13290 14720
rect 13398 14680 13407 14720
rect 13447 14680 13456 14720
rect 13498 14680 13507 14720
rect 13547 14680 13556 14720
rect 13675 14680 13684 14720
rect 13748 14680 13864 14720
rect 13987 14680 13996 14720
rect 14036 14680 14167 14720
rect 14224 14680 14233 14720
rect 14273 14680 14282 14720
rect 14537 14680 14668 14720
rect 14708 14680 14717 14720
rect 14896 14680 14905 14720
rect 14945 14680 15340 14720
rect 15380 14680 15389 14720
rect 15811 14680 15820 14720
rect 15860 14680 16216 14720
rect 16256 14680 16265 14720
rect 16387 14680 16396 14720
rect 16436 14680 16492 14720
rect 16532 14680 16567 14720
rect 16684 14680 16709 14720
rect 16749 14680 16820 14720
rect 16867 14680 16876 14720
rect 16916 14680 16963 14720
rect 17059 14680 17068 14720
rect 17108 14680 17117 14720
rect 17164 14680 17243 14720
rect 17283 14680 17292 14720
rect 17360 14680 17369 14720
rect 17409 14680 17418 14720
rect 17530 14711 17588 14720
rect 4291 14596 4300 14636
rect 4340 14596 4436 14636
rect 4483 14596 4492 14636
rect 4532 14596 4676 14636
rect 4396 14468 4436 14596
rect 4775 14552 4815 14661
rect 6067 14636 6107 14680
rect 6316 14636 6356 14680
rect 6508 14636 6548 14680
rect 7377 14636 7417 14680
rect 5443 14596 5452 14636
rect 5492 14596 5972 14636
rect 6067 14596 6124 14636
rect 6164 14596 6173 14636
rect 6316 14596 6412 14636
rect 6452 14596 6461 14636
rect 6508 14596 6892 14636
rect 6932 14596 7417 14636
rect 7564 14636 7604 14680
rect 8044 14636 8084 14680
rect 13516 14636 13556 14680
rect 14242 14636 14282 14680
rect 16684 14636 16724 14680
rect 16876 14636 16916 14680
rect 17164 14636 17204 14680
rect 17530 14671 17539 14711
rect 17579 14671 17588 14711
rect 17634 14680 17643 14720
rect 17683 14680 17731 14720
rect 17803 14680 17812 14720
rect 17876 14680 17992 14720
rect 18313 14680 18322 14720
rect 18362 14680 18520 14720
rect 18569 14680 18700 14720
rect 18740 14680 18749 14720
rect 18793 14680 18802 14720
rect 18842 14680 18892 14720
rect 18932 14680 18982 14720
rect 19363 14680 19372 14720
rect 19412 14680 19421 14720
rect 19505 14680 19564 14720
rect 19604 14680 19627 14720
rect 19667 14680 19676 14720
rect 19738 14680 19747 14720
rect 19787 14680 19796 14720
rect 19852 14680 20995 14720
rect 21035 14680 21044 14720
rect 21091 14680 21100 14720
rect 21140 14680 21149 14720
rect 21449 14680 21580 14720
rect 21620 14680 21629 14720
rect 22435 14680 22444 14720
rect 22484 14680 22548 14720
rect 22588 14680 22615 14720
rect 22915 14680 22924 14720
rect 22964 14680 23308 14720
rect 23348 14680 23357 14720
rect 23849 14680 23980 14720
rect 24020 14680 24029 14720
rect 24093 14680 24102 14720
rect 24142 14680 24151 14720
rect 24197 14713 24212 14753
rect 24556 14720 24596 14848
rect 26668 14804 26708 14848
rect 24643 14764 24652 14804
rect 24692 14764 24823 14804
rect 25193 14764 25228 14804
rect 25268 14764 25324 14804
rect 25364 14764 25373 14804
rect 25546 14795 26708 14804
rect 25546 14755 25555 14795
rect 25595 14764 26708 14795
rect 26851 14764 26860 14804
rect 26900 14764 26909 14804
rect 26956 14764 27148 14804
rect 27188 14764 27197 14804
rect 25595 14755 25604 14764
rect 25546 14754 25604 14755
rect 26860 14720 26900 14764
rect 26956 14720 26996 14764
rect 28108 14720 28148 15268
rect 28780 14972 28820 15520
rect 30403 15436 30412 15476
rect 30452 15436 30461 15476
rect 28867 15268 28876 15308
rect 28916 15268 28972 15308
rect 29012 15268 29047 15308
rect 29225 15268 29356 15308
rect 29396 15268 29405 15308
rect 28378 14932 28387 14972
rect 28427 14932 28820 14972
rect 28876 14932 30836 14972
rect 28876 14888 28916 14932
rect 28579 14848 28588 14888
rect 28628 14848 28916 14888
rect 30691 14848 30700 14888
rect 30740 14848 30749 14888
rect 30700 14804 30740 14848
rect 28393 14764 28402 14804
rect 28442 14764 30740 14804
rect 30796 14720 30836 14932
rect 30953 14848 31084 14888
rect 31124 14848 31133 14888
rect 24252 14713 24500 14720
rect 24197 14680 24500 14713
rect 24547 14680 24556 14720
rect 24596 14680 24605 14720
rect 24655 14680 24748 14720
rect 24817 14680 24835 14720
rect 24886 14680 24895 14720
rect 24935 14680 24940 14720
rect 24980 14680 25075 14720
rect 25289 14680 25420 14720
rect 25460 14680 25469 14720
rect 25642 14680 25651 14720
rect 25691 14680 25700 14720
rect 26580 14680 26668 14720
rect 26708 14680 26711 14720
rect 26751 14680 26760 14720
rect 26813 14711 26900 14720
rect 26813 14680 26851 14711
rect 17530 14670 17588 14671
rect 7564 14596 7660 14636
rect 7700 14596 7709 14636
rect 8044 14596 8236 14636
rect 8276 14596 8285 14636
rect 8873 14596 9004 14636
rect 9044 14596 9053 14636
rect 9100 14596 12980 14636
rect 13516 14596 14132 14636
rect 14179 14596 14188 14636
rect 14228 14596 14282 14636
rect 14476 14596 15916 14636
rect 15956 14596 15965 14636
rect 16099 14596 16108 14636
rect 16148 14596 16724 14636
rect 16867 14596 16876 14636
rect 16916 14596 16925 14636
rect 16972 14596 17204 14636
rect 17548 14636 17588 14670
rect 19372 14636 19412 14680
rect 19852 14636 19892 14680
rect 21100 14636 21140 14680
rect 17548 14596 17644 14636
rect 17684 14596 17693 14636
rect 18008 14596 18017 14636
rect 18057 14596 18494 14636
rect 18534 14596 19084 14636
rect 19124 14596 19133 14636
rect 19372 14596 19660 14636
rect 19700 14596 19892 14636
rect 20419 14596 20428 14636
rect 20468 14596 21140 14636
rect 22060 14636 22100 14680
rect 24099 14636 24139 14680
rect 24460 14636 24500 14680
rect 25651 14636 25691 14680
rect 26842 14671 26851 14680
rect 26891 14671 26900 14711
rect 26947 14680 26956 14720
rect 26996 14680 27005 14720
rect 27113 14680 27244 14720
rect 27284 14680 27293 14720
rect 27427 14680 27436 14720
rect 27476 14680 27532 14720
rect 27572 14680 27607 14720
rect 27689 14680 27820 14720
rect 27860 14680 27869 14720
rect 27994 14680 28003 14720
rect 28043 14680 28148 14720
rect 28361 14680 28492 14720
rect 28532 14680 28541 14720
rect 28841 14680 28972 14720
rect 29012 14680 29021 14720
rect 30377 14680 30508 14720
rect 30548 14680 30557 14720
rect 30691 14680 30700 14720
rect 30740 14680 30836 14720
rect 30883 14680 30892 14720
rect 30932 14680 30941 14720
rect 26842 14670 26900 14671
rect 30892 14636 30932 14680
rect 22060 14596 24020 14636
rect 24099 14596 24268 14636
rect 24308 14596 24317 14636
rect 24460 14596 26764 14636
rect 26804 14596 26813 14636
rect 27052 14596 29356 14636
rect 29396 14596 29405 14636
rect 29635 14596 29644 14636
rect 29684 14596 30932 14636
rect 5932 14552 5972 14596
rect 9100 14552 9140 14596
rect 4775 14512 5204 14552
rect 5705 14512 5827 14552
rect 5876 14512 5885 14552
rect 5932 14512 9140 14552
rect 4396 14428 4820 14468
rect 4780 14384 4820 14428
rect 5164 14384 5204 14512
rect 12940 14468 12980 14596
rect 14092 14552 14132 14596
rect 14476 14552 14516 14596
rect 16972 14552 17012 14596
rect 23980 14552 24020 14596
rect 27052 14552 27092 14596
rect 13385 14512 13507 14552
rect 13556 14512 13565 14552
rect 13769 14512 13804 14552
rect 13844 14512 13900 14552
rect 13940 14512 13949 14552
rect 14092 14512 14516 14552
rect 14563 14512 14572 14552
rect 14612 14512 14621 14552
rect 15900 14512 16012 14552
rect 16091 14512 16100 14552
rect 16387 14512 16396 14552
rect 16436 14512 16588 14552
rect 16628 14512 16637 14552
rect 16963 14512 16972 14552
rect 17012 14512 17021 14552
rect 17609 14512 17731 14552
rect 17780 14512 17789 14552
rect 17923 14512 17932 14552
rect 17972 14512 18220 14552
rect 18260 14512 18269 14552
rect 18595 14512 18604 14552
rect 18644 14512 22732 14552
rect 22772 14512 22781 14552
rect 23299 14512 23308 14552
rect 23348 14512 23452 14552
rect 23492 14512 23501 14552
rect 23980 14512 27092 14552
rect 29827 14512 29836 14552
rect 29876 14512 29885 14552
rect 14572 14468 14612 14512
rect 5923 14428 5932 14468
rect 5972 14428 11692 14468
rect 11732 14428 11741 14468
rect 11980 14428 12596 14468
rect 12940 14428 14612 14468
rect 16060 14468 16100 14512
rect 16060 14428 24364 14468
rect 24404 14428 24413 14468
rect 11980 14384 12020 14428
rect 12556 14384 12596 14428
rect 4343 14344 4352 14384
rect 4720 14344 4729 14384
rect 4780 14344 5068 14384
rect 5108 14344 5117 14384
rect 5164 14344 6892 14384
rect 6932 14344 6941 14384
rect 7555 14344 7564 14384
rect 7604 14344 12020 14384
rect 12117 14344 12126 14384
rect 12494 14344 12503 14384
rect 12556 14344 19660 14384
rect 19700 14344 19709 14384
rect 19891 14344 19900 14384
rect 20268 14344 20277 14384
rect 27665 14344 27674 14384
rect 28042 14344 28051 14384
rect 29836 14300 29876 14512
rect 4876 14260 7468 14300
rect 7508 14260 7517 14300
rect 10339 14260 10348 14300
rect 10388 14260 10540 14300
rect 10580 14260 10589 14300
rect 11068 14260 14092 14300
rect 14132 14260 14141 14300
rect 14563 14260 14572 14300
rect 14612 14260 15244 14300
rect 15284 14260 15293 14300
rect 18211 14260 18220 14300
rect 18260 14260 22292 14300
rect 4876 14216 4916 14260
rect 652 14176 1612 14216
rect 1652 14176 1661 14216
rect 1786 14176 1795 14216
rect 1835 14176 1844 14216
rect 1891 14176 1900 14216
rect 1940 14176 2380 14216
rect 2420 14176 2429 14216
rect 3706 14176 3715 14216
rect 3755 14176 4244 14216
rect 4867 14176 4876 14216
rect 4916 14176 4925 14216
rect 4972 14176 5452 14216
rect 5492 14176 5501 14216
rect 5626 14176 5635 14216
rect 5684 14176 5815 14216
rect 6178 14176 7276 14216
rect 7316 14176 9428 14216
rect 9955 14176 9964 14216
rect 10004 14176 10444 14216
rect 10484 14176 10493 14216
rect 10627 14176 10636 14216
rect 10676 14176 10807 14216
rect 0 13964 400 13984
rect 652 13964 692 14176
rect 4972 14132 5012 14176
rect 0 13924 692 13964
rect 748 14092 1123 14132
rect 1163 14092 1172 14132
rect 2001 14092 2010 14132
rect 2050 14092 2659 14132
rect 2699 14092 2708 14132
rect 2755 14092 2764 14132
rect 2804 14092 5012 14132
rect 5068 14092 5836 14132
rect 5876 14092 5885 14132
rect 0 13904 400 13924
rect 0 13544 400 13564
rect 0 13504 652 13544
rect 692 13504 701 13544
rect 0 13484 400 13504
rect 748 13292 788 14092
rect 5068 14048 5108 14092
rect 5548 14048 5588 14092
rect 6178 14048 6218 14176
rect 9388 14132 9428 14176
rect 11068 14132 11108 14260
rect 22252 14216 22292 14260
rect 24652 14260 27148 14300
rect 27188 14260 27197 14300
rect 28204 14260 29876 14300
rect 24652 14216 24692 14260
rect 14179 14176 14188 14216
rect 14228 14176 14237 14216
rect 14633 14176 14755 14216
rect 14804 14176 14813 14216
rect 15209 14176 15340 14216
rect 15380 14176 15389 14216
rect 16195 14176 16204 14216
rect 16244 14176 16483 14216
rect 16523 14176 16532 14216
rect 18883 14176 18892 14216
rect 18932 14176 19372 14216
rect 19412 14176 19421 14216
rect 20044 14176 20428 14216
rect 20468 14176 20477 14216
rect 21283 14176 21292 14216
rect 21332 14176 21812 14216
rect 22234 14176 22243 14216
rect 22283 14176 22292 14216
rect 23788 14176 24692 14216
rect 24809 14176 24940 14216
rect 24980 14176 24989 14216
rect 25219 14176 25228 14216
rect 25268 14176 25612 14216
rect 25652 14176 25661 14216
rect 25961 14176 26092 14216
rect 26132 14176 26141 14216
rect 26921 14176 26956 14216
rect 26996 14176 27052 14216
rect 27092 14176 27101 14216
rect 27235 14176 27244 14216
rect 27284 14176 27415 14216
rect 14188 14132 14228 14176
rect 6316 14092 9004 14132
rect 9044 14092 9053 14132
rect 9379 14092 9388 14132
rect 9428 14092 10196 14132
rect 10531 14092 10540 14132
rect 10580 14092 11108 14132
rect 11203 14092 11212 14132
rect 11252 14092 11732 14132
rect 14188 14092 14860 14132
rect 14900 14092 14909 14132
rect 15139 14092 15148 14132
rect 15188 14092 15447 14132
rect 15487 14092 15496 14132
rect 16762 14123 17644 14132
rect 6316 14048 6356 14092
rect 10156 14048 10196 14092
rect 11068 14048 11108 14092
rect 1027 14008 1036 14048
rect 1076 14008 1085 14048
rect 1132 14008 1208 14048
rect 1248 14008 1257 14048
rect 1315 14008 1324 14048
rect 1364 14008 1495 14048
rect 1690 14008 1699 14048
rect 1748 14008 1879 14048
rect 2179 14008 2188 14048
rect 2228 14008 2323 14048
rect 2363 14008 2372 14048
rect 2509 14008 2518 14048
rect 2558 14008 3292 14048
rect 3332 14008 3341 14048
rect 3521 14008 3530 14048
rect 3570 14008 3619 14048
rect 3715 14008 3724 14048
rect 3764 14008 3895 14048
rect 4963 14008 4972 14048
rect 5012 14008 5021 14048
rect 5068 14008 5091 14048
rect 5131 14008 5140 14048
rect 5200 14008 5209 14048
rect 5249 14008 5492 14048
rect 5539 14008 5548 14048
rect 5588 14008 5597 14048
rect 5801 14008 5932 14048
rect 5972 14008 5981 14048
rect 6160 14008 6169 14048
rect 6209 14008 6218 14048
rect 6307 14008 6316 14048
rect 6356 14008 6403 14048
rect 6499 14008 6508 14048
rect 6548 14008 6557 14048
rect 7747 14008 7756 14048
rect 7796 14008 10060 14048
rect 10100 14008 10109 14048
rect 10156 14008 10297 14048
rect 10337 14008 10348 14048
rect 10388 14008 10397 14048
rect 10601 14008 10732 14048
rect 10772 14008 10781 14048
rect 10960 14008 10969 14048
rect 11009 14008 11108 14048
rect 11194 14008 11203 14048
rect 11243 14008 11308 14048
rect 11348 14008 11383 14048
rect 835 13840 844 13880
rect 884 13840 893 13880
rect 163 13252 172 13292
rect 212 13252 500 13292
rect 643 13252 652 13292
rect 692 13252 788 13292
rect 844 13272 884 13840
rect 1036 13796 1076 14008
rect 1132 13964 1172 14008
rect 1132 13924 1228 13964
rect 1268 13924 1277 13964
rect 1036 13756 1612 13796
rect 1652 13756 2764 13796
rect 2804 13756 2813 13796
rect 2956 13460 2996 14008
rect 3532 13964 3572 14008
rect 3523 13924 3532 13964
rect 3572 13924 3581 13964
rect 3103 13588 3112 13628
rect 3480 13588 3489 13628
rect 2947 13420 2956 13460
rect 2996 13420 3005 13460
rect 3689 13420 3724 13460
rect 3764 13420 3820 13460
rect 3860 13420 3869 13460
rect 4972 13292 5012 14008
rect 5452 13964 5492 14008
rect 6316 13964 6356 14008
rect 6508 13964 6548 14008
rect 11692 13964 11732 14092
rect 16762 14083 16771 14123
rect 16811 14092 17644 14123
rect 17684 14092 17693 14132
rect 18892 14092 19316 14132
rect 16811 14083 16820 14092
rect 16762 14082 16820 14083
rect 18892 14048 18932 14092
rect 19276 14048 19316 14092
rect 20044 14048 20084 14176
rect 20131 14092 20140 14132
rect 20180 14092 21044 14132
rect 21449 14092 21484 14132
rect 21524 14092 21580 14132
rect 21620 14092 21629 14132
rect 21004 14048 21044 14092
rect 21772 14048 21812 14176
rect 23788 14132 23828 14176
rect 22243 14092 22252 14132
rect 22292 14092 23692 14132
rect 23732 14092 23828 14132
rect 23875 14092 23884 14132
rect 23924 14092 23933 14132
rect 23884 14048 23924 14092
rect 23980 14048 24020 14176
rect 24652 14132 24692 14176
rect 24163 14092 24172 14132
rect 24212 14092 24237 14132
rect 24425 14092 24460 14132
rect 24500 14092 24556 14132
rect 24596 14092 24605 14132
rect 24652 14092 24663 14132
rect 24703 14092 25268 14132
rect 24197 14048 24237 14092
rect 25228 14048 25268 14092
rect 12451 14008 12460 14048
rect 12500 14008 12652 14048
rect 12692 14008 12701 14048
rect 12835 14008 12844 14048
rect 12884 14008 12893 14048
rect 14100 14008 14188 14048
rect 14228 14008 14231 14048
rect 14271 14008 14280 14048
rect 14362 14039 14420 14048
rect 12844 13964 12884 14008
rect 14362 13999 14371 14039
rect 14411 13999 14420 14039
rect 14467 14008 14476 14048
rect 14516 14008 14525 14048
rect 14648 14008 14657 14048
rect 14708 14008 14828 14048
rect 14956 14039 14996 14048
rect 14362 13998 14420 13999
rect 5443 13924 5452 13964
rect 5492 13924 5501 13964
rect 5827 13924 5836 13964
rect 5876 13924 5885 13964
rect 6019 13924 6028 13964
rect 6091 13924 6199 13964
rect 6307 13924 6316 13964
rect 6356 13924 6365 13964
rect 6508 13924 6892 13964
rect 6932 13924 8332 13964
rect 8372 13924 8908 13964
rect 8948 13924 8957 13964
rect 10147 13924 10156 13964
rect 10219 13924 10327 13964
rect 10540 13924 10851 13964
rect 10891 13924 10900 13964
rect 11683 13924 11692 13964
rect 11732 13924 11741 13964
rect 12643 13924 12652 13964
rect 12692 13924 12884 13964
rect 12931 13924 12940 13964
rect 12980 13924 13111 13964
rect 5155 13756 5164 13796
rect 5204 13756 5356 13796
rect 5396 13756 5405 13796
rect 5836 13628 5876 13924
rect 10540 13880 10580 13924
rect 6281 13840 6316 13880
rect 6356 13840 6412 13880
rect 6452 13840 6461 13880
rect 7843 13840 7852 13880
rect 7892 13840 8140 13880
rect 8180 13840 9964 13880
rect 10004 13840 10580 13880
rect 11166 13840 11175 13880
rect 11215 13840 11404 13880
rect 11444 13840 11453 13880
rect 10540 13796 10580 13840
rect 14380 13796 14420 13998
rect 14476 13880 14516 14008
rect 15130 14008 15139 14048
rect 15179 14008 15188 14048
rect 15235 14008 15244 14048
rect 15284 14008 15415 14048
rect 16474 14008 16483 14048
rect 16523 14008 16532 14048
rect 14956 13964 14996 13999
rect 15148 13964 15188 14008
rect 16492 13964 16532 14008
rect 14956 13924 15052 13964
rect 15092 13924 15101 13964
rect 15148 13924 15340 13964
rect 15380 13924 15389 13964
rect 16300 13924 16532 13964
rect 16588 14039 16628 14048
rect 16858 14008 16867 14048
rect 16907 14008 16916 14048
rect 17035 14008 17044 14048
rect 17084 14008 17740 14048
rect 17780 14008 17789 14048
rect 18787 14008 18796 14048
rect 18836 14008 18892 14048
rect 18932 14008 18967 14048
rect 19075 14008 19084 14048
rect 19124 14008 19133 14048
rect 19267 14008 19276 14048
rect 19316 14008 19325 14048
rect 19459 14008 19468 14048
rect 19508 14008 20084 14048
rect 20227 14008 20236 14048
rect 20289 14008 20407 14048
rect 20515 14008 20524 14048
rect 20564 14008 20573 14048
rect 20681 14008 20812 14048
rect 20852 14008 20861 14048
rect 20986 14008 20995 14048
rect 21035 14008 21148 14048
rect 21188 14008 21204 14048
rect 21475 14008 21484 14048
rect 21524 14008 21593 14048
rect 21633 14008 21655 14048
rect 21772 14008 21868 14048
rect 21908 14008 21917 14048
rect 22435 14008 22444 14048
rect 22484 14008 22531 14048
rect 22571 14008 22615 14048
rect 23177 14008 23277 14048
rect 23348 14008 23357 14048
rect 23722 14008 23731 14048
rect 23771 14008 23924 14048
rect 23971 14008 23980 14048
rect 24020 14008 24029 14048
rect 24188 14008 24197 14048
rect 24237 14008 24259 14048
rect 24346 14008 24355 14048
rect 24395 14008 24404 14048
rect 24451 14008 24460 14048
rect 24500 14008 24652 14048
rect 24692 14008 24701 14048
rect 24809 14008 24940 14048
rect 24980 14008 24989 14048
rect 25125 14008 25137 14048
rect 25177 14008 25186 14048
rect 25228 14008 25276 14048
rect 25316 14008 25325 14048
rect 25507 14024 25516 14048
rect 15148 13880 15188 13924
rect 16300 13880 16340 13924
rect 16588 13880 16628 13999
rect 16876 13964 16916 14008
rect 16771 13924 16780 13964
rect 16820 13924 17548 13964
rect 17588 13924 17597 13964
rect 19084 13880 19124 14008
rect 20524 13964 20564 14008
rect 23404 13966 23432 14006
rect 23472 13966 23481 14006
rect 20524 13924 20620 13964
rect 20660 13924 20669 13964
rect 21004 13924 22147 13964
rect 22187 13924 22196 13964
rect 22714 13924 22723 13964
rect 22763 13924 22772 13964
rect 21004 13880 21044 13924
rect 14476 13840 15188 13880
rect 16291 13840 16300 13880
rect 16340 13840 16349 13880
rect 16540 13840 16628 13880
rect 17923 13840 17932 13880
rect 17972 13840 19028 13880
rect 19084 13840 20852 13880
rect 20986 13840 20995 13880
rect 21035 13840 21044 13880
rect 16540 13796 16580 13840
rect 18988 13796 19028 13840
rect 20812 13796 20852 13840
rect 10540 13756 11395 13796
rect 11435 13756 11596 13796
rect 11636 13756 11645 13796
rect 11923 13756 11932 13796
rect 11972 13756 13804 13796
rect 13844 13756 13853 13796
rect 14380 13756 14572 13796
rect 14612 13756 14621 13796
rect 14755 13756 14764 13796
rect 14804 13756 17164 13796
rect 17204 13756 17213 13796
rect 18883 13756 18892 13796
rect 18932 13756 18941 13796
rect 18988 13756 19852 13796
rect 19892 13756 19901 13796
rect 20812 13756 21484 13796
rect 21524 13756 21533 13796
rect 18892 13712 18932 13756
rect 8995 13672 9004 13712
rect 9044 13672 12748 13712
rect 12788 13672 16876 13712
rect 16916 13672 16925 13712
rect 18892 13672 19124 13712
rect 5452 13588 5876 13628
rect 6115 13588 6124 13628
rect 6164 13588 6173 13628
rect 10877 13588 10886 13628
rect 11254 13588 11263 13628
rect 18651 13588 18660 13628
rect 19028 13588 19037 13628
rect 5452 13292 5492 13588
rect 6124 13460 6164 13588
rect 7939 13504 7948 13544
rect 7988 13504 9196 13544
rect 9236 13504 9524 13544
rect 9667 13504 9676 13544
rect 9716 13504 12460 13544
rect 12500 13504 15724 13544
rect 15764 13504 15773 13544
rect 17068 13504 17260 13544
rect 17300 13504 17309 13544
rect 9484 13460 9524 13504
rect 5731 13420 5740 13460
rect 5780 13420 5904 13460
rect 5539 13336 5548 13376
rect 5588 13336 5719 13376
rect 5864 13292 5904 13420
rect 6028 13420 6604 13460
rect 6644 13420 6653 13460
rect 7459 13420 7468 13460
rect 7508 13420 9332 13460
rect 6028 13292 6068 13420
rect 9292 13376 9332 13420
rect 6115 13336 6124 13376
rect 6164 13336 6295 13376
rect 6665 13336 6700 13376
rect 6740 13336 6796 13376
rect 6836 13336 6845 13376
rect 7843 13336 7852 13376
rect 7892 13336 8276 13376
rect 8803 13336 8812 13376
rect 8852 13336 8908 13376
rect 8948 13336 8983 13376
rect 9274 13336 9283 13376
rect 9323 13336 9332 13376
rect 9484 13420 10636 13460
rect 10676 13420 11308 13460
rect 11348 13420 11357 13460
rect 8236 13292 8276 13336
rect 2563 13252 2572 13292
rect 2612 13252 2621 13292
rect 4649 13252 4771 13292
rect 4820 13252 4829 13292
rect 4963 13252 4972 13292
rect 5012 13252 5021 13292
rect 5452 13252 5588 13292
rect 5635 13252 5644 13292
rect 5684 13252 5815 13292
rect 5864 13252 5924 13292
rect 6019 13252 6028 13292
rect 6068 13252 6077 13292
rect 6403 13252 6412 13292
rect 6452 13252 6596 13292
rect 6761 13252 6892 13292
rect 6932 13252 6941 13292
rect 7555 13252 7564 13292
rect 7604 13252 7712 13292
rect 0 13124 400 13144
rect 460 13124 500 13252
rect 1018 13168 1027 13208
rect 1067 13168 1420 13208
rect 1460 13168 1469 13208
rect 0 13084 500 13124
rect 0 13064 400 13084
rect 2572 13040 2612 13252
rect 5548 13208 5588 13252
rect 5884 13208 5924 13252
rect 6556 13208 6596 13252
rect 7672 13208 7712 13252
rect 7804 13252 7948 13292
rect 7988 13252 7997 13292
rect 8218 13252 8227 13292
rect 8267 13252 8276 13292
rect 8515 13252 8524 13292
rect 8564 13252 8716 13292
rect 8756 13252 8765 13292
rect 7804 13219 7844 13252
rect 3331 13168 3340 13208
rect 3380 13168 3619 13208
rect 3659 13168 3668 13208
rect 3715 13168 3724 13208
rect 3764 13168 3895 13208
rect 4642 13168 4651 13208
rect 4691 13168 4700 13208
rect 4867 13168 4876 13208
rect 4916 13168 5047 13208
rect 5478 13168 5487 13208
rect 5527 13168 5588 13208
rect 5770 13168 5779 13208
rect 5819 13168 5828 13208
rect 5875 13168 5884 13208
rect 5924 13168 5933 13208
rect 6054 13168 6124 13208
rect 6164 13168 6185 13208
rect 6225 13168 6234 13208
rect 6547 13168 6556 13208
rect 6596 13168 6605 13208
rect 6691 13168 6700 13208
rect 6761 13168 6871 13208
rect 6953 13168 7027 13208
rect 7067 13168 7084 13208
rect 7124 13168 7133 13208
rect 7337 13168 7439 13208
rect 7508 13168 7517 13208
rect 7560 13168 7569 13208
rect 7609 13168 7618 13208
rect 7663 13168 7672 13208
rect 7712 13168 7721 13208
rect 7784 13179 7793 13219
rect 7833 13179 7844 13219
rect 9484 13208 9524 13420
rect 10156 13336 10828 13376
rect 10868 13336 10877 13376
rect 10156 13208 10196 13336
rect 10339 13252 10348 13292
rect 10411 13252 10519 13292
rect 10627 13252 10636 13292
rect 10676 13252 10732 13292
rect 10772 13252 10807 13292
rect 11308 13208 11348 13420
rect 12077 13292 12117 13504
rect 17068 13460 17108 13504
rect 14371 13420 14380 13460
rect 14420 13420 14476 13460
rect 14516 13420 14551 13460
rect 15031 13420 15532 13460
rect 15572 13420 15581 13460
rect 16291 13420 16300 13460
rect 16340 13420 16483 13460
rect 16523 13420 16532 13460
rect 17050 13420 17059 13460
rect 17099 13420 17108 13460
rect 17346 13420 17452 13460
rect 17492 13420 17960 13460
rect 12556 13336 13132 13376
rect 13172 13336 13181 13376
rect 13315 13336 13324 13376
rect 13364 13336 13703 13376
rect 13743 13336 13752 13376
rect 13795 13336 13804 13376
rect 13844 13336 13853 13376
rect 14755 13336 14764 13376
rect 14804 13336 14880 13376
rect 11395 13252 11404 13292
rect 11444 13252 11636 13292
rect 12077 13252 12115 13292
rect 12155 13252 12164 13292
rect 11596 13208 11636 13252
rect 12556 13208 12596 13336
rect 13804 13292 13844 13336
rect 14764 13292 14804 13336
rect 12666 13252 12675 13292
rect 12715 13252 12748 13292
rect 12788 13252 12846 13292
rect 12931 13252 12940 13292
rect 12980 13252 13036 13292
rect 13076 13252 13111 13292
rect 13203 13252 13604 13292
rect 13797 13252 13806 13292
rect 13846 13252 14860 13292
rect 14900 13252 14909 13292
rect 13203 13208 13243 13252
rect 13564 13250 13604 13252
rect 13564 13210 13612 13250
rect 13652 13210 13661 13250
rect 15031 13208 15071 13420
rect 17506 13376 17546 13420
rect 15235 13336 15244 13376
rect 15284 13336 15532 13376
rect 15572 13336 15581 13376
rect 15628 13336 17546 13376
rect 17602 13336 17740 13376
rect 17780 13336 17789 13376
rect 15628 13292 15668 13336
rect 15497 13252 15628 13292
rect 15668 13252 15677 13292
rect 16876 13252 16972 13292
rect 17012 13252 17021 13292
rect 17155 13252 17164 13292
rect 17204 13252 17213 13292
rect 17347 13252 17356 13292
rect 17396 13252 17492 13292
rect 16876 13208 16916 13252
rect 17164 13208 17204 13252
rect 17452 13208 17492 13252
rect 17602 13208 17642 13336
rect 17920 13292 17960 13420
rect 17920 13252 17972 13292
rect 17932 13208 17972 13252
rect 18094 13252 18220 13292
rect 18260 13252 18269 13292
rect 18094 13208 18134 13252
rect 18988 13208 19028 13217
rect 19084 13208 19124 13672
rect 20812 13504 22636 13544
rect 22676 13504 22685 13544
rect 20131 13420 20140 13460
rect 20180 13420 20716 13460
rect 20756 13420 20765 13460
rect 20812 13376 20852 13504
rect 22732 13460 22772 13924
rect 23404 13544 23444 13966
rect 24364 13964 24404 14008
rect 23587 13924 23596 13964
rect 23636 13924 23980 13964
rect 24020 13924 24029 13964
rect 24090 13924 24099 13964
rect 24139 13924 24148 13964
rect 24259 13924 24268 13964
rect 24308 13924 24404 13964
rect 24099 13880 24139 13924
rect 24460 13880 24500 14008
rect 25125 13964 25165 14008
rect 25409 13984 25466 14024
rect 25506 14008 25516 14024
rect 25556 14008 25565 14048
rect 25506 13984 25556 14008
rect 25612 13964 25652 14176
rect 27244 14132 27284 14176
rect 25804 14092 26708 14132
rect 25804 14048 25844 14092
rect 26668 14048 26708 14092
rect 27016 14092 27284 14132
rect 27331 14092 27340 14132
rect 27380 14092 27572 14132
rect 27016 14048 27056 14092
rect 27532 14048 27572 14092
rect 28204 14048 28244 14260
rect 25795 14008 25804 14048
rect 25844 14008 25975 14048
rect 26134 14008 26143 14048
rect 26183 14008 26188 14048
rect 26228 14008 26323 14048
rect 26659 14008 26668 14048
rect 26708 14008 26717 14048
rect 26998 14008 27007 14048
rect 27047 14008 27052 14048
rect 27092 14008 27216 14048
rect 27316 14027 27380 14048
rect 27514 14039 27572 14048
rect 27316 13987 27405 14027
rect 27445 13987 27454 14027
rect 27514 13999 27523 14039
rect 27563 13999 27572 14039
rect 27619 14008 27628 14048
rect 27672 14008 27799 14048
rect 28195 14008 28204 14048
rect 28244 14008 28253 14048
rect 28457 14008 28588 14048
rect 28628 14008 28637 14048
rect 30595 14008 30604 14048
rect 30644 14008 30883 14048
rect 30932 14008 30941 14048
rect 27514 13998 27572 13999
rect 27316 13964 27356 13987
rect 25125 13924 25268 13964
rect 25612 13924 26026 13964
rect 26066 13924 26075 13964
rect 26851 13924 26860 13964
rect 26930 13924 27031 13964
rect 27139 13924 27148 13964
rect 27188 13924 27356 13964
rect 28963 13924 28972 13964
rect 29012 13924 29347 13964
rect 29387 13924 29396 13964
rect 31075 13924 31084 13964
rect 31124 13924 31133 13964
rect 31258 13924 31267 13964
rect 31307 13924 31316 13964
rect 23491 13840 23500 13880
rect 23540 13840 23671 13880
rect 24099 13840 24500 13880
rect 25228 13880 25268 13924
rect 25228 13840 25324 13880
rect 25364 13840 25940 13880
rect 26275 13840 26284 13880
rect 26324 13840 26668 13880
rect 26708 13840 26764 13880
rect 26804 13840 26839 13880
rect 28771 13840 28780 13880
rect 28820 13840 28828 13880
rect 28868 13840 28951 13880
rect 25900 13796 25940 13840
rect 25891 13756 25900 13796
rect 25940 13756 27340 13796
rect 27380 13756 27389 13796
rect 27619 13756 27628 13796
rect 27668 13756 28972 13796
rect 29012 13756 30508 13796
rect 30548 13756 30557 13796
rect 26425 13588 26434 13628
rect 26802 13588 26811 13628
rect 23404 13504 24500 13544
rect 24460 13460 24500 13504
rect 21955 13420 21964 13460
rect 22004 13420 22772 13460
rect 23674 13420 23683 13460
rect 23723 13420 24268 13460
rect 24308 13420 24317 13460
rect 24451 13420 24460 13460
rect 24500 13420 24509 13460
rect 25769 13420 25804 13460
rect 25844 13420 25900 13460
rect 25940 13420 25949 13460
rect 26825 13420 26956 13460
rect 26996 13420 27005 13460
rect 19529 13336 19660 13376
rect 19700 13336 19709 13376
rect 20140 13336 20852 13376
rect 25219 13336 25228 13376
rect 25268 13336 25556 13376
rect 26755 13336 26764 13376
rect 26804 13336 27244 13376
rect 27284 13336 27293 13376
rect 29801 13336 29932 13376
rect 29972 13336 29981 13376
rect 20140 13292 20180 13336
rect 7936 13168 7945 13208
rect 7985 13168 7994 13208
rect 4660 13124 4700 13168
rect 5338 13126 5347 13166
rect 5387 13126 5396 13166
rect 5356 13124 5396 13126
rect 5788 13124 5828 13168
rect 6298 13126 6307 13166
rect 6347 13126 6356 13166
rect 6316 13124 6356 13126
rect 7569 13124 7609 13168
rect 7954 13124 7994 13168
rect 8044 13168 8087 13208
rect 8127 13168 8136 13208
rect 8201 13168 8332 13208
rect 8372 13168 8381 13208
rect 9034 13168 9043 13208
rect 9083 13168 9100 13208
rect 9140 13168 9223 13208
rect 9283 13168 9292 13208
rect 9332 13168 9341 13208
rect 9475 13168 9484 13208
rect 9524 13168 9533 13208
rect 10156 13168 10252 13208
rect 10292 13168 10301 13208
rect 10444 13168 10469 13208
rect 10509 13168 10518 13208
rect 10564 13168 10588 13208
rect 10628 13168 10637 13208
rect 10877 13168 10903 13208
rect 10943 13168 10964 13208
rect 11011 13168 11020 13208
rect 11083 13168 11191 13208
rect 11299 13168 11308 13208
rect 11348 13168 11357 13208
rect 11587 13168 11596 13208
rect 11636 13168 11645 13208
rect 12268 13168 12280 13208
rect 12320 13168 12329 13208
rect 12547 13168 12556 13208
rect 12596 13168 12605 13208
rect 12748 13168 12773 13208
rect 12813 13168 12822 13208
rect 12880 13168 12892 13208
rect 12932 13168 12941 13208
rect 13062 13168 13132 13208
rect 13172 13168 13193 13208
rect 13233 13168 13243 13208
rect 13420 13168 13468 13208
rect 13508 13168 13517 13208
rect 14249 13168 14380 13208
rect 14420 13168 14429 13208
rect 14563 13168 14572 13208
rect 14612 13168 14621 13208
rect 14722 13168 14731 13208
rect 14804 13168 14911 13208
rect 15022 13168 15031 13208
rect 15071 13168 15080 13208
rect 15462 13168 15471 13208
rect 15511 13168 15532 13208
rect 15572 13168 15642 13208
rect 15715 13168 15724 13208
rect 15789 13168 15895 13208
rect 16003 13168 16012 13208
rect 16052 13168 16300 13208
rect 16340 13168 16349 13208
rect 16457 13168 16483 13208
rect 16523 13168 16588 13208
rect 16628 13168 16684 13208
rect 16724 13168 16733 13208
rect 16867 13168 16876 13208
rect 16916 13168 16925 13208
rect 17050 13168 17059 13208
rect 17099 13168 17108 13208
rect 17164 13168 17177 13208
rect 17217 13168 17251 13208
rect 17328 13168 17337 13208
rect 17377 13168 17386 13208
rect 17434 13168 17443 13208
rect 17483 13168 17492 13208
rect 17580 13168 17589 13208
rect 17629 13168 17642 13208
rect 17705 13168 17827 13208
rect 17876 13168 17885 13208
rect 17932 13168 17982 13208
rect 18022 13168 18031 13208
rect 18076 13168 18085 13208
rect 18125 13168 18134 13208
rect 18202 13168 18211 13208
rect 18251 13168 18260 13208
rect 18307 13168 18316 13208
rect 18385 13168 18487 13208
rect 19028 13168 19124 13208
rect 19180 13252 20180 13292
rect 20227 13252 20236 13292
rect 20276 13252 21236 13292
rect 21283 13252 21292 13292
rect 21332 13252 21484 13292
rect 21524 13252 22004 13292
rect 22650 13252 22659 13292
rect 22699 13252 23308 13292
rect 23348 13252 23357 13292
rect 23980 13252 24500 13292
rect 24643 13252 24652 13292
rect 24692 13252 25460 13292
rect 4660 13084 5164 13124
rect 5204 13084 5213 13124
rect 5356 13084 5548 13124
rect 5588 13084 5597 13124
rect 5788 13084 6028 13124
rect 6068 13084 6077 13124
rect 6316 13084 7609 13124
rect 7907 13084 7948 13124
rect 7988 13084 7997 13124
rect 6412 13040 6452 13084
rect 7564 13040 7604 13084
rect 2572 13000 6452 13040
rect 6499 13000 6508 13040
rect 6548 13000 7459 13040
rect 7499 13000 7508 13040
rect 7555 13000 7564 13040
rect 7604 13000 7680 13040
rect 8044 12956 8084 13168
rect 8554 13126 8563 13166
rect 8603 13126 8660 13166
rect 8871 13126 8880 13166
rect 8920 13126 8948 13166
rect 8620 13040 8660 13126
rect 8908 13040 8948 13126
rect 8410 13000 8419 13040
rect 8459 13000 8620 13040
rect 8660 13000 8669 13040
rect 8899 13000 8908 13040
rect 8948 13000 8957 13040
rect 9292 12956 9332 13168
rect 10444 13124 10484 13168
rect 10025 13084 10156 13124
rect 10196 13084 10205 13124
rect 10422 13084 10444 13124
rect 10484 13084 10493 13124
rect 10564 13040 10604 13168
rect 10924 13124 10964 13168
rect 12268 13124 12308 13168
rect 12748 13124 12788 13168
rect 10915 13084 10924 13124
rect 10964 13084 10973 13124
rect 11395 13084 11404 13124
rect 11444 13084 12404 13124
rect 12451 13084 12460 13124
rect 12500 13084 12556 13124
rect 12596 13084 12631 13124
rect 12726 13084 12748 13124
rect 12788 13084 12797 13124
rect 12364 13040 12404 13084
rect 12880 13040 12920 13168
rect 13306 13126 13315 13166
rect 13355 13126 13364 13166
rect 13324 13124 13364 13126
rect 13420 13124 13460 13168
rect 13925 13126 13939 13166
rect 13979 13126 13988 13166
rect 13925 13124 13965 13126
rect 14572 13124 14612 13168
rect 15130 13126 15139 13166
rect 15179 13126 15188 13166
rect 15322 13126 15331 13166
rect 15371 13126 15380 13166
rect 13324 13084 13420 13124
rect 13460 13084 13482 13124
rect 13900 13084 13965 13124
rect 14083 13084 14092 13124
rect 14132 13084 14612 13124
rect 13900 13040 13940 13084
rect 14938 13042 14947 13082
rect 14987 13042 14996 13082
rect 9475 13000 9484 13040
rect 9524 13000 12308 13040
rect 12364 13000 13228 13040
rect 13268 13000 13277 13040
rect 13900 13000 14764 13040
rect 14804 13000 14813 13040
rect 12268 12956 12308 13000
rect 13900 12956 13940 13000
rect 3619 12916 3628 12956
rect 3668 12916 4820 12956
rect 7363 12916 7372 12956
rect 7412 12916 8428 12956
rect 8468 12916 8477 12956
rect 9292 12916 10156 12956
rect 10196 12916 11404 12956
rect 11444 12916 11453 12956
rect 12268 12916 13940 12956
rect 4780 12872 4820 12916
rect 14956 12872 14996 13042
rect 15148 13040 15188 13126
rect 15340 13040 15380 13126
rect 17067 13124 17107 13168
rect 16771 13084 16780 13124
rect 16820 13084 17107 13124
rect 17337 13124 17377 13168
rect 17602 13124 17642 13168
rect 18220 13124 18260 13168
rect 18988 13159 19028 13168
rect 17337 13084 17452 13124
rect 17492 13084 17501 13124
rect 17548 13084 17642 13124
rect 17731 13084 17740 13124
rect 17780 13084 18260 13124
rect 18680 13084 18689 13124
rect 18729 13084 18892 13124
rect 18932 13084 18941 13124
rect 15148 13000 15244 13040
rect 15284 13000 15380 13040
rect 17548 12956 17588 13084
rect 19180 13040 19220 13252
rect 21004 13208 21044 13252
rect 19747 13168 19756 13208
rect 19796 13199 20084 13208
rect 19796 13168 20044 13199
rect 20323 13168 20332 13208
rect 20372 13168 20812 13208
rect 20852 13168 20861 13208
rect 20995 13168 21004 13208
rect 21044 13168 21053 13208
rect 21100 13199 21140 13208
rect 20044 13150 20084 13159
rect 19939 13084 19948 13124
rect 19988 13084 19997 13124
rect 17993 13000 18115 13040
rect 18164 13000 18173 13040
rect 18499 13000 18508 13040
rect 18548 13000 18787 13040
rect 18827 13000 18836 13040
rect 18883 13000 18892 13040
rect 18932 13000 19220 13040
rect 19948 13040 19988 13084
rect 21100 13040 21140 13159
rect 21196 13124 21236 13252
rect 21964 13208 22004 13252
rect 23212 13208 23252 13252
rect 23980 13208 24020 13252
rect 24460 13208 24500 13252
rect 25420 13208 25460 13252
rect 25516 13208 25556 13336
rect 26851 13252 26860 13292
rect 26900 13252 27109 13292
rect 27149 13252 27676 13292
rect 27716 13252 28108 13292
rect 28148 13252 28157 13292
rect 28387 13252 28396 13292
rect 28436 13252 29012 13292
rect 30665 13252 30700 13292
rect 30740 13252 30796 13292
rect 30836 13252 30845 13292
rect 28972 13208 29012 13252
rect 21379 13168 21388 13208
rect 21428 13168 21559 13208
rect 21955 13168 21964 13208
rect 22004 13168 22013 13208
rect 22121 13168 22252 13208
rect 22292 13168 22301 13208
rect 22409 13168 22540 13208
rect 22580 13168 22589 13208
rect 22636 13168 22757 13208
rect 22797 13168 22806 13208
rect 23194 13168 23203 13208
rect 23243 13168 23328 13208
rect 23404 13168 23678 13208
rect 23718 13168 23727 13208
rect 24163 13168 24172 13208
rect 24212 13168 24221 13208
rect 24298 13168 24307 13208
rect 24347 13168 24356 13208
rect 24412 13168 24421 13208
rect 24500 13168 24601 13208
rect 25097 13168 25228 13208
rect 25268 13168 25277 13208
rect 25402 13168 25411 13208
rect 25451 13168 25460 13208
rect 25507 13168 25516 13208
rect 25556 13168 25565 13208
rect 25699 13168 25708 13208
rect 25748 13168 25757 13208
rect 25891 13168 25900 13208
rect 25940 13168 26071 13208
rect 26921 13168 27017 13208
rect 27092 13168 27101 13208
rect 27331 13168 27340 13208
rect 27380 13168 27511 13208
rect 27562 13168 27571 13208
rect 27611 13168 27620 13208
rect 28649 13168 28780 13208
rect 28820 13168 28829 13208
rect 28963 13168 28972 13208
rect 29012 13168 29143 13208
rect 30115 13168 30124 13208
rect 30164 13168 30604 13208
rect 30644 13168 30653 13208
rect 21196 13084 22444 13124
rect 22484 13084 22493 13124
rect 22636 13040 22676 13168
rect 23404 13124 23444 13168
rect 23980 13159 24020 13168
rect 24172 13124 24212 13168
rect 24316 13124 24356 13168
rect 25708 13124 25748 13168
rect 27580 13124 27620 13168
rect 31276 13124 31316 13924
rect 23395 13084 23404 13124
rect 23444 13084 23453 13124
rect 23505 13084 23514 13124
rect 23554 13084 23692 13124
rect 23732 13084 23741 13124
rect 24134 13084 24172 13124
rect 24212 13084 24221 13124
rect 24316 13084 25315 13124
rect 25355 13084 25748 13124
rect 25795 13084 25804 13124
rect 25844 13084 27620 13124
rect 28867 13084 28876 13124
rect 28916 13084 31316 13124
rect 27580 13040 27620 13084
rect 19948 13000 20812 13040
rect 20852 13000 21140 13040
rect 21475 13000 21484 13040
rect 21524 13000 22676 13040
rect 23290 13000 23299 13040
rect 23339 13000 23348 13040
rect 23875 13000 23884 13040
rect 23924 13000 24268 13040
rect 24308 13000 24317 13040
rect 27580 13000 30556 13040
rect 30596 13000 30605 13040
rect 15427 12916 15436 12956
rect 15476 12916 17588 12956
rect 18892 12872 18932 13000
rect 23308 12956 23348 13000
rect 23308 12916 23788 12956
rect 23828 12916 23837 12956
rect 24547 12916 24556 12956
rect 24596 12916 25228 12956
rect 25268 12916 25277 12956
rect 4343 12832 4352 12872
rect 4720 12832 4729 12872
rect 4780 12832 10100 12872
rect 12117 12832 12126 12872
rect 12494 12832 12503 12872
rect 14956 12832 15340 12872
rect 15380 12832 15389 12872
rect 16963 12832 16972 12872
rect 17012 12832 17164 12872
rect 17204 12832 18932 12872
rect 19891 12832 19900 12872
rect 20268 12832 20277 12872
rect 23107 12832 23116 12872
rect 23156 12832 23165 12872
rect 23683 12832 23692 12872
rect 23732 12832 27620 12872
rect 27665 12832 27674 12872
rect 28042 12832 28051 12872
rect 10060 12788 10100 12832
rect 3715 12748 3724 12788
rect 3764 12748 5356 12788
rect 5396 12748 5684 12788
rect 0 12704 400 12724
rect 0 12664 940 12704
rect 980 12664 989 12704
rect 3209 12664 3340 12704
rect 3380 12664 3389 12704
rect 4073 12664 4204 12704
rect 4244 12664 4253 12704
rect 4492 12664 4876 12704
rect 4916 12664 4925 12704
rect 0 12644 400 12664
rect 4492 12620 4532 12664
rect 5644 12620 5684 12748
rect 7468 12748 7948 12788
rect 7988 12748 7997 12788
rect 9379 12748 9388 12788
rect 9428 12748 9437 12788
rect 10060 12748 13516 12788
rect 13556 12748 13565 12788
rect 14371 12748 14380 12788
rect 14420 12748 14996 12788
rect 16195 12748 16204 12788
rect 16244 12748 18124 12788
rect 18164 12748 18811 12788
rect 7468 12704 7508 12748
rect 5731 12664 5740 12704
rect 5780 12664 6028 12704
rect 6068 12664 6077 12704
rect 6691 12664 6700 12704
rect 6740 12664 6892 12704
rect 6932 12664 6941 12704
rect 7459 12664 7468 12704
rect 7508 12664 7517 12704
rect 7756 12664 8524 12704
rect 8564 12664 8573 12704
rect 8899 12664 8908 12704
rect 8948 12664 9004 12704
rect 9044 12664 9079 12704
rect 4483 12580 4492 12620
rect 4532 12580 4541 12620
rect 4876 12580 4972 12620
rect 5012 12580 5108 12620
rect 5644 12580 7372 12620
rect 7412 12580 7421 12620
rect 4492 12536 4532 12580
rect 4876 12536 4916 12580
rect 1193 12496 1324 12536
rect 1364 12496 1373 12536
rect 1507 12496 1516 12536
rect 1556 12496 1565 12536
rect 2275 12496 2284 12536
rect 2324 12496 2764 12536
rect 2804 12496 2860 12536
rect 2900 12496 2964 12536
rect 3139 12496 3148 12536
rect 3188 12496 3197 12536
rect 4291 12496 4300 12536
rect 4340 12496 4349 12536
rect 4492 12496 4517 12536
rect 4557 12496 4579 12536
rect 4664 12496 4673 12536
rect 4713 12496 4916 12536
rect 4972 12527 5012 12536
rect 1516 12452 1556 12496
rect 1516 12412 2668 12452
rect 2708 12412 2717 12452
rect 1769 12328 1900 12368
rect 1940 12328 1949 12368
rect 3148 12284 3188 12496
rect 4300 12368 4340 12496
rect 4972 12452 5012 12487
rect 4410 12412 4419 12452
rect 4459 12412 5012 12452
rect 5068 12452 5108 12580
rect 6051 12536 6091 12580
rect 7372 12536 7412 12580
rect 7756 12536 7796 12664
rect 8116 12580 8140 12620
rect 8180 12580 8189 12620
rect 8116 12536 8156 12580
rect 9388 12536 9428 12748
rect 14956 12704 14996 12748
rect 11273 12664 11308 12704
rect 11348 12664 11404 12704
rect 11444 12664 11453 12704
rect 13018 12664 13027 12704
rect 13076 12664 13207 12704
rect 14441 12664 14563 12704
rect 14612 12664 14621 12704
rect 14938 12664 14947 12704
rect 14987 12664 14996 12704
rect 17059 12664 17068 12704
rect 17108 12664 17836 12704
rect 17876 12664 17885 12704
rect 18403 12664 18412 12704
rect 18452 12664 18520 12704
rect 9475 12580 9484 12620
rect 9524 12580 10100 12620
rect 5705 12496 5836 12536
rect 5876 12496 5885 12536
rect 6044 12496 6053 12536
rect 6093 12496 6102 12536
rect 6892 12496 6988 12536
rect 7028 12496 7037 12536
rect 5068 12412 5644 12452
rect 5684 12412 5693 12452
rect 5962 12443 6316 12452
rect 4300 12328 4724 12368
rect 4684 12284 4724 12328
rect 1193 12244 1324 12284
rect 1364 12244 1373 12284
rect 1420 12244 3188 12284
rect 4666 12244 4675 12284
rect 4715 12244 4724 12284
rect 1420 12200 1460 12244
rect 1219 12160 1228 12200
rect 1268 12160 1460 12200
rect 2659 12160 2668 12200
rect 2708 12160 4700 12200
rect 3103 12076 3112 12116
rect 3480 12076 3489 12116
rect 1795 11908 1804 11948
rect 1844 11908 2764 11948
rect 2804 11908 3668 11948
rect 4361 11908 4483 11948
rect 4532 11908 4541 11948
rect 3235 11824 3244 11864
rect 3284 11824 3293 11864
rect 1891 11740 1900 11780
rect 1940 11740 1949 11780
rect 2729 11740 2860 11780
rect 2900 11740 2909 11780
rect 3244 11696 3284 11824
rect 3628 11780 3668 11908
rect 3628 11740 4498 11780
rect 4538 11740 4547 11780
rect 4660 11696 4700 12160
rect 4972 12116 5012 12412
rect 5962 12403 5971 12443
rect 6011 12412 6316 12443
rect 6356 12412 6365 12452
rect 6011 12403 6020 12412
rect 5962 12402 6020 12403
rect 6892 12284 6932 12496
rect 7234 12494 7316 12503
rect 7363 12496 7372 12536
rect 7412 12496 7421 12536
rect 7554 12496 7563 12536
rect 7603 12496 7700 12536
rect 7747 12496 7756 12536
rect 7796 12496 7805 12536
rect 7219 12454 7228 12494
rect 7268 12454 7316 12494
rect 6976 12412 7084 12452
rect 7147 12412 7156 12452
rect 7276 12368 7316 12454
rect 7267 12328 7276 12368
rect 7316 12328 7325 12368
rect 6892 12244 7468 12284
rect 7508 12244 7517 12284
rect 7660 12200 7700 12496
rect 7944 12491 7953 12531
rect 7993 12491 8002 12531
rect 8093 12496 8107 12536
rect 8147 12496 8156 12536
rect 8262 12496 8332 12536
rect 8372 12496 8393 12536
rect 8433 12496 8442 12536
rect 8515 12496 8524 12536
rect 8587 12496 8695 12536
rect 8969 12496 9100 12536
rect 9140 12496 9149 12536
rect 9328 12496 9337 12536
rect 9377 12496 9428 12536
rect 10060 12536 10100 12580
rect 10492 12580 12556 12620
rect 12596 12580 12605 12620
rect 12844 12580 13996 12620
rect 14036 12580 14045 12620
rect 14467 12580 14476 12620
rect 14516 12580 14525 12620
rect 14572 12580 14996 12620
rect 16867 12580 16876 12620
rect 16916 12580 17012 12620
rect 10492 12536 10532 12580
rect 10060 12496 10492 12536
rect 10532 12496 10541 12536
rect 10627 12496 10636 12536
rect 10697 12496 10807 12536
rect 10954 12496 10963 12536
rect 11003 12496 11116 12536
rect 11156 12496 11165 12536
rect 7954 12368 7994 12491
rect 10636 12452 10676 12496
rect 11248 12464 11257 12504
rect 11297 12464 11306 12504
rect 12617 12496 12715 12536
rect 12788 12496 12797 12536
rect 11266 12452 11306 12464
rect 12844 12452 12884 12580
rect 14476 12536 14516 12580
rect 14572 12536 14612 12580
rect 14956 12536 14996 12580
rect 16972 12536 17012 12580
rect 18480 12578 18520 12664
rect 18595 12580 18604 12620
rect 18644 12580 18667 12620
rect 18471 12538 18480 12578
rect 18520 12538 18529 12578
rect 18627 12536 18667 12580
rect 18771 12536 18811 12748
rect 23116 12704 23156 12832
rect 27580 12788 27620 12832
rect 24268 12748 25940 12788
rect 26371 12748 26380 12788
rect 26420 12748 27244 12788
rect 27284 12748 27293 12788
rect 27580 12748 28724 12788
rect 24268 12704 24308 12748
rect 25900 12704 25940 12748
rect 26620 12704 26660 12748
rect 19049 12664 19075 12704
rect 19115 12664 19180 12704
rect 19220 12664 19229 12704
rect 22042 12664 22051 12704
rect 22091 12664 22540 12704
rect 22580 12664 22589 12704
rect 23020 12664 23156 12704
rect 23753 12664 23836 12704
rect 23876 12664 23884 12704
rect 23924 12664 23933 12704
rect 24250 12664 24259 12704
rect 24299 12664 24308 12704
rect 24451 12664 24460 12704
rect 24500 12664 25420 12704
rect 25460 12664 25469 12704
rect 25673 12664 25708 12704
rect 25748 12664 25804 12704
rect 25844 12664 25853 12704
rect 25900 12664 26228 12704
rect 26275 12664 26284 12704
rect 26324 12664 26476 12704
rect 26516 12664 26525 12704
rect 26611 12664 26620 12704
rect 26660 12664 26669 12704
rect 26938 12664 26947 12704
rect 26996 12664 27127 12704
rect 27523 12664 27532 12704
rect 27572 12664 27724 12704
rect 27764 12664 27773 12704
rect 28457 12664 28492 12704
rect 28532 12664 28588 12704
rect 28628 12664 28637 12704
rect 23020 12620 23060 12664
rect 21187 12580 21196 12620
rect 21236 12580 21258 12620
rect 21218 12536 21258 12580
rect 21484 12580 22100 12620
rect 23011 12580 23020 12620
rect 23060 12580 23069 12620
rect 23500 12580 25420 12620
rect 25460 12580 25469 12620
rect 21484 12536 21524 12580
rect 22060 12536 22100 12580
rect 23500 12536 23540 12580
rect 26188 12536 26228 12664
rect 26334 12580 26860 12620
rect 26900 12580 26909 12620
rect 27043 12580 27052 12620
rect 27092 12580 27140 12620
rect 27235 12580 27244 12620
rect 27284 12580 27293 12620
rect 28012 12580 28108 12620
rect 28148 12580 28157 12620
rect 28335 12580 28396 12620
rect 28436 12580 28445 12620
rect 26334 12536 26374 12580
rect 27100 12536 27140 12580
rect 27244 12536 27284 12580
rect 28012 12536 28052 12580
rect 28335 12536 28375 12580
rect 12931 12496 12940 12536
rect 12980 12496 13324 12536
rect 13364 12496 13373 12536
rect 13603 12496 13612 12536
rect 13652 12496 13699 12536
rect 13739 12496 13783 12536
rect 14371 12496 14380 12536
rect 14420 12496 14516 12536
rect 14563 12496 14572 12536
rect 14612 12496 14621 12536
rect 14755 12496 14764 12536
rect 14804 12496 14813 12536
rect 14947 12496 14956 12536
rect 14996 12496 15340 12536
rect 15380 12496 15389 12536
rect 16483 12496 16492 12536
rect 16532 12496 16588 12536
rect 16628 12496 16663 12536
rect 16771 12496 16780 12536
rect 16820 12496 16829 12536
rect 16963 12496 16972 12536
rect 17012 12496 17021 12536
rect 17155 12496 17164 12536
rect 17204 12496 17335 12536
rect 18618 12496 18627 12536
rect 18667 12496 18691 12536
rect 18754 12496 18763 12536
rect 18803 12496 18812 12536
rect 18979 12496 18988 12536
rect 19028 12496 19037 12536
rect 20707 12496 20716 12536
rect 20756 12496 21100 12536
rect 21140 12496 21149 12536
rect 21200 12496 21209 12536
rect 21249 12496 21283 12536
rect 21353 12496 21484 12536
rect 21524 12496 21533 12536
rect 21859 12496 21868 12536
rect 21908 12496 21917 12536
rect 22051 12496 22060 12536
rect 22100 12496 22109 12536
rect 23107 12496 23116 12536
rect 23156 12496 23212 12536
rect 23252 12496 23287 12536
rect 23491 12496 23500 12536
rect 23540 12496 23549 12536
rect 23683 12496 23692 12536
rect 23732 12496 23863 12536
rect 23971 12496 23980 12536
rect 24020 12496 24029 12536
rect 24163 12496 24172 12536
rect 24212 12496 24221 12536
rect 24329 12496 24460 12536
rect 24500 12496 24652 12536
rect 24692 12496 24701 12536
rect 25315 12496 25324 12536
rect 25364 12496 25373 12536
rect 25507 12496 25516 12536
rect 25556 12496 25565 12536
rect 25699 12496 25708 12536
rect 25748 12496 25757 12536
rect 25891 12496 25900 12536
rect 25940 12496 25949 12536
rect 26083 12496 26092 12536
rect 26132 12496 26141 12536
rect 26188 12496 26214 12536
rect 26254 12496 26263 12536
rect 26316 12496 26325 12536
rect 26365 12496 26374 12536
rect 26431 12527 26476 12536
rect 14764 12452 14804 12496
rect 8227 12412 8236 12452
rect 8276 12412 8285 12452
rect 8611 12412 8620 12452
rect 8660 12412 9219 12452
rect 9259 12412 9268 12452
rect 9667 12412 9676 12452
rect 9716 12412 10676 12452
rect 10819 12412 10828 12452
rect 10868 12412 10999 12452
rect 11266 12412 11788 12452
rect 11828 12412 11837 12452
rect 12826 12412 12835 12452
rect 12875 12412 12884 12452
rect 12931 12412 12940 12452
rect 12980 12412 14804 12452
rect 16780 12452 16820 12496
rect 17164 12452 17204 12496
rect 18124 12454 18172 12494
rect 18212 12454 18221 12494
rect 18124 12452 18164 12454
rect 16780 12412 17204 12452
rect 17836 12412 18164 12452
rect 18307 12412 18316 12452
rect 18356 12412 18365 12452
rect 18412 12412 18883 12452
rect 18923 12412 18932 12452
rect 7939 12328 7948 12368
rect 7988 12328 7997 12368
rect 8236 12284 8276 12412
rect 8323 12328 8332 12368
rect 8372 12328 8908 12368
rect 8948 12328 8957 12368
rect 10601 12328 10732 12368
rect 10772 12328 10781 12368
rect 11266 12284 11306 12412
rect 7843 12244 7852 12284
rect 7892 12244 8140 12284
rect 8180 12244 8189 12284
rect 8236 12244 8332 12284
rect 8372 12244 8381 12284
rect 8707 12244 8716 12284
rect 8756 12244 11306 12284
rect 12844 12200 12884 12412
rect 13027 12328 13036 12368
rect 13076 12328 13744 12368
rect 13784 12328 13793 12368
rect 13507 12244 13516 12284
rect 13556 12244 13612 12284
rect 13652 12244 13687 12284
rect 16457 12244 16588 12284
rect 16628 12244 16637 12284
rect 6979 12160 6988 12200
rect 7028 12160 10348 12200
rect 10388 12160 12884 12200
rect 13507 12160 13516 12200
rect 13556 12160 15724 12200
rect 15764 12160 15773 12200
rect 4972 12076 5164 12116
rect 5204 12076 9524 12116
rect 10877 12076 10886 12116
rect 11254 12076 11263 12116
rect 13123 12076 13132 12116
rect 13172 12076 16492 12116
rect 16532 12076 16541 12116
rect 5980 11992 7372 12032
rect 7412 11992 7421 12032
rect 7555 11992 7564 12032
rect 7604 11992 7988 12032
rect 8227 11992 8236 12032
rect 8276 11992 8285 12032
rect 5692 11824 5740 11864
rect 5780 11824 5789 11864
rect 4963 11740 4972 11780
rect 5012 11740 5251 11780
rect 5291 11740 5300 11780
rect 5692 11707 5732 11824
rect 5827 11740 5836 11780
rect 5876 11740 5923 11780
rect 1289 11656 1315 11696
rect 1355 11656 1420 11696
rect 1460 11656 1469 11696
rect 3244 11656 4108 11696
rect 4148 11656 4157 11696
rect 4579 11656 4588 11696
rect 4628 11656 4700 11696
rect 4867 11656 4876 11696
rect 4916 11656 5111 11696
rect 5151 11656 5160 11696
rect 5251 11656 5260 11696
rect 5300 11656 5356 11696
rect 5396 11656 5431 11696
rect 5683 11667 5692 11707
rect 5732 11667 5741 11707
rect 5836 11696 5876 11740
rect 5980 11696 6020 11992
rect 7948 11948 7988 11992
rect 8236 11948 8276 11992
rect 9484 11948 9524 12076
rect 17836 12032 17876 12412
rect 18316 12284 18356 12412
rect 18412 12368 18452 12412
rect 18403 12328 18412 12368
rect 18452 12328 18461 12368
rect 18316 12244 18508 12284
rect 18548 12244 18557 12284
rect 18988 12200 19028 12496
rect 21868 12452 21908 12496
rect 23347 12454 23356 12494
rect 23396 12454 23444 12494
rect 21868 12412 22060 12452
rect 22100 12412 22109 12452
rect 23212 12412 23235 12452
rect 23275 12412 23284 12452
rect 20681 12328 20812 12368
rect 20852 12328 20861 12368
rect 20131 12244 20140 12284
rect 20180 12244 22636 12284
rect 22676 12244 22685 12284
rect 10627 11992 10636 12032
rect 10676 11992 12212 12032
rect 12547 11992 12556 12032
rect 12596 11992 14476 12032
rect 14516 11992 16108 12032
rect 16148 11992 16157 12032
rect 16780 11992 17876 12032
rect 6844 11908 7172 11948
rect 6844 11864 6884 11908
rect 5818 11656 5827 11696
rect 5867 11656 5876 11696
rect 5962 11656 5971 11696
rect 6011 11656 6020 11696
rect 6067 11824 6884 11864
rect 6979 11824 6988 11864
rect 7028 11824 7037 11864
rect 6067 11705 6107 11824
rect 6348 11740 6700 11780
rect 6740 11740 6749 11780
rect 6067 11696 6116 11705
rect 6348 11696 6388 11740
rect 6844 11738 6884 11824
rect 6988 11780 7028 11824
rect 7132 11780 7172 11908
rect 7372 11908 7593 11948
rect 7372 11864 7412 11908
rect 7553 11906 7593 11908
rect 7948 11908 8276 11948
rect 9466 11908 9475 11948
rect 9515 11908 10444 11948
rect 10484 11908 10493 11948
rect 7553 11866 7564 11906
rect 7604 11866 7613 11906
rect 7363 11824 7372 11864
rect 7412 11824 7421 11864
rect 6970 11740 6979 11780
rect 7019 11740 7075 11780
rect 7132 11740 7468 11780
rect 7508 11740 7517 11780
rect 7651 11740 7660 11780
rect 7700 11740 7785 11780
rect 6835 11698 6844 11738
rect 6884 11698 6893 11738
rect 6067 11656 6076 11696
rect 6202 11656 6211 11696
rect 6251 11656 6260 11696
rect 6348 11656 6407 11696
rect 6447 11656 6456 11696
rect 6589 11656 6598 11696
rect 6638 11656 6788 11696
rect 6953 11656 7084 11696
rect 7124 11656 7133 11696
rect 7267 11656 7276 11696
rect 7316 11656 7324 11696
rect 7364 11656 7447 11696
rect 7494 11656 7564 11696
rect 7604 11656 7625 11696
rect 7665 11656 7674 11696
rect 6067 11647 6116 11656
rect 6067 11612 6107 11647
rect 922 11572 931 11612
rect 971 11572 1132 11612
rect 1172 11572 1181 11612
rect 2851 11572 2860 11612
rect 2900 11572 6107 11612
rect 6220 11612 6260 11656
rect 6748 11612 6788 11656
rect 7745 11654 7785 11740
rect 7948 11696 7988 11908
rect 8094 11824 8140 11864
rect 8180 11824 8225 11864
rect 8265 11824 8274 11864
rect 10147 11824 10156 11864
rect 10196 11824 10348 11864
rect 10388 11824 10397 11864
rect 10531 11824 10540 11864
rect 10580 11824 10924 11864
rect 10964 11824 10973 11864
rect 11020 11780 11060 11992
rect 12172 11948 12212 11992
rect 11491 11908 11500 11948
rect 11540 11908 11549 11948
rect 12163 11908 12172 11948
rect 12212 11908 12652 11948
rect 12692 11908 12701 11948
rect 12905 11908 13027 11948
rect 13076 11908 13085 11948
rect 11500 11864 11540 11908
rect 11395 11824 11404 11864
rect 11444 11824 11540 11864
rect 11587 11824 11596 11864
rect 11636 11824 13132 11864
rect 13172 11824 13181 11864
rect 8035 11740 8044 11780
rect 8084 11740 8093 11780
rect 8995 11740 9004 11780
rect 9044 11740 9676 11780
rect 9716 11740 9725 11780
rect 9955 11740 9964 11780
rect 10004 11740 10532 11780
rect 10915 11740 10924 11780
rect 10964 11740 11060 11780
rect 11369 11740 11500 11780
rect 11540 11740 11549 11780
rect 12652 11740 12748 11780
rect 12788 11740 12797 11780
rect 7906 11656 7915 11696
rect 7955 11656 7988 11696
rect 7738 11614 7747 11654
rect 7787 11614 7796 11654
rect 8044 11612 8084 11740
rect 8400 11698 8587 11738
rect 8400 11696 8440 11698
rect 8362 11656 8371 11696
rect 8411 11656 8440 11696
rect 8547 11696 8587 11698
rect 9484 11696 9524 11740
rect 10492 11696 10532 11740
rect 12652 11696 12692 11740
rect 12844 11696 12884 11824
rect 13372 11780 13412 11992
rect 16780 11948 16820 11992
rect 13795 11908 13804 11948
rect 13844 11908 16204 11948
rect 16244 11908 16253 11948
rect 16483 11908 16492 11948
rect 16532 11908 16541 11948
rect 16762 11908 16771 11948
rect 16811 11908 16820 11948
rect 13865 11824 13996 11864
rect 14036 11824 14045 11864
rect 14633 11824 14764 11864
rect 14804 11824 14813 11864
rect 15206 11824 15244 11864
rect 15284 11824 15293 11864
rect 12931 11740 12940 11780
rect 12980 11740 13322 11780
rect 13372 11740 13460 11780
rect 13769 11740 13900 11780
rect 13940 11740 13949 11780
rect 14563 11740 14572 11780
rect 14612 11740 15114 11780
rect 13282 11696 13322 11740
rect 13420 11696 13460 11740
rect 15074 11696 15114 11740
rect 15206 11696 15246 11824
rect 16012 11780 16052 11908
rect 16099 11824 16108 11864
rect 16148 11824 16196 11864
rect 16265 11824 16396 11864
rect 16436 11824 16445 11864
rect 15293 11740 15340 11780
rect 15380 11740 15389 11780
rect 15715 11740 15724 11780
rect 15764 11740 15895 11780
rect 16012 11740 16100 11780
rect 15340 11696 15380 11740
rect 16060 11696 16100 11740
rect 16156 11696 16196 11824
rect 16492 11780 16532 11908
rect 17836 11864 17876 11992
rect 18508 12160 19028 12200
rect 18508 11948 18548 12160
rect 18651 12076 18660 12116
rect 19028 12076 19037 12116
rect 18298 11908 18307 11948
rect 18347 11908 18548 11948
rect 18595 11908 18604 11948
rect 18644 11908 22964 11948
rect 16579 11824 16588 11864
rect 16628 11824 16820 11864
rect 17836 11855 18116 11864
rect 17836 11824 18076 11855
rect 16476 11740 16485 11780
rect 16525 11740 16534 11780
rect 16780 11696 16820 11824
rect 21283 11824 21292 11864
rect 21332 11824 22292 11864
rect 18076 11806 18116 11815
rect 22252 11780 22292 11824
rect 16924 11740 17740 11780
rect 17780 11740 17789 11780
rect 20323 11740 20332 11780
rect 20372 11740 20620 11780
rect 20660 11740 20669 11780
rect 21955 11740 21964 11780
rect 22004 11740 22013 11780
rect 22252 11740 22388 11780
rect 22531 11740 22540 11780
rect 22580 11740 22636 11780
rect 22676 11740 22711 11780
rect 22803 11740 22828 11780
rect 22868 11740 22877 11780
rect 16924 11696 16964 11740
rect 19852 11696 19892 11705
rect 21964 11696 22004 11740
rect 22348 11738 22388 11740
rect 22348 11698 22376 11738
rect 22416 11698 22425 11738
rect 22803 11696 22843 11740
rect 22924 11696 22964 11908
rect 23212 11780 23252 12412
rect 23404 11948 23444 12454
rect 23980 12452 24020 12496
rect 23875 12412 23884 12452
rect 23924 12412 24020 12452
rect 24172 12452 24212 12496
rect 24172 12412 24556 12452
rect 24596 12412 24605 12452
rect 25324 12284 25364 12496
rect 25516 12368 25556 12496
rect 25708 12452 25748 12496
rect 25699 12412 25708 12452
rect 25748 12412 25795 12452
rect 25900 12368 25940 12496
rect 26092 12452 26132 12496
rect 26471 12496 26476 12527
rect 26516 12496 26602 12536
rect 26755 12496 26764 12536
rect 26804 12496 26935 12536
rect 27091 12496 27100 12536
rect 27140 12496 27149 12536
rect 27242 12496 27251 12536
rect 27291 12496 27331 12536
rect 27427 12496 27436 12536
rect 27476 12496 27767 12536
rect 27807 12496 27816 12536
rect 27898 12527 27956 12536
rect 26431 12478 26471 12487
rect 26764 12452 26804 12496
rect 27898 12487 27907 12527
rect 27947 12487 27956 12527
rect 28003 12496 28012 12536
rect 28052 12496 28061 12536
rect 28157 12496 28201 12536
rect 28241 12496 28250 12536
rect 28317 12496 28326 12536
rect 28366 12496 28375 12536
rect 27898 12486 27956 12487
rect 27898 12452 27938 12486
rect 28204 12452 28244 12496
rect 28435 12478 28444 12518
rect 28484 12478 28493 12518
rect 26092 12412 26188 12452
rect 26228 12412 26237 12452
rect 26764 12412 27820 12452
rect 27860 12412 27938 12452
rect 28195 12412 28204 12452
rect 28244 12412 28253 12452
rect 27898 12368 27938 12412
rect 28444 12368 28484 12478
rect 28684 12452 28724 12748
rect 30473 12496 30595 12536
rect 30644 12496 30653 12536
rect 28684 12412 29059 12452
rect 29099 12412 29108 12452
rect 29923 12412 29932 12452
rect 29972 12412 29981 12452
rect 30970 12412 30979 12452
rect 31019 12412 31028 12452
rect 25516 12328 25804 12368
rect 25844 12328 25853 12368
rect 25900 12328 27724 12368
rect 27764 12328 27773 12368
rect 27898 12328 28492 12368
rect 28532 12328 28644 12368
rect 25900 12284 25940 12328
rect 23491 12244 23500 12284
rect 23540 12244 23587 12284
rect 23971 12244 23980 12284
rect 24020 12244 24172 12284
rect 24212 12244 24221 12284
rect 25324 12244 25940 12284
rect 28675 12244 28684 12284
rect 28724 12244 28733 12284
rect 23500 12200 23540 12244
rect 28684 12200 28724 12244
rect 23491 12160 23500 12200
rect 23540 12160 23549 12200
rect 23683 12160 23692 12200
rect 23732 12160 24268 12200
rect 24308 12160 24317 12200
rect 28684 12160 30700 12200
rect 30740 12160 30749 12200
rect 26425 12076 26434 12116
rect 26802 12076 26811 12116
rect 26179 11992 26188 12032
rect 26228 11992 26420 12032
rect 26380 11948 26420 11992
rect 30988 11948 31028 12412
rect 23299 11908 23308 11948
rect 23348 11908 23444 11948
rect 25577 11908 25612 11948
rect 25652 11908 25708 11948
rect 25748 11908 25757 11948
rect 26083 11908 26092 11948
rect 26132 11908 26188 11948
rect 26228 11908 26263 11948
rect 26371 11908 26380 11948
rect 26420 11908 26429 11948
rect 28003 11908 28012 11948
rect 28052 11908 28061 11948
rect 29731 11908 29740 11948
rect 29780 11908 31028 11948
rect 28012 11864 28052 11908
rect 28012 11824 31276 11864
rect 31316 11824 31325 11864
rect 23107 11740 23116 11780
rect 23156 11740 23252 11780
rect 23308 11740 23596 11780
rect 23636 11740 23645 11780
rect 24931 11740 24940 11780
rect 24980 11740 25420 11780
rect 25460 11740 26132 11780
rect 26179 11740 26188 11780
rect 26228 11740 26516 11780
rect 23308 11696 23348 11740
rect 25455 11696 25495 11740
rect 26092 11696 26132 11740
rect 26476 11696 26516 11740
rect 27724 11740 28204 11780
rect 28244 11740 28419 11780
rect 28459 11740 28468 11780
rect 28963 11740 28972 11780
rect 29012 11740 30356 11780
rect 27724 11696 27764 11740
rect 29932 11696 29972 11740
rect 30316 11696 30356 11740
rect 8547 11656 8908 11696
rect 8948 11656 8957 11696
rect 9065 11656 9142 11696
rect 9182 11656 9196 11696
rect 9236 11656 9245 11696
rect 9475 11656 9484 11696
rect 9524 11656 9533 11696
rect 9582 11656 9591 11696
rect 9631 11656 9772 11696
rect 9812 11656 9821 11696
rect 10060 11656 10156 11696
rect 10196 11656 10327 11696
rect 10409 11656 10483 11696
rect 10523 11656 10540 11696
rect 10580 11656 10589 11696
rect 11011 11656 11020 11696
rect 11060 11656 11107 11696
rect 11147 11656 11212 11696
rect 11252 11656 11261 11696
rect 11771 11656 11780 11696
rect 11820 11656 11829 11696
rect 12643 11656 12652 11696
rect 12692 11656 12701 11696
rect 12826 11656 12835 11696
rect 12875 11656 12884 11696
rect 13018 11656 13027 11696
rect 13067 11656 13076 11696
rect 13174 11656 13183 11696
rect 13223 11656 13232 11696
rect 13276 11656 13285 11696
rect 13325 11656 13334 11696
rect 13397 11656 13406 11696
rect 13446 11656 13460 11696
rect 13507 11656 13516 11696
rect 13585 11656 13687 11696
rect 13747 11656 13756 11696
rect 13796 11656 13805 11696
rect 13961 11656 14071 11696
rect 14132 11656 14141 11696
rect 14218 11656 14227 11696
rect 14267 11656 14284 11696
rect 14324 11656 14407 11696
rect 14563 11656 14572 11696
rect 14612 11656 14621 11696
rect 14755 11656 14764 11696
rect 14804 11656 14947 11696
rect 14987 11656 14996 11696
rect 15056 11656 15065 11696
rect 15105 11656 15114 11696
rect 15188 11656 15197 11696
rect 15237 11656 15246 11696
rect 15322 11656 15331 11696
rect 15371 11656 15380 11696
rect 15427 11656 15436 11696
rect 15505 11656 15607 11696
rect 15689 11656 15820 11696
rect 15860 11656 15869 11696
rect 15946 11687 16004 11696
rect 8199 11614 8208 11654
rect 8248 11614 8265 11654
rect 6220 11572 6508 11612
rect 6548 11572 6557 11612
rect 6748 11572 6988 11612
rect 7028 11572 7679 11612
rect 7639 11570 7679 11572
rect 7852 11572 8084 11612
rect 8225 11612 8265 11614
rect 10060 11612 10100 11656
rect 11788 11612 11828 11656
rect 13036 11612 13076 11656
rect 8225 11572 8397 11612
rect 8515 11572 8524 11612
rect 8564 11572 8947 11612
rect 8987 11572 10100 11612
rect 11395 11572 11404 11612
rect 11444 11572 11596 11612
rect 11636 11572 11645 11612
rect 11742 11572 11788 11612
rect 11828 11572 11837 11612
rect 12739 11572 12748 11612
rect 12788 11572 13076 11612
rect 13192 11612 13232 11656
rect 13756 11612 13796 11656
rect 13192 11572 13228 11612
rect 13268 11572 13277 11612
rect 13516 11572 13796 11612
rect 14572 11612 14612 11656
rect 15946 11647 15955 11687
rect 15995 11647 16004 11687
rect 16051 11656 16060 11696
rect 16100 11656 16109 11696
rect 16154 11656 16163 11696
rect 16203 11656 16265 11696
rect 16326 11656 16335 11696
rect 16375 11656 16413 11696
rect 16482 11656 16588 11696
rect 16653 11656 16662 11696
rect 16762 11656 16771 11696
rect 16811 11656 16820 11696
rect 16906 11656 16915 11696
rect 16955 11656 16964 11696
rect 17150 11656 17163 11696
rect 17203 11656 17212 11696
rect 17321 11656 17332 11696
rect 17372 11656 17452 11696
rect 17492 11656 17501 11696
rect 17993 11656 18115 11696
rect 18164 11656 18173 11696
rect 19354 11656 19363 11696
rect 19403 11656 19700 11696
rect 15946 11646 16004 11647
rect 14572 11572 15532 11612
rect 15572 11572 15581 11612
rect 7852 11570 7892 11572
rect 7639 11530 7892 11570
rect 3427 11488 3436 11528
rect 3476 11488 3607 11528
rect 3811 11488 3820 11528
rect 3860 11488 5108 11528
rect 5251 11488 5260 11528
rect 5300 11488 5443 11528
rect 5483 11488 5492 11528
rect 5609 11488 5731 11528
rect 5780 11488 5789 11528
rect 7162 11488 7171 11528
rect 7211 11488 7220 11528
rect 5068 11444 5108 11488
rect 7180 11444 7220 11488
rect 8357 11444 8397 11572
rect 13516 11528 13556 11572
rect 15964 11528 16004 11646
rect 16225 11528 16265 11656
rect 16373 11612 16413 11656
rect 17050 11645 17108 11654
rect 17050 11612 17059 11645
rect 16373 11572 16396 11612
rect 16436 11605 17059 11612
rect 17099 11605 17108 11645
rect 16436 11604 17108 11605
rect 16436 11572 17093 11604
rect 17150 11528 17190 11656
rect 19660 11528 19700 11656
rect 20297 11656 20428 11696
rect 20468 11656 20477 11696
rect 20681 11656 20716 11696
rect 20756 11656 20812 11696
rect 20852 11656 20861 11696
rect 20921 11656 20930 11696
rect 20970 11656 21388 11696
rect 21428 11656 21437 11696
rect 21737 11656 21868 11696
rect 21908 11656 21917 11696
rect 21964 11656 22051 11696
rect 22091 11656 22100 11696
rect 22156 11656 22204 11696
rect 22244 11656 22253 11696
rect 22530 11656 22540 11696
rect 22580 11656 22661 11696
rect 22701 11656 22710 11696
rect 22781 11656 22803 11696
rect 22843 11656 22852 11696
rect 22906 11656 22915 11696
rect 22955 11656 22964 11696
rect 23011 11656 23020 11696
rect 23060 11656 23069 11696
rect 23299 11656 23308 11696
rect 23348 11656 23357 11696
rect 23600 11656 23609 11696
rect 23649 11656 23980 11696
rect 24020 11656 24460 11696
rect 24500 11656 24509 11696
rect 25193 11656 25324 11696
rect 25364 11656 25373 11696
rect 25437 11656 25446 11696
rect 25486 11656 25495 11696
rect 25555 11656 25564 11696
rect 25604 11656 25613 11696
rect 25987 11656 25996 11696
rect 26036 11656 26045 11696
rect 26092 11656 26380 11696
rect 26420 11656 26429 11696
rect 26476 11656 26577 11696
rect 26617 11656 26626 11696
rect 26729 11656 26860 11696
rect 26900 11656 26909 11696
rect 27523 11656 27532 11696
rect 27572 11656 27715 11696
rect 27755 11656 27764 11696
rect 27811 11656 27820 11696
rect 27860 11656 27991 11696
rect 28169 11656 28300 11696
rect 28340 11656 28349 11696
rect 28483 11656 28492 11696
rect 28557 11656 28663 11696
rect 28771 11656 28780 11696
rect 28820 11656 28876 11696
rect 28916 11656 28951 11696
rect 29539 11656 29548 11696
rect 29588 11656 29740 11696
rect 29780 11656 29789 11696
rect 29923 11656 29932 11696
rect 29972 11656 29981 11696
rect 30115 11656 30124 11696
rect 30164 11656 30173 11696
rect 30307 11656 30316 11696
rect 30356 11656 30365 11696
rect 30569 11656 30691 11696
rect 30740 11656 30749 11696
rect 19852 11612 19892 11656
rect 22156 11612 22196 11656
rect 23020 11612 23060 11656
rect 19852 11572 21580 11612
rect 21620 11572 21629 11612
rect 21955 11572 21964 11612
rect 22004 11572 22196 11612
rect 22540 11572 23060 11612
rect 23203 11572 23212 11612
rect 23252 11572 23500 11612
rect 23540 11572 24172 11612
rect 24212 11572 24221 11612
rect 22540 11570 22580 11572
rect 22449 11530 22458 11570
rect 22498 11530 22580 11570
rect 24460 11528 24500 11656
rect 25564 11612 25604 11656
rect 25507 11572 25516 11612
rect 25556 11572 25604 11612
rect 25996 11612 26036 11656
rect 30124 11612 30164 11656
rect 25996 11572 26476 11612
rect 26516 11572 26525 11612
rect 28017 11572 28026 11612
rect 28066 11572 28204 11612
rect 28244 11572 28253 11612
rect 28675 11572 28684 11612
rect 28724 11572 30164 11612
rect 30211 11572 30220 11612
rect 30260 11572 31180 11612
rect 31220 11572 31229 11612
rect 8611 11488 8620 11528
rect 8660 11488 13412 11528
rect 13498 11488 13507 11528
rect 13547 11488 13556 11528
rect 14345 11488 14467 11528
rect 14516 11488 14525 11528
rect 15305 11488 15427 11528
rect 15476 11488 15485 11528
rect 15964 11488 16012 11528
rect 16052 11488 16061 11528
rect 16225 11488 17190 11528
rect 19049 11488 19180 11528
rect 19220 11488 19229 11528
rect 19660 11488 21484 11528
rect 21524 11488 21533 11528
rect 23779 11488 23788 11528
rect 23828 11488 23884 11528
rect 23924 11488 23959 11528
rect 24460 11488 25891 11528
rect 25931 11488 25940 11528
rect 27331 11488 27340 11528
rect 27380 11488 27532 11528
rect 27572 11488 27581 11528
rect 28579 11488 28588 11528
rect 28628 11488 30892 11528
rect 30932 11488 30941 11528
rect 13372 11444 13412 11488
rect 4003 11404 4012 11444
rect 4052 11404 5012 11444
rect 5068 11404 6604 11444
rect 6644 11404 6653 11444
rect 7180 11404 8236 11444
rect 8276 11404 8285 11444
rect 8357 11404 8468 11444
rect 9955 11404 9964 11444
rect 10004 11404 13268 11444
rect 13372 11404 19508 11444
rect 4343 11320 4352 11360
rect 4720 11320 4729 11360
rect 4972 11192 5012 11404
rect 8428 11360 8468 11404
rect 13228 11360 13268 11404
rect 5539 11320 5548 11360
rect 5588 11320 8332 11360
rect 8372 11320 8381 11360
rect 8428 11320 8716 11360
rect 8756 11320 8765 11360
rect 12117 11320 12126 11360
rect 12494 11320 12503 11360
rect 12739 11320 12748 11360
rect 12788 11320 13036 11360
rect 13076 11320 13085 11360
rect 13228 11320 14420 11360
rect 14380 11276 14420 11320
rect 15820 11320 16396 11360
rect 16436 11320 16445 11360
rect 15820 11276 15860 11320
rect 6499 11236 6508 11276
rect 6548 11236 13556 11276
rect 14380 11236 15860 11276
rect 16099 11236 16108 11276
rect 16148 11236 19220 11276
rect 13516 11192 13556 11236
rect 19180 11192 19220 11236
rect 19468 11192 19508 11404
rect 4073 11152 4195 11192
rect 4244 11152 4253 11192
rect 4649 11152 4771 11192
rect 4820 11152 4829 11192
rect 4972 11152 5164 11192
rect 5204 11152 5213 11192
rect 6857 11152 6940 11192
rect 6980 11152 6988 11192
rect 7028 11152 7037 11192
rect 7145 11152 7180 11192
rect 7220 11152 7276 11192
rect 7316 11152 7325 11192
rect 7913 11152 8044 11192
rect 8084 11152 8093 11192
rect 8419 11152 8428 11192
rect 8468 11152 8852 11192
rect 8899 11152 8908 11192
rect 8948 11152 9100 11192
rect 9140 11152 9149 11192
rect 10531 11152 10540 11192
rect 10595 11152 10711 11192
rect 11369 11152 11395 11192
rect 11435 11152 11500 11192
rect 11540 11152 11549 11192
rect 11657 11152 11692 11192
rect 11732 11152 11788 11192
rect 11828 11152 11837 11192
rect 12595 11152 12604 11192
rect 12644 11152 12940 11192
rect 12980 11152 12989 11192
rect 13507 11152 13516 11192
rect 13556 11152 13565 11192
rect 13891 11152 13900 11192
rect 13940 11152 14371 11192
rect 14411 11152 14420 11192
rect 15610 11152 15619 11192
rect 15659 11152 15820 11192
rect 15860 11152 15869 11192
rect 16553 11152 16684 11192
rect 16724 11152 16733 11192
rect 16867 11152 16876 11192
rect 16916 11152 17836 11192
rect 17876 11152 17885 11192
rect 19171 11152 19180 11192
rect 19220 11152 19229 11192
rect 19459 11152 19468 11192
rect 19508 11152 19517 11192
rect 8812 11108 8852 11152
rect 1315 11068 1324 11108
rect 1364 11068 1373 11108
rect 1603 11068 1612 11108
rect 1652 11068 1728 11108
rect 3898 11068 3907 11108
rect 3947 11068 4300 11108
rect 4340 11068 4349 11108
rect 6211 11068 6220 11108
rect 6260 11068 8754 11108
rect 8812 11068 9301 11108
rect 10147 11068 10156 11108
rect 10196 11068 11540 11108
rect 11587 11068 11596 11108
rect 11636 11068 12172 11108
rect 12212 11068 12221 11108
rect 12940 11068 14860 11108
rect 14900 11068 14909 11108
rect 15139 11068 15148 11108
rect 15188 11068 15476 11108
rect 1324 11024 1364 11068
rect 1612 11024 1652 11068
rect 8714 11024 8754 11068
rect 1123 10984 1132 11024
rect 1172 10984 1181 11024
rect 1248 10984 1257 11024
rect 1297 10984 1364 11024
rect 1411 10984 1420 11024
rect 1460 10984 2092 11024
rect 2132 10984 2141 11024
rect 2572 10984 2860 11024
rect 2900 10984 2956 11024
rect 2996 10984 3005 11024
rect 3427 10984 3436 11024
rect 3488 10984 3607 11024
rect 4099 10984 4108 11024
rect 4148 10984 4157 11024
rect 4298 10984 4396 11024
rect 4460 10984 4478 11024
rect 4540 10984 4557 11024
rect 4597 10984 4606 11024
rect 4687 10984 4696 11024
rect 4736 10984 4745 11024
rect 4828 10984 4862 11024
rect 4902 10984 4911 11024
rect 4954 10984 4963 11024
rect 5003 11003 5012 11024
rect 5003 10984 5019 11003
rect 5129 10984 5260 11024
rect 5300 10984 5309 11024
rect 5417 10984 5497 11024
rect 5537 10984 5548 11024
rect 5588 10984 5597 11024
rect 6115 10984 6124 11024
rect 6164 10984 6412 11024
rect 6452 10984 6461 11024
rect 6586 10984 6595 11024
rect 6635 10984 6644 11024
rect 7075 10984 7084 11024
rect 7124 10984 7133 11024
rect 7241 10984 7372 11024
rect 7412 10984 7421 11024
rect 7529 10984 7609 11024
rect 7649 10984 7660 11024
rect 7700 10984 7709 11024
rect 8009 10984 8140 11024
rect 8180 10984 8189 11024
rect 8323 10984 8332 11024
rect 8397 10984 8503 11024
rect 8611 10984 8620 11024
rect 8660 10984 8669 11024
rect 8714 10984 8742 11024
rect 8782 10984 8791 11024
rect 8860 10984 8869 11024
rect 8948 10984 9049 11024
rect 9261 11015 9301 11068
rect 11500 11024 11540 11068
rect 1132 10940 1172 10984
rect 2572 10940 2612 10984
rect 1132 10900 1268 10940
rect 1315 10900 1324 10940
rect 1364 10900 2612 10940
rect 2659 10900 2668 10940
rect 2708 10900 3283 10940
rect 3323 10900 3332 10940
rect 1001 10816 1132 10856
rect 1172 10816 1181 10856
rect 1228 10436 1268 10900
rect 1507 10732 1516 10772
rect 1556 10732 2284 10772
rect 2324 10732 2333 10772
rect 4108 10688 4148 10984
rect 4540 10940 4580 10984
rect 4696 10940 4736 10984
rect 4828 10940 4868 10984
rect 4972 10963 5019 10984
rect 4540 10900 4588 10940
rect 4628 10900 4637 10940
rect 4684 10900 4736 10940
rect 4780 10900 4868 10940
rect 4684 10856 4724 10900
rect 4675 10816 4684 10856
rect 4724 10816 4733 10856
rect 4780 10772 4820 10900
rect 4979 10856 5019 10963
rect 6604 10940 6644 10984
rect 5386 10931 5740 10940
rect 5386 10891 5395 10931
rect 5435 10900 5740 10931
rect 5780 10900 5789 10940
rect 6307 10900 6316 10940
rect 6356 10900 6644 10940
rect 7084 10940 7124 10984
rect 7084 10900 7276 10940
rect 7316 10900 7325 10940
rect 7498 10931 7852 10940
rect 5435 10891 5444 10900
rect 5386 10890 5444 10891
rect 7498 10891 7507 10931
rect 7547 10900 7852 10931
rect 7892 10900 7901 10940
rect 8227 10900 8236 10940
rect 8299 10900 8407 10940
rect 7547 10891 7556 10900
rect 7498 10890 7556 10891
rect 4867 10816 4876 10856
rect 4916 10816 5019 10856
rect 4195 10732 4204 10772
rect 4244 10732 4820 10772
rect 5404 10688 5444 10890
rect 8620 10856 8660 10984
rect 9261 10966 9301 10975
rect 9370 11015 9428 11024
rect 9370 10975 9379 11015
rect 9419 10975 9428 11015
rect 9480 10984 9489 11024
rect 9529 10984 9964 11024
rect 10004 10984 10013 11024
rect 10205 10984 10252 11024
rect 10292 11015 10376 11024
rect 10292 10984 10336 11015
rect 9370 10974 9428 10975
rect 9388 10940 9428 10974
rect 10426 10984 10435 11024
rect 10484 10984 10615 11024
rect 11011 10984 11020 11024
rect 11060 10984 11063 11024
rect 11103 10984 11191 11024
rect 11297 10984 11306 11024
rect 11346 10984 11444 11024
rect 11500 10984 11596 11024
rect 11636 10984 11645 11024
rect 11753 10984 11788 11024
rect 11828 10984 11884 11024
rect 11924 10984 11933 11024
rect 10336 10966 10376 10975
rect 11404 10940 11444 10984
rect 12940 10940 12980 11068
rect 15436 11024 15476 11068
rect 16012 11068 16108 11108
rect 16148 11068 16157 11108
rect 16780 11068 17260 11108
rect 17300 11068 17309 11108
rect 17602 11068 17644 11108
rect 17684 11068 17693 11108
rect 16012 11066 16052 11068
rect 15964 11026 16052 11066
rect 13123 10984 13132 11024
rect 13172 10984 13243 11024
rect 13292 10984 13301 11024
rect 13341 10984 13350 11024
rect 13795 10984 13804 11024
rect 13869 10984 13975 11024
rect 14188 10984 14270 11024
rect 14310 10984 14319 11024
rect 14467 10984 14476 11024
rect 14516 10984 14525 11024
rect 14572 11015 14612 11024
rect 9388 10900 9772 10940
rect 9812 10900 10156 10940
rect 10196 10900 10205 10940
rect 11194 10900 11203 10940
rect 11243 10900 11252 10940
rect 11404 10900 11500 10940
rect 11540 10900 11549 10940
rect 11779 10900 11788 10940
rect 11828 10900 12364 10940
rect 12404 10900 12413 10940
rect 12460 10900 12980 10940
rect 11212 10856 11252 10900
rect 8620 10816 9100 10856
rect 9140 10816 9149 10856
rect 9571 10816 9580 10856
rect 9620 10816 10051 10856
rect 10091 10816 10100 10856
rect 10339 10816 10348 10856
rect 10388 10816 11252 10856
rect 6586 10732 6595 10772
rect 6644 10732 6775 10772
rect 8899 10732 8908 10772
rect 8948 10732 11692 10772
rect 11732 10732 11741 10772
rect 12460 10688 12500 10900
rect 13203 10856 13243 10984
rect 13294 10940 13334 10984
rect 13481 10942 13612 10982
rect 13652 10942 13661 10982
rect 13294 10900 13324 10940
rect 13364 10900 13374 10940
rect 13722 10900 13731 10940
rect 13771 10900 13996 10940
rect 14036 10900 14045 10940
rect 14188 10856 14228 10984
rect 14476 10940 14516 10984
rect 14275 10900 14284 10940
rect 14324 10900 14516 10940
rect 14825 10984 14956 11024
rect 14996 10984 15005 11024
rect 15113 10984 15193 11024
rect 15233 10984 15244 11024
rect 15284 10984 15293 11024
rect 15418 10984 15427 11024
rect 15467 10984 15476 11024
rect 15763 10984 15772 11024
rect 15812 10984 15821 11024
rect 13203 10816 13516 10856
rect 13556 10816 13565 10856
rect 13996 10816 14228 10856
rect 13996 10772 14036 10816
rect 14572 10772 14612 10975
rect 15772 10940 15812 10984
rect 15964 10940 16004 11026
rect 16780 11024 16820 11068
rect 17602 11024 17642 11068
rect 19660 11024 19700 11488
rect 19891 11320 19900 11360
rect 20268 11320 20277 11360
rect 24547 11320 24556 11360
rect 24596 11320 26996 11360
rect 27665 11320 27674 11360
rect 28042 11320 28051 11360
rect 19747 11236 19756 11276
rect 19796 11236 26132 11276
rect 21859 11152 21868 11192
rect 21908 11152 23980 11192
rect 24020 11152 24029 11192
rect 16234 10984 16243 11024
rect 16283 10984 16300 11024
rect 16340 10984 16423 11024
rect 16771 10984 16780 11024
rect 16820 10984 16829 11024
rect 17008 10984 17017 11024
rect 17057 10984 17164 11024
rect 17204 10984 17213 11024
rect 17347 10984 17356 11024
rect 17396 10984 17405 11024
rect 17584 10984 17593 11024
rect 17633 10984 17642 11024
rect 17731 10984 17740 11024
rect 17780 10984 17789 11024
rect 17923 10984 17932 11024
rect 17972 10984 18103 11024
rect 18682 10984 18691 11024
rect 18731 10984 18740 11024
rect 18953 10984 19084 11024
rect 19124 10984 19133 11024
rect 19180 10984 19276 11024
rect 19316 10984 19325 11024
rect 19642 10984 19651 11024
rect 19691 10984 19700 11024
rect 20140 11068 20620 11108
rect 20660 11068 20669 11108
rect 20812 11068 21196 11108
rect 21236 11068 21484 11108
rect 21524 11068 21533 11108
rect 22121 11068 22252 11108
rect 22292 11068 22301 11108
rect 22732 11068 23404 11108
rect 23444 11068 23453 11108
rect 24076 11068 24172 11108
rect 24212 11068 25036 11108
rect 25076 11068 25085 11108
rect 20140 11015 20180 11068
rect 20812 11024 20852 11068
rect 22732 11024 22772 11068
rect 24076 11024 24116 11068
rect 16090 10942 16099 10982
rect 16139 10942 16148 10982
rect 15082 10931 15340 10940
rect 15082 10891 15091 10931
rect 15131 10900 15340 10931
rect 15380 10900 15389 10940
rect 15436 10900 15812 10940
rect 15907 10900 15916 10940
rect 15956 10900 16004 10940
rect 15131 10891 15140 10900
rect 15082 10890 15140 10891
rect 15436 10856 15476 10900
rect 16108 10856 16148 10942
rect 16841 10931 16972 10940
rect 16841 10900 16915 10931
rect 16906 10891 16915 10900
rect 16955 10900 16972 10931
rect 17012 10900 17021 10940
rect 16955 10891 16964 10900
rect 16906 10890 16964 10891
rect 15390 10816 15399 10856
rect 15476 10816 15570 10856
rect 15881 10816 16012 10856
rect 16052 10816 16061 10856
rect 16108 10816 16396 10856
rect 16436 10816 16445 10856
rect 17356 10772 17396 10984
rect 17740 10940 17780 10984
rect 17482 10931 17644 10940
rect 17482 10891 17491 10931
rect 17531 10900 17644 10931
rect 17684 10900 17780 10940
rect 17827 10900 17836 10940
rect 17876 10900 18307 10940
rect 18347 10900 18356 10940
rect 17531 10891 17540 10900
rect 17482 10890 17540 10891
rect 18700 10856 18740 10984
rect 19180 10940 19220 10984
rect 20611 10984 20620 11024
rect 20660 10984 20852 11024
rect 20969 10984 21100 11024
rect 21140 10984 21149 11024
rect 21209 10984 21218 11024
rect 21258 10984 21388 11024
rect 21428 10984 21437 11024
rect 21763 10984 21772 11024
rect 21812 10984 21821 11024
rect 21946 10984 21955 11024
rect 22004 10984 22156 11024
rect 22196 10984 22205 11024
rect 22339 10984 22348 11024
rect 22388 10984 22397 11024
rect 22714 10984 22723 11024
rect 22763 10984 22772 11024
rect 22819 10984 22828 11024
rect 22868 10984 22999 11024
rect 23177 10984 23212 11024
rect 23252 10984 23308 11024
rect 23348 10984 23357 11024
rect 23482 10984 23491 11024
rect 23540 10984 23671 11024
rect 23753 10984 23884 11024
rect 23924 10984 23933 11024
rect 24058 10984 24067 11024
rect 24107 10984 24116 11024
rect 24268 11012 24460 11024
rect 20140 10966 20180 10975
rect 21772 10940 21812 10984
rect 22348 10940 22388 10984
rect 24169 10972 24178 11012
rect 24218 10984 24460 11012
rect 24500 10984 24509 11024
rect 24730 10984 24739 11024
rect 24779 10984 25996 11024
rect 26036 10984 26045 11024
rect 24218 10972 24308 10984
rect 26092 10940 26132 11236
rect 26956 11192 26996 11320
rect 26659 11152 26668 11192
rect 26708 11152 26860 11192
rect 26900 11152 26909 11192
rect 26956 11152 26995 11192
rect 27035 11152 27044 11192
rect 27907 11152 27916 11192
rect 27956 11152 28780 11192
rect 28820 11152 28829 11192
rect 26947 11068 26956 11108
rect 26996 11068 28588 11108
rect 28628 11068 28637 11108
rect 31145 11068 31267 11108
rect 31316 11068 31325 11108
rect 27628 11024 27668 11068
rect 27181 10984 27190 11024
rect 27230 10984 27340 11024
rect 27380 10984 27389 11024
rect 27514 10984 27523 11024
rect 27563 10984 27572 11024
rect 27619 10984 27628 11024
rect 27668 10984 27677 11024
rect 27977 10984 28108 11024
rect 28148 10984 29356 11024
rect 29396 10984 29405 11024
rect 30761 10984 30883 11024
rect 30932 10984 30941 11024
rect 27532 10940 27572 10984
rect 18874 10900 18883 10940
rect 18932 10900 19063 10940
rect 19171 10900 19180 10940
rect 19220 10900 19229 10940
rect 20585 10900 20716 10940
rect 20756 10900 20765 10940
rect 21772 10900 24116 10940
rect 24355 10900 24364 10940
rect 24404 10900 24413 10940
rect 25411 10900 25420 10940
rect 25460 10900 25469 10940
rect 26092 10900 26284 10940
rect 26324 10900 26333 10940
rect 27532 10900 29548 10940
rect 29588 10900 29597 10940
rect 30979 10900 30988 10940
rect 31028 10900 31037 10940
rect 18394 10816 18403 10856
rect 18443 10816 18452 10856
rect 18412 10772 18452 10816
rect 13306 10732 13315 10772
rect 13355 10732 13364 10772
rect 13987 10732 13996 10772
rect 14036 10732 14045 10772
rect 14572 10732 16108 10772
rect 16148 10732 16157 10772
rect 17356 10732 17932 10772
rect 17972 10732 18452 10772
rect 18700 10816 19948 10856
rect 19988 10816 19997 10856
rect 4108 10648 5444 10688
rect 6787 10648 6796 10688
rect 6836 10648 7316 10688
rect 7276 10604 7316 10648
rect 9196 10648 12500 10688
rect 9196 10604 9236 10648
rect 3103 10564 3112 10604
rect 3480 10564 3489 10604
rect 7276 10564 9236 10604
rect 10877 10564 10886 10604
rect 11254 10564 11263 10604
rect 8131 10480 8140 10520
rect 8180 10480 8620 10520
rect 8660 10480 8669 10520
rect 643 10396 652 10436
rect 692 10396 3724 10436
rect 3764 10396 3773 10436
rect 4841 10396 4876 10436
rect 4916 10396 4972 10436
rect 5012 10396 5021 10436
rect 5722 10396 5731 10436
rect 5771 10396 6740 10436
rect 7267 10396 7276 10436
rect 7316 10396 7325 10436
rect 9283 10396 9292 10436
rect 9332 10396 9475 10436
rect 9515 10396 9524 10436
rect 10636 10396 12748 10436
rect 12788 10396 12797 10436
rect 2362 10312 2371 10352
rect 2411 10312 2420 10352
rect 2380 10268 2420 10312
rect 3052 10312 6356 10352
rect 6595 10312 6604 10352
rect 6644 10312 6653 10352
rect 3052 10268 3092 10312
rect 1564 10228 2284 10268
rect 2324 10228 2333 10268
rect 2380 10228 2612 10268
rect 3043 10228 3052 10268
rect 3092 10228 3101 10268
rect 4469 10228 4492 10268
rect 4532 10228 4541 10268
rect 4673 10228 4684 10268
rect 4724 10228 4733 10268
rect 6089 10228 6220 10268
rect 6260 10228 6269 10268
rect 1564 10184 1604 10228
rect 2572 10184 2612 10228
rect 4307 10184 4316 10195
rect 835 10144 844 10184
rect 884 10144 1036 10184
rect 1076 10144 1085 10184
rect 1289 10144 1324 10184
rect 1364 10144 1420 10184
rect 1460 10144 1469 10184
rect 1546 10144 1555 10184
rect 1595 10144 1604 10184
rect 1708 10144 1996 10184
rect 2036 10144 2083 10184
rect 2123 10144 2132 10184
rect 2179 10144 2188 10184
rect 2228 10144 2359 10184
rect 2572 10144 2711 10184
rect 2751 10144 2760 10184
rect 2842 10144 2851 10184
rect 2891 10144 2900 10184
rect 2947 10144 2956 10184
rect 2996 10144 3127 10184
rect 3523 10144 3532 10184
rect 3572 10144 3716 10184
rect 3785 10144 3916 10184
rect 3956 10144 3965 10184
rect 4156 10155 4316 10184
rect 4356 10155 4365 10195
rect 4492 10184 4532 10228
rect 4673 10184 4713 10228
rect 4948 10184 5012 10189
rect 6316 10184 6356 10312
rect 6604 10268 6644 10312
rect 6442 10259 6644 10268
rect 6442 10219 6451 10259
rect 6491 10228 6644 10259
rect 6700 10268 6740 10396
rect 7049 10312 7180 10352
rect 7220 10312 7229 10352
rect 6700 10228 6915 10268
rect 6955 10228 6964 10268
rect 7075 10228 7084 10268
rect 7124 10228 7220 10268
rect 6491 10219 6500 10228
rect 6442 10218 6500 10219
rect 7180 10184 7220 10228
rect 7276 10184 7316 10396
rect 10636 10352 10676 10396
rect 7939 10312 7948 10352
rect 7988 10312 8468 10352
rect 8515 10312 8524 10352
rect 8564 10312 9004 10352
rect 9044 10312 10676 10352
rect 10723 10312 10732 10352
rect 10772 10312 10891 10352
rect 8428 10268 8468 10312
rect 7363 10228 7372 10268
rect 7412 10228 7651 10268
rect 7691 10228 7700 10268
rect 7747 10228 7756 10268
rect 7796 10228 7852 10268
rect 7892 10228 7927 10268
rect 8044 10228 8236 10268
rect 8276 10228 8285 10268
rect 8419 10228 8428 10268
rect 8468 10228 8477 10268
rect 8611 10228 8620 10268
rect 8660 10228 10540 10268
rect 10580 10228 10755 10268
rect 10795 10228 10804 10268
rect 8044 10184 8084 10228
rect 10851 10184 10891 10312
rect 10972 10226 11012 10396
rect 11068 10312 11116 10352
rect 11156 10312 11165 10352
rect 11779 10312 11788 10352
rect 11828 10312 12268 10352
rect 12308 10312 12317 10352
rect 12556 10312 13228 10352
rect 13268 10312 13277 10352
rect 11068 10268 11108 10312
rect 11068 10228 11093 10268
rect 11133 10228 11142 10268
rect 11299 10228 11308 10268
rect 11348 10228 11404 10268
rect 11444 10228 11479 10268
rect 11849 10228 11884 10268
rect 11924 10228 11980 10268
rect 12020 10228 12029 10268
rect 12233 10228 12364 10268
rect 12404 10228 12413 10268
rect 12556 10226 12596 10312
rect 13324 10268 13364 10732
rect 18700 10688 18740 10816
rect 24076 10772 24116 10900
rect 24364 10856 24404 10900
rect 24163 10816 24172 10856
rect 24212 10816 24404 10856
rect 28483 10816 28492 10856
rect 28532 10816 29492 10856
rect 29452 10772 29492 10816
rect 23002 10732 23011 10772
rect 23051 10732 23500 10772
rect 23540 10732 23549 10772
rect 24076 10732 24844 10772
rect 24884 10732 24893 10772
rect 28771 10732 28780 10772
rect 28820 10732 28829 10772
rect 28937 10732 28972 10772
rect 29012 10732 29068 10772
rect 29108 10732 29117 10772
rect 29225 10732 29356 10772
rect 29396 10732 29405 10772
rect 29452 10732 30412 10772
rect 30452 10732 30461 10772
rect 17452 10648 18740 10688
rect 17452 10604 17492 10648
rect 13603 10564 13612 10604
rect 13652 10564 13900 10604
rect 13940 10564 17492 10604
rect 18651 10564 18660 10604
rect 19028 10564 19037 10604
rect 19084 10564 20428 10604
rect 20468 10564 21292 10604
rect 21332 10564 21341 10604
rect 26425 10564 26434 10604
rect 26802 10564 26811 10604
rect 19084 10520 19124 10564
rect 28780 10520 28820 10732
rect 18700 10480 19124 10520
rect 19180 10480 20620 10520
rect 20660 10480 20669 10520
rect 21379 10480 21388 10520
rect 21428 10480 25132 10520
rect 25172 10480 27188 10520
rect 28780 10480 30164 10520
rect 18700 10436 18740 10480
rect 14825 10396 14947 10436
rect 14996 10396 15005 10436
rect 17251 10396 17260 10436
rect 17300 10396 18740 10436
rect 14659 10312 14668 10352
rect 14708 10312 15188 10352
rect 13306 10228 13315 10268
rect 13355 10228 13364 10268
rect 13507 10228 13516 10268
rect 13556 10228 14092 10268
rect 14132 10228 14141 10268
rect 14410 10228 14419 10268
rect 14459 10228 14572 10268
rect 14612 10228 14621 10268
rect 14740 10228 14860 10268
rect 14900 10228 14909 10268
rect 10963 10186 10972 10226
rect 11012 10186 11021 10226
rect 12490 10186 12499 10226
rect 12539 10186 12596 10226
rect 14428 10184 14468 10228
rect 14740 10184 14780 10228
rect 15148 10184 15188 10312
rect 16780 10312 16876 10352
rect 16916 10312 16925 10352
rect 17164 10312 17548 10352
rect 17588 10312 17597 10352
rect 16780 10268 16820 10312
rect 15305 10228 15340 10268
rect 15380 10228 15436 10268
rect 15476 10228 15485 10268
rect 15658 10259 15820 10268
rect 15658 10219 15667 10259
rect 15707 10228 15820 10259
rect 15860 10228 15869 10268
rect 16387 10228 16396 10268
rect 16436 10228 16492 10268
rect 16532 10228 16567 10268
rect 16714 10259 16820 10268
rect 15707 10219 15716 10228
rect 15658 10218 15716 10219
rect 16714 10219 16723 10259
rect 16763 10228 16820 10259
rect 17164 10268 17204 10312
rect 17164 10228 17187 10268
rect 17227 10228 17236 10268
rect 17443 10228 17452 10268
rect 17492 10228 17534 10268
rect 16763 10219 16772 10228
rect 16714 10218 16772 10219
rect 17447 10184 17487 10228
rect 18700 10184 18740 10396
rect 18787 10312 18796 10352
rect 18836 10312 19084 10352
rect 19124 10312 19133 10352
rect 19180 10268 19220 10480
rect 27148 10436 27188 10480
rect 19555 10396 19564 10436
rect 19604 10396 21100 10436
rect 21140 10396 21149 10436
rect 22435 10396 22444 10436
rect 22484 10396 23212 10436
rect 23252 10396 23261 10436
rect 24451 10396 24460 10436
rect 24500 10396 24652 10436
rect 24692 10396 24748 10436
rect 24788 10396 25804 10436
rect 25844 10396 25853 10436
rect 27139 10396 27148 10436
rect 27188 10396 27197 10436
rect 29539 10396 29548 10436
rect 29588 10396 29932 10436
rect 29972 10396 29981 10436
rect 18892 10228 19220 10268
rect 19276 10312 20716 10352
rect 20756 10312 20765 10352
rect 20899 10312 20908 10352
rect 20948 10312 21100 10352
rect 21140 10312 21716 10352
rect 23683 10312 23692 10352
rect 23732 10312 24076 10352
rect 24116 10312 25036 10352
rect 25076 10312 25085 10352
rect 25289 10312 25420 10352
rect 25460 10312 25469 10352
rect 27523 10312 27532 10352
rect 27572 10312 28387 10352
rect 28427 10312 28436 10352
rect 18892 10184 18932 10228
rect 19276 10184 19316 10312
rect 20044 10228 21580 10268
rect 21620 10228 21629 10268
rect 20044 10184 20084 10228
rect 21676 10184 21716 10312
rect 30124 10268 30164 10480
rect 21955 10228 21964 10268
rect 22004 10228 24556 10268
rect 24596 10228 24605 10268
rect 28291 10228 28300 10268
rect 28340 10228 30068 10268
rect 30124 10228 30260 10268
rect 30595 10228 30604 10268
rect 30644 10228 31036 10268
rect 31076 10228 31085 10268
rect 24556 10184 24596 10228
rect 28588 10184 28628 10228
rect 30028 10184 30068 10228
rect 30220 10184 30260 10228
rect 4156 10144 4354 10155
rect 4492 10144 4507 10184
rect 4547 10144 4556 10184
rect 4618 10144 4627 10184
rect 4667 10144 4713 10184
rect 4757 10144 4766 10184
rect 4806 10144 4815 10184
rect 4858 10144 4867 10184
rect 4907 10144 4972 10184
rect 5012 10144 5037 10184
rect 5321 10144 5356 10184
rect 5396 10144 5443 10184
rect 5483 10144 5492 10184
rect 5539 10144 5548 10184
rect 5588 10144 5719 10184
rect 6307 10144 6316 10184
rect 6356 10144 6365 10184
rect 6531 10144 6547 10184
rect 6587 10144 6596 10184
rect 6665 10144 6796 10184
rect 6836 10144 6845 10184
rect 7024 10144 7033 10184
rect 7073 10144 7082 10184
rect 7171 10144 7180 10184
rect 7220 10144 7229 10184
rect 7276 10144 7377 10184
rect 7417 10144 7426 10184
rect 7522 10144 7531 10184
rect 7571 10144 7604 10184
rect 7747 10144 7756 10184
rect 7796 10144 7852 10184
rect 7892 10144 7927 10184
rect 8035 10144 8044 10184
rect 8084 10144 8093 10184
rect 8140 10144 8236 10184
rect 8276 10144 8285 10184
rect 8332 10144 8524 10184
rect 8564 10144 8573 10184
rect 8620 10144 8643 10184
rect 8683 10144 8692 10184
rect 8752 10144 8761 10184
rect 8801 10144 8908 10184
rect 8948 10144 8957 10184
rect 9229 10144 9238 10184
rect 9278 10144 9868 10184
rect 9908 10144 9917 10184
rect 10505 10144 10636 10184
rect 10676 10144 10685 10184
rect 10851 10144 10867 10184
rect 10907 10144 10916 10184
rect 11196 10144 11205 10184
rect 11245 10144 11273 10184
rect 11534 10144 11543 10184
rect 11583 10144 11592 10184
rect 11674 10144 11683 10184
rect 11723 10144 11732 10184
rect 11779 10144 11788 10184
rect 11828 10144 11959 10184
rect 12036 10144 12045 10184
rect 12085 10144 12116 10184
rect 12163 10144 12172 10184
rect 12233 10144 12343 10184
rect 13194 10144 13203 10184
rect 13243 10144 13252 10184
rect 13315 10144 13324 10184
rect 13364 10144 13420 10184
rect 13460 10144 13495 10184
rect 13891 10144 13900 10184
rect 13940 10144 14468 10184
rect 14605 10144 14614 10184
rect 14654 10144 14780 10184
rect 14825 10175 14956 10184
rect 14825 10144 14851 10175
rect 1708 10016 1748 10144
rect 2668 10016 2708 10144
rect 2860 10100 2900 10144
rect 2755 10060 2764 10100
rect 2804 10060 2900 10100
rect 3676 10100 3716 10144
rect 4156 10100 4196 10144
rect 4775 10100 4815 10144
rect 6531 10100 6571 10144
rect 3676 10060 4052 10100
rect 4147 10060 4156 10100
rect 4196 10060 4205 10100
rect 4579 10060 4588 10100
rect 4628 10060 4815 10100
rect 6499 10060 6508 10100
rect 6548 10060 6571 10100
rect 7042 10100 7082 10144
rect 7564 10100 7604 10144
rect 8140 10100 8180 10144
rect 7042 10060 7124 10100
rect 7488 10060 7564 10100
rect 7604 10060 7613 10100
rect 8092 10060 8180 10100
rect 8332 10100 8372 10144
rect 8332 10060 8468 10100
rect 4012 10016 4052 10060
rect 7084 10016 7124 10060
rect 8092 10016 8132 10060
rect 8428 10016 8468 10060
rect 922 9976 931 10016
rect 971 9976 980 10016
rect 1699 9976 1708 10016
rect 1748 9976 1757 10016
rect 2668 9976 3052 10016
rect 3092 9976 3101 10016
rect 4012 9976 5068 10016
rect 5108 9976 5117 10016
rect 5705 9976 5836 10016
rect 5876 9976 5885 10016
rect 6595 9976 6604 10016
rect 6644 9976 6700 10016
rect 6740 9976 6775 10016
rect 7084 9976 7948 10016
rect 7988 9976 7997 10016
rect 8044 9976 8132 10016
rect 8218 9976 8227 10016
rect 8267 9976 8468 10016
rect 940 9848 980 9976
rect 940 9808 2572 9848
rect 2612 9808 2621 9848
rect 4204 9764 4244 9976
rect 8044 9932 8084 9976
rect 8620 9932 8660 10144
rect 11233 10100 11273 10144
rect 9034 10060 9043 10100
rect 9083 10060 9196 10100
rect 9236 10060 9245 10100
rect 10531 10060 10540 10100
rect 10580 10060 11273 10100
rect 11543 10100 11583 10144
rect 11692 10100 11732 10144
rect 12076 10100 12116 10144
rect 13200 10100 13240 10144
rect 14842 10135 14851 10144
rect 14891 10144 14956 10175
rect 14996 10144 15005 10184
rect 15139 10144 15148 10184
rect 15188 10144 15197 10184
rect 15401 10144 15532 10184
rect 15572 10144 15581 10184
rect 15760 10144 15769 10184
rect 15809 10144 16108 10184
rect 16148 10144 16157 10184
rect 16457 10144 16588 10184
rect 16628 10144 16637 10184
rect 16816 10144 16825 10184
rect 16865 10144 16916 10184
rect 17059 10144 17068 10184
rect 17108 10144 17117 10184
rect 17296 10144 17305 10184
rect 17345 10144 17354 10184
rect 17438 10144 17447 10184
rect 17487 10144 17496 10184
rect 17626 10144 17635 10184
rect 17684 10144 17815 10184
rect 18473 10144 18604 10184
rect 18644 10144 18653 10184
rect 18700 10144 18719 10184
rect 18759 10144 18768 10184
rect 18883 10144 18892 10184
rect 18932 10144 18941 10184
rect 18994 10144 19003 10184
rect 19043 10144 19084 10184
rect 19124 10144 19174 10184
rect 19267 10144 19276 10184
rect 19316 10144 19325 10184
rect 19817 10144 19948 10184
rect 19988 10144 19997 10184
rect 20201 10144 20320 10184
rect 20372 10144 20381 10184
rect 20524 10144 21148 10184
rect 21188 10144 21197 10184
rect 21283 10144 21292 10184
rect 21332 10144 21388 10184
rect 21428 10144 21463 10184
rect 21676 10144 21772 10184
rect 21812 10144 21821 10184
rect 22505 10144 22636 10184
rect 22676 10144 22685 10184
rect 23369 10144 23500 10184
rect 23540 10144 23549 10184
rect 24547 10144 24556 10184
rect 24596 10144 24605 10184
rect 24809 10144 24940 10184
rect 24980 10144 24989 10184
rect 25315 10144 25324 10184
rect 25364 10144 26668 10184
rect 26708 10144 26717 10184
rect 26851 10144 26860 10184
rect 26900 10144 27052 10184
rect 27092 10144 27436 10184
rect 27476 10144 27485 10184
rect 27977 10144 28108 10184
rect 28148 10144 28157 10184
rect 28387 10144 28396 10184
rect 28436 10144 28445 10184
rect 28579 10144 28588 10184
rect 28628 10144 28637 10184
rect 28937 10144 29068 10184
rect 29108 10144 29117 10184
rect 29164 10144 29932 10184
rect 29972 10144 29981 10184
rect 30028 10144 30047 10184
rect 30087 10144 30096 10184
rect 30211 10144 30220 10184
rect 30260 10144 30269 10184
rect 30316 10144 30355 10184
rect 30395 10144 30404 10184
rect 30499 10144 30508 10184
rect 30548 10144 30850 10184
rect 30890 10144 30899 10184
rect 14891 10135 14900 10144
rect 14842 10134 14900 10135
rect 11543 10060 11636 10100
rect 11692 10060 11980 10100
rect 12020 10060 12029 10100
rect 12076 10060 14380 10100
rect 14420 10060 14429 10100
rect 11596 9932 11636 10060
rect 15148 9932 15188 10144
rect 16876 10100 16916 10144
rect 17067 10100 17107 10144
rect 16841 10060 16876 10100
rect 16916 10060 16972 10100
rect 17012 10060 17021 10100
rect 17067 10060 17164 10100
rect 17204 10060 17267 10100
rect 17067 10016 17107 10060
rect 17314 10016 17354 10144
rect 20044 10135 20084 10144
rect 20524 10100 20564 10144
rect 17827 10060 17836 10100
rect 17876 10060 19180 10100
rect 19220 10060 19229 10100
rect 19651 10060 19660 10100
rect 19700 10060 19742 10100
rect 19782 10060 19831 10100
rect 20419 10060 20428 10100
rect 20468 10060 20476 10100
rect 20516 10060 20599 10100
rect 26668 10016 26708 10144
rect 28396 10100 28436 10144
rect 29164 10100 29204 10144
rect 30316 10100 30356 10144
rect 26755 10060 26764 10100
rect 26804 10060 29204 10100
rect 29731 10060 29740 10100
rect 29780 10060 30356 10100
rect 30403 10060 30412 10100
rect 30452 10060 30556 10100
rect 30596 10060 30605 10100
rect 15811 9976 15820 10016
rect 15860 9976 17107 10016
rect 17260 9976 17354 10016
rect 17417 9976 17548 10016
rect 17588 9976 17597 10016
rect 19721 9976 19843 10016
rect 19892 9976 19901 10016
rect 23261 9976 23308 10016
rect 23348 9976 23357 10016
rect 23779 9976 23788 10016
rect 23828 9976 24172 10016
rect 24212 9976 24221 10016
rect 24442 9976 24451 10016
rect 24491 9976 24844 10016
rect 24884 9976 24893 10016
rect 26668 9976 27052 10016
rect 27092 9976 27101 10016
rect 27305 9976 27340 10016
rect 27380 9976 27436 10016
rect 27476 9976 27485 10016
rect 17260 9932 17300 9976
rect 23308 9932 23348 9976
rect 8035 9892 8044 9932
rect 8084 9892 8093 9932
rect 8620 9892 10388 9932
rect 10435 9892 10444 9932
rect 10484 9892 14284 9932
rect 14324 9892 14333 9932
rect 15148 9892 17260 9932
rect 17300 9892 17309 9932
rect 19756 9892 20428 9932
rect 20468 9892 20477 9932
rect 20707 9892 20716 9932
rect 20756 9892 23252 9932
rect 23299 9892 23308 9932
rect 23348 9892 23357 9932
rect 24364 9892 29356 9932
rect 29396 9892 29405 9932
rect 10348 9848 10388 9892
rect 19756 9848 19796 9892
rect 23212 9848 23252 9892
rect 24364 9848 24404 9892
rect 4343 9808 4352 9848
rect 4720 9808 4729 9848
rect 7564 9808 9044 9848
rect 9379 9808 9388 9848
rect 9428 9808 10196 9848
rect 10348 9808 11596 9848
rect 11636 9808 11645 9848
rect 12117 9808 12126 9848
rect 12494 9808 12503 9848
rect 17443 9808 17452 9848
rect 17492 9808 19796 9848
rect 19891 9808 19900 9848
rect 20268 9808 20277 9848
rect 20611 9808 20620 9848
rect 20660 9808 23060 9848
rect 23212 9808 24404 9848
rect 24451 9808 24460 9848
rect 24500 9808 25612 9848
rect 25652 9808 26612 9848
rect 27665 9808 27674 9848
rect 28042 9808 28051 9848
rect 7564 9764 7604 9808
rect 1708 9724 3628 9764
rect 3668 9724 3677 9764
rect 4204 9724 4340 9764
rect 1594 9640 1603 9680
rect 1643 9640 1652 9680
rect 1027 9472 1036 9512
rect 1076 9472 1123 9512
rect 1163 9472 1207 9512
rect 1385 9472 1420 9512
rect 1460 9472 1516 9512
rect 1556 9472 1565 9512
rect 1612 9428 1652 9640
rect 1708 9512 1748 9724
rect 4300 9680 4340 9724
rect 6149 9724 7564 9764
rect 7604 9724 7613 9764
rect 7756 9724 8564 9764
rect 1891 9640 1900 9680
rect 1940 9640 2188 9680
rect 2228 9640 2237 9680
rect 2842 9640 2851 9680
rect 2891 9640 3052 9680
rect 3092 9640 3101 9680
rect 4291 9640 4300 9680
rect 4340 9640 4349 9680
rect 5801 9640 5836 9680
rect 5876 9640 5932 9680
rect 5972 9640 5981 9680
rect 2188 9596 2228 9640
rect 2188 9556 2324 9596
rect 2947 9556 2956 9596
rect 2996 9556 3127 9596
rect 2284 9512 2324 9556
rect 6149 9512 6189 9724
rect 6394 9640 6403 9680
rect 6443 9640 7220 9680
rect 7337 9640 7459 9680
rect 7508 9640 7517 9680
rect 7180 9596 7220 9640
rect 7756 9596 7796 9724
rect 8524 9680 8564 9724
rect 7843 9640 7852 9680
rect 7892 9640 8419 9680
rect 8459 9640 8468 9680
rect 8515 9640 8524 9680
rect 8564 9640 8573 9680
rect 8777 9640 8908 9680
rect 8948 9640 8957 9680
rect 6487 9556 6618 9596
rect 6658 9556 6667 9596
rect 6883 9556 6892 9596
rect 6932 9556 7124 9596
rect 7180 9556 7852 9596
rect 7892 9556 7901 9596
rect 8201 9556 8321 9596
rect 8372 9556 8381 9596
rect 7084 9512 7124 9556
rect 9004 9512 9044 9808
rect 10156 9764 10196 9808
rect 10156 9724 15572 9764
rect 16003 9724 16012 9764
rect 16052 9724 21676 9764
rect 21716 9724 21725 9764
rect 15532 9680 15572 9724
rect 23020 9680 23060 9808
rect 9187 9640 9196 9680
rect 9236 9640 10348 9680
rect 10388 9640 10483 9680
rect 10523 9640 10532 9680
rect 10819 9640 10828 9680
rect 10868 9640 11107 9680
rect 11147 9640 11404 9680
rect 11444 9640 11453 9680
rect 11587 9640 11596 9680
rect 11636 9640 11779 9680
rect 11819 9640 11828 9680
rect 11875 9640 11884 9680
rect 11924 9640 12364 9680
rect 12404 9640 12413 9680
rect 13588 9640 13597 9680
rect 13637 9640 13687 9680
rect 14419 9640 14428 9680
rect 14468 9640 14956 9680
rect 14996 9640 15005 9680
rect 15523 9640 15532 9680
rect 15572 9640 15581 9680
rect 15955 9640 15964 9680
rect 16004 9640 17164 9680
rect 17204 9640 17213 9680
rect 17746 9640 18316 9680
rect 18356 9640 18365 9680
rect 18499 9640 18508 9680
rect 18548 9640 18835 9680
rect 18875 9640 18884 9680
rect 19241 9640 19372 9680
rect 19412 9640 19421 9680
rect 19468 9640 19700 9680
rect 19843 9640 19852 9680
rect 19892 9640 20276 9680
rect 20515 9640 20524 9680
rect 20564 9640 22636 9680
rect 22676 9640 22685 9680
rect 23020 9640 25612 9680
rect 25652 9640 25661 9680
rect 13647 9596 13687 9640
rect 17746 9596 17786 9640
rect 19468 9596 19508 9640
rect 19660 9596 19700 9640
rect 10531 9556 10540 9596
rect 10580 9556 11212 9596
rect 11252 9556 11261 9596
rect 11308 9556 11932 9596
rect 11972 9556 11981 9596
rect 13507 9556 13516 9596
rect 13556 9556 13687 9596
rect 14620 9556 17786 9596
rect 18691 9556 18700 9596
rect 18740 9556 19508 9596
rect 19555 9556 19564 9596
rect 19604 9556 19613 9596
rect 19660 9556 19892 9596
rect 20009 9556 20131 9596
rect 20180 9556 20189 9596
rect 1699 9472 1708 9512
rect 1748 9472 1757 9512
rect 2050 9472 2059 9512
rect 2099 9472 2188 9512
rect 2228 9472 2237 9512
rect 2284 9472 2345 9512
rect 2385 9472 2394 9512
rect 2506 9472 2515 9512
rect 2555 9472 2612 9512
rect 2659 9472 2668 9512
rect 2708 9472 2755 9512
rect 2795 9472 2839 9512
rect 2903 9472 3063 9512
rect 3103 9472 5644 9512
rect 5684 9472 5693 9512
rect 5801 9472 5932 9512
rect 5972 9472 5981 9512
rect 6140 9472 6149 9512
rect 6189 9472 6198 9512
rect 6298 9472 6307 9512
rect 6347 9472 6356 9512
rect 6403 9472 6412 9512
rect 6452 9472 6796 9512
rect 6836 9472 6845 9512
rect 6970 9472 6979 9512
rect 7019 9472 7028 9512
rect 7084 9472 7127 9512
rect 7167 9472 7176 9512
rect 7363 9472 7372 9512
rect 7412 9472 7543 9512
rect 7817 9472 7948 9512
rect 7988 9472 7997 9512
rect 8065 9472 8140 9512
rect 8180 9472 8182 9512
rect 8222 9472 8243 9512
rect 8620 9503 8756 9512
rect 2572 9428 2612 9472
rect 2903 9428 2943 9472
rect 6316 9428 6356 9472
rect 1612 9388 1804 9428
rect 1844 9388 1853 9428
rect 1987 9388 1996 9428
rect 2036 9388 2188 9428
rect 2228 9388 2237 9428
rect 2563 9388 2572 9428
rect 2612 9388 2621 9428
rect 2851 9388 2860 9428
rect 2900 9388 2943 9428
rect 5827 9388 5836 9428
rect 5876 9388 6051 9428
rect 6091 9388 6100 9428
rect 6211 9388 6220 9428
rect 6260 9388 6356 9428
rect 6988 9428 7028 9472
rect 8140 9471 8228 9472
rect 8660 9472 8756 9503
rect 8803 9472 8812 9512
rect 8852 9472 8861 9512
rect 8995 9472 9004 9512
rect 9044 9472 10444 9512
rect 10484 9472 10493 9512
rect 10627 9472 10636 9512
rect 10688 9472 10807 9512
rect 10915 9472 10924 9512
rect 10964 9472 11006 9512
rect 11046 9472 11095 9512
rect 11308 9503 11348 9556
rect 8620 9454 8660 9463
rect 8716 9428 8756 9472
rect 6988 9388 7084 9428
rect 7124 9388 7133 9428
rect 7258 9388 7267 9428
rect 7307 9388 7756 9428
rect 7796 9388 7805 9428
rect 8074 9419 8132 9428
rect 8074 9379 8083 9419
rect 8123 9379 8132 9419
rect 8707 9388 8716 9428
rect 8756 9388 8765 9428
rect 8074 9378 8132 9379
rect 8092 9344 8132 9378
rect 2275 9304 2284 9344
rect 2324 9304 5260 9344
rect 5300 9304 5309 9344
rect 8092 9304 8180 9344
rect 8140 9260 8180 9304
rect 8812 9260 8852 9472
rect 11395 9472 11404 9512
rect 11444 9472 11447 9512
rect 11487 9472 11575 9512
rect 11683 9472 11692 9512
rect 11732 9472 11863 9512
rect 12067 9472 12076 9512
rect 12116 9472 12247 9512
rect 12809 9472 12844 9512
rect 12884 9472 12940 9512
rect 12980 9472 12989 9512
rect 13219 9472 13228 9512
rect 13268 9472 13399 9512
rect 13577 9472 13612 9512
rect 13652 9472 13699 9512
rect 13739 9472 13757 9512
rect 13804 9503 13900 9512
rect 11308 9454 11348 9463
rect 13844 9472 13900 9503
rect 13940 9472 14004 9512
rect 14153 9503 14284 9512
rect 14153 9472 14275 9503
rect 14324 9472 14333 9512
rect 13804 9428 13844 9463
rect 14266 9463 14275 9472
rect 14315 9463 14324 9472
rect 14266 9462 14324 9463
rect 11578 9388 11587 9428
rect 11627 9388 11884 9428
rect 11924 9388 11933 9428
rect 13027 9388 13036 9428
rect 13076 9388 13844 9428
rect 14620 9344 14660 9556
rect 16695 9512 16735 9556
rect 14729 9503 14860 9512
rect 14729 9472 14755 9503
rect 14746 9463 14755 9472
rect 14795 9472 14860 9503
rect 14900 9472 14909 9512
rect 15305 9472 15436 9512
rect 15476 9472 15485 9512
rect 15610 9472 15619 9512
rect 15659 9472 15668 9512
rect 14795 9463 14804 9472
rect 14746 9462 14804 9463
rect 14899 9388 14908 9428
rect 14948 9388 14956 9428
rect 14996 9388 15079 9428
rect 13219 9304 13228 9344
rect 13268 9304 14660 9344
rect 15628 9344 15668 9472
rect 15802 9503 15820 9512
rect 15802 9463 15811 9503
rect 15860 9472 15991 9512
rect 16099 9472 16108 9512
rect 16148 9472 16588 9512
rect 16628 9472 16637 9512
rect 16694 9472 16703 9512
rect 16743 9472 16752 9512
rect 16867 9472 16876 9512
rect 16916 9472 17452 9512
rect 17492 9472 17501 9512
rect 17548 9472 17591 9512
rect 17631 9472 17640 9512
rect 17827 9472 17836 9512
rect 17876 9472 18007 9512
rect 19021 9472 19030 9512
rect 19070 9472 19220 9512
rect 19267 9472 19276 9512
rect 19316 9472 19468 9512
rect 19508 9472 19517 9512
rect 15851 9463 15860 9472
rect 15802 9462 15860 9463
rect 16588 9428 16628 9472
rect 17548 9428 17588 9472
rect 19180 9428 19220 9472
rect 19564 9428 19604 9556
rect 19852 9512 19892 9556
rect 19810 9472 19819 9512
rect 19859 9472 19892 9512
rect 20028 9472 20037 9512
rect 20077 9472 20180 9512
rect 19699 9430 19708 9470
rect 19748 9430 19757 9470
rect 16588 9388 16724 9428
rect 17251 9388 17260 9428
rect 17300 9388 17588 9428
rect 17635 9388 17644 9428
rect 17684 9388 17731 9428
rect 17771 9388 17815 9428
rect 17923 9388 17932 9428
rect 17972 9388 18316 9428
rect 18356 9388 18365 9428
rect 19049 9388 19180 9428
rect 19220 9388 19468 9428
rect 19508 9388 19517 9428
rect 19564 9388 19587 9428
rect 19627 9388 19636 9428
rect 16684 9344 16724 9388
rect 15628 9304 16588 9344
rect 16628 9304 16637 9344
rect 16684 9304 18700 9344
rect 18740 9304 18749 9344
rect 1289 9220 1324 9260
rect 1364 9220 1420 9260
rect 1460 9220 1469 9260
rect 3619 9220 3628 9260
rect 3668 9220 5588 9260
rect 5923 9220 5932 9260
rect 5972 9220 6604 9260
rect 6644 9220 6653 9260
rect 8140 9220 8332 9260
rect 8372 9220 8852 9260
rect 13459 9220 13468 9260
rect 13508 9220 13612 9260
rect 13652 9220 13661 9260
rect 14083 9220 14092 9260
rect 14132 9220 14380 9260
rect 14420 9220 14429 9260
rect 5548 9092 5588 9220
rect 6019 9136 6028 9176
rect 6068 9136 13228 9176
rect 13268 9136 13277 9176
rect 259 9052 268 9092
rect 308 9052 500 9092
rect 3103 9052 3112 9092
rect 3480 9052 3489 9092
rect 5548 9052 9772 9092
rect 9812 9052 9821 9092
rect 10877 9052 10886 9092
rect 11254 9052 11263 9092
rect 18651 9052 18660 9092
rect 19028 9052 19037 9092
rect 0 8924 400 8944
rect 460 8924 500 9052
rect 8572 8968 9196 9008
rect 9236 8968 11404 9008
rect 11444 8968 11453 9008
rect 0 8884 500 8924
rect 1097 8884 1219 8924
rect 1268 8884 1277 8924
rect 1987 8884 1996 8924
rect 2036 8884 2572 8924
rect 2612 8884 2621 8924
rect 3785 8884 3907 8924
rect 3956 8884 3965 8924
rect 4012 8884 4876 8924
rect 4916 8884 4925 8924
rect 5626 8884 5635 8924
rect 5675 8884 8084 8924
rect 8201 8884 8323 8924
rect 8372 8884 8381 8924
rect 0 8864 400 8884
rect 2188 8800 2380 8840
rect 2420 8800 2429 8840
rect 2572 8800 2764 8840
rect 2804 8800 2813 8840
rect 2188 8672 2228 8800
rect 2572 8756 2612 8800
rect 4012 8756 4052 8884
rect 2275 8716 2284 8756
rect 2324 8716 2420 8756
rect 2554 8716 2563 8756
rect 2603 8716 2612 8756
rect 2755 8716 2764 8756
rect 2804 8716 3668 8756
rect 2380 8672 2420 8716
rect 2956 8672 2996 8716
rect 3628 8672 3668 8716
rect 3724 8716 4052 8756
rect 4660 8800 7028 8840
rect 3724 8672 3764 8716
rect 1603 8632 1612 8672
rect 1652 8632 2092 8672
rect 2132 8632 2228 8672
rect 2275 8632 2284 8672
rect 2324 8632 2333 8672
rect 2380 8632 2423 8672
rect 2463 8632 2472 8672
rect 2659 8632 2668 8672
rect 2708 8632 2717 8672
rect 2938 8632 2947 8672
rect 2987 8632 3072 8672
rect 3235 8632 3244 8672
rect 3284 8632 3476 8672
rect 3610 8632 3619 8672
rect 3659 8632 3668 8672
rect 3715 8632 3724 8672
rect 3764 8632 3773 8672
rect 3907 8632 3916 8672
rect 3956 8632 4195 8672
rect 4235 8632 4244 8672
rect 4291 8632 4300 8672
rect 4340 8632 4471 8672
rect 2284 8588 2324 8632
rect 1795 8548 1804 8588
rect 1844 8548 2380 8588
rect 2420 8548 2484 8588
rect 0 8504 400 8524
rect 2668 8504 2708 8632
rect 3436 8588 3476 8632
rect 3724 8588 3764 8632
rect 3436 8548 3764 8588
rect 3820 8548 4503 8588
rect 4543 8548 4552 8588
rect 3820 8504 3860 8548
rect 4660 8504 4700 8800
rect 4969 8716 4978 8756
rect 5018 8716 5164 8756
rect 5204 8716 5213 8756
rect 6988 8672 7028 8800
rect 8044 8672 8084 8884
rect 8572 8672 8612 8968
rect 19714 8924 19754 9430
rect 19852 9388 19925 9428
rect 19965 9388 19974 9428
rect 19852 9344 19892 9388
rect 20140 9344 20180 9472
rect 19852 9304 19948 9344
rect 19988 9304 19997 9344
rect 20131 9304 20140 9344
rect 20180 9304 20189 9344
rect 20236 9092 20276 9640
rect 22444 9556 24211 9596
rect 24251 9556 24844 9596
rect 24884 9556 24893 9596
rect 25795 9556 25804 9596
rect 25844 9556 26132 9596
rect 22444 9512 22484 9556
rect 26092 9512 26132 9556
rect 26572 9512 26612 9808
rect 27043 9724 27052 9764
rect 27092 9724 27572 9764
rect 27532 9680 27572 9724
rect 28204 9724 29012 9764
rect 26764 9640 27436 9680
rect 27476 9640 27485 9680
rect 27532 9640 27619 9680
rect 27659 9640 27668 9680
rect 27715 9640 27724 9680
rect 27764 9640 28108 9680
rect 28148 9640 28157 9680
rect 26764 9512 26804 9640
rect 28204 9596 28244 9724
rect 28972 9680 29012 9724
rect 28649 9640 28684 9680
rect 28724 9640 28780 9680
rect 28820 9640 28829 9680
rect 28963 9640 28972 9680
rect 29012 9640 29021 9680
rect 26851 9556 26860 9596
rect 26900 9556 28244 9596
rect 28291 9556 28300 9596
rect 28340 9556 28724 9596
rect 30211 9556 30220 9596
rect 30260 9556 30508 9596
rect 30548 9556 30557 9596
rect 31171 9556 31180 9596
rect 31220 9556 31267 9596
rect 31307 9556 31351 9596
rect 27388 9512 27428 9556
rect 28684 9512 28724 9556
rect 22426 9472 22435 9512
rect 22475 9472 22484 9512
rect 23299 9472 23308 9512
rect 23348 9472 23416 9512
rect 23456 9472 23479 9512
rect 23587 9472 23596 9512
rect 23636 9472 23645 9512
rect 23770 9472 23779 9512
rect 23828 9472 23959 9512
rect 24355 9472 24364 9512
rect 24416 9472 24535 9512
rect 24940 9485 25036 9512
rect 20419 9388 20428 9428
rect 20468 9388 20899 9428
rect 20948 9388 20957 9428
rect 21763 9388 21772 9428
rect 21812 9388 21821 9428
rect 22810 9388 22819 9428
rect 22859 9388 23060 9428
rect 23242 9388 23251 9428
rect 23291 9388 23500 9428
rect 23540 9388 23549 9428
rect 23020 9344 23060 9388
rect 23596 9344 23636 9472
rect 24846 9445 24855 9485
rect 24895 9472 25036 9485
rect 25076 9472 25085 9512
rect 25769 9472 25804 9512
rect 25844 9472 25900 9512
rect 25940 9472 25949 9512
rect 26083 9472 26092 9512
rect 26132 9472 26141 9512
rect 26188 9472 26214 9512
rect 26254 9472 26263 9512
rect 26332 9472 26341 9512
rect 26381 9472 26420 9512
rect 26563 9472 26572 9512
rect 26612 9472 26621 9512
rect 26746 9472 26755 9512
rect 26795 9472 26804 9512
rect 26851 9472 26860 9512
rect 26900 9472 27244 9512
rect 27284 9472 27293 9512
rect 27370 9472 27379 9512
rect 27419 9472 27428 9512
rect 27514 9472 27523 9512
rect 27572 9472 27703 9512
rect 27825 9472 27834 9512
rect 27874 9472 28108 9512
rect 28148 9472 28157 9512
rect 24895 9445 24980 9472
rect 25036 9428 25076 9472
rect 26188 9428 26228 9472
rect 26380 9428 26420 9472
rect 28472 9445 28481 9485
rect 28521 9445 28530 9485
rect 28618 9472 28627 9512
rect 28667 9472 28724 9512
rect 30403 9472 30412 9512
rect 30452 9472 30883 9512
rect 30932 9472 30941 9512
rect 24623 9388 24652 9428
rect 24692 9388 24754 9428
rect 24794 9388 24803 9428
rect 25036 9388 26228 9428
rect 26275 9388 26284 9428
rect 26324 9388 26420 9428
rect 27043 9388 27052 9428
rect 27092 9388 27187 9428
rect 27227 9388 27236 9428
rect 28478 9344 28518 9445
rect 29225 9388 29347 9428
rect 29396 9388 29405 9428
rect 31075 9388 31084 9428
rect 31124 9388 31133 9428
rect 23020 9304 23308 9344
rect 23348 9304 23357 9344
rect 23596 9304 24460 9344
rect 24500 9304 24509 9344
rect 26371 9304 26380 9344
rect 26420 9304 26956 9344
rect 26996 9304 28300 9344
rect 28340 9304 28349 9344
rect 28478 9304 28972 9344
rect 29012 9304 29021 9344
rect 23657 9220 23779 9260
rect 23828 9220 23837 9260
rect 24643 9220 24652 9260
rect 24692 9220 24701 9260
rect 26729 9220 26860 9260
rect 26900 9220 26909 9260
rect 20419 9136 20428 9176
rect 20468 9136 21964 9176
rect 22004 9136 22013 9176
rect 20236 9052 23692 9092
rect 23732 9052 23741 9092
rect 19939 8968 19948 9008
rect 19988 8968 21292 9008
rect 21332 8968 21341 9008
rect 21571 8968 21580 9008
rect 21620 8968 23060 9008
rect 23020 8924 23060 8968
rect 12643 8884 12652 8924
rect 12692 8884 12844 8924
rect 12884 8884 12893 8924
rect 13699 8884 13708 8924
rect 13748 8884 13900 8924
rect 13940 8884 13949 8924
rect 14458 8884 14467 8924
rect 14507 8884 14516 8924
rect 14563 8884 14572 8924
rect 14612 8884 16684 8924
rect 16724 8884 16733 8924
rect 17452 8884 19604 8924
rect 19714 8884 20035 8924
rect 20075 8884 20084 8924
rect 23020 8884 23452 8924
rect 23492 8884 23501 8924
rect 14476 8840 14516 8884
rect 11194 8800 11203 8840
rect 11243 8800 12076 8840
rect 12116 8800 12125 8840
rect 14476 8800 15668 8840
rect 9091 8716 9100 8756
rect 9140 8716 9196 8756
rect 9236 8716 9271 8756
rect 10924 8716 11212 8756
rect 11252 8716 11261 8756
rect 11395 8716 11404 8756
rect 11444 8716 11587 8756
rect 11627 8716 11636 8756
rect 11779 8716 11788 8756
rect 11828 8716 12404 8756
rect 13603 8716 13612 8756
rect 13652 8716 13661 8756
rect 13708 8716 14572 8756
rect 14612 8716 14621 8756
rect 15043 8716 15052 8756
rect 15092 8716 15532 8756
rect 15572 8716 15581 8756
rect 9772 8672 9812 8681
rect 10924 8672 10964 8716
rect 12364 8714 12404 8716
rect 12364 8705 12408 8714
rect 12364 8674 12368 8705
rect 5059 8632 5068 8672
rect 5108 8632 6028 8672
rect 6068 8632 6077 8672
rect 6874 8632 6883 8672
rect 6923 8632 6932 8672
rect 6979 8632 6988 8672
rect 7028 8632 7084 8672
rect 7124 8632 7188 8672
rect 8026 8632 8035 8672
rect 8075 8632 8084 8672
rect 8131 8632 8140 8672
rect 8180 8632 8612 8672
rect 8698 8632 8707 8672
rect 8747 8632 8756 8672
rect 8803 8632 8812 8672
rect 8852 8632 9004 8672
rect 9044 8632 9053 8672
rect 9161 8632 9292 8672
rect 9332 8632 9341 8672
rect 9641 8632 9772 8672
rect 9812 8632 9821 8672
rect 10217 8632 10291 8672
rect 10331 8632 10348 8672
rect 10388 8632 10397 8672
rect 10906 8632 10915 8672
rect 10955 8632 10964 8672
rect 11011 8632 11020 8672
rect 11060 8632 11069 8672
rect 11369 8632 11467 8672
rect 11540 8632 11549 8672
rect 11683 8632 11692 8672
rect 11732 8632 11863 8672
rect 12137 8632 12259 8672
rect 12308 8632 12317 8672
rect 13612 8672 13652 8716
rect 13708 8672 13748 8716
rect 14764 8672 14804 8681
rect 15628 8672 15668 8800
rect 17452 8756 17492 8884
rect 17539 8800 17548 8840
rect 17588 8831 17828 8840
rect 17588 8800 17788 8831
rect 18115 8800 18124 8840
rect 18164 8800 19220 8840
rect 17788 8782 17828 8791
rect 15715 8716 15724 8756
rect 15787 8716 15895 8756
rect 16012 8716 16108 8756
rect 16148 8716 16157 8756
rect 16444 8716 16876 8756
rect 16916 8716 17108 8756
rect 16012 8672 16052 8716
rect 12368 8656 12408 8665
rect 12451 8632 12460 8672
rect 12500 8632 13508 8672
rect 13565 8632 13603 8672
rect 13643 8632 13652 8672
rect 13699 8632 13708 8672
rect 13748 8632 13757 8672
rect 14633 8632 14764 8672
rect 14804 8632 14813 8672
rect 15031 8632 15040 8672
rect 15080 8632 15436 8672
rect 15476 8632 15485 8672
rect 15619 8632 15628 8672
rect 15668 8632 15677 8672
rect 15856 8632 15865 8672
rect 15905 8632 16052 8672
rect 16108 8632 16195 8672
rect 16235 8632 16244 8672
rect 16291 8643 16300 8683
rect 16340 8643 16349 8683
rect 16444 8672 16484 8716
rect 17068 8672 17108 8716
rect 17194 8747 17492 8756
rect 17194 8707 17203 8747
rect 17243 8716 17492 8747
rect 18019 8716 18028 8756
rect 18068 8716 18220 8756
rect 18260 8716 18269 8756
rect 18442 8747 18508 8756
rect 17243 8707 17252 8716
rect 17194 8706 17252 8707
rect 18442 8707 18451 8747
rect 18491 8716 18508 8747
rect 18548 8716 18631 8756
rect 18491 8707 18500 8716
rect 18442 8706 18500 8707
rect 18307 8672 18316 8693
rect 6892 8588 6932 8632
rect 8716 8588 8756 8632
rect 9772 8623 9812 8632
rect 11020 8588 11060 8632
rect 13468 8588 13508 8632
rect 13708 8588 13748 8632
rect 14764 8623 14804 8632
rect 16108 8588 16148 8632
rect 16300 8588 16340 8643
rect 16436 8632 16445 8672
rect 16485 8632 16494 8672
rect 16566 8632 16575 8672
rect 16615 8632 16628 8672
rect 16675 8632 16684 8672
rect 16753 8632 16855 8672
rect 17059 8632 17068 8672
rect 17108 8632 17117 8672
rect 17296 8632 17305 8672
rect 17345 8632 17396 8672
rect 17818 8632 17827 8672
rect 17867 8632 18315 8672
rect 18356 8653 18365 8693
rect 19180 8672 19220 8800
rect 19564 8756 19604 8884
rect 19843 8800 19852 8840
rect 19892 8800 20524 8840
rect 20564 8800 20573 8840
rect 21641 8800 21772 8840
rect 21812 8800 21821 8840
rect 23020 8800 24556 8840
rect 24596 8800 24605 8840
rect 23020 8756 23060 8800
rect 19564 8716 23060 8756
rect 23299 8716 23308 8756
rect 23348 8716 24404 8756
rect 24451 8716 24460 8756
rect 24500 8716 24542 8756
rect 18355 8632 18364 8653
rect 18544 8632 18553 8672
rect 18593 8632 18644 8672
rect 19171 8632 19180 8672
rect 19220 8632 19229 8672
rect 19450 8632 19459 8672
rect 19499 8632 19508 8672
rect 19555 8632 19564 8672
rect 19604 8632 20236 8672
rect 20276 8632 20285 8672
rect 20329 8632 20338 8672
rect 20378 8632 23404 8672
rect 23444 8632 23453 8672
rect 23779 8632 23788 8672
rect 23828 8632 23924 8672
rect 23971 8632 23980 8672
rect 24020 8632 24076 8672
rect 24116 8632 24151 8672
rect 16588 8588 16628 8632
rect 17356 8588 17396 8632
rect 18604 8588 18644 8632
rect 19468 8588 19508 8632
rect 23884 8588 23924 8632
rect 24364 8588 24404 8716
rect 24460 8672 24500 8716
rect 24652 8714 24692 9220
rect 26425 9052 26434 9092
rect 26802 9052 26811 9092
rect 27091 8884 27100 8924
rect 27140 8884 27532 8924
rect 27572 8884 27581 8924
rect 28841 8884 28972 8924
rect 29012 8884 29021 8924
rect 29923 8884 29932 8924
rect 29972 8884 29981 8924
rect 29932 8840 29972 8884
rect 24835 8800 24844 8840
rect 24884 8800 25996 8840
rect 26036 8800 26045 8840
rect 26441 8800 26572 8840
rect 26612 8800 26621 8840
rect 26668 8800 29972 8840
rect 30953 8800 30988 8840
rect 31028 8800 31084 8840
rect 31124 8800 31133 8840
rect 24634 8674 24643 8714
rect 24683 8674 24692 8714
rect 24844 8672 24884 8800
rect 26668 8756 26708 8800
rect 24931 8716 24940 8756
rect 24980 8716 26708 8756
rect 26764 8716 28876 8756
rect 28916 8716 28925 8756
rect 29993 8716 30034 8756
rect 30074 8716 30124 8756
rect 30164 8716 30173 8756
rect 26764 8672 26804 8716
rect 24446 8632 24455 8672
rect 24495 8632 24504 8672
rect 24835 8632 24844 8672
rect 24884 8632 24893 8672
rect 25036 8632 26804 8672
rect 26947 8632 26956 8672
rect 26996 8632 27127 8672
rect 27977 8632 28108 8672
rect 28148 8632 28157 8672
rect 29347 8632 29356 8672
rect 29396 8632 29644 8672
rect 29684 8632 29693 8672
rect 29827 8632 29836 8672
rect 29876 8632 30124 8672
rect 30164 8632 30173 8672
rect 30499 8632 30508 8672
rect 30587 8632 30679 8672
rect 5609 8548 5731 8588
rect 5780 8548 5789 8588
rect 6892 8548 6988 8588
rect 7028 8548 7037 8588
rect 8716 8548 8812 8588
rect 8852 8548 8916 8588
rect 11020 8548 12980 8588
rect 13468 8548 13748 8588
rect 13836 8548 13914 8588
rect 13954 8548 13996 8588
rect 14036 8548 14465 8588
rect 14505 8548 14514 8588
rect 15196 8548 16148 8588
rect 16291 8548 16300 8588
rect 16340 8548 16376 8588
rect 16588 8548 16876 8588
rect 16916 8548 16925 8588
rect 17155 8548 17164 8588
rect 17204 8548 17396 8588
rect 18019 8548 18028 8588
rect 18068 8548 18316 8588
rect 18356 8548 18365 8588
rect 18508 8548 18644 8588
rect 19075 8548 19084 8588
rect 19124 8548 19508 8588
rect 19555 8548 19564 8588
rect 19604 8548 19613 8588
rect 19747 8548 19756 8588
rect 19796 8548 20030 8588
rect 20070 8548 20079 8588
rect 23875 8548 23884 8588
rect 23924 8548 24055 8588
rect 24364 8548 24556 8588
rect 24596 8548 24605 8588
rect 0 8464 748 8504
rect 788 8464 797 8504
rect 2266 8464 2275 8504
rect 2315 8464 2708 8504
rect 3139 8464 3148 8504
rect 3188 8464 3860 8504
rect 4387 8464 4396 8504
rect 4436 8464 4700 8504
rect 7145 8464 7276 8504
rect 7316 8464 7325 8504
rect 0 8444 400 8464
rect 8716 8420 8756 8548
rect 11500 8504 11540 8548
rect 10313 8464 10444 8504
rect 10484 8464 10493 8504
rect 11491 8464 11500 8504
rect 11540 8464 11549 8504
rect 11980 8495 12212 8504
rect 11980 8464 12163 8495
rect 1795 8380 1804 8420
rect 1844 8380 8756 8420
rect 4343 8296 4352 8336
rect 4720 8296 4729 8336
rect 7468 8296 11924 8336
rect 1036 8212 3820 8252
rect 3860 8212 3869 8252
rect 0 8084 400 8104
rect 1036 8084 1076 8212
rect 7468 8168 7508 8296
rect 11884 8168 11924 8296
rect 11980 8252 12020 8464
rect 12154 8455 12163 8464
rect 12203 8455 12212 8495
rect 12154 8454 12212 8455
rect 12940 8420 12980 8548
rect 14284 8420 14324 8548
rect 15196 8504 15236 8548
rect 17356 8504 17396 8548
rect 18508 8504 18548 8548
rect 14371 8464 14380 8504
rect 14420 8464 14668 8504
rect 14708 8464 14717 8504
rect 15187 8464 15196 8504
rect 15236 8464 15245 8504
rect 16666 8464 16675 8504
rect 16715 8464 16724 8504
rect 16771 8464 16780 8504
rect 16820 8464 16972 8504
rect 17012 8464 17021 8504
rect 17356 8464 17836 8504
rect 17876 8464 18548 8504
rect 19564 8504 19604 8548
rect 19564 8464 19796 8504
rect 15196 8420 15236 8464
rect 12940 8380 13940 8420
rect 14284 8380 15236 8420
rect 16684 8420 16724 8464
rect 16684 8380 17068 8420
rect 17108 8380 17117 8420
rect 12117 8296 12126 8336
rect 12494 8296 12503 8336
rect 11980 8212 12308 8252
rect 12268 8168 12308 8212
rect 13900 8168 13940 8380
rect 17923 8296 17932 8336
rect 17972 8296 19276 8336
rect 19316 8296 19325 8336
rect 14947 8212 14956 8252
rect 14996 8212 18164 8252
rect 18403 8212 18412 8252
rect 18452 8212 18461 8252
rect 18124 8168 18164 8212
rect 18412 8168 18452 8212
rect 19756 8168 19796 8464
rect 23980 8420 24020 8548
rect 25036 8420 25076 8632
rect 28649 8464 28780 8504
rect 28820 8464 28829 8504
rect 30403 8464 30412 8504
rect 30452 8464 30748 8504
rect 30788 8464 30797 8504
rect 23980 8380 25076 8420
rect 19891 8296 19900 8336
rect 20268 8296 20277 8336
rect 27665 8296 27674 8336
rect 28042 8296 28051 8336
rect 19852 8212 25036 8252
rect 25076 8212 25460 8252
rect 19852 8168 19892 8212
rect 25420 8168 25460 8212
rect 2467 8128 2476 8168
rect 2516 8128 2764 8168
rect 2804 8128 2813 8168
rect 3226 8128 3235 8168
rect 3275 8128 3532 8168
rect 3572 8128 3581 8168
rect 4099 8128 4108 8168
rect 4148 8128 4195 8168
rect 4235 8128 4279 8168
rect 4483 8128 4492 8168
rect 4532 8128 4541 8168
rect 5033 8128 5164 8168
rect 5204 8128 5395 8168
rect 5435 8128 5444 8168
rect 6857 8128 6988 8168
rect 7028 8128 7037 8168
rect 7450 8128 7459 8168
rect 7499 8128 7508 8168
rect 11866 8128 11875 8168
rect 11915 8128 11924 8168
rect 12250 8128 12259 8168
rect 12299 8128 12308 8168
rect 12460 8128 13324 8168
rect 13364 8128 13373 8168
rect 13891 8128 13900 8168
rect 13940 8128 13949 8168
rect 16553 8128 16588 8168
rect 16628 8128 16684 8168
rect 16724 8128 16733 8168
rect 16867 8128 16876 8168
rect 16916 8128 17047 8168
rect 17347 8128 17356 8168
rect 17396 8128 18019 8168
rect 18059 8128 18068 8168
rect 18115 8128 18124 8168
rect 18164 8128 18295 8168
rect 18403 8128 18412 8168
rect 18452 8128 18499 8168
rect 19075 8128 19084 8168
rect 19124 8128 19363 8168
rect 19403 8128 19412 8168
rect 19459 8128 19468 8168
rect 19508 8128 19639 8168
rect 19738 8128 19747 8168
rect 19787 8128 19796 8168
rect 19843 8128 19852 8168
rect 19892 8128 19901 8168
rect 22051 8128 22060 8168
rect 22100 8128 23116 8168
rect 23156 8128 23165 8168
rect 25411 8128 25420 8168
rect 25460 8128 25469 8168
rect 27907 8128 27916 8168
rect 27956 8128 28108 8168
rect 28148 8128 28157 8168
rect 28780 8128 28876 8168
rect 28916 8128 28925 8168
rect 29155 8128 29164 8168
rect 29204 8128 29836 8168
rect 29876 8128 29885 8168
rect 29993 8128 30124 8168
rect 30164 8128 30173 8168
rect 4204 8084 4244 8128
rect 4492 8084 4532 8128
rect 0 8044 1076 8084
rect 1132 8044 2420 8084
rect 2467 8044 2476 8084
rect 2516 8044 2525 8084
rect 4204 8044 4436 8084
rect 4492 8044 5684 8084
rect 0 8024 400 8044
rect 1132 8000 1172 8044
rect 2380 8000 2420 8044
rect 2476 8000 2516 8044
rect 4396 8000 4436 8044
rect 931 7960 940 8000
rect 980 7960 989 8000
rect 1123 7960 1132 8000
rect 1172 7960 1181 8000
rect 1498 7960 1507 8000
rect 1547 7960 1556 8000
rect 1603 7960 1612 8000
rect 1652 7960 1748 8000
rect 2249 7960 2380 8000
rect 2420 7960 2429 8000
rect 2476 7960 2564 8000
rect 0 7664 400 7684
rect 940 7664 980 7960
rect 1516 7916 1556 7960
rect 1507 7876 1516 7916
rect 1556 7876 1603 7916
rect 1708 7832 1748 7960
rect 2524 7958 2564 7960
rect 2668 7960 2903 8000
rect 2943 7960 2952 8000
rect 3043 7960 3052 8000
rect 3092 7960 3148 8000
rect 3188 7960 3223 8000
rect 4291 7960 4300 8000
rect 4340 7960 4349 8000
rect 4396 7960 4684 8000
rect 4724 7960 4733 8000
rect 5059 7960 5068 8000
rect 5108 7960 5348 8000
rect 5417 7960 5539 8000
rect 5588 7960 5597 8000
rect 5644 7991 5684 8044
rect 6604 8044 6892 8084
rect 6932 8044 7276 8084
rect 7316 8044 7325 8084
rect 7372 8044 7756 8084
rect 7796 8044 7805 8084
rect 12081 8044 12090 8084
rect 12130 8044 12364 8084
rect 12404 8044 12413 8084
rect 6604 8000 6644 8044
rect 7372 8000 7412 8044
rect 12460 8000 12500 8128
rect 12547 8044 12556 8084
rect 12596 8044 12980 8084
rect 12940 8000 12980 8044
rect 16684 8044 17356 8084
rect 17396 8044 17405 8084
rect 17801 8044 17921 8084
rect 17972 8044 17981 8084
rect 18220 8044 21428 8084
rect 16684 8000 16724 8044
rect 2524 7918 2563 7958
rect 2603 7918 2612 7958
rect 1027 7792 1036 7832
rect 1076 7792 1708 7832
rect 1748 7792 1757 7832
rect 2668 7748 2708 7960
rect 4300 7916 4340 7960
rect 5308 7916 5348 7960
rect 6586 7960 6595 8000
rect 6635 7960 6644 8000
rect 6691 7960 6700 8000
rect 6740 7960 6871 8000
rect 7075 7960 7084 8000
rect 7124 7960 7127 8000
rect 7167 7960 7255 8000
rect 7363 7960 7372 8000
rect 7412 7960 7421 8000
rect 7651 7960 7660 8000
rect 7700 7960 7709 8000
rect 7843 7960 7852 8000
rect 7892 7960 8908 8000
rect 8948 7960 8957 8000
rect 9571 7960 9580 8000
rect 9620 7960 9676 8000
rect 9716 7960 9751 8000
rect 11770 7960 11779 8000
rect 11819 7960 11828 8000
rect 11875 7960 11884 8000
rect 11924 7960 11933 8000
rect 12436 7960 12445 8000
rect 12485 7960 12500 8000
rect 12547 7960 12556 8000
rect 12596 7960 12605 8000
rect 12940 7960 13036 8000
rect 13076 7960 13085 8000
rect 5644 7942 5684 7951
rect 3034 7876 3043 7916
rect 3083 7876 3092 7916
rect 4300 7876 5348 7916
rect 3052 7832 3092 7876
rect 3052 7792 3532 7832
rect 3572 7792 3581 7832
rect 5308 7748 5348 7876
rect 6604 7832 6644 7960
rect 7660 7916 7700 7960
rect 7258 7876 7267 7916
rect 7307 7876 7316 7916
rect 7363 7876 7372 7916
rect 7412 7876 7700 7916
rect 7276 7832 7316 7876
rect 11788 7832 11828 7960
rect 11884 7916 11924 7960
rect 12556 7916 12596 7960
rect 13169 7928 13178 7968
rect 13218 7928 13240 7968
rect 13961 7960 14092 8000
rect 14132 7960 14141 8000
rect 14659 7960 14668 8000
rect 14708 7960 14717 8000
rect 14851 7960 14860 8000
rect 14900 7960 15628 8000
rect 15668 7960 15677 8000
rect 16099 7960 16108 8000
rect 16148 7960 16492 8000
rect 16532 7960 16541 8000
rect 16666 7960 16675 8000
rect 16715 7960 16724 8000
rect 16867 7960 16876 8000
rect 16916 7960 16925 8000
rect 17059 7960 17068 8000
rect 17108 7960 17260 8000
rect 17300 7960 17309 8000
rect 17443 7960 17452 8000
rect 17492 7960 17501 8000
rect 18220 7991 18260 8044
rect 11884 7876 12596 7916
rect 13200 7832 13240 7928
rect 14668 7916 14708 7960
rect 16876 7916 16916 7960
rect 17459 7916 17499 7960
rect 18403 7960 18412 8000
rect 18452 7960 18508 8000
rect 18548 7960 18583 8000
rect 19256 7960 19265 8000
rect 19316 7960 19436 8000
rect 19564 7991 19604 8000
rect 18220 7942 18260 7951
rect 18739 7918 18748 7958
rect 18788 7918 18797 7958
rect 20035 7960 20044 8000
rect 20084 7960 20428 8000
rect 20468 7960 20477 8000
rect 14668 7876 15148 7916
rect 15188 7876 15197 7916
rect 15331 7876 15340 7916
rect 15380 7876 17499 7916
rect 18496 7876 18604 7916
rect 18667 7876 18676 7916
rect 5923 7792 5932 7832
rect 5972 7792 6644 7832
rect 7267 7792 7276 7832
rect 7316 7792 7363 7832
rect 11788 7792 12748 7832
rect 12788 7792 13240 7832
rect 17459 7832 17499 7876
rect 18754 7832 18794 7918
rect 19564 7916 19604 7951
rect 19459 7876 19468 7916
rect 19508 7876 19604 7916
rect 19945 7876 19954 7916
rect 19994 7876 20564 7916
rect 17459 7792 18220 7832
rect 18260 7792 18269 7832
rect 18403 7792 18412 7832
rect 18452 7792 18794 7832
rect 1786 7708 1795 7748
rect 1835 7708 2764 7748
rect 2804 7708 2813 7748
rect 5308 7708 7084 7748
rect 7124 7708 7133 7748
rect 9427 7708 9436 7748
rect 9476 7708 9484 7748
rect 9524 7708 9607 7748
rect 12067 7708 12076 7748
rect 12116 7708 12980 7748
rect 14755 7708 14764 7748
rect 14804 7708 14956 7748
rect 14996 7708 15005 7748
rect 12940 7664 12980 7708
rect 0 7624 460 7664
rect 500 7624 509 7664
rect 940 7624 1804 7664
rect 1844 7624 1853 7664
rect 12940 7624 14284 7664
rect 14324 7624 14333 7664
rect 0 7604 400 7624
rect 3103 7540 3112 7580
rect 3480 7540 3489 7580
rect 10877 7540 10886 7580
rect 11254 7540 11263 7580
rect 18651 7540 18660 7580
rect 19028 7540 19037 7580
rect 748 7456 1612 7496
rect 1652 7456 1661 7496
rect 17059 7456 17068 7496
rect 17108 7456 19652 7496
rect 0 7244 400 7264
rect 748 7244 788 7456
rect 1385 7372 1507 7412
rect 1556 7372 1565 7412
rect 2947 7372 2956 7412
rect 2996 7372 3148 7412
rect 3188 7372 3197 7412
rect 4099 7372 4108 7412
rect 4148 7372 4972 7412
rect 5012 7372 5021 7412
rect 6874 7372 6883 7412
rect 6923 7372 7276 7412
rect 7316 7372 7325 7412
rect 7852 7372 8852 7412
rect 8899 7372 8908 7412
rect 8948 7372 9964 7412
rect 10004 7372 10013 7412
rect 11971 7372 11980 7412
rect 12020 7372 12364 7412
rect 12404 7372 12413 7412
rect 12617 7372 12739 7412
rect 12788 7372 12797 7412
rect 14746 7372 14755 7412
rect 14795 7372 15724 7412
rect 15764 7372 15773 7412
rect 18211 7372 18220 7412
rect 18260 7372 18412 7412
rect 18452 7372 18461 7412
rect 0 7204 788 7244
rect 1516 7244 1556 7372
rect 2092 7288 7124 7328
rect 2092 7244 2132 7288
rect 7084 7244 7124 7288
rect 1516 7204 1891 7244
rect 1931 7204 1940 7244
rect 2083 7204 2092 7244
rect 2132 7204 2141 7244
rect 2755 7204 2764 7244
rect 2804 7204 2996 7244
rect 4361 7235 4492 7244
rect 4361 7204 4435 7235
rect 0 7184 400 7204
rect 2956 7160 2996 7204
rect 4426 7195 4435 7204
rect 4475 7204 4492 7235
rect 4532 7204 4541 7244
rect 4748 7204 4780 7244
rect 4820 7204 4829 7244
rect 7084 7204 7220 7244
rect 4475 7195 4484 7204
rect 4426 7194 4484 7195
rect 4748 7193 4788 7204
rect 1210 7120 1219 7160
rect 1259 7120 1268 7160
rect 1315 7120 1324 7160
rect 1364 7120 1516 7160
rect 1556 7120 1565 7160
rect 1699 7120 1708 7160
rect 1748 7120 1751 7160
rect 1791 7120 1879 7160
rect 1987 7120 1996 7160
rect 2036 7120 2045 7160
rect 2179 7120 2188 7160
rect 2228 7120 2284 7160
rect 2324 7120 2359 7160
rect 2467 7120 2476 7160
rect 2516 7120 2525 7160
rect 2668 7120 2851 7160
rect 2891 7120 2900 7160
rect 2947 7120 2956 7160
rect 2996 7120 3005 7160
rect 3052 7120 3532 7160
rect 3572 7120 3581 7160
rect 4099 7120 4108 7160
rect 4148 7120 4300 7160
rect 4340 7120 4349 7160
rect 4525 7120 4534 7160
rect 4574 7120 4583 7160
rect 4677 7153 4686 7193
rect 4726 7153 4788 7193
rect 7180 7160 7220 7204
rect 7852 7160 7892 7372
rect 8122 7288 8131 7328
rect 8171 7288 8180 7328
rect 8140 7244 8180 7288
rect 8812 7244 8852 7372
rect 19612 7328 19652 7456
rect 20524 7412 20564 7876
rect 20297 7372 20419 7412
rect 20468 7372 20477 7412
rect 20524 7372 21292 7412
rect 21332 7372 21341 7412
rect 21388 7328 21428 8044
rect 21772 8044 22828 8084
rect 22868 8044 22877 8084
rect 23098 8044 23107 8084
rect 23147 8044 23788 8084
rect 23828 8044 23837 8084
rect 25594 8044 25603 8084
rect 25643 8044 26860 8084
rect 26900 8044 26909 8084
rect 21772 8000 21812 8044
rect 28780 8000 28820 8128
rect 28876 8044 29932 8084
rect 29972 8044 30644 8084
rect 28876 8000 28916 8044
rect 30604 8000 30644 8044
rect 21545 7960 21676 8000
rect 21716 7960 21725 8000
rect 21772 7991 21827 8000
rect 21772 7960 21787 7991
rect 21676 7942 21716 7951
rect 21787 7942 21827 7951
rect 21898 7991 21964 8000
rect 21898 7951 21907 7991
rect 21947 7960 21964 7991
rect 22004 7960 22339 8000
rect 22379 7960 22388 8000
rect 22627 7960 22636 8000
rect 22676 7960 22732 8000
rect 22772 7960 22807 8000
rect 23482 7960 23491 8000
rect 23531 7960 23980 8000
rect 24020 7960 24029 8000
rect 25978 7960 25987 8000
rect 26036 7960 26167 8000
rect 28762 7960 28771 8000
rect 28811 7960 28820 8000
rect 28867 7960 28876 8000
rect 28916 7960 28925 8000
rect 29722 7960 29731 8000
rect 29771 7960 29780 8000
rect 29829 7960 29838 8000
rect 29878 7960 30028 8000
rect 30068 7960 30077 8000
rect 30307 7960 30316 8000
rect 30356 7960 30499 8000
rect 30539 7960 30548 8000
rect 30595 7960 30604 8000
rect 30644 7960 30653 8000
rect 21947 7951 21956 7960
rect 21898 7950 21956 7951
rect 29740 7916 29780 7960
rect 24643 7876 24652 7916
rect 24692 7876 24701 7916
rect 26563 7876 26572 7916
rect 26612 7876 26621 7916
rect 27523 7876 27532 7916
rect 27572 7876 28396 7916
rect 28436 7876 28445 7916
rect 29740 7876 29836 7916
rect 29876 7876 29885 7916
rect 30953 7792 31084 7832
rect 31124 7792 31133 7832
rect 21475 7708 21484 7748
rect 21524 7708 25036 7748
rect 25076 7708 25085 7748
rect 30569 7708 30604 7748
rect 30644 7708 30700 7748
rect 30740 7708 30749 7748
rect 26425 7540 26434 7580
rect 26802 7540 26811 7580
rect 21475 7372 21484 7412
rect 21524 7372 22060 7412
rect 22100 7372 22109 7412
rect 23491 7372 23500 7412
rect 23540 7372 28396 7412
rect 28436 7372 29031 7412
rect 30019 7372 30028 7412
rect 30068 7372 30508 7412
rect 30548 7372 30557 7412
rect 9475 7288 9484 7328
rect 9524 7288 10411 7328
rect 19450 7288 19459 7328
rect 19499 7288 19508 7328
rect 19603 7288 19612 7328
rect 19652 7288 20756 7328
rect 21388 7288 23060 7328
rect 24521 7288 24652 7328
rect 24692 7288 24701 7328
rect 28745 7288 28876 7328
rect 28916 7288 28925 7328
rect 8105 7204 8236 7244
rect 8276 7204 8564 7244
rect 8812 7204 8908 7244
rect 8948 7204 8957 7244
rect 9475 7204 9484 7244
rect 9524 7204 9533 7244
rect 8524 7160 8564 7204
rect 4963 7120 4972 7160
rect 5023 7120 5143 7160
rect 6569 7120 6700 7160
rect 6740 7120 6749 7160
rect 6874 7120 6883 7160
rect 6932 7120 7063 7160
rect 7180 7120 7843 7160
rect 7883 7120 7892 7160
rect 7939 7120 7948 7160
rect 7988 7120 7997 7160
rect 8131 7120 8140 7160
rect 8180 7120 8375 7160
rect 8415 7120 8424 7160
rect 8506 7120 8515 7160
rect 8555 7120 8564 7160
rect 8611 7120 8620 7160
rect 8660 7120 8791 7160
rect 9082 7120 9091 7160
rect 9131 7120 9140 7160
rect 1228 7076 1268 7120
rect 1996 7076 2036 7120
rect 1181 7036 1228 7076
rect 1268 7036 1277 7076
rect 1996 7036 2380 7076
rect 2420 7036 2429 7076
rect 1228 6908 1268 7036
rect 1507 6952 1516 6992
rect 1556 6952 1996 6992
rect 2036 6952 2188 6992
rect 2228 6952 2237 6992
rect 2476 6908 2516 7120
rect 1228 6868 2516 6908
rect 0 6824 400 6844
rect 0 6784 1900 6824
rect 1940 6784 1949 6824
rect 0 6764 400 6784
rect 2668 6656 2708 7120
rect 2860 7076 2900 7120
rect 3052 7076 3092 7120
rect 4531 7076 4571 7120
rect 7948 7076 7988 7120
rect 9100 7076 9140 7120
rect 2860 7036 3092 7076
rect 3148 7036 3159 7076
rect 3199 7036 3208 7076
rect 4003 7036 4012 7076
rect 4052 7036 4204 7076
rect 4244 7036 4253 7076
rect 4531 7036 4820 7076
rect 3148 6992 3188 7036
rect 4780 6992 4820 7036
rect 2851 6952 2860 6992
rect 2900 6952 3188 6992
rect 4762 6952 4771 6992
rect 4811 6952 4820 6992
rect 4343 6784 4352 6824
rect 4720 6784 4729 6824
rect 4780 6740 4820 6952
rect 7468 7036 9140 7076
rect 9257 7036 9388 7076
rect 9428 7036 9437 7076
rect 2755 6700 2764 6740
rect 2804 6700 3532 6740
rect 3572 6700 3581 6740
rect 3820 6700 4628 6740
rect 1891 6616 1900 6656
rect 1940 6616 1949 6656
rect 2179 6616 2188 6656
rect 2228 6616 2237 6656
rect 2659 6616 2668 6656
rect 2708 6616 2717 6656
rect 1900 6488 1940 6616
rect 2188 6572 2228 6616
rect 3820 6572 3860 6700
rect 3907 6616 3916 6656
rect 3956 6616 3965 6656
rect 2188 6532 2996 6572
rect 2956 6488 2996 6532
rect 3148 6532 3628 6572
rect 3668 6532 3860 6572
rect 3148 6488 3188 6532
rect 3916 6488 3956 6616
rect 4588 6572 4628 6700
rect 4684 6700 4820 6740
rect 4963 6700 4972 6740
rect 5012 6700 6751 6740
rect 4684 6656 4724 6700
rect 4675 6616 4684 6656
rect 4724 6616 4733 6656
rect 6089 6616 6211 6656
rect 6260 6616 6269 6656
rect 6711 6572 6751 6700
rect 7468 6656 7508 7036
rect 8585 6952 8707 6992
rect 8756 6952 8765 6992
rect 9484 6656 9524 7204
rect 10147 7162 10156 7202
rect 10196 7162 10327 7202
rect 10036 7120 10045 7160
rect 10085 7120 10100 7160
rect 10156 7144 10196 7153
rect 10371 7160 10411 7288
rect 12460 7244 12499 7272
rect 11116 7204 11348 7244
rect 11116 7160 11156 7204
rect 10371 7120 10967 7160
rect 11007 7120 11016 7160
rect 11098 7120 11107 7160
rect 11147 7120 11156 7160
rect 11203 7120 11212 7160
rect 11252 7120 11261 7160
rect 7459 6616 7468 6656
rect 7508 6616 7517 6656
rect 8026 6616 8035 6656
rect 8075 6616 8620 6656
rect 8660 6616 8669 6656
rect 9283 6616 9292 6656
rect 9332 6616 9524 6656
rect 10060 6656 10100 7120
rect 11212 7076 11252 7120
rect 11020 7036 11252 7076
rect 11308 7076 11348 7204
rect 12172 7232 12499 7244
rect 12539 7232 12548 7272
rect 19468 7244 19508 7288
rect 12172 7204 12500 7232
rect 12940 7204 13556 7244
rect 14275 7204 14284 7244
rect 14324 7204 14612 7244
rect 12172 7160 12212 7204
rect 11779 7120 11788 7160
rect 11828 7120 12172 7160
rect 12212 7120 12221 7160
rect 12425 7120 12547 7160
rect 12596 7120 12605 7160
rect 12940 7076 12980 7204
rect 13027 7120 13036 7160
rect 13076 7120 13228 7160
rect 13268 7120 13277 7160
rect 13414 7120 13423 7160
rect 13463 7120 13474 7160
rect 13434 7076 13474 7120
rect 11308 7036 12980 7076
rect 13389 7036 13420 7076
rect 13460 7036 13474 7076
rect 11020 6656 11060 7036
rect 11290 6952 11299 6992
rect 11339 6952 11788 6992
rect 11828 6952 11837 6992
rect 12250 6952 12259 6992
rect 12299 6952 12556 6992
rect 12596 6952 12605 6992
rect 13402 6952 13411 6992
rect 13451 6952 13460 6992
rect 12117 6784 12126 6824
rect 12494 6784 12503 6824
rect 10060 6616 10156 6656
rect 10196 6616 10205 6656
rect 10819 6616 10828 6656
rect 10868 6616 11060 6656
rect 11884 6616 12547 6656
rect 12587 6616 12596 6656
rect 10156 6572 10196 6616
rect 4588 6532 5108 6572
rect 5068 6488 5108 6532
rect 6124 6532 6604 6572
rect 6644 6532 6653 6572
rect 6702 6532 6711 6572
rect 6751 6532 7412 6572
rect 8009 6532 8140 6572
rect 8180 6532 8189 6572
rect 8995 6532 9004 6572
rect 9044 6532 10060 6572
rect 10100 6532 10109 6572
rect 10156 6532 10676 6572
rect 6124 6488 6164 6532
rect 7372 6488 7412 6532
rect 10060 6488 10100 6532
rect 10636 6488 10676 6532
rect 11884 6488 11924 6616
rect 12748 6532 12940 6572
rect 12980 6532 12989 6572
rect 12748 6488 12788 6532
rect 13420 6488 13460 6952
rect 13516 6908 13556 7204
rect 14572 7160 14612 7204
rect 18028 7204 18499 7244
rect 18539 7204 18548 7244
rect 18691 7204 18700 7244
rect 18740 7204 19084 7244
rect 19124 7204 19133 7244
rect 19468 7204 20372 7244
rect 18028 7160 18068 7204
rect 20332 7160 20372 7204
rect 20716 7160 20756 7288
rect 23020 7244 23060 7288
rect 22156 7204 22388 7244
rect 23020 7204 26764 7244
rect 26804 7204 26813 7244
rect 27523 7204 27532 7244
rect 27611 7204 27703 7244
rect 28771 7204 28780 7244
rect 28820 7204 28829 7244
rect 22156 7160 22196 7204
rect 22348 7160 22388 7204
rect 28780 7160 28820 7204
rect 28991 7160 29031 7372
rect 29609 7288 29644 7328
rect 29684 7288 29740 7328
rect 29780 7288 29972 7328
rect 29932 7244 29972 7288
rect 29914 7204 29923 7244
rect 29963 7204 29972 7244
rect 30115 7204 30124 7244
rect 30164 7204 30316 7244
rect 30356 7204 30365 7244
rect 30595 7204 30604 7244
rect 30650 7204 30775 7244
rect 29588 7193 29636 7202
rect 14458 7120 14467 7160
rect 14507 7120 14516 7160
rect 14563 7120 14572 7160
rect 14612 7120 14621 7160
rect 15065 7120 15148 7160
rect 15188 7120 15196 7160
rect 15236 7120 15245 7160
rect 15331 7120 15340 7160
rect 15380 7120 15628 7160
rect 15668 7120 15677 7160
rect 17923 7120 17932 7160
rect 17972 7120 18013 7160
rect 18053 7120 18103 7160
rect 18350 7120 18359 7160
rect 18399 7120 18408 7160
rect 18595 7120 18604 7160
rect 18644 7120 18775 7160
rect 19267 7120 19276 7160
rect 19316 7120 19325 7160
rect 19450 7120 19459 7160
rect 19499 7120 19948 7160
rect 19988 7120 20044 7160
rect 20084 7120 20093 7160
rect 20227 7120 20236 7160
rect 20276 7120 20285 7160
rect 20332 7120 20414 7160
rect 20454 7120 20463 7160
rect 21209 7120 21292 7160
rect 21332 7120 21340 7160
rect 21380 7120 21389 7160
rect 21475 7120 21484 7160
rect 21524 7120 21655 7160
rect 22132 7120 22141 7160
rect 22181 7120 22196 7160
rect 22243 7120 22252 7160
rect 22292 7120 22301 7160
rect 22348 7120 23060 7160
rect 23107 7120 23116 7160
rect 23156 7120 23308 7160
rect 23348 7120 23357 7160
rect 23491 7120 23500 7160
rect 23540 7120 23671 7160
rect 23767 7120 23776 7160
rect 23816 7120 23825 7160
rect 24259 7120 24268 7160
rect 24308 7120 24788 7160
rect 24905 7120 25024 7160
rect 25076 7120 25085 7160
rect 25132 7120 25180 7160
rect 25220 7120 26284 7160
rect 26324 7120 26333 7160
rect 27757 7120 27766 7160
rect 27806 7120 28108 7160
rect 28148 7120 28157 7160
rect 28579 7120 28588 7160
rect 28628 7120 28820 7160
rect 28867 7120 28876 7160
rect 28916 7120 28925 7160
rect 28982 7120 28991 7160
rect 29031 7120 29040 7160
rect 29155 7120 29164 7160
rect 29204 7120 29213 7160
rect 29347 7120 29356 7160
rect 29396 7120 29405 7160
rect 29469 7120 29478 7160
rect 29518 7120 29527 7160
rect 29588 7153 29596 7193
rect 29636 7160 29684 7193
rect 29636 7153 29644 7160
rect 29596 7144 29644 7153
rect 29635 7120 29644 7144
rect 29684 7120 29709 7160
rect 29774 7120 29783 7160
rect 29823 7120 29832 7160
rect 30019 7120 30028 7160
rect 30068 7120 30199 7160
rect 30691 7120 30700 7160
rect 30740 7120 30871 7160
rect 14476 7076 14516 7120
rect 18359 7076 18399 7120
rect 19276 7076 19316 7120
rect 20236 7076 20276 7120
rect 20716 7111 20756 7120
rect 14476 7036 14860 7076
rect 14900 7036 15092 7076
rect 15052 6992 15092 7036
rect 18125 7036 18399 7076
rect 18508 7036 19220 7076
rect 19276 7036 20524 7076
rect 20564 7036 20573 7076
rect 18125 6992 18165 7036
rect 18508 6992 18548 7036
rect 15034 6952 15043 6992
rect 15083 6952 15092 6992
rect 17914 6952 17923 6992
rect 17963 6952 18165 6992
rect 18403 6952 18412 6992
rect 18452 6952 18548 6992
rect 13516 6868 17932 6908
rect 17972 6868 17981 6908
rect 16204 6700 17786 6740
rect 16204 6656 16244 6700
rect 13507 6616 13516 6656
rect 13556 6616 15148 6656
rect 15188 6616 15197 6656
rect 15820 6616 16204 6656
rect 16244 6616 16253 6656
rect 16841 6616 16972 6656
rect 17012 6616 17021 6656
rect 13708 6532 14092 6572
rect 14132 6532 14141 6572
rect 15034 6532 15043 6572
rect 15083 6532 15340 6572
rect 15380 6532 15389 6572
rect 13708 6488 13748 6532
rect 15820 6488 15860 6616
rect 15916 6532 17492 6572
rect 15916 6488 15956 6532
rect 17452 6488 17492 6532
rect 17746 6488 17786 6700
rect 18125 6656 18165 6952
rect 19180 6908 19220 7036
rect 22252 6992 22292 7120
rect 23020 7076 23060 7120
rect 23785 7076 23825 7120
rect 24748 7076 24788 7120
rect 25132 7076 25172 7120
rect 28876 7076 28916 7120
rect 23020 7036 23203 7076
rect 23243 7036 23252 7076
rect 23785 7036 24364 7076
rect 24404 7036 24413 7076
rect 24748 7036 25172 7076
rect 28073 7036 28195 7076
rect 28244 7036 28253 7076
rect 28771 7036 28780 7076
rect 28820 7036 28916 7076
rect 29164 7076 29204 7120
rect 29164 7036 29260 7076
rect 29300 7036 29309 7076
rect 29356 6992 29396 7120
rect 29487 7076 29527 7120
rect 29783 7076 29823 7120
rect 29487 7036 29548 7076
rect 29588 7036 29597 7076
rect 29783 7036 30124 7076
rect 30164 7036 30173 7076
rect 20489 6952 20620 6992
rect 20660 6952 20669 6992
rect 22252 6952 23212 6992
rect 23252 6952 23261 6992
rect 23340 6952 23404 6992
rect 23444 6952 23500 6992
rect 23540 6952 23596 6992
rect 23636 6952 23645 6992
rect 23849 6952 23932 6992
rect 23972 6952 23980 6992
rect 24020 6952 24029 6992
rect 24259 6952 24268 6992
rect 24308 6952 24364 6992
rect 24404 6952 24439 6992
rect 29155 6952 29164 6992
rect 29204 6952 29396 6992
rect 24268 6908 24308 6952
rect 19180 6868 23732 6908
rect 23875 6868 23884 6908
rect 23924 6868 24308 6908
rect 19891 6784 19900 6824
rect 20268 6784 20277 6824
rect 21772 6784 23596 6824
rect 23636 6784 23645 6824
rect 18211 6700 18220 6740
rect 18260 6700 20180 6740
rect 20515 6700 20524 6740
rect 20564 6700 21620 6740
rect 20140 6656 20180 6700
rect 21580 6656 21620 6700
rect 18125 6616 18211 6656
rect 18251 6616 18260 6656
rect 20140 6616 20620 6656
rect 20660 6616 20669 6656
rect 21562 6616 21571 6656
rect 21611 6616 21620 6656
rect 21772 6572 21812 6784
rect 23692 6656 23732 6868
rect 27665 6784 27674 6824
rect 28042 6784 28051 6824
rect 22409 6616 22492 6656
rect 22532 6616 22540 6656
rect 22580 6616 22589 6656
rect 23491 6616 23500 6656
rect 23540 6616 23549 6656
rect 23674 6616 23683 6656
rect 23723 6616 23732 6656
rect 26633 6616 26755 6656
rect 26804 6616 26813 6656
rect 28771 6616 28780 6656
rect 28820 6616 29539 6656
rect 29588 6616 29597 6656
rect 23500 6572 23540 6616
rect 17923 6532 17932 6572
rect 17972 6532 21812 6572
rect 23116 6532 23404 6572
rect 23444 6532 23453 6572
rect 23500 6532 24020 6572
rect 23116 6488 23156 6532
rect 23980 6488 24020 6532
rect 25228 6532 26132 6572
rect 28387 6532 28396 6572
rect 28436 6532 28959 6572
rect 29155 6532 29164 6572
rect 29204 6532 29251 6572
rect 29291 6532 29335 6572
rect 29443 6532 29452 6572
rect 29492 6532 29751 6572
rect 29791 6532 29800 6572
rect 25228 6488 25268 6532
rect 26092 6488 26132 6532
rect 28396 6488 28436 6532
rect 28919 6488 28959 6532
rect 29260 6488 29300 6532
rect 1498 6448 1507 6488
rect 1547 6448 1556 6488
rect 1603 6448 1612 6488
rect 1652 6448 1783 6488
rect 1900 6448 2188 6488
rect 2228 6448 2237 6488
rect 2345 6448 2476 6488
rect 2516 6448 2900 6488
rect 2947 6448 2956 6488
rect 2996 6448 3005 6488
rect 3139 6448 3148 6488
rect 3188 6448 3197 6488
rect 3514 6448 3523 6488
rect 3563 6448 3572 6488
rect 3619 6448 3628 6488
rect 3668 6448 3677 6488
rect 3916 6448 4204 6488
rect 4244 6448 4291 6488
rect 4331 6448 4340 6488
rect 4387 6448 4396 6488
rect 4436 6448 4567 6488
rect 4867 6448 4876 6488
rect 4916 6448 4925 6488
rect 5059 6448 5068 6488
rect 5108 6448 5117 6488
rect 6115 6448 6124 6488
rect 6164 6448 6173 6488
rect 6394 6448 6403 6488
rect 6443 6448 6452 6488
rect 6499 6448 6508 6488
rect 6548 6448 6557 6488
rect 6979 6448 6988 6488
rect 7028 6448 7037 6488
rect 7084 6448 7276 6488
rect 7316 6448 7325 6488
rect 7372 6448 7934 6488
rect 7974 6448 7983 6488
rect 8105 6448 8236 6488
rect 8276 6448 8285 6488
rect 9065 6448 9196 6488
rect 9236 6448 9245 6488
rect 9353 6448 9388 6488
rect 9428 6448 9484 6488
rect 9524 6448 9533 6488
rect 9667 6448 9676 6488
rect 9716 6448 9847 6488
rect 9955 6448 9964 6488
rect 10004 6448 10013 6488
rect 10060 6448 10540 6488
rect 10580 6448 10589 6488
rect 10636 6448 10679 6488
rect 10719 6448 10728 6488
rect 11866 6448 11875 6488
rect 11915 6448 11924 6488
rect 11971 6448 11980 6488
rect 12020 6448 12151 6488
rect 12739 6448 12748 6488
rect 12788 6448 12797 6488
rect 13027 6448 13036 6488
rect 13076 6448 13085 6488
rect 13420 6448 13612 6488
rect 13652 6448 13661 6488
rect 13708 6448 13731 6488
rect 13771 6448 13780 6488
rect 13840 6448 13849 6488
rect 13889 6448 13940 6488
rect 13987 6448 13996 6488
rect 14036 6448 14045 6488
rect 14170 6448 14179 6488
rect 14219 6448 14228 6488
rect 14275 6448 14284 6488
rect 14324 6448 14711 6488
rect 14751 6448 14760 6488
rect 14947 6448 14956 6488
rect 14996 6448 15127 6488
rect 15802 6448 15811 6488
rect 15851 6448 15860 6488
rect 15907 6448 15916 6488
rect 15956 6448 15965 6488
rect 16387 6448 16396 6488
rect 16436 6448 16673 6488
rect 16713 6448 16722 6488
rect 16810 6448 16819 6488
rect 16859 6448 16905 6488
rect 17417 6448 17443 6488
rect 17483 6448 17548 6488
rect 17588 6448 17597 6488
rect 17731 6448 17740 6488
rect 17780 6448 17789 6488
rect 18115 6448 18124 6488
rect 18165 6448 18295 6488
rect 19049 6448 19084 6488
rect 19124 6448 19180 6488
rect 19220 6448 19229 6488
rect 20201 6448 20323 6488
rect 20372 6448 20381 6488
rect 21763 6448 21772 6488
rect 21812 6448 21821 6488
rect 21929 6448 22060 6488
rect 22100 6448 22109 6488
rect 22217 6448 22348 6488
rect 22388 6448 22397 6488
rect 23098 6448 23107 6488
rect 23147 6448 23156 6488
rect 23203 6448 23212 6488
rect 23252 6448 23500 6488
rect 23540 6448 23549 6488
rect 23971 6448 23980 6488
rect 24020 6448 24029 6488
rect 25097 6448 25219 6488
rect 25268 6448 25277 6488
rect 25324 6448 25948 6488
rect 25988 6448 25997 6488
rect 26083 6448 26092 6488
rect 26132 6448 26141 6488
rect 27043 6448 27052 6488
rect 27092 6448 27476 6488
rect 27689 6448 27820 6488
rect 27860 6448 27869 6488
rect 28012 6448 28060 6488
rect 28100 6448 28109 6488
rect 28169 6448 28300 6488
rect 28340 6448 28349 6488
rect 28396 6448 28444 6488
rect 28484 6448 28493 6488
rect 28579 6448 28588 6488
rect 28628 6448 28780 6488
rect 28820 6448 28829 6488
rect 28910 6448 28919 6488
rect 28959 6448 28968 6488
rect 29155 6448 29164 6488
rect 29204 6448 29213 6488
rect 29260 6448 29443 6488
rect 29483 6448 29492 6488
rect 30595 6448 30604 6488
rect 30644 6448 30775 6488
rect 0 6404 400 6424
rect 1516 6404 1556 6448
rect 2860 6404 2900 6448
rect 3532 6404 3572 6448
rect 3628 6404 3668 6448
rect 0 6364 556 6404
rect 596 6364 605 6404
rect 1516 6364 2284 6404
rect 2324 6364 2764 6404
rect 2804 6364 2813 6404
rect 2860 6364 3052 6404
rect 3092 6364 3101 6404
rect 3485 6364 3532 6404
rect 3572 6364 3581 6404
rect 3628 6364 3916 6404
rect 3956 6364 3965 6404
rect 0 6344 400 6364
rect 4876 6320 4916 6448
rect 5875 6406 5884 6446
rect 5924 6406 5933 6446
rect 5884 6320 5924 6406
rect 6412 6404 6452 6448
rect 6010 6364 6019 6404
rect 6068 6364 6452 6404
rect 6508 6320 6548 6448
rect 6988 6320 7028 6448
rect 7084 6404 7124 6448
rect 8236 6430 8276 6439
rect 7075 6364 7084 6404
rect 7124 6364 7133 6404
rect 9676 6320 9716 6448
rect 9964 6404 10004 6448
rect 9964 6364 11500 6404
rect 11540 6364 11549 6404
rect 13036 6320 13076 6448
rect 13900 6404 13940 6448
rect 13891 6364 13900 6404
rect 13940 6364 13949 6404
rect 13996 6320 14036 6448
rect 14188 6404 14228 6448
rect 16865 6404 16905 6448
rect 17740 6404 17780 6448
rect 17875 6406 17884 6446
rect 17924 6406 17933 6446
rect 14141 6364 14188 6404
rect 14228 6364 14237 6404
rect 14729 6364 14851 6404
rect 14900 6364 14909 6404
rect 16483 6364 16492 6404
rect 16532 6364 16905 6404
rect 17635 6364 17644 6404
rect 17684 6364 17780 6404
rect 17879 6320 17919 6406
rect 21772 6404 21812 6448
rect 25324 6404 25364 6448
rect 27436 6404 27476 6448
rect 28012 6404 28052 6448
rect 28300 6404 28340 6448
rect 29164 6404 29204 6448
rect 18010 6364 18019 6404
rect 18059 6364 18068 6404
rect 21772 6364 22252 6404
rect 22292 6364 22301 6404
rect 23881 6364 23890 6404
rect 23930 6364 24172 6404
rect 24212 6364 24221 6404
rect 24876 6364 24940 6404
rect 24980 6364 25036 6404
rect 25076 6364 25364 6404
rect 25481 6364 25612 6404
rect 25652 6364 25661 6404
rect 26953 6364 26962 6404
rect 27002 6364 27340 6404
rect 27380 6364 27389 6404
rect 27436 6364 27475 6404
rect 27515 6364 27524 6404
rect 28003 6364 28012 6404
rect 28052 6364 28061 6404
rect 28300 6364 29059 6404
rect 29099 6364 29108 6404
rect 29164 6364 29260 6404
rect 29300 6364 29309 6404
rect 30499 6364 30508 6404
rect 30554 6364 30679 6404
rect 2851 6280 2860 6320
rect 2900 6280 4916 6320
rect 5801 6280 5932 6320
rect 5972 6280 6548 6320
rect 6595 6280 6604 6320
rect 6644 6280 9716 6320
rect 12154 6280 12163 6320
rect 12203 6280 12556 6320
rect 12596 6280 12605 6320
rect 13036 6280 13420 6320
rect 13460 6280 14036 6320
rect 16771 6280 16780 6320
rect 16820 6280 17919 6320
rect 13036 6236 13076 6280
rect 18028 6236 18068 6364
rect 20131 6280 20140 6320
rect 20180 6280 22828 6320
rect 22868 6280 22877 6320
rect 25385 6280 25516 6320
rect 25556 6280 25565 6320
rect 26668 6280 30452 6320
rect 4291 6196 4300 6236
rect 4340 6196 4972 6236
rect 5012 6196 5021 6236
rect 10060 6196 13076 6236
rect 15977 6196 16099 6236
rect 16148 6196 16157 6236
rect 17731 6196 17740 6236
rect 17780 6196 18068 6236
rect 18403 6196 18412 6236
rect 18452 6196 18691 6236
rect 18731 6196 18740 6236
rect 20585 6196 20716 6236
rect 20756 6196 20765 6236
rect 25865 6196 25987 6236
rect 26036 6196 26045 6236
rect 10060 6152 10100 6196
rect 26668 6152 26708 6280
rect 30412 6236 30452 6280
rect 29731 6196 29740 6236
rect 29780 6196 29789 6236
rect 30403 6196 30412 6236
rect 30452 6196 30461 6236
rect 29740 6152 29780 6196
rect 67 6112 76 6152
rect 116 6112 500 6152
rect 6787 6112 6796 6152
rect 6836 6112 10100 6152
rect 18499 6112 18508 6152
rect 18548 6112 26708 6152
rect 28771 6112 28780 6152
rect 28820 6112 29260 6152
rect 29300 6112 29309 6152
rect 29740 6112 30892 6152
rect 30932 6112 30941 6152
rect 0 5984 400 6004
rect 460 5984 500 6112
rect 3103 6028 3112 6068
rect 3480 6028 3489 6068
rect 6499 6028 6508 6068
rect 6548 6028 7084 6068
rect 7124 6028 7220 6068
rect 10877 6028 10886 6068
rect 11254 6028 11263 6068
rect 18651 6028 18660 6068
rect 19028 6028 19037 6068
rect 26425 6028 26434 6068
rect 26802 6028 26811 6068
rect 7180 5984 7220 6028
rect 0 5944 500 5984
rect 2860 5944 6700 5984
rect 6740 5944 6749 5984
rect 7180 5944 17740 5984
rect 17780 5944 17789 5984
rect 17923 5944 17932 5984
rect 17972 5944 21964 5984
rect 22004 5944 22013 5984
rect 27756 5944 27820 5984
rect 27860 5944 29644 5984
rect 29684 5944 30260 5984
rect 0 5924 400 5944
rect 2860 5900 2900 5944
rect 27916 5900 27956 5944
rect 2668 5860 2900 5900
rect 4265 5860 4348 5900
rect 4388 5860 4396 5900
rect 4436 5860 4820 5900
rect 2668 5732 2708 5860
rect 4553 5776 4684 5816
rect 4724 5776 4733 5816
rect 1036 5692 1228 5732
rect 1268 5692 1277 5732
rect 2345 5692 2467 5732
rect 2516 5692 2525 5732
rect 2659 5692 2668 5732
rect 2708 5692 2717 5732
rect 3052 5692 3532 5732
rect 3572 5692 3581 5732
rect 4195 5692 4204 5732
rect 4244 5692 4588 5732
rect 4628 5692 4637 5732
rect 1036 5648 1076 5692
rect 3052 5648 3092 5692
rect 521 5608 652 5648
rect 692 5608 701 5648
rect 1027 5608 1036 5648
rect 1076 5608 1085 5648
rect 1132 5608 1603 5648
rect 1643 5608 1652 5648
rect 1699 5608 1708 5648
rect 1748 5608 1879 5648
rect 2179 5608 2188 5648
rect 2228 5608 2327 5648
rect 2367 5608 2376 5648
rect 2563 5608 2572 5648
rect 2612 5608 2621 5648
rect 2729 5608 2860 5648
rect 2900 5608 2909 5648
rect 3043 5608 3052 5648
rect 3092 5608 3101 5648
rect 3427 5608 3436 5648
rect 3476 5608 3485 5648
rect 1132 5480 1172 5608
rect 2572 5564 2612 5608
rect 2572 5524 2956 5564
rect 2996 5524 3005 5564
rect 1123 5440 1132 5480
rect 1172 5440 1181 5480
rect 1987 5440 1996 5480
rect 2036 5440 2668 5480
rect 2708 5440 2717 5480
rect 3436 5396 3476 5608
rect 3532 5564 3572 5692
rect 4780 5690 4820 5860
rect 6988 5860 12980 5900
rect 16361 5860 16483 5900
rect 16532 5860 16541 5900
rect 20419 5860 20428 5900
rect 20468 5860 20908 5900
rect 20948 5860 20957 5900
rect 21353 5860 21475 5900
rect 21524 5860 21533 5900
rect 21580 5860 25228 5900
rect 25268 5860 25277 5900
rect 25402 5860 25411 5900
rect 25451 5860 25612 5900
rect 25652 5860 25661 5900
rect 27898 5860 27907 5900
rect 27947 5860 27956 5900
rect 29251 5860 29260 5900
rect 29300 5860 30028 5900
rect 30068 5860 30077 5900
rect 5731 5776 5740 5816
rect 5780 5807 6892 5816
rect 5780 5776 6268 5807
rect 6308 5776 6892 5807
rect 6932 5776 6941 5816
rect 6268 5758 6308 5767
rect 6988 5732 7028 5860
rect 12940 5816 12980 5860
rect 21580 5816 21620 5860
rect 7267 5776 7276 5816
rect 7316 5776 7988 5816
rect 9571 5776 9580 5816
rect 9620 5776 9629 5816
rect 10051 5776 10060 5816
rect 10100 5776 10868 5816
rect 12940 5776 14228 5816
rect 17635 5776 17644 5816
rect 17684 5776 17693 5816
rect 18220 5776 18412 5816
rect 18452 5776 18461 5816
rect 18892 5776 21620 5816
rect 21964 5776 22051 5816
rect 22091 5776 22100 5816
rect 22339 5776 22348 5816
rect 22388 5776 23116 5816
rect 23156 5776 23165 5816
rect 28876 5776 29164 5816
rect 29204 5776 29213 5816
rect 29827 5776 29836 5816
rect 29876 5776 29972 5816
rect 7948 5732 7988 5776
rect 9580 5732 9620 5776
rect 10828 5732 10868 5776
rect 14188 5732 14228 5776
rect 17644 5732 17684 5776
rect 18220 5732 18260 5776
rect 18892 5732 18932 5776
rect 21964 5732 22004 5776
rect 6403 5692 6412 5732
rect 6452 5692 6787 5732
rect 6827 5692 6836 5732
rect 6979 5692 6988 5732
rect 7028 5692 7037 5732
rect 7948 5692 9100 5732
rect 9140 5692 9332 5732
rect 9475 5692 9484 5732
rect 9524 5692 9533 5732
rect 9580 5692 10252 5732
rect 10292 5692 10301 5732
rect 10828 5692 10867 5732
rect 10907 5692 10916 5732
rect 11068 5692 11308 5732
rect 11348 5692 12556 5732
rect 12596 5692 12605 5732
rect 13027 5692 13036 5732
rect 13076 5692 13228 5732
rect 13268 5692 13277 5732
rect 14188 5692 15380 5732
rect 4762 5650 4771 5690
rect 4811 5650 4820 5690
rect 9292 5690 9332 5692
rect 9292 5650 9340 5690
rect 9380 5650 9389 5690
rect 3619 5608 3628 5648
rect 3668 5608 3724 5648
rect 3764 5608 3799 5648
rect 4169 5608 4204 5648
rect 4244 5608 4300 5648
rect 4340 5608 4349 5648
rect 4867 5608 4876 5648
rect 4939 5608 5047 5648
rect 5443 5608 5452 5648
rect 5492 5608 5501 5648
rect 5609 5608 5740 5648
rect 5780 5608 6124 5648
rect 6164 5608 6173 5648
rect 6269 5608 6307 5648
rect 6347 5608 6356 5648
rect 4396 5566 4435 5606
rect 4475 5566 4484 5606
rect 4396 5564 4436 5566
rect 5452 5564 5492 5608
rect 6316 5564 6356 5608
rect 6412 5608 6647 5648
rect 6687 5608 6696 5648
rect 6883 5608 6892 5648
rect 6932 5608 6941 5648
rect 7075 5608 7084 5648
rect 7124 5608 7180 5648
rect 7220 5608 7255 5648
rect 7372 5608 7852 5648
rect 7892 5608 7901 5648
rect 8227 5608 8236 5648
rect 8276 5608 8285 5648
rect 8633 5608 8716 5648
rect 8756 5608 8764 5648
rect 8804 5608 8813 5648
rect 8899 5608 8908 5648
rect 8948 5608 9044 5648
rect 3532 5524 4436 5564
rect 4675 5524 4684 5564
rect 4724 5524 6068 5564
rect 6307 5524 6316 5564
rect 6356 5524 6365 5564
rect 6028 5480 6068 5524
rect 6412 5480 6452 5608
rect 6892 5564 6932 5608
rect 6499 5524 6508 5564
rect 6548 5524 6932 5564
rect 7372 5480 7412 5608
rect 8236 5564 8276 5608
rect 9004 5564 9044 5608
rect 8236 5524 8660 5564
rect 8899 5524 8908 5564
rect 8948 5524 9044 5564
rect 8620 5480 8660 5524
rect 9484 5480 9524 5692
rect 11068 5648 11108 5692
rect 12748 5648 12788 5657
rect 12844 5648 12932 5651
rect 14188 5648 14228 5692
rect 15340 5648 15380 5692
rect 16314 5692 16396 5732
rect 16436 5692 16780 5732
rect 16820 5692 16829 5732
rect 17644 5692 17727 5732
rect 18019 5692 18028 5732
rect 18068 5692 18260 5732
rect 18307 5692 18316 5732
rect 18356 5692 18691 5732
rect 18731 5692 18740 5732
rect 18883 5692 18892 5732
rect 18932 5692 18941 5732
rect 20428 5692 20756 5732
rect 21481 5692 21490 5732
rect 21530 5692 22004 5732
rect 24460 5692 25268 5732
rect 16314 5690 16354 5692
rect 16300 5681 16354 5690
rect 9802 5608 9811 5648
rect 9851 5608 10060 5648
rect 10100 5608 10109 5648
rect 11050 5608 11059 5648
rect 11099 5608 11108 5648
rect 11194 5608 11203 5648
rect 11252 5608 11383 5648
rect 12329 5608 12449 5648
rect 12500 5608 12509 5648
rect 12617 5608 12748 5648
rect 12788 5608 12797 5648
rect 12844 5608 12892 5648
rect 12932 5608 12941 5648
rect 13018 5608 13027 5648
rect 13067 5608 13076 5648
rect 13123 5608 13132 5648
rect 13172 5608 13228 5648
rect 13268 5608 13303 5648
rect 13987 5608 13996 5648
rect 14036 5608 14045 5648
rect 14188 5608 14284 5648
rect 14324 5608 14333 5648
rect 14489 5608 14572 5648
rect 14612 5608 14620 5648
rect 14660 5608 14669 5648
rect 14755 5608 14764 5648
rect 14804 5608 14860 5648
rect 14900 5608 14935 5648
rect 15226 5608 15235 5648
rect 15275 5608 15284 5648
rect 15331 5608 15340 5648
rect 15380 5608 15389 5648
rect 15436 5608 15956 5648
rect 16186 5608 16195 5648
rect 16235 5608 16244 5648
rect 16340 5650 16354 5681
rect 17687 5690 17727 5692
rect 17687 5681 17732 5690
rect 17687 5650 17692 5681
rect 16300 5632 16340 5641
rect 17417 5608 17548 5648
rect 17588 5608 17597 5648
rect 18220 5648 18260 5692
rect 20428 5648 20468 5692
rect 20716 5648 20756 5692
rect 22060 5681 22376 5690
rect 22060 5650 22336 5681
rect 17692 5632 17732 5641
rect 17827 5608 17836 5648
rect 17876 5608 18124 5648
rect 18164 5608 18173 5648
rect 18220 5608 18263 5648
rect 18303 5608 18312 5648
rect 18354 5608 18551 5648
rect 18591 5608 18600 5648
rect 18787 5608 18796 5648
rect 18836 5608 18845 5648
rect 20131 5608 20140 5648
rect 20180 5608 20372 5648
rect 20419 5608 20428 5648
rect 20468 5608 20477 5648
rect 20602 5608 20611 5648
rect 20651 5608 20660 5648
rect 20707 5608 20716 5648
rect 20756 5608 20765 5648
rect 21571 5608 21580 5648
rect 21620 5608 21964 5648
rect 22004 5608 22013 5648
rect 9639 5566 9648 5606
rect 9688 5566 9716 5606
rect 12748 5599 12788 5608
rect 3610 5440 3619 5480
rect 3659 5440 3668 5480
rect 3715 5440 3724 5480
rect 3764 5440 4876 5480
rect 4916 5440 4925 5480
rect 5801 5440 5932 5480
rect 5972 5440 5981 5480
rect 6028 5440 6452 5480
rect 6691 5440 6700 5480
rect 6740 5440 7412 5480
rect 8131 5440 8140 5480
rect 8180 5440 8332 5480
rect 8372 5440 8381 5480
rect 8602 5440 8611 5480
rect 8651 5440 9524 5480
rect 2860 5356 3476 5396
rect 2860 5228 2900 5356
rect 1219 5188 1228 5228
rect 1268 5188 2900 5228
rect 3628 5228 3668 5440
rect 7372 5396 7412 5440
rect 9676 5396 9716 5566
rect 7372 5356 9716 5396
rect 11116 5524 11511 5564
rect 11551 5524 11560 5564
rect 11875 5524 11884 5564
rect 11924 5524 12547 5564
rect 12587 5524 12596 5564
rect 4343 5272 4352 5312
rect 4720 5272 4729 5312
rect 6883 5272 6892 5312
rect 6932 5272 8716 5312
rect 8756 5272 8765 5312
rect 3628 5188 4340 5228
rect 1577 5020 1708 5060
rect 1748 5020 1757 5060
rect 2860 4976 2900 5188
rect 3235 5104 3244 5144
rect 3284 5104 3293 5144
rect 3523 5104 3532 5144
rect 3572 5104 3860 5144
rect 3907 5104 3916 5144
rect 3956 5104 4108 5144
rect 4148 5104 4157 5144
rect 3244 5060 3284 5104
rect 3244 5020 3764 5060
rect 3724 4976 3764 5020
rect 3820 4976 3860 5104
rect 4300 4976 4340 5188
rect 11116 5144 11156 5524
rect 12844 5480 12884 5608
rect 13036 5564 13076 5608
rect 13996 5564 14036 5608
rect 15244 5564 15284 5608
rect 15436 5564 15476 5608
rect 13036 5524 13844 5564
rect 13996 5524 15284 5564
rect 15427 5524 15436 5564
rect 15476 5524 15485 5564
rect 15532 5524 15543 5564
rect 15583 5524 15592 5564
rect 13036 5480 13076 5524
rect 13804 5480 13844 5524
rect 14476 5480 14516 5524
rect 11290 5440 11299 5480
rect 11339 5440 11348 5480
rect 11395 5440 11404 5480
rect 11444 5440 11575 5480
rect 12556 5440 12652 5480
rect 12692 5440 12884 5480
rect 12931 5440 12940 5480
rect 12980 5440 13076 5480
rect 13786 5440 13795 5480
rect 13835 5440 13844 5480
rect 14458 5440 14467 5480
rect 14507 5440 14516 5480
rect 5731 5104 5740 5144
rect 5780 5104 6028 5144
rect 6068 5104 6077 5144
rect 7468 5104 8044 5144
rect 8084 5104 8093 5144
rect 9763 5104 9772 5144
rect 9812 5104 10196 5144
rect 10531 5104 10540 5144
rect 10580 5104 10589 5144
rect 11002 5104 11011 5144
rect 11051 5104 11156 5144
rect 4474 5020 4483 5060
rect 4523 5020 5356 5060
rect 5396 5020 5405 5060
rect 5356 4976 5396 5020
rect 7468 4976 7508 5104
rect 7642 5020 7651 5060
rect 7691 5020 7838 5060
rect 7878 5020 7887 5060
rect 8044 5020 8620 5060
rect 8660 5020 8669 5060
rect 8044 4976 8084 5020
rect 10156 4976 10196 5104
rect 10540 5060 10580 5104
rect 11308 5060 11348 5440
rect 12117 5272 12126 5312
rect 12494 5272 12503 5312
rect 12556 5228 12596 5440
rect 12739 5356 12748 5396
rect 12788 5356 14572 5396
rect 14612 5356 14621 5396
rect 12268 5188 12596 5228
rect 12739 5188 12748 5228
rect 12788 5188 14476 5228
rect 14516 5188 14525 5228
rect 12268 5144 12308 5188
rect 12259 5104 12268 5144
rect 12308 5104 12317 5144
rect 12442 5104 12451 5144
rect 12491 5104 12884 5144
rect 14458 5104 14467 5144
rect 14507 5104 14516 5144
rect 12460 5060 12500 5104
rect 10540 5020 11348 5060
rect 12067 5020 12076 5060
rect 12116 5020 12500 5060
rect 10732 4976 10772 5020
rect 12844 4976 12884 5104
rect 1481 4936 1516 4976
rect 1556 4936 1612 4976
rect 1652 4936 1661 4976
rect 1795 4936 1804 4976
rect 1844 4936 1975 4976
rect 2371 4936 2380 4976
rect 2420 4936 2851 4976
rect 2891 4936 2900 4976
rect 2947 4936 2956 4976
rect 2996 4936 3005 4976
rect 3401 4936 3436 4976
rect 3476 4936 3532 4976
rect 3572 4936 3581 4976
rect 3715 4936 3724 4976
rect 3764 4936 3773 4976
rect 3820 4936 4151 4976
rect 4191 4936 4200 4976
rect 4300 4936 4396 4976
rect 4436 4936 4445 4976
rect 5338 4936 5347 4976
rect 5387 4936 5396 4976
rect 5443 4936 5452 4976
rect 5492 4936 5623 4976
rect 7241 4936 7339 4976
rect 7412 4936 7508 4976
rect 7555 4936 7564 4976
rect 7604 4936 8084 4976
rect 8140 4967 8180 4976
rect 2956 4892 2996 4936
rect 3724 4892 3764 4936
rect 8681 4936 8812 4976
rect 8852 4936 8861 4976
rect 8995 4936 9004 4976
rect 9044 4936 9379 4976
rect 9419 4936 9428 4976
rect 9475 4936 9484 4976
rect 9524 4936 9655 4976
rect 10138 4936 10147 4976
rect 10187 4936 10196 4976
rect 10243 4936 10252 4976
rect 10292 4936 10423 4976
rect 10656 4936 10699 4976
rect 10739 4936 10772 4976
rect 10915 4936 10924 4976
rect 10964 4936 11095 4976
rect 11866 4936 11875 4976
rect 11915 4936 11924 4976
rect 11971 4936 11980 4976
rect 12026 4936 12151 4976
rect 12473 4936 12556 4976
rect 12596 4936 12604 4976
rect 12644 4936 12653 4976
rect 12739 4936 12748 4976
rect 12788 4936 12797 4976
rect 12844 4936 13175 4976
rect 13215 4936 13224 4976
rect 13411 4936 13420 4976
rect 13460 4936 13591 4976
rect 8140 4892 8180 4927
rect 11884 4892 11924 4936
rect 12748 4892 12788 4936
rect 14476 4892 14516 5104
rect 14572 4976 14612 5356
rect 15532 5144 15572 5524
rect 15916 5396 15956 5608
rect 16204 5564 16244 5608
rect 18354 5564 18394 5608
rect 18796 5564 18836 5608
rect 16099 5524 16108 5564
rect 16148 5524 16244 5564
rect 17836 5524 18124 5564
rect 18164 5524 18173 5564
rect 18220 5524 18394 5564
rect 18700 5524 18836 5564
rect 20332 5564 20372 5608
rect 20620 5564 20660 5608
rect 20332 5524 20660 5564
rect 20908 5524 20919 5564
rect 20959 5524 20968 5564
rect 17836 5480 17876 5524
rect 17827 5440 17836 5480
rect 17876 5440 17885 5480
rect 18220 5396 18260 5524
rect 18700 5480 18740 5524
rect 18403 5440 18412 5480
rect 18452 5440 18740 5480
rect 19930 5440 19939 5480
rect 19979 5440 19988 5480
rect 19948 5396 19988 5440
rect 15916 5356 18124 5396
rect 18164 5356 18260 5396
rect 18316 5356 19988 5396
rect 18316 5312 18356 5356
rect 15619 5272 15628 5312
rect 15668 5272 18356 5312
rect 19891 5272 19900 5312
rect 20268 5272 20277 5312
rect 20332 5228 20372 5524
rect 20585 5440 20707 5480
rect 20756 5440 20765 5480
rect 14755 5104 14764 5144
rect 14804 5104 15572 5144
rect 15628 5188 16492 5228
rect 16532 5188 16541 5228
rect 18403 5188 18412 5228
rect 18452 5188 19508 5228
rect 15628 5060 15668 5188
rect 15715 5104 15724 5144
rect 15764 5104 16148 5144
rect 16483 5104 16492 5144
rect 16532 5104 17356 5144
rect 17396 5104 17405 5144
rect 18403 5104 18412 5144
rect 18452 5104 19276 5144
rect 19316 5104 19325 5144
rect 15340 5020 15668 5060
rect 15340 4976 15380 5020
rect 16108 4976 16148 5104
rect 16553 5020 16588 5060
rect 16628 5020 16684 5060
rect 16724 5020 16733 5060
rect 17011 4976 17051 5104
rect 17242 5020 17251 5060
rect 17291 5020 17356 5060
rect 17396 5020 17431 5060
rect 18028 5020 18316 5060
rect 18356 5020 18365 5060
rect 18700 5020 18796 5060
rect 18836 5020 18845 5060
rect 18028 4976 18068 5020
rect 18700 4976 18740 5020
rect 18892 4976 18932 5104
rect 19468 5060 19508 5188
rect 20140 5188 20372 5228
rect 20140 5144 20180 5188
rect 20908 5144 20948 5524
rect 22060 5144 22100 5650
rect 24460 5648 24500 5692
rect 25228 5648 25268 5692
rect 28876 5648 28916 5776
rect 29932 5732 29972 5776
rect 29609 5692 29731 5732
rect 29780 5692 29789 5732
rect 29923 5692 29932 5732
rect 29972 5692 29981 5732
rect 30220 5690 30260 5944
rect 30473 5860 30595 5900
rect 30644 5860 30653 5900
rect 30220 5681 30303 5690
rect 30220 5650 30263 5681
rect 22336 5632 22376 5641
rect 22426 5608 22435 5648
rect 22475 5608 22540 5648
rect 22580 5608 22615 5648
rect 24067 5608 24076 5648
rect 24116 5608 24460 5648
rect 24500 5608 24509 5648
rect 24739 5608 24748 5648
rect 24788 5608 24797 5648
rect 25219 5608 25228 5648
rect 25268 5608 25277 5648
rect 25402 5608 25411 5648
rect 25451 5608 25460 5648
rect 25795 5608 25804 5648
rect 25844 5608 25853 5648
rect 25902 5608 25911 5648
rect 25951 5608 25996 5648
rect 26036 5608 26082 5648
rect 27139 5608 27148 5648
rect 27188 5608 27619 5648
rect 27659 5608 27668 5648
rect 27715 5608 27724 5648
rect 27764 5608 28108 5648
rect 28148 5608 28157 5648
rect 28474 5608 28483 5648
rect 28523 5608 28972 5648
rect 29012 5608 29021 5648
rect 29085 5608 29094 5648
rect 29134 5608 29143 5648
rect 29212 5608 29221 5648
rect 29261 5608 29452 5648
rect 29492 5608 29501 5648
rect 29582 5608 29591 5648
rect 29631 5608 29644 5648
rect 29684 5608 29762 5648
rect 29828 5608 29837 5648
rect 29877 5608 29886 5648
rect 29993 5608 30124 5648
rect 30164 5608 30173 5648
rect 30892 5648 30932 5657
rect 30263 5632 30303 5641
rect 30761 5608 30892 5648
rect 30932 5608 30941 5648
rect 24748 5564 24788 5608
rect 25420 5564 25460 5608
rect 23020 5524 25460 5564
rect 22243 5440 22252 5480
rect 22292 5440 22555 5480
rect 22595 5440 22604 5480
rect 23020 5312 23060 5524
rect 24809 5440 24940 5480
rect 24980 5440 24989 5480
rect 25594 5440 25603 5480
rect 25643 5440 25652 5480
rect 25612 5396 25652 5440
rect 24547 5356 24556 5396
rect 24596 5356 25652 5396
rect 20131 5104 20140 5144
rect 20180 5104 20189 5144
rect 20410 5104 20419 5144
rect 20459 5104 20468 5144
rect 20707 5104 20716 5144
rect 20756 5104 20948 5144
rect 21449 5104 21571 5144
rect 21620 5104 21629 5144
rect 21859 5104 21868 5144
rect 21908 5104 22100 5144
rect 22156 5272 23060 5312
rect 20428 5060 20468 5104
rect 22156 5060 22196 5272
rect 23203 5188 23212 5228
rect 23252 5188 24596 5228
rect 22793 5104 22915 5144
rect 22964 5104 22973 5144
rect 24041 5104 24172 5144
rect 24212 5104 24221 5144
rect 24346 5104 24355 5144
rect 24395 5104 24404 5144
rect 24364 5060 24404 5104
rect 18979 5020 18988 5060
rect 19028 5020 19171 5060
rect 19211 5020 19220 5060
rect 19468 5020 20468 5060
rect 20707 5020 20716 5060
rect 20756 5020 22196 5060
rect 23788 5020 24404 5060
rect 24556 5060 24596 5188
rect 25804 5144 25844 5608
rect 29103 5564 29143 5608
rect 28785 5524 28794 5564
rect 28834 5524 28876 5564
rect 28916 5524 28965 5564
rect 29103 5524 29548 5564
rect 29588 5524 29597 5564
rect 29836 5480 29876 5608
rect 30892 5599 30932 5608
rect 30307 5524 30316 5564
rect 30356 5524 30590 5564
rect 30630 5524 30639 5564
rect 28570 5440 28579 5480
rect 28619 5440 28628 5480
rect 28675 5440 28684 5480
rect 28724 5440 29876 5480
rect 30403 5440 30412 5480
rect 30452 5440 30796 5480
rect 30836 5440 30845 5480
rect 28588 5396 28628 5440
rect 28588 5356 29452 5396
rect 29492 5356 29501 5396
rect 27665 5272 27674 5312
rect 28042 5272 28051 5312
rect 28588 5228 28628 5356
rect 27523 5188 27532 5228
rect 27572 5188 27581 5228
rect 28012 5188 28628 5228
rect 27532 5144 27572 5188
rect 28012 5144 28052 5188
rect 25786 5104 25795 5144
rect 25835 5104 25844 5144
rect 26650 5104 26659 5144
rect 26699 5104 26708 5144
rect 26668 5060 26708 5104
rect 24556 5020 25844 5060
rect 19468 4976 19508 5020
rect 23788 4976 23828 5020
rect 24556 4976 24596 5020
rect 14563 4936 14572 4976
rect 14612 4936 14621 4976
rect 15322 4936 15331 4976
rect 15371 4936 15380 4976
rect 15427 4936 15436 4976
rect 15476 4936 15820 4976
rect 15860 4936 15869 4976
rect 15948 4936 16012 4976
rect 16052 4936 16099 4976
rect 16139 4936 16148 4976
rect 16195 4936 16204 4976
rect 16244 4936 16253 4976
rect 16649 4936 16780 4976
rect 16820 4936 16829 4976
rect 17002 4936 17011 4976
rect 17051 4936 17060 4976
rect 17144 4936 17153 4976
rect 17204 4936 17324 4976
rect 17449 4936 17458 4976
rect 17498 4936 17644 4976
rect 17684 4936 17693 4976
rect 18010 4936 18019 4976
rect 18059 4936 18068 4976
rect 18115 4936 18124 4976
rect 18164 4936 18295 4976
rect 18691 4936 18700 4976
rect 18740 4936 18749 4976
rect 18892 4936 18917 4976
rect 18957 4936 18966 4976
rect 19037 4936 19073 4976
rect 19113 4936 19124 4976
rect 15436 4892 15476 4936
rect 16204 4892 16244 4936
rect 17460 4892 17500 4936
rect 19084 4892 19124 4936
rect 19372 4967 19412 4976
rect 19468 4936 19660 4976
rect 19700 4936 19709 4976
rect 20035 4936 20044 4976
rect 20084 4936 20524 4976
rect 20564 4936 20573 4976
rect 21545 4936 21676 4976
rect 21716 4936 21725 4976
rect 23107 4936 23116 4976
rect 23156 4936 23287 4976
rect 23369 4936 23443 4976
rect 23483 4936 23500 4976
rect 23540 4936 23549 4976
rect 23770 4936 23779 4976
rect 23819 4936 23828 4976
rect 23875 4936 23884 4976
rect 23924 4936 24055 4976
rect 24532 4936 24541 4976
rect 24581 4936 24596 4976
rect 24643 4936 24652 4976
rect 24692 4936 25708 4976
rect 25748 4936 25757 4976
rect 19372 4892 19412 4927
rect 25804 4892 25844 5020
rect 25996 5020 26708 5060
rect 26860 5104 27572 5144
rect 28003 5104 28012 5144
rect 28052 5104 28061 5144
rect 28378 5104 28387 5144
rect 28427 5104 30164 5144
rect 30307 5104 30316 5144
rect 30356 5104 30365 5144
rect 30490 5104 30499 5144
rect 30548 5104 30679 5144
rect 25996 4976 26036 5020
rect 26860 4976 26900 5104
rect 27235 5020 27244 5060
rect 27284 5020 27293 5060
rect 27523 5020 27532 5060
rect 27572 5020 28492 5060
rect 28532 5020 28541 5060
rect 29356 5020 30068 5060
rect 27244 4976 27284 5020
rect 29356 4976 29396 5020
rect 30028 4976 30068 5020
rect 30124 4976 30164 5104
rect 30316 5060 30356 5104
rect 30316 5020 30836 5060
rect 30796 4976 30836 5020
rect 25972 4936 25981 4976
rect 26021 4936 26036 4976
rect 26083 4936 26092 4976
rect 26132 4936 26263 4976
rect 26851 4936 26860 4976
rect 26900 4936 26909 4976
rect 27017 4936 27148 4976
rect 27188 4936 27197 4976
rect 27244 4936 27811 4976
rect 27851 4936 27860 4976
rect 27977 4936 28012 4976
rect 28052 4936 28108 4976
rect 28148 4936 28157 4976
rect 28280 4936 28289 4976
rect 28340 4936 28460 4976
rect 28588 4967 28628 4976
rect 28958 4936 29068 4976
rect 29120 4936 29138 4976
rect 29225 4936 29356 4976
rect 29396 4936 29405 4976
rect 29530 4936 29539 4976
rect 29579 4936 29923 4976
rect 29963 4936 29972 4976
rect 30019 4936 30028 4976
rect 30068 4936 30077 4976
rect 30124 4936 30508 4976
rect 30548 4936 30652 4976
rect 30692 4936 30701 4976
rect 30787 4936 30796 4976
rect 30836 4936 30845 4976
rect 28588 4892 28628 4927
rect 2956 4852 3628 4892
rect 3668 4852 3677 4892
rect 3724 4852 4291 4892
rect 4331 4852 4340 4892
rect 7337 4852 7459 4892
rect 7508 4852 8180 4892
rect 10627 4852 10636 4892
rect 10676 4852 10819 4892
rect 10859 4852 11212 4892
rect 11252 4852 11261 4892
rect 11837 4852 11884 4892
rect 11924 4852 11933 4892
rect 12748 4852 12980 4892
rect 13027 4852 13036 4892
rect 13076 4852 13315 4892
rect 13355 4852 13364 4892
rect 13507 4852 13516 4892
rect 13556 4852 13565 4892
rect 14476 4852 15476 4892
rect 15907 4852 15916 4892
rect 15956 4852 16244 4892
rect 16906 4883 17500 4892
rect 12940 4808 12980 4852
rect 12940 4768 13228 4808
rect 13268 4768 13277 4808
rect 7747 4684 7756 4724
rect 7796 4684 7843 4724
rect 7883 4684 7927 4724
rect 8947 4684 8956 4724
rect 8996 4684 10060 4724
rect 10100 4684 10109 4724
rect 10156 4684 13132 4724
rect 13172 4684 13181 4724
rect 10156 4640 10196 4684
rect 8803 4600 8812 4640
rect 8852 4600 10196 4640
rect 3103 4516 3112 4556
rect 3480 4516 3489 4556
rect 10877 4516 10886 4556
rect 11254 4516 11263 4556
rect 13516 4472 13556 4852
rect 16906 4843 16915 4883
rect 16955 4852 17500 4883
rect 18595 4852 18604 4892
rect 18644 4852 18653 4892
rect 18796 4852 18819 4892
rect 18859 4852 18868 4892
rect 19075 4852 19084 4892
rect 19124 4852 19133 4892
rect 19372 4852 24844 4892
rect 24884 4852 24893 4892
rect 25804 4852 27956 4892
rect 28457 4852 28588 4892
rect 28628 4852 28915 4892
rect 28955 4852 28964 4892
rect 16955 4843 16964 4852
rect 16906 4842 16964 4843
rect 18604 4808 18644 4852
rect 17251 4768 17260 4808
rect 17300 4768 18644 4808
rect 18796 4808 18836 4852
rect 19372 4808 19412 4852
rect 27916 4808 27956 4852
rect 29932 4808 29972 4936
rect 18796 4768 19412 4808
rect 23491 4768 23500 4808
rect 23540 4768 24076 4808
rect 24116 4768 24125 4808
rect 27916 4768 28492 4808
rect 28532 4768 30452 4808
rect 17059 4684 17068 4724
rect 17108 4684 19084 4724
rect 19124 4684 19133 4724
rect 20515 4684 20524 4724
rect 20564 4684 23060 4724
rect 23107 4684 23116 4724
rect 23156 4684 27244 4724
rect 27284 4684 27293 4724
rect 29530 4684 29539 4724
rect 29579 4684 30316 4724
rect 30356 4684 30365 4724
rect 23020 4640 23060 4684
rect 23020 4600 28204 4640
rect 28244 4600 28253 4640
rect 18651 4516 18660 4556
rect 19028 4516 19037 4556
rect 26425 4516 26434 4556
rect 26802 4516 26811 4556
rect 9388 4432 11884 4472
rect 11924 4432 13036 4472
rect 13076 4432 13085 4472
rect 13516 4432 24884 4472
rect 1795 4348 1804 4388
rect 1844 4348 2900 4388
rect 3427 4348 3436 4388
rect 3476 4348 3532 4388
rect 3572 4348 3607 4388
rect 7241 4348 7372 4388
rect 7412 4348 7421 4388
rect 8515 4348 8524 4388
rect 8564 4348 9100 4388
rect 9140 4348 9149 4388
rect 556 4264 1612 4304
rect 1652 4264 1661 4304
rect 556 4136 596 4264
rect 1612 4220 1652 4264
rect 1420 4180 2228 4220
rect 1420 4136 1460 4180
rect 2188 4136 2228 4180
rect 2860 4136 2900 4348
rect 9388 4304 9428 4432
rect 9475 4348 9484 4388
rect 9524 4348 11596 4388
rect 11636 4348 12748 4388
rect 12788 4348 12797 4388
rect 13123 4348 13132 4388
rect 13172 4348 13420 4388
rect 13460 4348 13469 4388
rect 16265 4348 16300 4388
rect 16340 4348 16396 4388
rect 16436 4348 16445 4388
rect 18307 4348 18316 4388
rect 18356 4348 18412 4388
rect 18452 4348 18487 4388
rect 18700 4348 20716 4388
rect 20756 4348 20765 4388
rect 21182 4348 21676 4388
rect 21716 4348 21725 4388
rect 5059 4264 5068 4304
rect 5108 4264 5117 4304
rect 5338 4264 5347 4304
rect 5387 4264 9428 4304
rect 5068 4220 5108 4264
rect 5068 4180 5251 4220
rect 5291 4180 5300 4220
rect 5347 4180 5356 4220
rect 5396 4180 5500 4220
rect 5540 4180 5549 4220
rect 6604 4180 6892 4220
rect 6932 4180 6941 4220
rect 7180 4180 7843 4220
rect 7883 4180 7892 4220
rect 9193 4180 9202 4220
rect 9242 4180 10004 4220
rect 6604 4136 6644 4180
rect 7180 4136 7220 4180
rect 9964 4136 10004 4180
rect 10156 4136 10196 4348
rect 10627 4264 10636 4304
rect 10676 4264 10964 4304
rect 13891 4264 13900 4304
rect 13940 4264 15052 4304
rect 15092 4264 18028 4304
rect 18068 4264 18077 4304
rect 10924 4220 10964 4264
rect 10243 4180 10252 4220
rect 10292 4180 10772 4220
rect 10906 4180 10915 4220
rect 10955 4180 10964 4220
rect 11491 4180 11500 4220
rect 11540 4180 12556 4220
rect 12596 4180 13076 4220
rect 10732 4136 10772 4180
rect 13036 4136 13076 4180
rect 14476 4136 14516 4264
rect 18700 4220 18740 4348
rect 21182 4220 21222 4348
rect 24844 4304 24884 4432
rect 25900 4432 28012 4472
rect 28052 4432 29684 4472
rect 25900 4388 25940 4432
rect 25882 4348 25891 4388
rect 25931 4348 25940 4388
rect 26083 4348 26092 4388
rect 26132 4348 26659 4388
rect 26699 4348 26708 4388
rect 27322 4348 27331 4388
rect 27371 4348 29527 4388
rect 21274 4264 21283 4304
rect 21323 4264 21332 4304
rect 16492 4180 17635 4220
rect 17675 4180 18740 4220
rect 19657 4180 19666 4220
rect 19706 4180 21222 4220
rect 21292 4220 21332 4264
rect 24844 4264 26996 4304
rect 21292 4180 21778 4220
rect 21818 4180 21827 4220
rect 16492 4136 16532 4180
rect 24844 4136 24884 4264
rect 25981 4220 26021 4264
rect 25981 4180 26068 4220
rect 556 4096 748 4136
rect 788 4096 797 4136
rect 922 4096 931 4136
rect 971 4096 1132 4136
rect 1172 4096 1181 4136
rect 1420 4096 1432 4136
rect 1472 4096 1481 4136
rect 1524 4096 1612 4136
rect 1652 4096 1655 4136
rect 1695 4096 1704 4136
rect 1786 4096 1795 4136
rect 1835 4096 1844 4136
rect 1891 4096 1900 4136
rect 1940 4096 1949 4136
rect 2057 4096 2188 4136
rect 2228 4096 2237 4136
rect 2371 4096 2380 4136
rect 2420 4096 2551 4136
rect 2860 4096 3340 4136
rect 3380 4096 3389 4136
rect 3523 4096 3532 4136
rect 3572 4096 3581 4136
rect 4841 4096 4876 4136
rect 4916 4096 4972 4136
rect 5012 4096 5021 4136
rect 5443 4096 5452 4136
rect 5492 4096 5635 4136
rect 5675 4096 5684 4136
rect 6211 4096 6220 4136
rect 6260 4096 6269 4136
rect 6595 4096 6604 4136
rect 6644 4096 6653 4136
rect 6700 4096 7171 4136
rect 7211 4096 7220 4136
rect 7267 4096 7276 4136
rect 7316 4096 7703 4136
rect 7743 4096 7752 4136
rect 7939 4096 7948 4136
rect 7988 4096 7997 4136
rect 8393 4096 8515 4136
rect 8564 4096 8573 4136
rect 8803 4096 8812 4136
rect 8852 4096 9292 4136
rect 9332 4096 9341 4136
rect 9833 4096 9964 4136
rect 10004 4096 10013 4136
rect 10156 4096 10339 4136
rect 10379 4096 10388 4136
rect 10627 4096 10636 4136
rect 10676 4096 10685 4136
rect 10732 4096 10775 4136
rect 10815 4096 10824 4136
rect 11011 4096 11020 4136
rect 11060 4096 11308 4136
rect 11348 4096 11357 4136
rect 11404 4096 11452 4136
rect 11492 4096 11501 4136
rect 11587 4096 11596 4136
rect 11636 4096 12364 4136
rect 12404 4096 12413 4136
rect 12460 4096 12506 4136
rect 12546 4096 12980 4136
rect 13027 4096 13036 4136
rect 13076 4096 13085 4136
rect 13219 4096 13228 4136
rect 13268 4096 13420 4136
rect 13460 4096 14092 4136
rect 14132 4096 14141 4136
rect 14467 4096 14476 4136
rect 14516 4096 14525 4136
rect 15881 4096 16003 4136
rect 16052 4096 16061 4136
rect 16361 4096 16492 4136
rect 16532 4096 16541 4136
rect 16675 4096 16684 4136
rect 16724 4096 16855 4136
rect 17417 4096 17515 4136
rect 17588 4096 17597 4136
rect 17644 4096 17740 4136
rect 17780 4096 17789 4136
rect 18019 4096 18028 4136
rect 18068 4096 18211 4136
rect 18251 4096 18260 4136
rect 18307 4096 18316 4136
rect 18356 4096 18487 4136
rect 19747 4096 19756 4136
rect 19796 4096 19805 4136
rect 20986 4096 20995 4136
rect 21035 4096 21044 4136
rect 21091 4096 21100 4136
rect 21140 4096 21271 4136
rect 21859 4096 21868 4136
rect 21908 4096 22924 4136
rect 22964 4096 22973 4136
rect 23491 4096 23500 4136
rect 23540 4096 23549 4136
rect 23683 4096 23692 4136
rect 23732 4096 24172 4136
rect 24212 4096 24221 4136
rect 24844 4096 24940 4136
rect 24980 4096 24989 4136
rect 25289 4096 25324 4136
rect 25364 4096 25420 4136
rect 25460 4096 25469 4136
rect 25866 4107 25875 4147
rect 25915 4107 25924 4147
rect 26028 4136 26068 4180
rect 26350 4180 26380 4220
rect 26420 4180 26429 4220
rect 26350 4136 26390 4180
rect 26956 4136 26996 4264
rect 27820 4264 28204 4304
rect 28244 4264 28300 4304
rect 28340 4264 28349 4304
rect 27113 4180 27148 4220
rect 27188 4180 27197 4220
rect 1804 4052 1844 4096
rect 835 4012 844 4052
rect 884 4012 1844 4052
rect 1900 4052 1940 4096
rect 3532 4052 3572 4096
rect 6220 4052 6260 4096
rect 1900 4012 2284 4052
rect 2324 4012 2333 4052
rect 2851 4012 2860 4052
rect 2900 4012 3572 4052
rect 3907 4012 3916 4052
rect 3956 4012 6604 4052
rect 6644 4012 6653 4052
rect 6700 3968 6740 4096
rect 7948 4052 7988 4096
rect 9964 4052 10004 4096
rect 10636 4052 10676 4096
rect 11404 4052 11444 4096
rect 12460 4052 12500 4096
rect 7852 4012 7988 4052
rect 8817 4012 8826 4052
rect 8866 4012 9763 4052
rect 9803 4012 9812 4052
rect 9964 4012 11444 4052
rect 11875 4012 11884 4052
rect 11924 4012 12500 4052
rect 12940 4052 12980 4096
rect 12940 4012 13900 4052
rect 13940 4012 13949 4052
rect 16305 4012 16314 4052
rect 16354 4012 16588 4052
rect 16628 4012 16637 4052
rect 643 3928 652 3968
rect 692 3928 1267 3968
rect 1307 3928 1516 3968
rect 1556 3928 1565 3968
rect 1978 3928 1987 3968
rect 2027 3928 2036 3968
rect 4745 3928 4771 3968
rect 4811 3928 4876 3968
rect 4916 3928 4925 3968
rect 6691 3928 6700 3968
rect 6740 3928 6749 3968
rect 1996 3884 2036 3928
rect 1996 3844 5644 3884
rect 5684 3844 5693 3884
rect 4343 3760 4352 3800
rect 4720 3760 4729 3800
rect 2179 3676 2188 3716
rect 2228 3676 3916 3716
rect 3956 3676 3965 3716
rect 7852 3632 7892 4012
rect 17644 3968 17684 4096
rect 19756 4052 19796 4096
rect 17818 4012 17827 4052
rect 17867 4012 19796 4052
rect 8026 3928 8035 3968
rect 8075 3928 8611 3968
rect 8651 3928 8660 3968
rect 8707 3928 8716 3968
rect 8756 3928 8887 3968
rect 9929 3928 10051 3968
rect 10100 3928 10109 3968
rect 11098 3928 11107 3968
rect 11147 3928 11156 3968
rect 11290 3928 11299 3968
rect 11348 3928 11479 3968
rect 12521 3928 12556 3968
rect 12596 3928 12652 3968
rect 12692 3928 12701 3968
rect 14563 3928 14572 3968
rect 14612 3928 14621 3968
rect 15907 3928 15916 3968
rect 15956 3928 16099 3968
rect 16139 3928 16148 3968
rect 16675 3928 16684 3968
rect 16724 3928 17684 3968
rect 19337 3928 19459 3968
rect 19508 3928 19517 3968
rect 8620 3884 8660 3928
rect 8620 3844 9620 3884
rect 4867 3592 4876 3632
rect 4916 3592 5452 3632
rect 5492 3592 5501 3632
rect 5635 3592 5644 3632
rect 5684 3592 5740 3632
rect 5780 3592 5815 3632
rect 5897 3592 5923 3632
rect 5963 3592 6028 3632
rect 6068 3592 6796 3632
rect 6836 3592 6845 3632
rect 7738 3592 7747 3632
rect 7787 3592 7892 3632
rect 1411 3508 1420 3548
rect 1460 3508 1844 3548
rect 3811 3508 3820 3548
rect 3860 3508 8812 3548
rect 8852 3508 8861 3548
rect 1804 3464 1844 3508
rect 9580 3464 9620 3844
rect 9859 3592 9868 3632
rect 9908 3592 10676 3632
rect 10723 3592 10732 3632
rect 10772 3592 11020 3632
rect 11060 3592 11069 3632
rect 10636 3464 10676 3592
rect 1001 3424 1132 3464
rect 1172 3424 1181 3464
rect 1786 3424 1795 3464
rect 1835 3424 1996 3464
rect 2036 3424 2045 3464
rect 4387 3424 4396 3464
rect 4436 3424 4445 3464
rect 4553 3424 4684 3464
rect 4724 3424 4733 3464
rect 4867 3424 4876 3464
rect 4916 3424 5164 3464
rect 5204 3424 5213 3464
rect 5539 3424 5548 3464
rect 5588 3424 5597 3464
rect 5993 3424 6028 3464
rect 6068 3424 6124 3464
rect 6164 3424 6508 3464
rect 6548 3424 6557 3464
rect 7546 3424 7555 3464
rect 7595 3424 7700 3464
rect 8515 3424 8524 3464
rect 8564 3424 9475 3464
rect 9515 3424 9524 3464
rect 9571 3424 9580 3464
rect 9620 3424 9629 3464
rect 10618 3424 10627 3464
rect 10667 3424 10676 3464
rect 10723 3424 10732 3464
rect 10772 3424 10903 3464
rect 4396 3380 4436 3424
rect 4876 3380 4916 3424
rect 1267 3340 1276 3380
rect 1316 3340 1420 3380
rect 1460 3340 1469 3380
rect 2467 3340 2476 3380
rect 2516 3340 2525 3380
rect 4396 3340 4916 3380
rect 5548 3380 5588 3424
rect 7660 3380 7700 3424
rect 5548 3340 6932 3380
rect 6892 3296 6932 3340
rect 7660 3340 10156 3380
rect 10196 3340 10205 3380
rect 4675 3256 4684 3296
rect 4724 3256 4972 3296
rect 5012 3256 6124 3296
rect 6164 3256 6173 3296
rect 6883 3256 6892 3296
rect 6932 3256 7527 3296
rect 7567 3256 7576 3296
rect 3331 3172 3340 3212
rect 3380 3172 3389 3212
rect 3523 3172 3532 3212
rect 3572 3172 3724 3212
rect 3764 3172 3773 3212
rect 6211 3172 6220 3212
rect 6260 3172 7084 3212
rect 7124 3172 7133 3212
rect 3340 3128 3380 3172
rect 7660 3128 7700 3340
rect 11116 3212 11156 3928
rect 12117 3760 12126 3800
rect 12494 3760 12503 3800
rect 11971 3592 11980 3632
rect 12020 3592 12029 3632
rect 12643 3592 12652 3632
rect 12692 3592 13036 3632
rect 13076 3592 13085 3632
rect 13193 3592 13315 3632
rect 13364 3592 13373 3632
rect 13987 3592 13996 3632
rect 14036 3592 14275 3632
rect 14315 3592 14324 3632
rect 11980 3548 12020 3592
rect 11596 3508 11884 3548
rect 11924 3508 11933 3548
rect 11980 3508 12500 3548
rect 11596 3464 11636 3508
rect 12460 3464 12500 3508
rect 13034 3464 13074 3592
rect 14572 3548 14612 3928
rect 21004 3884 21044 4096
rect 23500 4052 23540 4096
rect 25876 4052 25916 4107
rect 26010 4096 26019 4136
rect 26059 4096 26068 4136
rect 26306 4096 26315 4136
rect 26355 4096 26390 4136
rect 26443 4096 26452 4136
rect 26516 4096 26632 4136
rect 27148 4136 27188 4180
rect 27820 4136 27860 4264
rect 28003 4180 28012 4220
rect 28052 4180 28061 4220
rect 28012 4136 28052 4180
rect 28396 4136 28436 4348
rect 29347 4264 29356 4304
rect 29396 4264 29405 4304
rect 29356 4136 29396 4264
rect 29487 4178 29527 4348
rect 29644 4220 29684 4432
rect 30412 4304 30452 4768
rect 30089 4264 30220 4304
rect 30260 4264 30269 4304
rect 30412 4264 30932 4304
rect 29626 4180 29635 4220
rect 29675 4180 29684 4220
rect 30569 4180 30700 4220
rect 30740 4180 30749 4220
rect 29487 4138 29500 4178
rect 29540 4138 29549 4178
rect 30892 4136 30932 4264
rect 27148 4096 27160 4136
rect 27200 4096 27209 4136
rect 27330 4096 27339 4136
rect 27379 4096 27436 4136
rect 27476 4096 27510 4136
rect 27675 4096 27684 4136
rect 27724 4096 27733 4136
rect 27811 4096 27820 4136
rect 27860 4096 27869 4136
rect 27965 4096 27998 4136
rect 28038 4096 28052 4136
rect 28128 4096 28137 4136
rect 28177 4096 28186 4136
rect 28291 4096 28300 4136
rect 28340 4096 28436 4136
rect 29347 4096 29356 4136
rect 29396 4096 29405 4136
rect 29731 4096 29740 4136
rect 29780 4096 29911 4136
rect 30228 4096 30316 4136
rect 30356 4096 30359 4136
rect 30399 4096 30408 4136
rect 30490 4096 30499 4136
rect 30539 4096 30548 4136
rect 30595 4096 30604 4136
rect 30644 4096 30653 4136
rect 30883 4096 30892 4136
rect 30932 4096 30941 4136
rect 31075 4096 31084 4136
rect 31124 4096 31133 4136
rect 23500 4012 23828 4052
rect 25795 4012 25804 4052
rect 25844 4012 25916 4052
rect 26170 4085 26228 4094
rect 26956 4087 26996 4096
rect 26170 4045 26179 4085
rect 26219 4045 26228 4085
rect 27693 4052 27733 4096
rect 28146 4052 28186 4096
rect 30508 4052 30548 4096
rect 30604 4052 30644 4096
rect 26170 4044 26228 4045
rect 23465 3928 23596 3968
rect 23636 3928 23645 3968
rect 21004 3844 21524 3884
rect 19891 3760 19900 3800
rect 20268 3760 20277 3800
rect 16204 3676 17588 3716
rect 17635 3676 17644 3716
rect 17684 3676 19796 3716
rect 16204 3548 16244 3676
rect 17548 3632 17588 3676
rect 19756 3632 19796 3676
rect 16457 3592 16588 3632
rect 16628 3592 16637 3632
rect 17225 3592 17356 3632
rect 17396 3592 17405 3632
rect 17539 3592 17548 3632
rect 17588 3592 17971 3632
rect 18011 3592 18020 3632
rect 19162 3592 19171 3632
rect 19211 3592 19220 3632
rect 19738 3592 19747 3632
rect 19787 3592 19796 3632
rect 19852 3676 20524 3716
rect 20564 3676 20573 3716
rect 14476 3508 14612 3548
rect 14860 3508 15332 3548
rect 14476 3464 14516 3508
rect 14860 3464 14900 3508
rect 15292 3506 15332 3508
rect 16108 3508 16244 3548
rect 16588 3548 16628 3592
rect 19180 3548 19220 3592
rect 19852 3548 19892 3676
rect 21484 3632 21524 3844
rect 16588 3508 17204 3548
rect 18307 3508 18316 3548
rect 18356 3508 19220 3548
rect 15292 3466 15312 3506
rect 15352 3466 15361 3506
rect 16108 3464 16148 3508
rect 17164 3464 17204 3508
rect 11578 3424 11587 3464
rect 11627 3424 11636 3464
rect 11683 3424 11692 3464
rect 11732 3424 11788 3464
rect 11828 3424 11863 3464
rect 12041 3424 12172 3464
rect 12212 3424 12221 3464
rect 12329 3424 12460 3464
rect 12500 3424 12509 3464
rect 12994 3424 13003 3464
rect 13043 3424 13074 3464
rect 13219 3424 13228 3464
rect 13268 3424 13399 3464
rect 13784 3424 13793 3464
rect 13844 3424 13964 3464
rect 14092 3455 14284 3464
rect 14132 3424 14284 3455
rect 14324 3424 14333 3464
rect 14452 3424 14461 3464
rect 14501 3424 14516 3464
rect 14563 3424 14572 3464
rect 14612 3424 14900 3464
rect 15010 3424 15019 3464
rect 15092 3424 15199 3464
rect 15466 3424 15475 3464
rect 15515 3424 15820 3464
rect 15860 3424 15869 3464
rect 16099 3424 16108 3464
rect 16148 3424 16157 3464
rect 16361 3424 16492 3464
rect 16532 3424 16541 3464
rect 16867 3424 16876 3464
rect 16916 3424 16925 3464
rect 17155 3424 17164 3464
rect 17204 3424 17213 3464
rect 18014 3424 18124 3464
rect 18176 3424 18185 3464
rect 18298 3424 18307 3464
rect 18347 3424 18356 3464
rect 18473 3424 18508 3464
rect 18548 3424 18604 3464
rect 18644 3424 18653 3464
rect 14092 3406 14132 3415
rect 14476 3380 14516 3424
rect 16876 3380 16916 3424
rect 13085 3340 13123 3380
rect 13163 3340 13172 3380
rect 14476 3340 15148 3380
rect 15188 3340 15197 3380
rect 15244 3340 16396 3380
rect 16436 3340 16916 3380
rect 13132 3296 13172 3340
rect 15244 3296 15284 3340
rect 18316 3296 18356 3424
rect 19180 3380 19220 3508
rect 19276 3508 19892 3548
rect 20236 3592 20515 3632
rect 20555 3592 20564 3632
rect 21466 3592 21475 3632
rect 21515 3592 21524 3632
rect 22121 3592 22243 3632
rect 22292 3592 22301 3632
rect 22819 3592 22828 3632
rect 22868 3592 22915 3632
rect 22955 3592 22999 3632
rect 23674 3592 23683 3632
rect 23723 3592 23732 3632
rect 19276 3464 19316 3508
rect 20236 3464 20276 3592
rect 23692 3464 23732 3592
rect 19267 3424 19276 3464
rect 19316 3424 19447 3464
rect 19651 3424 19660 3464
rect 19700 3424 19852 3464
rect 19892 3424 19901 3464
rect 20131 3424 20140 3464
rect 20180 3424 20236 3464
rect 20276 3424 20311 3464
rect 20515 3424 20524 3464
rect 20564 3424 20620 3464
rect 20660 3424 20695 3464
rect 20995 3424 21004 3464
rect 21044 3424 21140 3464
rect 21545 3424 21676 3464
rect 21716 3424 21725 3464
rect 21833 3424 21964 3464
rect 22004 3424 22013 3464
rect 22339 3424 22348 3464
rect 22388 3424 22397 3464
rect 22601 3424 22636 3464
rect 22676 3424 22732 3464
rect 22772 3424 22781 3464
rect 23203 3424 23212 3464
rect 23252 3424 23732 3464
rect 21100 3380 21140 3424
rect 19180 3340 21140 3380
rect 21676 3380 21716 3424
rect 22348 3380 22388 3424
rect 23788 3380 23828 4012
rect 24713 3928 24835 3968
rect 24884 3928 24893 3968
rect 26183 3884 26223 4044
rect 26523 4012 26572 4052
rect 26612 4012 26654 4052
rect 26694 4012 26703 4052
rect 27331 4012 27340 4052
rect 27380 4012 27572 4052
rect 27693 4012 28052 4052
rect 28146 4012 28204 4052
rect 28244 4012 28253 4052
rect 28300 4012 29827 4052
rect 29867 4012 29876 4052
rect 30461 4012 30508 4052
rect 30548 4012 30557 4052
rect 30604 4012 30988 4052
rect 31028 4012 31037 4052
rect 27532 3968 27572 4012
rect 26851 3928 26860 3968
rect 26900 3928 26909 3968
rect 27514 3928 27523 3968
rect 27563 3928 27572 3968
rect 28012 3968 28052 4012
rect 28300 3968 28340 4012
rect 31084 3968 31124 4096
rect 28012 3928 28340 3968
rect 28675 3928 28684 3968
rect 28724 3928 28780 3968
rect 28820 3928 28855 3968
rect 30220 3928 31124 3968
rect 26860 3884 26900 3928
rect 25411 3844 25420 3884
rect 25460 3844 26900 3884
rect 27665 3760 27674 3800
rect 28042 3760 28051 3800
rect 24460 3676 25324 3716
rect 25364 3676 26380 3716
rect 26420 3676 27148 3716
rect 27188 3676 27197 3716
rect 27820 3676 28204 3716
rect 28244 3676 29740 3716
rect 29780 3676 29789 3716
rect 24460 3464 24500 3676
rect 27820 3632 27860 3676
rect 30220 3632 30260 3928
rect 25289 3592 25420 3632
rect 25460 3592 25469 3632
rect 25690 3592 25699 3632
rect 25739 3592 25748 3632
rect 25795 3592 25804 3632
rect 25844 3592 25996 3632
rect 26036 3592 26572 3632
rect 26612 3592 26621 3632
rect 27811 3592 27820 3632
rect 27860 3592 27869 3632
rect 28963 3592 28972 3632
rect 29012 3592 29356 3632
rect 29396 3592 30260 3632
rect 25708 3548 25748 3592
rect 24940 3508 25748 3548
rect 27436 3508 28588 3548
rect 28628 3508 28637 3548
rect 28867 3508 28876 3548
rect 28916 3508 31267 3548
rect 31307 3508 31316 3548
rect 24940 3464 24980 3508
rect 27436 3464 27476 3508
rect 23971 3424 23980 3464
rect 24020 3424 24172 3464
rect 24212 3424 24460 3464
rect 24500 3424 24509 3464
rect 24643 3424 24652 3464
rect 24692 3424 24701 3464
rect 24809 3424 24940 3464
rect 24980 3424 24989 3464
rect 25315 3424 25324 3464
rect 25364 3424 25804 3464
rect 25844 3424 27052 3464
rect 27092 3424 27101 3464
rect 27418 3424 27427 3464
rect 27467 3424 27476 3464
rect 27523 3424 27532 3464
rect 27572 3424 27703 3464
rect 28195 3424 28204 3464
rect 28244 3424 28396 3464
rect 28436 3424 28445 3464
rect 28649 3424 28780 3464
rect 28820 3424 28829 3464
rect 30403 3424 30412 3464
rect 30452 3424 30883 3464
rect 30923 3424 30932 3464
rect 24652 3380 24692 3424
rect 27436 3380 27476 3424
rect 21676 3340 22388 3380
rect 23113 3340 23122 3380
rect 23162 3340 23212 3380
rect 23252 3340 23293 3380
rect 23404 3340 23890 3380
rect 23930 3340 27476 3380
rect 13123 3256 13132 3296
rect 13172 3256 13181 3296
rect 13647 3256 14572 3296
rect 14612 3256 14621 3296
rect 15235 3256 15244 3296
rect 15284 3256 15293 3296
rect 17635 3256 17644 3296
rect 17684 3256 18356 3296
rect 13647 3212 13687 3256
rect 21100 3212 21140 3340
rect 22348 3296 22388 3340
rect 23404 3296 23444 3340
rect 27532 3296 27572 3424
rect 30211 3340 30220 3380
rect 30260 3340 30269 3380
rect 22348 3256 23444 3296
rect 25699 3256 25708 3296
rect 25748 3256 27572 3296
rect 11116 3172 13687 3212
rect 13786 3172 13795 3212
rect 13835 3172 13844 3212
rect 14345 3172 14467 3212
rect 14516 3172 14525 3212
rect 18595 3172 18604 3212
rect 18644 3172 19276 3212
rect 19316 3172 19325 3212
rect 19459 3172 19468 3212
rect 19508 3172 20236 3212
rect 20276 3172 20285 3212
rect 21100 3172 22964 3212
rect 23779 3172 23788 3212
rect 23828 3172 24556 3212
rect 24596 3172 24605 3212
rect 28147 3172 28156 3212
rect 28196 3172 28780 3212
rect 28820 3172 28829 3212
rect 29225 3172 29356 3212
rect 29396 3172 29405 3212
rect 13804 3128 13844 3172
rect 22924 3128 22964 3172
rect 3340 3088 7700 3128
rect 8707 3088 8716 3128
rect 8756 3088 12172 3128
rect 12212 3088 12221 3128
rect 13804 3088 14860 3128
rect 14900 3088 14909 3128
rect 18211 3088 18220 3128
rect 18260 3088 21004 3128
rect 21044 3088 21053 3128
rect 22915 3088 22924 3128
rect 22964 3088 24940 3128
rect 24980 3088 24989 3128
rect 3103 3004 3112 3044
rect 3480 3004 3489 3044
rect 10877 3004 10886 3044
rect 11254 3004 11263 3044
rect 18651 3004 18660 3044
rect 19028 3004 19037 3044
rect 26425 3004 26434 3044
rect 26802 3004 26811 3044
rect 1891 2836 1900 2876
rect 1940 2836 1949 2876
rect 3785 2836 3916 2876
rect 3956 2836 3965 2876
rect 6316 2836 6836 2876
rect 7354 2836 7363 2876
rect 7403 2836 7468 2876
rect 7508 2836 7543 2876
rect 9466 2836 9475 2876
rect 9515 2836 10636 2876
rect 10676 2836 10685 2876
rect 13219 2836 13228 2876
rect 13268 2836 13420 2876
rect 13460 2836 13469 2876
rect 13699 2836 13708 2876
rect 13748 2836 17068 2876
rect 17108 2836 17117 2876
rect 18377 2836 18508 2876
rect 18548 2836 18557 2876
rect 20227 2836 20236 2876
rect 20276 2836 21044 2876
rect 21091 2836 21100 2876
rect 21140 2836 21187 2876
rect 21227 2836 21271 2876
rect 22540 2836 22772 2876
rect 22819 2836 22828 2876
rect 22868 2836 23164 2876
rect 23204 2836 24548 2876
rect 24835 2836 24844 2876
rect 24884 2836 27092 2876
rect 28745 2836 28771 2876
rect 28811 2836 28876 2876
rect 28916 2836 28925 2876
rect 1900 2792 1940 2836
rect 1228 2752 1940 2792
rect 2345 2752 2476 2792
rect 2516 2752 2525 2792
rect 4579 2752 4588 2792
rect 4628 2752 4876 2792
rect 4916 2752 4925 2792
rect 1001 2668 1132 2708
rect 1172 2668 1181 2708
rect 1228 2624 1268 2752
rect 1315 2668 1324 2708
rect 1387 2668 1652 2708
rect 1612 2624 1652 2668
rect 3052 2668 3628 2708
rect 3668 2668 4724 2708
rect 3052 2624 3092 2668
rect 4684 2624 4724 2668
rect 6316 2624 6356 2836
rect 6796 2792 6836 2836
rect 21004 2792 21044 2836
rect 22540 2792 22580 2836
rect 6569 2752 6700 2792
rect 6740 2752 6749 2792
rect 6796 2752 6892 2792
rect 6932 2752 7796 2792
rect 6892 2668 7084 2708
rect 7124 2668 7700 2708
rect 6892 2666 6932 2668
rect 1219 2584 1228 2624
rect 1268 2584 1277 2624
rect 1456 2584 1465 2624
rect 1505 2584 1514 2624
rect 1594 2584 1603 2624
rect 1643 2584 1652 2624
rect 1699 2584 1708 2624
rect 1748 2584 2900 2624
rect 3043 2584 3052 2624
rect 3092 2584 3101 2624
rect 3235 2584 3244 2624
rect 3284 2584 3293 2624
rect 3401 2584 3523 2624
rect 3572 2584 3581 2624
rect 4457 2584 4588 2624
rect 4628 2584 4637 2624
rect 4684 2584 4894 2624
rect 4934 2584 4943 2624
rect 5827 2584 5836 2624
rect 5876 2584 6028 2624
rect 6068 2584 6077 2624
rect 6298 2584 6307 2624
rect 6347 2584 6356 2624
rect 6424 2657 6932 2666
rect 6464 2626 6932 2657
rect 7660 2624 7700 2668
rect 7756 2666 7796 2752
rect 12652 2752 15916 2792
rect 15956 2752 15965 2792
rect 16108 2752 16204 2792
rect 16244 2752 16253 2792
rect 16300 2752 17356 2792
rect 17396 2752 17405 2792
rect 19267 2752 19276 2792
rect 19316 2752 20468 2792
rect 21004 2752 22580 2792
rect 22627 2752 22636 2792
rect 22676 2752 22685 2792
rect 12652 2708 12692 2752
rect 16108 2708 16148 2752
rect 9196 2668 9388 2708
rect 9428 2668 9859 2708
rect 9899 2668 9908 2708
rect 12329 2668 12451 2708
rect 12500 2668 12509 2708
rect 12643 2668 12652 2708
rect 12692 2668 12701 2708
rect 14755 2668 14764 2708
rect 14804 2668 14956 2708
rect 14996 2668 15005 2708
rect 15907 2668 15916 2708
rect 15956 2668 16148 2708
rect 7756 2657 7839 2666
rect 7756 2626 7799 2657
rect 6424 2608 6464 2617
rect 7066 2584 7075 2624
rect 7115 2584 7124 2624
rect 7171 2584 7180 2624
rect 7220 2584 7229 2624
rect 7651 2584 7660 2624
rect 7700 2584 7709 2624
rect 9196 2624 9236 2668
rect 16300 2666 16340 2752
rect 16387 2668 16396 2708
rect 16436 2668 16445 2708
rect 17635 2668 17644 2708
rect 17684 2668 17746 2708
rect 17786 2668 17815 2708
rect 18601 2668 18610 2708
rect 18650 2668 19180 2708
rect 19220 2668 19229 2708
rect 16243 2626 16252 2666
rect 16292 2626 16340 2666
rect 16396 2624 16436 2668
rect 17164 2624 17204 2633
rect 7799 2608 7839 2617
rect 8410 2584 8419 2624
rect 8459 2584 8468 2624
rect 8515 2584 8524 2624
rect 8564 2584 8908 2624
rect 8948 2584 8957 2624
rect 9178 2584 9187 2624
rect 9227 2584 9236 2624
rect 9283 2584 9292 2624
rect 9332 2584 9719 2624
rect 9759 2584 9768 2624
rect 9955 2584 9964 2624
rect 10004 2584 10013 2624
rect 10723 2584 10732 2624
rect 10772 2584 11500 2624
rect 11540 2584 11549 2624
rect 12163 2584 12172 2624
rect 12212 2584 12311 2624
rect 12351 2584 12360 2624
rect 12547 2584 12556 2624
rect 12596 2584 12727 2624
rect 13001 2584 13123 2624
rect 13172 2584 13181 2624
rect 13425 2584 13434 2624
rect 13474 2584 13708 2624
rect 13748 2584 13757 2624
rect 14467 2584 14476 2624
rect 14516 2584 14615 2624
rect 14655 2584 14664 2624
rect 14746 2584 14755 2624
rect 14795 2584 14804 2624
rect 14851 2584 14860 2624
rect 14900 2584 15031 2624
rect 16003 2584 16012 2624
rect 16052 2584 16061 2624
rect 16122 2584 16131 2624
rect 16171 2584 16180 2624
rect 16396 2584 16435 2624
rect 16475 2584 16484 2624
rect 16529 2584 16538 2624
rect 16578 2584 16587 2624
rect 17033 2584 17164 2624
rect 17204 2584 17588 2624
rect 17827 2584 17836 2624
rect 17876 2584 18508 2624
rect 18548 2584 18557 2624
rect 18691 2584 18700 2624
rect 18740 2584 19604 2624
rect 19651 2584 19660 2624
rect 19700 2584 19939 2624
rect 19979 2584 19988 2624
rect 20116 2584 20236 2624
rect 20287 2584 20296 2624
rect 1474 2540 1514 2584
rect 1708 2540 1748 2584
rect 2860 2540 2900 2584
rect 3244 2540 3284 2584
rect 1385 2500 1516 2540
rect 1556 2500 1748 2540
rect 1905 2500 1914 2540
rect 1954 2500 2092 2540
rect 2132 2500 2141 2540
rect 2851 2500 2860 2540
rect 2900 2500 3380 2540
rect 4649 2500 4684 2540
rect 4724 2500 4780 2540
rect 4820 2500 4829 2540
rect 3340 2456 3380 2500
rect 7084 2456 7124 2584
rect 7180 2540 7220 2584
rect 7180 2500 7988 2540
rect 7948 2456 7988 2500
rect 8428 2456 8468 2584
rect 9292 2540 9332 2584
rect 9964 2540 10004 2584
rect 14764 2540 14804 2584
rect 8812 2500 9332 2540
rect 9484 2500 10004 2540
rect 13027 2500 13036 2540
rect 13076 2500 13228 2540
rect 13268 2500 13277 2540
rect 14275 2500 14284 2540
rect 14324 2500 14804 2540
rect 8812 2456 8852 2500
rect 3226 2416 3235 2456
rect 3275 2416 3284 2456
rect 3340 2416 4780 2456
rect 4820 2416 4829 2456
rect 5059 2416 5068 2456
rect 5108 2416 5117 2456
rect 5347 2416 5356 2456
rect 5396 2416 5405 2456
rect 5731 2416 5740 2456
rect 5780 2447 7124 2456
rect 5780 2416 6211 2447
rect 3244 2204 3284 2416
rect 4343 2248 4352 2288
rect 4720 2248 4729 2288
rect 3244 2164 4340 2204
rect 1228 2080 2092 2120
rect 2132 2080 2141 2120
rect 2860 2080 4195 2120
rect 4235 2080 4244 2120
rect 1228 1952 1268 2080
rect 2860 2036 2900 2080
rect 1315 1996 1324 2036
rect 1364 1996 1603 2036
rect 1643 1996 1652 2036
rect 1708 1996 2900 2036
rect 1708 1952 1748 1996
rect 4300 1952 4340 2164
rect 1219 1912 1228 1952
rect 1268 1912 1277 1952
rect 1402 1912 1411 1952
rect 1451 1912 1748 1952
rect 1978 1912 1987 1952
rect 2036 1912 2167 1952
rect 4291 1912 4300 1952
rect 4340 1912 4396 1952
rect 4436 1912 4500 1952
rect 4649 1912 4684 1952
rect 4724 1912 4780 1952
rect 4820 1912 4829 1952
rect 5068 1868 5108 2416
rect 5356 2288 5396 2416
rect 6202 2407 6211 2416
rect 6251 2416 7124 2447
rect 7939 2416 7948 2456
rect 7988 2416 7997 2456
rect 8428 2416 8756 2456
rect 8803 2416 8812 2456
rect 8852 2416 8861 2456
rect 6251 2407 6260 2416
rect 6202 2406 6260 2407
rect 5164 2248 5396 2288
rect 5164 1952 5204 2248
rect 5260 2164 7124 2204
rect 5260 2120 5300 2164
rect 5251 2080 5260 2120
rect 5300 2080 5309 2120
rect 6761 2080 6796 2120
rect 6836 2080 6892 2120
rect 6932 2080 6941 2120
rect 6019 1996 6028 2036
rect 6068 1996 7028 2036
rect 6988 1952 7028 1996
rect 5164 1912 5452 1952
rect 5492 1912 5501 1952
rect 6281 1912 6412 1952
rect 6452 1912 6461 1952
rect 6970 1912 6979 1952
rect 7019 1912 7028 1952
rect 7084 1952 7124 2164
rect 8716 2036 8756 2416
rect 9484 2120 9524 2500
rect 10042 2416 10051 2456
rect 10091 2416 10100 2456
rect 10618 2416 10627 2456
rect 10667 2416 10676 2456
rect 10915 2416 10924 2456
rect 10964 2416 11308 2456
rect 11348 2416 11357 2456
rect 10060 2204 10100 2416
rect 10636 2372 10676 2416
rect 16012 2372 16052 2584
rect 16131 2540 16171 2584
rect 16547 2540 16587 2584
rect 17164 2575 17204 2584
rect 16131 2500 16204 2540
rect 16244 2500 16253 2540
rect 16547 2500 16588 2540
rect 16628 2500 16637 2540
rect 16856 2500 16865 2540
rect 16905 2500 17068 2540
rect 17108 2500 17117 2540
rect 17548 2456 17588 2584
rect 16553 2416 16684 2456
rect 16724 2416 16733 2456
rect 16954 2416 16963 2456
rect 17003 2416 17012 2456
rect 17059 2416 17068 2456
rect 17108 2416 17356 2456
rect 17396 2416 17405 2456
rect 17530 2416 17539 2456
rect 17579 2416 17588 2456
rect 16972 2372 17012 2416
rect 10147 2332 10156 2372
rect 10196 2332 11596 2372
rect 11636 2332 11645 2372
rect 16012 2332 17012 2372
rect 19564 2372 19604 2584
rect 20428 2540 20468 2752
rect 21484 2624 21524 2633
rect 22636 2624 22676 2752
rect 22732 2708 22772 2836
rect 22819 2752 22828 2792
rect 22868 2752 24212 2792
rect 22732 2668 23212 2708
rect 23252 2668 23587 2708
rect 23627 2668 23636 2708
rect 23753 2668 23788 2708
rect 23828 2668 23884 2708
rect 23924 2668 23933 2708
rect 23980 2668 24076 2708
rect 24116 2668 24125 2708
rect 23980 2624 24020 2668
rect 24172 2624 24212 2752
rect 24508 2624 24548 2836
rect 24652 2752 25564 2792
rect 25604 2752 25613 2792
rect 26729 2752 26860 2792
rect 26900 2752 26909 2792
rect 24652 2624 24692 2752
rect 24748 2668 25460 2708
rect 20611 2584 20620 2624
rect 20660 2584 21484 2624
rect 21667 2584 21676 2624
rect 21716 2584 21964 2624
rect 22004 2584 22013 2624
rect 22147 2584 22156 2624
rect 22196 2584 22540 2624
rect 22580 2584 22589 2624
rect 22636 2584 22662 2624
rect 22702 2584 22711 2624
rect 22780 2584 22789 2624
rect 22829 2584 22924 2624
rect 22964 2584 23028 2624
rect 23212 2584 23308 2624
rect 23348 2584 23357 2624
rect 23458 2584 23467 2624
rect 23507 2584 23516 2624
rect 23683 2584 23692 2624
rect 23732 2584 23788 2624
rect 23828 2584 23863 2624
rect 23971 2584 23980 2624
rect 24020 2584 24029 2624
rect 24154 2584 24163 2624
rect 24203 2584 24364 2624
rect 24404 2584 24413 2624
rect 24499 2584 24508 2624
rect 24548 2584 24557 2624
rect 24643 2584 24652 2624
rect 24692 2584 24701 2624
rect 21484 2575 21524 2584
rect 22828 2540 22868 2584
rect 20009 2500 20044 2540
rect 20084 2500 20140 2540
rect 20180 2500 20189 2540
rect 20428 2500 21182 2540
rect 21222 2500 21231 2540
rect 21859 2500 21868 2540
rect 21908 2500 22868 2540
rect 21379 2416 21388 2456
rect 21428 2416 21580 2456
rect 21620 2416 21629 2456
rect 22217 2416 22348 2456
rect 22388 2416 22397 2456
rect 22627 2416 22636 2456
rect 22676 2416 22828 2456
rect 22868 2416 22877 2456
rect 19564 2332 19756 2372
rect 19796 2332 22540 2372
rect 22580 2332 22589 2372
rect 12117 2248 12126 2288
rect 12494 2248 12503 2288
rect 13795 2248 13804 2288
rect 13844 2248 14516 2288
rect 19891 2248 19900 2288
rect 20268 2248 20277 2288
rect 14476 2204 14516 2248
rect 10060 2164 14420 2204
rect 14476 2164 18412 2204
rect 18452 2164 18461 2204
rect 18700 2164 22156 2204
rect 22196 2164 22205 2204
rect 8995 2080 9004 2120
rect 9044 2080 9524 2120
rect 10339 2080 10348 2120
rect 10388 2080 10397 2120
rect 10601 2080 10723 2120
rect 10772 2080 10781 2120
rect 12259 2080 12268 2120
rect 12308 2080 12317 2120
rect 13001 2080 13132 2120
rect 13172 2080 13181 2120
rect 13420 2080 13747 2120
rect 13787 2080 13804 2120
rect 13844 2080 13853 2120
rect 10348 2036 10388 2080
rect 8716 1996 9236 2036
rect 9196 1952 9236 1996
rect 9868 1996 10156 2036
rect 10196 1996 10205 2036
rect 10348 1996 10636 2036
rect 10676 1996 11252 2036
rect 9868 1952 9908 1996
rect 11212 1952 11252 1996
rect 7084 1912 8908 1952
rect 8948 1912 9004 1952
rect 9044 1912 9079 1952
rect 9187 1912 9196 1952
rect 9236 1912 9245 1952
rect 9859 1912 9868 1952
rect 9908 1912 9917 1952
rect 10243 1912 10252 1952
rect 10292 1912 10301 1952
rect 10723 1912 10732 1952
rect 10772 1912 10828 1952
rect 10868 1912 10903 1952
rect 11203 1912 11212 1952
rect 11252 1912 11261 1952
rect 11657 1912 11788 1952
rect 11828 1912 11837 1952
rect 12041 1912 12172 1952
rect 12212 1912 12221 1952
rect 9196 1868 9236 1912
rect 10252 1868 10292 1912
rect 12268 1868 12308 2080
rect 13420 2036 13460 2080
rect 12355 1996 12364 2036
rect 12404 1996 13460 2036
rect 13900 1952 13940 2164
rect 14380 2120 14420 2164
rect 13987 2080 13996 2120
rect 14036 2080 14045 2120
rect 14153 2080 14275 2120
rect 14324 2080 14333 2120
rect 14380 2080 14899 2120
rect 14939 2080 14948 2120
rect 15811 2080 15820 2120
rect 15860 2080 16204 2120
rect 16244 2080 18019 2120
rect 18059 2080 18068 2120
rect 18307 2080 18316 2120
rect 18356 2080 18604 2120
rect 18644 2080 18653 2120
rect 13996 2036 14036 2080
rect 18316 2036 18356 2080
rect 13996 1996 15188 2036
rect 18225 1996 18234 2036
rect 18274 1996 18356 2036
rect 12547 1912 12556 1952
rect 12596 1912 12739 1952
rect 12779 1912 12788 1952
rect 12835 1912 12844 1952
rect 12884 1912 13036 1952
rect 13076 1912 13085 1952
rect 13193 1912 13324 1952
rect 13364 1912 13373 1952
rect 13507 1912 13516 1952
rect 13556 1912 13804 1952
rect 13844 1912 13853 1952
rect 13900 1912 14380 1952
rect 14420 1912 14429 1952
rect 14755 1912 14764 1952
rect 14804 1912 15043 1952
rect 15083 1912 15092 1952
rect 15148 1943 15188 1996
rect 18700 1952 18740 2164
rect 23212 2120 23252 2584
rect 23476 2540 23516 2584
rect 24748 2540 24788 2668
rect 25420 2624 25460 2668
rect 27052 2624 27092 2836
rect 30185 2752 30316 2792
rect 30356 2752 30365 2792
rect 28396 2668 29356 2708
rect 29396 2668 29405 2708
rect 28396 2624 28436 2668
rect 25193 2584 25228 2624
rect 25268 2584 25324 2624
rect 25364 2584 25373 2624
rect 25673 2584 25756 2624
rect 25796 2584 25804 2624
rect 25844 2584 25853 2624
rect 27052 2584 28204 2624
rect 28244 2584 28253 2624
rect 28387 2584 28396 2624
rect 28436 2584 28445 2624
rect 28579 2584 28588 2624
rect 28628 2584 28637 2624
rect 28762 2584 28771 2624
rect 28811 2584 28820 2624
rect 28954 2584 28963 2624
rect 29003 2584 29012 2624
rect 29251 2584 29260 2624
rect 29300 2584 29443 2624
rect 29483 2584 29492 2624
rect 30115 2584 30124 2624
rect 30164 2584 30173 2624
rect 25420 2540 25460 2584
rect 28588 2540 28628 2584
rect 28780 2540 28820 2584
rect 23476 2500 23596 2540
rect 23636 2500 23645 2540
rect 24067 2500 24076 2540
rect 24116 2500 24788 2540
rect 25112 2500 25121 2540
rect 25161 2500 25364 2540
rect 25420 2500 25996 2540
rect 26036 2500 26045 2540
rect 28204 2500 28628 2540
rect 28771 2500 28780 2540
rect 28820 2500 28867 2540
rect 25210 2416 25219 2456
rect 25259 2416 25268 2456
rect 25228 2372 25268 2416
rect 24163 2332 24172 2372
rect 24212 2332 25268 2372
rect 25324 2372 25364 2500
rect 28204 2372 28244 2500
rect 28291 2416 28300 2456
rect 28340 2416 28349 2456
rect 25324 2332 28244 2372
rect 25324 2288 25364 2332
rect 24259 2248 24268 2288
rect 24308 2248 25364 2288
rect 27665 2248 27674 2288
rect 28042 2248 28051 2288
rect 21475 2080 21484 2120
rect 21524 2080 21964 2120
rect 22004 2080 22013 2120
rect 22636 2080 23116 2120
rect 23156 2080 23165 2120
rect 23212 2080 24652 2120
rect 24692 2080 24701 2120
rect 27523 2080 27532 2120
rect 27572 2080 28108 2120
rect 28148 2080 28157 2120
rect 22636 2036 22676 2080
rect 19564 1996 22676 2036
rect 23116 2036 23156 2080
rect 23116 1996 23980 2036
rect 24020 1996 26228 2036
rect 19564 1952 19604 1996
rect 14764 1868 14804 1912
rect 16291 1912 16300 1952
rect 16340 1912 16780 1952
rect 16820 1912 16829 1952
rect 17914 1912 17923 1952
rect 17963 1912 17972 1952
rect 18019 1912 18028 1952
rect 18068 1912 18595 1952
rect 18635 1912 18644 1952
rect 18691 1912 18700 1952
rect 18740 1912 18749 1952
rect 19546 1912 19555 1952
rect 19595 1912 19604 1952
rect 21737 1912 21811 1952
rect 21851 1912 21868 1952
rect 21908 1912 21917 1952
rect 21997 1912 22006 1952
rect 22046 1912 22348 1952
rect 22388 1912 22397 1952
rect 22714 1912 22723 1952
rect 22763 1912 22772 1952
rect 22818 1914 22827 1954
rect 22867 1914 22876 1954
rect 26188 1952 26228 1996
rect 15148 1894 15188 1903
rect 17932 1868 17972 1912
rect 18700 1868 18740 1912
rect 22732 1868 22772 1912
rect 22828 1868 22868 1914
rect 23299 1912 23308 1952
rect 23348 1912 23357 1952
rect 23491 1912 23500 1952
rect 23540 1912 23549 1952
rect 24041 1912 24163 1952
rect 24212 1912 24221 1952
rect 24329 1912 24460 1952
rect 24500 1912 24509 1952
rect 25193 1912 25324 1952
rect 25364 1912 25373 1952
rect 26170 1912 26179 1952
rect 26219 1912 26228 1952
rect 28204 1952 28244 2332
rect 28300 2036 28340 2416
rect 28972 2120 29012 2584
rect 29155 2416 29164 2456
rect 29204 2416 29213 2456
rect 28570 2080 28579 2120
rect 28619 2080 29012 2120
rect 29164 2036 29204 2416
rect 30124 2120 30164 2584
rect 30124 2080 31084 2120
rect 31124 2080 31133 2120
rect 28300 1996 28628 2036
rect 28675 1996 28684 2036
rect 28724 1996 28916 2036
rect 29164 1996 30164 2036
rect 28588 1952 28628 1996
rect 28204 1912 28478 1952
rect 28518 1912 28527 1952
rect 28588 1943 28820 1952
rect 28588 1912 28780 1943
rect 23308 1868 23348 1912
rect 23500 1868 23540 1912
rect 2659 1828 2668 1868
rect 2708 1828 2717 1868
rect 3523 1828 3532 1868
rect 3572 1828 3820 1868
rect 3860 1828 3869 1868
rect 5068 1828 9044 1868
rect 9196 1828 11500 1868
rect 11540 1828 11549 1868
rect 12268 1828 14804 1868
rect 15436 1828 17644 1868
rect 17684 1828 17693 1868
rect 17932 1828 18740 1868
rect 19049 1828 19180 1868
rect 19220 1828 19229 1868
rect 20832 1828 20908 1868
rect 20948 1828 20957 1868
rect 22627 1828 22636 1868
rect 22676 1828 22772 1868
rect 22819 1828 22828 1868
rect 22868 1828 22912 1868
rect 23020 1828 23348 1868
rect 23491 1828 23500 1868
rect 23540 1828 24268 1868
rect 24308 1828 24317 1868
rect 25795 1828 25804 1868
rect 25844 1828 25853 1868
rect 26851 1828 26860 1868
rect 26900 1828 26909 1868
rect 27715 1828 27724 1868
rect 27764 1828 28108 1868
rect 28148 1828 28157 1868
rect 3907 1744 3916 1784
rect 3956 1744 5836 1784
rect 5876 1744 5885 1784
rect 6115 1744 6124 1784
rect 6164 1744 7024 1784
rect 7064 1744 7073 1784
rect 7433 1744 7564 1784
rect 7604 1744 7613 1784
rect 9004 1700 9044 1828
rect 15436 1784 15476 1828
rect 12940 1744 13556 1784
rect 15427 1744 15436 1784
rect 15476 1744 15485 1784
rect 16649 1744 16780 1784
rect 16820 1744 16829 1784
rect 12940 1700 12980 1744
rect 13516 1700 13556 1744
rect 17932 1700 17972 1828
rect 23020 1784 23060 1828
rect 25804 1784 25844 1828
rect 20995 1744 21004 1784
rect 21044 1744 21100 1784
rect 21140 1744 21175 1784
rect 23002 1744 23011 1784
rect 23051 1744 23060 1784
rect 23657 1744 23788 1784
rect 23828 1744 23837 1784
rect 24451 1744 24460 1784
rect 24500 1744 25844 1784
rect 28780 1784 28820 1903
rect 28876 1868 28916 1996
rect 30124 1952 30164 1996
rect 29705 1912 29836 1952
rect 29876 1912 29885 1952
rect 30115 1912 30124 1952
rect 30164 1912 30173 1952
rect 30857 1912 30988 1952
rect 31028 1912 31037 1952
rect 31171 1912 31180 1952
rect 31220 1912 31229 1952
rect 31180 1868 31220 1912
rect 28876 1828 29155 1868
rect 29195 1828 31220 1868
rect 28780 1744 30988 1784
rect 31028 1744 31037 1784
rect 4771 1660 4780 1700
rect 4820 1660 5059 1700
rect 5099 1660 5108 1700
rect 5609 1660 5740 1700
rect 5780 1660 5789 1700
rect 9004 1660 12980 1700
rect 13289 1660 13420 1700
rect 13460 1660 13469 1700
rect 13516 1660 14764 1700
rect 14804 1660 17972 1700
rect 18089 1660 18220 1700
rect 18260 1660 18269 1700
rect 18883 1660 18892 1700
rect 18932 1660 19084 1700
rect 19124 1660 19133 1700
rect 23177 1660 23308 1700
rect 23348 1660 23357 1700
rect 30665 1660 30796 1700
rect 30836 1660 30845 1700
rect 2083 1576 2092 1616
rect 2132 1576 5932 1616
rect 5972 1576 5981 1616
rect 6691 1576 6700 1616
rect 6740 1576 10732 1616
rect 10772 1576 10781 1616
rect 3103 1492 3112 1532
rect 3480 1492 3489 1532
rect 10877 1492 10886 1532
rect 11254 1492 11263 1532
rect 18651 1492 18660 1532
rect 19028 1492 19037 1532
rect 26425 1492 26434 1532
rect 26802 1492 26811 1532
rect 4867 1408 4876 1448
rect 4916 1408 5548 1448
rect 5588 1408 10388 1448
rect 13507 1408 13516 1448
rect 13556 1408 19660 1448
rect 19700 1408 19709 1448
rect 10348 1364 10388 1408
rect 8297 1324 8428 1364
rect 8468 1324 8477 1364
rect 10339 1324 10348 1364
rect 10388 1324 10397 1364
rect 11203 1324 11212 1364
rect 11252 1324 12556 1364
rect 12596 1324 12605 1364
rect 12713 1324 12844 1364
rect 12884 1324 12893 1364
rect 16867 1324 16876 1364
rect 16916 1324 17644 1364
rect 17684 1324 17693 1364
rect 19948 1324 23500 1364
rect 23540 1324 23549 1364
rect 24451 1324 24460 1364
rect 24500 1324 25228 1364
rect 25268 1324 25277 1364
rect 28483 1324 28492 1364
rect 28532 1324 29836 1364
rect 29876 1324 29885 1364
rect 2537 1240 2668 1280
rect 2708 1240 2717 1280
rect 4378 1240 4387 1280
rect 4427 1240 4436 1280
rect 4819 1240 4828 1280
rect 4868 1240 4972 1280
rect 5012 1240 5021 1280
rect 5155 1240 5164 1280
rect 5204 1240 6548 1280
rect 10531 1240 10540 1280
rect 10580 1240 11788 1280
rect 11828 1240 11837 1280
rect 13027 1240 13036 1280
rect 13076 1240 13324 1280
rect 13364 1240 15052 1280
rect 15092 1240 15101 1280
rect 18979 1240 18988 1280
rect 19028 1240 19180 1280
rect 19220 1240 19229 1280
rect 4396 1196 4436 1240
rect 6508 1196 6548 1240
rect 4396 1156 5059 1196
rect 5099 1156 5300 1196
rect 6499 1156 6508 1196
rect 6548 1156 6557 1196
rect 7555 1156 7564 1196
rect 7604 1156 7613 1196
rect 9100 1156 15860 1196
rect 16771 1156 16780 1196
rect 16820 1156 16829 1196
rect 18796 1156 19084 1196
rect 19124 1156 19133 1196
rect 5260 1112 5300 1156
rect 5827 1114 5836 1154
rect 5876 1145 6007 1154
rect 5876 1114 5923 1145
rect 3811 1072 3820 1112
rect 3860 1072 4204 1112
rect 4244 1072 4253 1112
rect 4378 1072 4387 1112
rect 4436 1072 4567 1112
rect 4675 1072 4684 1112
rect 4724 1072 4733 1112
rect 4788 1072 4876 1112
rect 4916 1072 4919 1112
rect 4959 1072 4968 1112
rect 5156 1072 5165 1112
rect 5205 1072 5214 1112
rect 5260 1072 5443 1112
rect 5483 1072 5492 1112
rect 5914 1105 5923 1114
rect 5963 1114 6007 1145
rect 5963 1105 5972 1114
rect 9100 1112 9140 1156
rect 5914 1104 5972 1105
rect 6874 1072 6883 1112
rect 6923 1072 8524 1112
rect 8564 1072 9140 1112
rect 9187 1072 9196 1112
rect 9236 1072 9245 1112
rect 9859 1072 9868 1112
rect 9908 1072 10147 1112
rect 10187 1072 10196 1112
rect 10723 1072 10732 1112
rect 10772 1072 10915 1112
rect 10955 1072 10964 1112
rect 11383 1072 11392 1112
rect 11432 1072 11444 1112
rect 11539 1072 11548 1112
rect 11588 1072 11596 1112
rect 11636 1072 12364 1112
rect 12404 1072 12413 1112
rect 12634 1072 12643 1112
rect 12683 1072 12692 1112
rect 12739 1072 12748 1112
rect 12788 1072 12940 1112
rect 12980 1072 12989 1112
rect 13036 1072 13175 1112
rect 13215 1072 13224 1112
rect 13306 1072 13315 1112
rect 13355 1072 13364 1112
rect 13411 1072 13420 1112
rect 13460 1072 13591 1112
rect 14275 1072 14284 1112
rect 14324 1072 14333 1112
rect 14458 1072 14467 1112
rect 14507 1072 14516 1112
rect 14681 1072 14764 1112
rect 14804 1072 14812 1112
rect 14852 1072 14861 1112
rect 14947 1072 14956 1112
rect 14996 1072 15052 1112
rect 15092 1072 15127 1112
rect 15820 1107 15860 1156
rect 18796 1112 18836 1156
rect 19948 1112 19988 1324
rect 20777 1240 20908 1280
rect 20948 1240 20957 1280
rect 21571 1240 21580 1280
rect 21620 1240 21676 1280
rect 21716 1240 21751 1280
rect 25027 1240 25036 1280
rect 25076 1240 25324 1280
rect 25364 1240 25373 1280
rect 23779 1156 23788 1196
rect 23828 1156 23837 1196
rect 24643 1156 24652 1196
rect 24692 1156 24701 1196
rect 25219 1156 25228 1196
rect 25268 1156 26851 1196
rect 26891 1156 26900 1196
rect 30307 1156 30316 1196
rect 30356 1156 30365 1196
rect 30778 1156 30787 1196
rect 30836 1156 30967 1196
rect 24652 1112 24692 1156
rect 26284 1112 26324 1156
rect 16012 1107 16099 1112
rect 15820 1072 16099 1107
rect 16139 1072 16148 1112
rect 18787 1072 18796 1112
rect 18836 1072 18845 1112
rect 18892 1072 18911 1112
rect 18951 1072 18960 1112
rect 19075 1072 19084 1112
rect 19124 1072 19988 1112
rect 20035 1072 20044 1112
rect 20084 1072 20093 1112
rect 20707 1072 20716 1112
rect 20756 1072 21475 1112
rect 21515 1072 21524 1112
rect 23098 1072 23107 1112
rect 23156 1072 23287 1112
rect 24067 1072 24076 1112
rect 24116 1072 24692 1112
rect 25843 1072 25852 1112
rect 25892 1072 25916 1112
rect 25961 1072 25996 1112
rect 26036 1072 26092 1112
rect 26132 1072 26141 1112
rect 26275 1072 26284 1112
rect 26324 1072 26333 1112
rect 27401 1072 27532 1112
rect 27572 1072 27581 1112
rect 30281 1072 30403 1112
rect 30452 1072 30461 1112
rect 4684 1028 4724 1072
rect 5164 1028 5204 1072
rect 4684 988 4820 1028
rect 5164 988 5644 1028
rect 5684 988 5693 1028
rect 5745 988 5754 1028
rect 5794 988 5932 1028
rect 5972 988 7220 1028
rect 4780 776 4820 988
rect 5242 904 5251 944
rect 5291 904 5300 944
rect 5417 904 5539 944
rect 5588 904 5597 944
rect 6019 904 6028 944
rect 6068 904 6076 944
rect 6116 904 6199 944
rect 5260 860 5300 904
rect 5260 820 6412 860
rect 6452 820 6461 860
rect 4343 736 4352 776
rect 4720 736 4729 776
rect 4780 736 5740 776
rect 5780 736 5789 776
rect 7180 692 7220 988
rect 9196 944 9236 1072
rect 10627 988 10636 1028
rect 10676 988 11020 1028
rect 11060 988 11069 1028
rect 11177 988 11226 1028
rect 11266 988 11308 1028
rect 11348 988 11357 1028
rect 8803 904 8812 944
rect 8852 904 9236 944
rect 9196 860 9236 904
rect 11404 860 11444 1072
rect 12652 1028 12692 1072
rect 12605 988 12652 1028
rect 12692 988 12701 1028
rect 13036 944 13076 1072
rect 13027 904 13036 944
rect 13076 904 13085 944
rect 13324 860 13364 1072
rect 13498 988 13507 1028
rect 13556 988 13687 1028
rect 9196 820 11444 860
rect 12547 820 12556 860
rect 12596 820 13364 860
rect 12117 736 12126 776
rect 12494 736 12503 776
rect 14284 692 14324 1072
rect 14476 1028 14516 1072
rect 15820 1067 16052 1072
rect 18892 1028 18932 1072
rect 20044 1028 20084 1072
rect 25876 1028 25916 1072
rect 14476 988 14708 1028
rect 14668 944 14708 988
rect 14371 904 14380 944
rect 14420 904 14429 944
rect 14650 904 14659 944
rect 14699 904 14708 944
rect 14956 988 15715 1028
rect 15755 988 15764 1028
rect 18211 988 18220 1028
rect 18260 988 18932 1028
rect 19747 988 19756 1028
rect 19796 988 20084 1028
rect 22714 988 22723 1028
rect 22763 988 23308 1028
rect 23348 988 23357 1028
rect 25876 988 26188 1028
rect 26228 988 26237 1028
rect 14380 860 14420 904
rect 14956 860 14996 988
rect 19756 944 19796 988
rect 18019 904 18028 944
rect 18068 904 19796 944
rect 21667 904 21676 944
rect 21716 904 21725 944
rect 21676 860 21716 904
rect 14380 820 14996 860
rect 15043 820 15052 860
rect 15092 820 21716 860
rect 19891 736 19900 776
rect 20268 736 20277 776
rect 27665 736 27674 776
rect 28042 736 28051 776
rect 7180 652 14324 692
<< via2 >>
rect 16396 28624 16436 28664
rect 13900 28540 13940 28580
rect 23308 28540 23348 28580
rect 30028 28540 30068 28580
rect 12364 28372 12404 28412
rect 17644 28372 17684 28412
rect 10060 28204 10100 28244
rect 20428 28204 20468 28244
rect 14668 28120 14708 28160
rect 21388 28120 21428 28160
rect 15436 28036 15476 28076
rect 20524 28036 20564 28076
rect 4352 27952 4720 27992
rect 12126 27952 12494 27992
rect 19900 27952 20268 27992
rect 27674 27952 28042 27992
rect 9292 27868 9332 27908
rect 11788 27868 11828 27908
rect 16204 27868 16244 27908
rect 21100 27868 21140 27908
rect 11596 27784 11636 27824
rect 17836 27784 17876 27824
rect 29260 27784 29300 27824
rect 8524 27700 8564 27740
rect 11692 27700 11732 27740
rect 23980 27700 24020 27740
rect 26956 27700 26996 27740
rect 28492 27700 28532 27740
rect 3628 27616 3659 27656
rect 3659 27616 3668 27656
rect 11596 27616 11627 27656
rect 11627 27616 11636 27656
rect 15148 27616 15188 27656
rect 17068 27616 17108 27656
rect 19084 27616 19124 27656
rect 20140 27616 20180 27656
rect 22732 27616 22763 27656
rect 22763 27616 22772 27656
rect 25612 27616 25652 27656
rect 25900 27616 25931 27656
rect 25931 27616 25940 27656
rect 3532 27532 3572 27572
rect 5740 27532 5780 27572
rect 6700 27532 6740 27572
rect 8236 27532 8276 27572
rect 9292 27532 9332 27572
rect 3148 27448 3188 27488
rect 15724 27532 15764 27572
rect 16780 27532 16811 27572
rect 16811 27532 16820 27572
rect 17740 27532 17780 27572
rect 24460 27532 24500 27572
rect 20812 27448 20852 27488
rect 27820 27532 27860 27572
rect 29356 27647 29396 27656
rect 29356 27616 29387 27647
rect 29387 27616 29396 27647
rect 28972 27532 29012 27572
rect 29452 27532 29492 27572
rect 29932 27532 29972 27572
rect 3724 27364 3764 27404
rect 7468 27364 7508 27404
rect 9676 27364 9716 27404
rect 10540 27364 10580 27404
rect 13324 27364 13364 27404
rect 13804 27364 13844 27404
rect 14476 27364 14516 27404
rect 14668 27364 14708 27404
rect 19660 27364 19700 27404
rect 30316 27448 30356 27488
rect 31084 27448 31124 27488
rect 25516 27364 25556 27404
rect 27148 27364 27188 27404
rect 28684 27364 28724 27404
rect 30412 27364 30452 27404
rect 20908 27280 20948 27320
rect 3112 27196 3480 27236
rect 10886 27196 11254 27236
rect 18660 27196 19028 27236
rect 8716 27112 8756 27152
rect 18124 27112 18164 27152
rect 24940 27112 24980 27152
rect 26434 27196 26802 27236
rect 3916 27028 3956 27068
rect 11692 27028 11732 27068
rect 17068 27028 17108 27068
rect 17740 27028 17780 27068
rect 20716 27028 20756 27068
rect 26956 27028 26996 27068
rect 30796 27028 30836 27068
rect 3532 26944 3572 26984
rect 3724 26944 3764 26984
rect 5548 26944 5588 26984
rect 6700 26944 6740 26984
rect 9292 26944 9332 26984
rect 13324 26944 13364 26984
rect 13708 26944 13748 26984
rect 15724 26944 15764 26984
rect 24460 26944 24500 26984
rect 26188 26944 26228 26984
rect 27820 26944 27860 26984
rect 8524 26860 8564 26900
rect 10828 26860 10868 26900
rect 12460 26860 12500 26900
rect 16780 26860 16820 26900
rect 19660 26860 19700 26900
rect 20812 26860 20852 26900
rect 23116 26860 23156 26900
rect 4876 26776 4916 26816
rect 6316 26776 6356 26816
rect 7468 26776 7508 26816
rect 12748 26776 12788 26816
rect 14380 26776 14420 26816
rect 16204 26776 16244 26816
rect 17068 26776 17108 26816
rect 20140 26776 20171 26816
rect 20171 26776 20180 26816
rect 24172 26776 24212 26816
rect 25516 26776 25556 26816
rect 26284 26776 26323 26816
rect 26323 26776 26324 26816
rect 27052 26776 27092 26816
rect 27436 26860 27476 26900
rect 28780 26860 28820 26900
rect 31084 26860 31124 26900
rect 27628 26776 27668 26816
rect 28492 26776 28532 26816
rect 30892 26776 30923 26816
rect 30923 26776 30932 26816
rect 4780 26692 4820 26732
rect 5452 26692 5492 26732
rect 6220 26692 6260 26732
rect 9196 26692 9236 26732
rect 7756 26608 7796 26648
rect 8620 26608 8660 26648
rect 4780 26524 4820 26564
rect 4352 26440 4720 26480
rect 3724 26188 3764 26228
rect 10252 26692 10292 26732
rect 12844 26608 12884 26648
rect 14668 26608 14708 26648
rect 10444 26524 10484 26564
rect 11404 26524 11444 26564
rect 23788 26692 23828 26732
rect 25708 26692 25739 26732
rect 25739 26692 25748 26732
rect 25996 26692 26036 26732
rect 27532 26692 27572 26732
rect 12126 26440 12494 26480
rect 12940 26440 12980 26480
rect 13804 26440 13844 26480
rect 16108 26440 16148 26480
rect 11980 26356 12020 26396
rect 16972 26356 17012 26396
rect 17164 26356 17204 26396
rect 18892 26356 18932 26396
rect 19276 26356 19316 26396
rect 23116 26608 23156 26648
rect 23596 26608 23635 26648
rect 23635 26608 23636 26648
rect 24076 26608 24116 26648
rect 19900 26440 20268 26480
rect 27340 26608 27380 26648
rect 25612 26524 25652 26564
rect 23404 26440 23444 26480
rect 27674 26440 28042 26480
rect 8236 26272 8276 26312
rect 8716 26272 8756 26312
rect 9676 26272 9707 26312
rect 9707 26272 9716 26312
rect 10156 26272 10196 26312
rect 11404 26272 11435 26312
rect 11435 26272 11444 26312
rect 11596 26272 11636 26312
rect 15148 26272 15188 26312
rect 17452 26272 17483 26312
rect 17483 26272 17492 26312
rect 18124 26272 18155 26312
rect 18155 26272 18164 26312
rect 19564 26272 19604 26312
rect 19948 26272 19988 26312
rect 23980 26272 24011 26312
rect 24011 26272 24020 26312
rect 26188 26272 26228 26312
rect 5836 26188 5876 26228
rect 9100 26188 9140 26228
rect 11884 26188 11924 26228
rect 12556 26188 12596 26228
rect 12844 26188 12875 26228
rect 12875 26188 12884 26228
rect 3628 26104 3659 26144
rect 3659 26104 3668 26144
rect 5068 26104 5108 26144
rect 5740 26104 5780 26144
rect 6220 26104 6260 26144
rect 8332 26104 8372 26144
rect 9196 26104 9197 26144
rect 9197 26104 9236 26144
rect 9964 26104 10004 26144
rect 17356 26188 17396 26228
rect 24076 26188 24116 26228
rect 24748 26188 24788 26228
rect 25996 26188 26036 26228
rect 26284 26188 26324 26228
rect 27052 26188 27092 26228
rect 10636 26104 10665 26144
rect 10665 26104 10676 26144
rect 11308 26104 11348 26144
rect 11980 26104 12020 26144
rect 12460 26104 12500 26144
rect 12652 26104 12691 26144
rect 12691 26104 12692 26144
rect 12940 26104 12980 26144
rect 14476 26104 14516 26144
rect 15820 26104 15860 26144
rect 16108 26104 16148 26144
rect 16588 26104 16595 26144
rect 16595 26104 16628 26144
rect 18028 26104 18068 26144
rect 18892 26135 18932 26144
rect 18892 26104 18932 26135
rect 5164 26020 5204 26060
rect 5548 26020 5588 26060
rect 8908 26020 8948 26060
rect 9292 26020 9332 26060
rect 11500 26020 11540 26060
rect 12844 26020 12884 26060
rect 13708 26020 13748 26060
rect 16204 26020 16244 26060
rect 9004 25936 9044 25976
rect 10060 25936 10100 25976
rect 10828 25936 10868 25976
rect 12748 25936 12788 25976
rect 16492 25936 16532 25976
rect 17548 25936 17588 25976
rect 18028 25936 18068 25976
rect 19468 26104 19508 26144
rect 19948 26104 19988 26144
rect 20716 26104 20756 26144
rect 21004 26104 21044 26144
rect 23884 26104 23913 26144
rect 23913 26104 23924 26144
rect 24172 26135 24212 26144
rect 24172 26104 24212 26135
rect 24652 26104 24692 26144
rect 25420 26104 25460 26144
rect 28684 26188 28724 26228
rect 20620 26020 20660 26060
rect 20812 26020 20835 26060
rect 20835 26020 20852 26060
rect 24844 26020 24884 26060
rect 25708 26020 25748 26060
rect 27628 26104 27668 26144
rect 28492 26104 28532 26144
rect 31180 26104 31220 26144
rect 26092 26020 26132 26060
rect 26956 26020 26996 26060
rect 27148 26020 27188 26060
rect 28012 26020 28052 26060
rect 30988 26020 31028 26060
rect 19852 25936 19892 25976
rect 22252 25936 22292 25976
rect 24940 25936 24980 25976
rect 25996 25936 26036 25976
rect 27244 25936 27284 25976
rect 27820 25936 27860 25976
rect 28780 25936 28820 25976
rect 30028 25936 30068 25976
rect 31084 25936 31124 25976
rect 8140 25852 8180 25892
rect 10444 25852 10484 25892
rect 11404 25852 11444 25892
rect 11980 25852 12020 25892
rect 19372 25852 19412 25892
rect 20140 25852 20180 25892
rect 26860 25852 26900 25892
rect 28396 25852 28427 25892
rect 28427 25852 28436 25892
rect 4204 25768 4244 25808
rect 11692 25768 11732 25808
rect 19180 25768 19220 25808
rect 27340 25768 27380 25808
rect 3112 25684 3480 25724
rect 8332 25684 8372 25724
rect 9868 25684 9908 25724
rect 10444 25684 10484 25724
rect 10886 25684 11254 25724
rect 15148 25684 15188 25724
rect 17068 25684 17108 25724
rect 18660 25684 19028 25724
rect 26434 25684 26802 25724
rect 26956 25684 26996 25724
rect 29932 25684 29972 25724
rect 17356 25600 17396 25640
rect 25804 25600 25844 25640
rect 28972 25600 29012 25640
rect 6316 25516 6356 25556
rect 10156 25516 10196 25556
rect 11308 25516 11348 25556
rect 12844 25516 12884 25556
rect 19564 25516 19604 25556
rect 19756 25516 19796 25556
rect 20332 25516 20372 25556
rect 23788 25516 23828 25556
rect 25612 25516 25652 25556
rect 26476 25516 26516 25556
rect 27244 25516 27284 25556
rect 5068 25432 5108 25472
rect 6892 25432 6932 25472
rect 10732 25432 10772 25472
rect 11500 25432 11540 25472
rect 13036 25432 13076 25472
rect 14668 25432 14708 25472
rect 19852 25432 19892 25472
rect 21196 25432 21236 25472
rect 23596 25432 23636 25472
rect 3052 25348 3092 25388
rect 5644 25348 5684 25388
rect 8908 25348 8948 25388
rect 9964 25348 10004 25388
rect 10540 25348 10580 25388
rect 11116 25348 11155 25388
rect 11155 25348 11156 25388
rect 2572 25264 2612 25304
rect 22252 25348 22292 25388
rect 23884 25348 23924 25388
rect 5260 25264 5300 25304
rect 5548 25264 5579 25304
rect 5579 25264 5588 25304
rect 5740 25264 5780 25304
rect 9004 25264 9044 25304
rect 9292 25264 9323 25304
rect 9323 25264 9332 25304
rect 10828 25264 10829 25304
rect 10829 25264 10868 25304
rect 11596 25264 11636 25304
rect 12652 25264 12663 25304
rect 12663 25264 12692 25304
rect 13324 25264 13364 25304
rect 14476 25264 14516 25304
rect 15340 25264 15380 25304
rect 16492 25264 16532 25304
rect 17356 25264 17387 25304
rect 17387 25264 17396 25304
rect 17548 25264 17588 25304
rect 18700 25264 18740 25304
rect 18892 25264 18932 25304
rect 19468 25264 19508 25304
rect 19852 25264 19892 25304
rect 20140 25264 20180 25304
rect 20620 25264 20651 25304
rect 20651 25264 20660 25304
rect 4780 25180 4820 25220
rect 4352 24928 4720 24968
rect 4780 24844 4820 24884
rect 5452 24844 5492 24884
rect 5836 25096 5876 25136
rect 6988 25096 7028 25136
rect 8140 25096 8171 25136
rect 8171 25096 8180 25136
rect 8524 25096 8564 25136
rect 25516 25432 25556 25472
rect 24556 25348 24596 25388
rect 22732 25264 22772 25304
rect 24748 25348 24788 25388
rect 24940 25348 24980 25388
rect 26092 25348 26132 25388
rect 26284 25348 26324 25388
rect 26668 25348 26708 25388
rect 26956 25348 26996 25388
rect 27820 25348 27860 25388
rect 28012 25348 28052 25388
rect 30316 25348 30356 25388
rect 25118 25299 25137 25304
rect 25137 25299 25158 25304
rect 25118 25264 25158 25299
rect 25900 25264 25940 25304
rect 26572 25264 26612 25304
rect 26860 25264 26900 25304
rect 28204 25264 28244 25304
rect 28684 25264 28724 25304
rect 30892 25264 30932 25304
rect 11980 25180 12020 25220
rect 16588 25180 16628 25220
rect 17932 25180 17972 25220
rect 18124 25180 18164 25220
rect 19276 25180 19316 25220
rect 23980 25180 24020 25220
rect 24940 25180 24980 25220
rect 25612 25180 25652 25220
rect 10156 25096 10196 25136
rect 11692 25096 11732 25136
rect 11884 25096 11924 25136
rect 16012 25096 16052 25136
rect 17644 25096 17684 25136
rect 18892 25096 18923 25136
rect 18923 25096 18932 25136
rect 9676 25012 9716 25052
rect 10924 25012 10964 25052
rect 11308 25012 11348 25052
rect 17356 25012 17396 25052
rect 18220 25012 18260 25052
rect 9868 24928 9908 24968
rect 11500 24928 11540 24968
rect 12126 24928 12494 24968
rect 14476 24928 14516 24968
rect 19900 24928 20268 24968
rect 4876 24676 4916 24716
rect 8332 24676 8372 24716
rect 8908 24676 8948 24716
rect 2188 24592 2228 24632
rect 4204 24592 4244 24632
rect 4396 24592 4436 24632
rect 4972 24592 5012 24632
rect 5164 24592 5195 24632
rect 5195 24592 5204 24632
rect 5644 24592 5675 24632
rect 5675 24592 5684 24632
rect 6220 24592 6251 24632
rect 6251 24592 6260 24632
rect 8716 24592 8741 24632
rect 8741 24592 8756 24632
rect 9004 24592 9044 24632
rect 10444 24760 10484 24800
rect 20332 24844 20372 24884
rect 15340 24760 15380 24800
rect 17548 24760 17588 24800
rect 18124 24760 18164 24800
rect 18892 24760 18932 24800
rect 20236 24760 20276 24800
rect 9964 24676 10004 24716
rect 10156 24676 10196 24716
rect 11596 24676 11636 24716
rect 18028 24676 18039 24716
rect 18039 24676 18068 24716
rect 18220 24676 18260 24716
rect 18988 24676 19028 24716
rect 9580 24592 9620 24632
rect 10924 24592 10955 24632
rect 10955 24592 10964 24632
rect 11404 24592 11444 24632
rect 11692 24592 11732 24632
rect 14380 24592 14420 24632
rect 14860 24592 14900 24632
rect 6892 24508 6932 24548
rect 8236 24508 8276 24548
rect 8524 24508 8564 24548
rect 9772 24508 9812 24548
rect 10252 24508 10292 24548
rect 10540 24508 10571 24548
rect 10571 24508 10580 24548
rect 1900 24424 1940 24464
rect 3052 24424 3092 24464
rect 5068 24424 5108 24464
rect 5644 24424 5684 24464
rect 5836 24424 5876 24464
rect 16108 24592 16148 24632
rect 16972 24592 16984 24632
rect 16984 24592 17012 24632
rect 17452 24592 17492 24632
rect 18412 24592 18452 24632
rect 19756 24592 19785 24632
rect 19785 24592 19796 24632
rect 20236 24592 20276 24632
rect 11116 24508 11147 24548
rect 11147 24508 11156 24548
rect 13036 24508 13076 24548
rect 15148 24508 15188 24548
rect 19084 24508 19124 24548
rect 19372 24508 19412 24548
rect 22828 25096 22868 25136
rect 24364 25096 24404 25136
rect 25132 25096 25172 25136
rect 25420 25096 25460 25136
rect 26284 25180 26324 25220
rect 26956 25180 26996 25220
rect 26476 25096 26516 25136
rect 26380 25012 26420 25052
rect 27674 24928 28042 24968
rect 26860 24844 26900 24884
rect 25036 24760 25076 24800
rect 21196 24676 21236 24716
rect 24940 24676 24980 24716
rect 25420 24676 25460 24716
rect 25804 24676 25844 24716
rect 22828 24592 22868 24632
rect 24364 24592 24373 24632
rect 24373 24592 24404 24632
rect 24556 24592 24596 24632
rect 24748 24592 24773 24632
rect 24773 24592 24788 24632
rect 25036 24592 25076 24632
rect 26380 24760 26420 24800
rect 26572 24760 26612 24800
rect 28684 24760 28724 24800
rect 26188 24676 26228 24716
rect 26764 24676 26804 24716
rect 27436 24676 27476 24716
rect 28396 24676 28436 24716
rect 25612 24592 25652 24632
rect 26956 24592 26996 24632
rect 27340 24592 27380 24632
rect 27724 24592 27764 24632
rect 29548 24592 29588 24632
rect 26668 24508 26708 24548
rect 28108 24508 28148 24548
rect 28396 24508 28436 24548
rect 31276 24508 31316 24548
rect 11500 24424 11540 24464
rect 11884 24424 11924 24464
rect 14188 24424 14228 24464
rect 17164 24424 17204 24464
rect 19180 24424 19220 24464
rect 22924 24424 22964 24464
rect 23212 24424 23252 24464
rect 24556 24424 24596 24464
rect 27532 24424 27572 24464
rect 29932 24424 29972 24464
rect 30604 24424 30644 24464
rect 3532 24340 3572 24380
rect 5356 24340 5396 24380
rect 10444 24340 10484 24380
rect 13900 24340 13940 24380
rect 15244 24340 15284 24380
rect 19084 24340 19124 24380
rect 21580 24340 21620 24380
rect 24652 24340 24692 24380
rect 25804 24340 25844 24380
rect 27148 24340 27179 24380
rect 27179 24340 27188 24380
rect 28780 24340 28820 24380
rect 3628 24256 3668 24296
rect 16972 24256 17012 24296
rect 22348 24256 22388 24296
rect 23212 24256 23252 24296
rect 24460 24256 24500 24296
rect 29452 24256 29492 24296
rect 3112 24172 3480 24212
rect 8620 24172 8660 24212
rect 10444 24172 10484 24212
rect 10886 24172 11254 24212
rect 1900 23836 1940 23876
rect 2572 23752 2603 23792
rect 2603 23752 2612 23792
rect 3532 23783 3572 23792
rect 3532 23752 3572 23783
rect 2188 23668 2228 23708
rect 3628 23584 3668 23624
rect 18660 24172 19028 24212
rect 24844 24172 24884 24212
rect 26434 24172 26802 24212
rect 5164 24088 5204 24128
rect 13420 24088 13460 24128
rect 20812 24088 20852 24128
rect 27340 24088 27380 24128
rect 5260 24004 5291 24044
rect 5291 24004 5300 24044
rect 10540 24004 10580 24044
rect 11692 24004 11732 24044
rect 16012 24004 16052 24044
rect 18412 24004 18452 24044
rect 19276 24004 19316 24044
rect 22732 24004 22772 24044
rect 26956 24004 26996 24044
rect 4396 23836 4436 23876
rect 7084 23920 7124 23960
rect 9100 23920 9140 23960
rect 9292 23920 9332 23960
rect 10828 23920 10868 23960
rect 4204 23752 4244 23792
rect 5548 23752 5588 23792
rect 7468 23752 7508 23792
rect 9004 23836 9044 23876
rect 10060 23836 10100 23876
rect 11884 23836 11924 23876
rect 12556 23836 12587 23876
rect 12587 23836 12596 23876
rect 18892 23951 18932 23960
rect 18892 23920 18900 23951
rect 18900 23920 18932 23951
rect 19084 23920 19124 23960
rect 19468 23920 19508 23960
rect 24556 23920 24596 23960
rect 25516 23920 25556 23960
rect 26572 23920 26612 23960
rect 27148 23920 27188 23960
rect 14380 23836 14420 23876
rect 15148 23836 15188 23876
rect 17164 23836 17204 23876
rect 20812 23836 20852 23876
rect 22924 23836 22964 23876
rect 9292 23752 9332 23792
rect 10444 23752 10484 23792
rect 10924 23752 10964 23792
rect 13900 23752 13940 23792
rect 14188 23752 14228 23792
rect 14860 23752 14900 23792
rect 15244 23752 15284 23792
rect 17932 23752 17972 23792
rect 18412 23752 18452 23792
rect 18988 23752 19028 23792
rect 19660 23752 19688 23792
rect 19688 23752 19700 23792
rect 22732 23752 22763 23792
rect 22763 23752 22772 23792
rect 24076 23752 24116 23792
rect 4780 23668 4820 23708
rect 4352 23416 4720 23456
rect 2188 23332 2228 23372
rect 4972 23668 5012 23708
rect 5356 23668 5396 23708
rect 8620 23668 8660 23708
rect 13612 23668 13652 23708
rect 20332 23668 20372 23708
rect 5260 23584 5300 23624
rect 8044 23584 8084 23624
rect 8332 23584 8372 23624
rect 8716 23584 8747 23624
rect 8747 23584 8756 23624
rect 10540 23584 10580 23624
rect 11212 23584 11252 23624
rect 12844 23584 12884 23624
rect 5260 23416 5300 23456
rect 11692 23416 11732 23456
rect 12126 23416 12494 23456
rect 4876 23164 4916 23204
rect 7852 23248 7892 23288
rect 10252 23248 10292 23288
rect 8908 23164 8948 23204
rect 10924 23248 10964 23288
rect 10540 23164 10580 23204
rect 11212 23164 11252 23204
rect 844 23080 884 23120
rect 3628 23080 3668 23120
rect 5932 23080 5963 23120
rect 5963 23080 5972 23120
rect 6220 23080 6260 23120
rect 7372 23080 7412 23120
rect 8044 23080 8084 23120
rect 8812 23080 8843 23120
rect 8843 23080 8852 23120
rect 11116 23080 11156 23120
rect 11500 23080 11540 23120
rect 12460 23164 12500 23204
rect 17932 23584 17972 23624
rect 19084 23584 19115 23624
rect 19115 23584 19124 23624
rect 22252 23584 22292 23624
rect 23308 23584 23339 23624
rect 23339 23584 23348 23624
rect 24940 23836 24980 23876
rect 28492 24004 28532 24044
rect 31276 24004 31316 24044
rect 28492 23836 28532 23876
rect 30028 23836 30068 23876
rect 24460 23752 24499 23792
rect 24499 23752 24500 23792
rect 24844 23752 24884 23792
rect 25804 23752 25844 23792
rect 26380 23752 26420 23792
rect 26860 23752 26900 23792
rect 27820 23752 27860 23792
rect 28300 23752 28340 23792
rect 28780 23752 28820 23792
rect 29356 23752 29387 23792
rect 29387 23752 29396 23792
rect 23596 23668 23636 23708
rect 23692 23584 23732 23624
rect 15820 23500 15860 23540
rect 22348 23500 22388 23540
rect 24556 23668 24596 23708
rect 25900 23668 25940 23708
rect 24652 23584 24692 23624
rect 26188 23584 26228 23624
rect 26572 23584 26603 23624
rect 26603 23584 26612 23624
rect 26860 23584 26900 23624
rect 27532 23584 27572 23624
rect 28684 23584 28724 23624
rect 19900 23416 20268 23456
rect 20428 23416 20468 23456
rect 25516 23416 25556 23456
rect 26092 23416 26132 23456
rect 27674 23416 28042 23456
rect 24076 23332 24116 23372
rect 24460 23332 24500 23372
rect 24940 23332 24980 23372
rect 16588 23248 16628 23288
rect 17932 23248 17972 23288
rect 20332 23248 20372 23288
rect 23596 23248 23636 23288
rect 26956 23248 26996 23288
rect 29356 23248 29396 23288
rect 30988 23248 31028 23288
rect 12940 23164 12980 23204
rect 16108 23164 16148 23204
rect 18892 23164 18932 23204
rect 19276 23164 19316 23204
rect 24364 23164 24404 23204
rect 25324 23164 25364 23204
rect 25996 23164 26036 23204
rect 27148 23164 27188 23204
rect 27436 23164 27476 23204
rect 30508 23164 30548 23204
rect 4300 22996 4340 23036
rect 5548 22996 5588 23036
rect 7084 22996 7124 23036
rect 7468 22996 7508 23036
rect 9100 22996 9140 23036
rect 10444 22996 10484 23036
rect 2092 22912 2132 22952
rect 7852 22912 7892 22952
rect 11020 22912 11060 22952
rect 11692 22912 11732 22952
rect 12556 23080 12557 23120
rect 12557 23080 12596 23120
rect 13612 23080 13643 23120
rect 13643 23080 13652 23120
rect 16012 23080 16052 23120
rect 16972 23080 17012 23120
rect 17356 23080 17396 23120
rect 17644 23111 17684 23120
rect 17644 23080 17675 23111
rect 17675 23080 17684 23111
rect 17932 23080 17972 23120
rect 18412 23080 18452 23120
rect 18988 23080 19028 23120
rect 19180 23080 19220 23120
rect 20332 23080 20372 23120
rect 20908 23080 20948 23120
rect 22252 23080 22292 23120
rect 23692 23080 23723 23120
rect 23723 23080 23732 23120
rect 24460 23080 24500 23120
rect 24652 23080 24683 23120
rect 24683 23080 24692 23120
rect 24940 23080 24980 23120
rect 25516 23080 25547 23120
rect 25547 23080 25556 23120
rect 11980 22996 12020 23036
rect 14668 22996 14708 23036
rect 19372 22996 19412 23036
rect 12460 22912 12500 22952
rect 26860 23080 26876 23120
rect 26876 23080 26900 23120
rect 29356 23080 29387 23120
rect 29387 23080 29396 23120
rect 21100 22996 21140 23036
rect 24556 22996 24596 23036
rect 24748 22912 24788 22952
rect 25996 22996 26036 23036
rect 26380 22996 26420 23036
rect 26668 22996 26708 23036
rect 27340 22996 27380 23036
rect 3628 22828 3668 22868
rect 8332 22828 8372 22868
rect 16780 22828 16820 22868
rect 19564 22828 19604 22868
rect 20332 22828 20372 22868
rect 21772 22828 21812 22868
rect 25228 22828 25268 22868
rect 10636 22744 10676 22784
rect 25804 22828 25844 22868
rect 27244 22828 27284 22868
rect 29932 22996 29972 23036
rect 28972 22744 29012 22784
rect 30796 22744 30836 22784
rect 3112 22660 3480 22700
rect 10886 22660 11254 22700
rect 18660 22660 19028 22700
rect 26434 22660 26802 22700
rect 30124 22660 30164 22700
rect 12076 22576 12116 22616
rect 14476 22576 14516 22616
rect 27628 22576 27668 22616
rect 28204 22576 28244 22616
rect 30220 22576 30260 22616
rect 844 22492 884 22532
rect 7660 22492 7700 22532
rect 12748 22492 12788 22532
rect 18604 22492 18644 22532
rect 19372 22492 19412 22532
rect 25228 22492 25268 22532
rect 6028 22408 6068 22448
rect 6508 22408 6548 22448
rect 9676 22408 9716 22448
rect 10636 22408 10676 22448
rect 11404 22408 11444 22448
rect 12844 22408 12884 22448
rect 19276 22408 19316 22448
rect 19756 22408 19796 22448
rect 2092 22324 2132 22364
rect 4300 22324 4340 22364
rect 8620 22324 8660 22364
rect 12076 22324 12116 22364
rect 12460 22324 12500 22364
rect 25324 22408 25364 22448
rect 27052 22408 27092 22448
rect 19084 22324 19124 22364
rect 21772 22324 21812 22364
rect 24844 22324 24884 22364
rect 26188 22324 26228 22364
rect 27532 22324 27572 22364
rect 28396 22324 28436 22364
rect 30220 22324 30260 22364
rect 30796 22324 30836 22364
rect 2572 22240 2612 22280
rect 3628 22240 3659 22280
rect 3659 22240 3668 22280
rect 4972 22240 5012 22280
rect 5548 22240 5588 22280
rect 6028 22240 6068 22280
rect 8044 22240 8084 22280
rect 8332 22240 8372 22280
rect 8716 22240 8756 22280
rect 11308 22240 11348 22280
rect 11788 22240 11828 22280
rect 12364 22240 12404 22280
rect 13324 22240 13364 22280
rect 15244 22240 15284 22280
rect 16108 22240 16139 22280
rect 16139 22240 16148 22280
rect 19180 22240 19220 22280
rect 21100 22240 21140 22280
rect 21964 22240 22004 22280
rect 22252 22240 22292 22280
rect 23692 22240 23732 22280
rect 24460 22240 24500 22280
rect 25132 22240 25172 22280
rect 26092 22240 26132 22280
rect 27724 22240 27764 22280
rect 28108 22240 28148 22280
rect 29452 22240 29492 22280
rect 30124 22240 30164 22280
rect 31084 22240 31124 22280
rect 8908 22156 8948 22196
rect 5644 22072 5684 22112
rect 9292 22072 9332 22112
rect 9964 22072 9995 22112
rect 9995 22072 10004 22112
rect 10156 22072 10196 22112
rect 12652 22156 12692 22196
rect 12844 22156 12884 22196
rect 13036 22156 13076 22196
rect 17644 22156 17684 22196
rect 20908 22156 20948 22196
rect 21484 22156 21524 22196
rect 22060 22156 22100 22196
rect 23980 22156 24020 22196
rect 25900 22156 25940 22196
rect 26188 22156 26228 22196
rect 27436 22156 27476 22196
rect 18604 22072 18635 22112
rect 18635 22072 18644 22112
rect 20620 22072 20660 22112
rect 22540 22072 22580 22112
rect 22924 22072 22964 22112
rect 23692 22072 23723 22112
rect 23723 22072 23732 22112
rect 25804 22072 25844 22112
rect 6412 21988 6452 22028
rect 13228 21988 13268 22028
rect 28780 22072 28820 22112
rect 23500 21988 23540 22028
rect 27340 21988 27380 22028
rect 31084 21988 31124 22028
rect 4352 21904 4720 21944
rect 12126 21904 12494 21944
rect 19900 21904 20268 21944
rect 25612 21904 25652 21944
rect 27674 21904 28042 21944
rect 28396 21904 28436 21944
rect 30412 21820 30452 21860
rect 364 21736 404 21776
rect 11692 21736 11732 21776
rect 12748 21736 12788 21776
rect 13132 21736 13172 21776
rect 17740 21736 17780 21776
rect 4972 21652 5012 21692
rect 5644 21652 5684 21692
rect 652 21568 692 21608
rect 2860 21568 2900 21608
rect 4108 21568 4148 21608
rect 4012 21484 4052 21524
rect 4684 21568 4724 21608
rect 8812 21568 8852 21608
rect 21964 21736 22004 21776
rect 22252 21736 22292 21776
rect 25228 21736 25268 21776
rect 26092 21736 26132 21776
rect 27340 21736 27380 21776
rect 28972 21736 29012 21776
rect 29452 21736 29492 21776
rect 30220 21736 30260 21776
rect 30892 21736 30932 21776
rect 19852 21652 19892 21692
rect 20140 21652 20180 21692
rect 23980 21652 24020 21692
rect 9388 21568 9428 21608
rect 11212 21568 11252 21608
rect 11500 21568 11540 21608
rect 4972 21484 5012 21524
rect 5356 21484 5396 21524
rect 6508 21484 6548 21524
rect 11692 21568 11732 21608
rect 13036 21568 13076 21608
rect 13324 21568 13364 21608
rect 13612 21568 13652 21608
rect 16108 21568 16148 21608
rect 17644 21568 17675 21608
rect 17675 21568 17684 21608
rect 18988 21568 19028 21608
rect 19276 21568 19316 21608
rect 19948 21568 19988 21608
rect 21580 21568 21620 21608
rect 22060 21568 22091 21608
rect 22091 21568 22100 21608
rect 22924 21568 22964 21608
rect 24652 21568 24692 21608
rect 26380 21652 26420 21692
rect 26860 21652 26900 21692
rect 28108 21652 28148 21692
rect 28492 21652 28532 21692
rect 30028 21652 30068 21692
rect 9964 21484 10004 21524
rect 10732 21484 10772 21524
rect 11308 21484 11348 21524
rect 16492 21484 16523 21524
rect 16523 21484 16532 21524
rect 17068 21484 17099 21524
rect 17099 21484 17108 21524
rect 17548 21484 17588 21524
rect 17836 21484 17867 21524
rect 17867 21484 17876 21524
rect 2668 21400 2708 21440
rect 5164 21400 5204 21440
rect 25516 21568 25556 21608
rect 22348 21484 22388 21524
rect 9004 21400 9044 21440
rect 10444 21400 10484 21440
rect 11404 21400 11444 21440
rect 11980 21400 12020 21440
rect 12364 21400 12404 21440
rect 14476 21400 14516 21440
rect 19756 21400 19796 21440
rect 22444 21400 22484 21440
rect 2764 21316 2804 21356
rect 7276 21316 7316 21356
rect 7948 21316 7988 21356
rect 8332 21316 8372 21356
rect 9388 21316 9428 21356
rect 9676 21316 9707 21356
rect 9707 21316 9716 21356
rect 16396 21316 16436 21356
rect 19180 21316 19220 21356
rect 21004 21316 21044 21356
rect 1996 21232 2036 21272
rect 24748 21232 24788 21272
rect 3112 21148 3480 21188
rect 4684 21148 4724 21188
rect 9004 21148 9044 21188
rect 10886 21148 11254 21188
rect 11404 21148 11444 21188
rect 16396 21148 16436 21188
rect 18660 21148 19028 21188
rect 4108 21064 4148 21104
rect 12364 21064 12404 21104
rect 24652 21064 24692 21104
rect 652 20980 692 21020
rect 25804 21400 25844 21440
rect 25708 21316 25748 21356
rect 27436 21568 27476 21608
rect 27628 21568 27668 21608
rect 28588 21568 28628 21608
rect 26284 21484 26324 21524
rect 26572 21484 26612 21524
rect 27340 21484 27380 21524
rect 27148 21400 27188 21440
rect 25996 21316 26036 21356
rect 28012 21316 28052 21356
rect 29644 21568 29684 21608
rect 30508 21568 30548 21608
rect 30988 21568 31028 21608
rect 28300 21484 28340 21524
rect 28780 21484 28820 21524
rect 30220 21400 30260 21440
rect 28780 21316 28820 21356
rect 27436 21232 27476 21272
rect 30124 21232 30164 21272
rect 26434 21148 26802 21188
rect 4972 20980 5012 21020
rect 11212 20980 11252 21020
rect 11500 20980 11540 21020
rect 13612 20980 13652 21020
rect 15052 20980 15092 21020
rect 16108 20980 16148 21020
rect 23404 20980 23444 21020
rect 26572 20980 26612 21020
rect 26764 20980 26804 21020
rect 27436 20980 27476 21020
rect 28204 20980 28244 21020
rect 28588 20980 28628 21020
rect 29644 20980 29684 21020
rect 11404 20896 11444 20936
rect 11980 20896 12020 20936
rect 16588 20896 16628 20936
rect 2668 20812 2708 20852
rect 5740 20812 5780 20852
rect 7180 20812 7220 20852
rect 7852 20812 7892 20852
rect 9004 20812 9044 20852
rect 11692 20812 11732 20852
rect 14476 20812 14516 20852
rect 15148 20812 15188 20852
rect 16492 20812 16532 20852
rect 17260 20812 17300 20852
rect 17548 20812 17588 20852
rect 19276 20812 19315 20852
rect 19315 20812 19316 20852
rect 20140 20812 20180 20852
rect 20524 20812 20564 20852
rect 21004 20812 21035 20852
rect 21035 20812 21044 20852
rect 2572 20728 2603 20768
rect 2603 20728 2612 20768
rect 2860 20728 2900 20768
rect 3148 20728 3188 20768
rect 3436 20728 3476 20768
rect 4204 20728 4244 20768
rect 4684 20728 4724 20768
rect 5260 20728 5300 20768
rect 5452 20728 5492 20768
rect 7276 20728 7316 20768
rect 8044 20728 8051 20768
rect 8051 20728 8084 20768
rect 10444 20728 10484 20768
rect 10732 20728 10772 20768
rect 11596 20728 11636 20768
rect 16396 20728 16436 20768
rect 17932 20728 17971 20768
rect 17971 20728 17972 20768
rect 19852 20728 19892 20768
rect 20428 20728 20468 20768
rect 1228 20644 1268 20684
rect 2956 20644 2987 20684
rect 2987 20644 2996 20684
rect 4300 20644 4331 20684
rect 4331 20644 4340 20684
rect 5164 20644 5204 20684
rect 6316 20644 6356 20684
rect 11020 20644 11060 20684
rect 12748 20644 12788 20684
rect 12940 20644 12980 20684
rect 14380 20644 14420 20684
rect 15916 20644 15956 20684
rect 22444 20812 22484 20852
rect 24940 20896 24980 20936
rect 26092 20896 26132 20936
rect 24172 20812 24212 20852
rect 25804 20812 25844 20852
rect 26476 20896 26516 20936
rect 27244 20812 27284 20852
rect 25516 20728 25556 20768
rect 25900 20728 25940 20768
rect 28012 20812 28052 20852
rect 28300 20812 28340 20852
rect 28588 20812 28628 20852
rect 28780 20812 28820 20852
rect 30604 20812 30644 20852
rect 26476 20728 26514 20768
rect 26514 20728 26516 20768
rect 17644 20644 17684 20684
rect 18988 20644 19028 20684
rect 19948 20644 19988 20684
rect 20620 20644 20660 20684
rect 20908 20644 20948 20684
rect 5548 20560 5588 20600
rect 8140 20560 8180 20600
rect 10924 20560 10955 20600
rect 10955 20560 10964 20600
rect 24556 20644 24596 20684
rect 27820 20728 27860 20768
rect 28492 20728 28532 20768
rect 30220 20728 30260 20768
rect 27436 20644 27476 20684
rect 14092 20560 14132 20600
rect 22636 20560 22676 20600
rect 25036 20560 25076 20600
rect 25612 20560 25652 20600
rect 25804 20560 25844 20600
rect 27052 20560 27092 20600
rect 27340 20560 27380 20600
rect 28300 20560 28340 20600
rect 11884 20476 11924 20516
rect 460 20392 500 20432
rect 4352 20392 4720 20432
rect 9004 20392 9044 20432
rect 12126 20392 12494 20432
rect 19900 20392 20268 20432
rect 27674 20392 28042 20432
rect 1324 20308 1364 20348
rect 4108 20308 4148 20348
rect 11980 20308 12020 20348
rect 19180 20308 19220 20348
rect 24556 20308 24596 20348
rect 24748 20308 24788 20348
rect 1420 20224 1460 20264
rect 10924 20224 10964 20264
rect 13420 20224 13451 20264
rect 13451 20224 13460 20264
rect 14476 20224 14516 20264
rect 17068 20224 17108 20264
rect 17260 20224 17300 20264
rect 17836 20224 17876 20264
rect 20908 20224 20948 20264
rect 25228 20308 25268 20348
rect 26764 20308 26804 20348
rect 27052 20308 27092 20348
rect 26668 20224 26708 20264
rect 27148 20224 27179 20264
rect 27179 20224 27188 20264
rect 27436 20224 27476 20264
rect 31180 20224 31220 20264
rect 940 20140 980 20180
rect 3436 20140 3476 20180
rect 3820 20140 3860 20180
rect 6700 20140 6740 20180
rect 8524 20140 8564 20180
rect 10060 20140 10100 20180
rect 13516 20140 13556 20180
rect 14380 20140 14411 20180
rect 14411 20140 14420 20180
rect 18988 20140 19028 20180
rect 23116 20140 23156 20180
rect 1804 20056 1844 20096
rect 2284 20056 2324 20096
rect 2668 20056 2708 20096
rect 2860 20056 2900 20096
rect 3628 20056 3668 20096
rect 3916 20056 3956 20096
rect 4300 20056 4340 20096
rect 4492 20056 4532 20096
rect 5164 20056 5195 20096
rect 5195 20056 5204 20096
rect 6988 20056 7028 20096
rect 7276 20056 7316 20096
rect 7756 20056 7787 20096
rect 7787 20056 7796 20096
rect 9004 20056 9035 20096
rect 9035 20056 9044 20096
rect 1708 19972 1748 20012
rect 3340 19972 3380 20012
rect 3724 19972 3764 20012
rect 4204 19972 4244 20012
rect 4972 19972 5012 20012
rect 5548 19972 5588 20012
rect 6796 19972 6836 20012
rect 7564 19972 7604 20012
rect 8140 19972 8180 20012
rect 8716 19972 8756 20012
rect 1228 19888 1268 19928
rect 2956 19888 2996 19928
rect 4876 19888 4916 19928
rect 1324 19804 1364 19844
rect 2380 19804 2420 19844
rect 5836 19888 5876 19928
rect 6124 19888 6164 19928
rect 10732 20056 10772 20096
rect 11020 20056 11051 20096
rect 11051 20056 11060 20096
rect 11212 20056 11252 20096
rect 13228 20056 13259 20096
rect 13259 20056 13268 20096
rect 15052 20056 15092 20096
rect 15820 20056 15860 20096
rect 16396 20056 16436 20096
rect 16588 20056 16619 20096
rect 16619 20056 16628 20096
rect 17107 20056 17147 20096
rect 17452 20056 17492 20096
rect 18124 20056 18164 20096
rect 18508 20087 18548 20096
rect 18508 20056 18539 20087
rect 18539 20056 18548 20087
rect 7180 19888 7220 19928
rect 8044 19888 8084 19928
rect 8428 19888 8468 19928
rect 11404 19972 11444 20012
rect 13708 19972 13748 20012
rect 10732 19888 10772 19928
rect 13804 19888 13844 19928
rect 6412 19804 6452 19844
rect 6988 19804 7028 19844
rect 11500 19804 11540 19844
rect 13036 19804 13076 19844
rect 748 19720 788 19760
rect 2860 19720 2900 19760
rect 4588 19720 4628 19760
rect 3112 19636 3480 19676
rect 844 19552 884 19592
rect 17356 19972 17387 20012
rect 17387 19972 17396 20012
rect 25996 20140 26036 20180
rect 27340 20140 27380 20180
rect 27628 20140 27668 20180
rect 28204 20140 28244 20180
rect 19276 20056 19316 20096
rect 19852 20056 19892 20096
rect 20428 20056 20468 20096
rect 20236 19972 20276 20012
rect 25036 20056 25067 20096
rect 25067 20056 25076 20096
rect 25324 20056 25355 20096
rect 25355 20056 25364 20096
rect 25708 20056 25739 20096
rect 25739 20056 25748 20096
rect 27532 20056 27572 20096
rect 29452 20056 29492 20096
rect 30316 20056 30356 20096
rect 30508 20087 30548 20096
rect 30508 20056 30539 20087
rect 30539 20056 30548 20087
rect 20524 19972 20564 20012
rect 20908 19972 20948 20012
rect 26572 19972 26612 20012
rect 27052 19972 27092 20012
rect 28876 19972 28916 20012
rect 30892 19972 30932 20012
rect 17260 19888 17300 19928
rect 19660 19888 19700 19928
rect 20716 19888 20756 19928
rect 17644 19804 17684 19844
rect 19468 19804 19508 19844
rect 20236 19804 20276 19844
rect 21100 19804 21140 19844
rect 17452 19720 17492 19760
rect 10886 19636 11254 19676
rect 11596 19636 11636 19676
rect 11980 19636 12020 19676
rect 16972 19636 17012 19676
rect 18660 19636 19028 19676
rect 25036 19888 25076 19928
rect 26284 19888 26324 19928
rect 24748 19804 24788 19844
rect 26434 19636 26802 19676
rect 2956 19468 2996 19508
rect 4204 19468 4244 19508
rect 5164 19468 5204 19508
rect 7276 19468 7316 19508
rect 7756 19468 7796 19508
rect 9772 19468 9812 19508
rect 11884 19468 11924 19508
rect 16396 19468 16436 19508
rect 17356 19468 17396 19508
rect 17644 19468 17675 19508
rect 17675 19468 17684 19508
rect 1324 19384 1364 19424
rect 1804 19384 1844 19424
rect 3628 19384 3668 19424
rect 4492 19384 4532 19424
rect 6988 19384 7028 19424
rect 1132 19300 1172 19340
rect 1708 19300 1748 19340
rect 3148 19300 3171 19340
rect 3171 19300 3188 19340
rect 3916 19300 3956 19340
rect 4780 19300 4820 19340
rect 5836 19300 5876 19340
rect 7660 19384 7700 19424
rect 10924 19384 10964 19424
rect 11980 19384 12020 19424
rect 14956 19384 14996 19424
rect 19660 19384 19700 19424
rect 6316 19300 6356 19340
rect 8140 19300 8180 19340
rect 8908 19300 8931 19340
rect 8931 19300 8948 19340
rect 9772 19300 9812 19340
rect 10732 19300 10772 19340
rect 11308 19300 11348 19340
rect 11500 19300 11540 19340
rect 13228 19300 13268 19340
rect 14860 19300 14900 19340
rect 17260 19300 17300 19340
rect 18508 19300 18548 19340
rect 2092 19216 2132 19256
rect 2764 19216 2804 19256
rect 4492 19216 4532 19256
rect 5740 19216 5780 19256
rect 6604 19216 6644 19256
rect 7852 19216 7883 19256
rect 7883 19216 7892 19256
rect 9292 19216 9320 19256
rect 9320 19216 9332 19256
rect 9964 19216 10004 19256
rect 11404 19216 11444 19256
rect 12460 19216 12500 19256
rect 13516 19216 13556 19256
rect 13804 19216 13844 19256
rect 14476 19216 14516 19256
rect 1516 19132 1556 19172
rect 1900 19132 1940 19172
rect 2188 19132 2228 19172
rect 2380 19132 2420 19172
rect 2860 19132 2900 19172
rect 3052 19132 3092 19172
rect 3340 19132 3380 19172
rect 3820 19132 3860 19172
rect 5548 19132 5588 19172
rect 6028 19132 6059 19172
rect 6059 19132 6068 19172
rect 1036 19048 1076 19088
rect 6700 19048 6740 19088
rect 1804 18964 1844 19004
rect 8716 19132 8756 19172
rect 9004 19132 9044 19172
rect 11980 19132 12020 19172
rect 12556 19132 12596 19172
rect 13132 19132 13172 19172
rect 7564 19048 7604 19088
rect 8812 19048 8852 19088
rect 6892 18964 6932 19004
rect 7276 18964 7316 19004
rect 1612 18880 1652 18920
rect 4352 18880 4720 18920
rect 9004 18880 9044 18920
rect 15820 19216 15860 19256
rect 15052 19132 15092 19172
rect 10924 19048 10964 19088
rect 14476 19048 14516 19088
rect 15148 19048 15188 19088
rect 15436 19048 15476 19088
rect 15724 19048 15764 19088
rect 19756 19300 19796 19340
rect 20524 19384 20564 19424
rect 21196 19384 21236 19424
rect 21868 19384 21908 19424
rect 24844 19384 24884 19424
rect 20812 19300 20852 19340
rect 21100 19300 21140 19340
rect 22828 19300 22868 19340
rect 23500 19300 23540 19340
rect 24652 19300 24692 19340
rect 17548 19216 17588 19256
rect 18220 19216 18260 19256
rect 19180 19216 19211 19256
rect 19211 19216 19220 19256
rect 19468 19216 19479 19256
rect 19479 19216 19508 19256
rect 20908 19216 20948 19256
rect 21388 19216 21428 19256
rect 23692 19216 23730 19256
rect 23730 19216 23732 19256
rect 24172 19216 24203 19256
rect 24203 19216 24212 19256
rect 25324 19216 25364 19256
rect 16876 19132 16916 19172
rect 17164 19132 17204 19172
rect 17356 19132 17396 19172
rect 18988 19132 19028 19172
rect 19372 19132 19412 19172
rect 28780 19804 28820 19844
rect 30316 19468 30356 19508
rect 28108 19300 28148 19340
rect 29836 19300 29876 19340
rect 30892 19216 30923 19256
rect 30923 19216 30932 19256
rect 25036 19132 25076 19172
rect 26092 19132 26132 19172
rect 27340 19132 27380 19172
rect 28300 19132 28340 19172
rect 28492 19132 28532 19172
rect 16108 19048 16148 19088
rect 16684 19048 16724 19088
rect 17452 19048 17492 19088
rect 17644 19048 17684 19088
rect 19276 19048 19307 19088
rect 19307 19048 19316 19088
rect 20908 19048 20948 19088
rect 23404 19048 23435 19088
rect 23435 19048 23444 19088
rect 24076 19079 24116 19088
rect 24076 19048 24107 19079
rect 24107 19048 24116 19079
rect 24748 19048 24779 19088
rect 24779 19048 24788 19088
rect 27436 19048 27476 19088
rect 28588 19048 28628 19088
rect 10828 18964 10868 19004
rect 11404 18964 11444 19004
rect 14572 18964 14612 19004
rect 11692 18880 11732 18920
rect 12126 18880 12494 18920
rect 19900 18880 20268 18920
rect 76 18796 116 18836
rect 2092 18796 2132 18836
rect 3148 18796 3188 18836
rect 1132 18712 1172 18752
rect 1900 18712 1931 18752
rect 1931 18712 1940 18752
rect 27052 18964 27092 19004
rect 27674 18880 28042 18920
rect 2764 18712 2804 18752
rect 4204 18712 4244 18752
rect 4972 18712 5012 18752
rect 5740 18712 5780 18752
rect 6892 18712 6932 18752
rect 8140 18712 8180 18752
rect 8908 18712 8939 18752
rect 8939 18712 8948 18752
rect 9292 18712 9332 18752
rect 11308 18712 11348 18752
rect 13420 18712 13460 18752
rect 14476 18712 14516 18752
rect 16684 18712 16724 18752
rect 17932 18712 17963 18752
rect 17963 18712 17972 18752
rect 18220 18712 18260 18752
rect 19372 18712 19403 18752
rect 19403 18712 19412 18752
rect 20236 18712 20276 18752
rect 27148 18712 27188 18752
rect 28492 18712 28532 18752
rect 29452 18712 29492 18752
rect 3724 18628 3764 18668
rect 4780 18628 4820 18668
rect 2092 18544 2132 18584
rect 1228 18460 1259 18500
rect 1259 18460 1268 18500
rect 5644 18628 5684 18668
rect 5932 18628 5972 18668
rect 7660 18628 7700 18668
rect 8812 18628 8838 18668
rect 8838 18628 8852 18668
rect 9004 18628 9044 18668
rect 10828 18628 10868 18668
rect 11980 18628 12020 18668
rect 16876 18628 16916 18668
rect 19468 18628 19508 18668
rect 20812 18628 20852 18668
rect 21388 18628 21428 18668
rect 23692 18628 23732 18668
rect 24460 18628 24491 18668
rect 24491 18628 24500 18668
rect 27436 18628 27476 18668
rect 28780 18628 28820 18668
rect 2668 18544 2708 18584
rect 2956 18544 2996 18584
rect 4300 18575 4340 18584
rect 4300 18544 4340 18575
rect 1708 18460 1739 18500
rect 1739 18460 1748 18500
rect 2284 18460 2307 18500
rect 2307 18460 2324 18500
rect 2764 18460 2804 18500
rect 4684 18460 4724 18500
rect 5068 18460 5099 18500
rect 5099 18460 5108 18500
rect 2092 18292 2132 18332
rect 4012 18292 4043 18332
rect 4043 18292 4052 18332
rect 2188 18208 2228 18248
rect 3112 18124 3480 18164
rect 6028 18460 6068 18500
rect 6604 18544 6644 18584
rect 6892 18544 6932 18584
rect 7180 18544 7220 18584
rect 7564 18544 7595 18584
rect 7595 18544 7604 18584
rect 8140 18544 8180 18584
rect 6220 18460 6260 18500
rect 6508 18460 6548 18500
rect 7372 18460 7412 18500
rect 11212 18544 11252 18584
rect 11788 18544 11828 18584
rect 13132 18544 13172 18584
rect 13708 18544 13748 18584
rect 14476 18544 14516 18584
rect 14860 18544 14900 18584
rect 16684 18544 16724 18584
rect 8812 18460 8852 18500
rect 9100 18460 9140 18500
rect 11404 18460 11444 18500
rect 11692 18460 11732 18500
rect 16108 18460 16148 18500
rect 7756 18376 7796 18416
rect 15916 18376 15956 18416
rect 6316 18292 6356 18332
rect 7660 18292 7700 18332
rect 6796 18208 6836 18248
rect 11020 18292 11060 18332
rect 13612 18292 13652 18332
rect 14764 18292 14804 18332
rect 13516 18208 13556 18248
rect 10886 18124 11254 18164
rect 4972 18040 5012 18080
rect 5164 18040 5204 18080
rect 12844 18040 12884 18080
rect 1420 17956 1451 17996
rect 1451 17956 1460 17996
rect 1708 17956 1748 17996
rect 17836 18544 17867 18584
rect 17867 18544 17876 18584
rect 18124 18544 18135 18584
rect 18135 18544 18164 18584
rect 16492 18460 16532 18500
rect 17068 18460 17108 18500
rect 17356 18460 17396 18500
rect 17548 18460 17588 18500
rect 18028 18460 18068 18500
rect 18988 18544 19028 18584
rect 20236 18544 20276 18584
rect 21004 18544 21044 18584
rect 23500 18544 23540 18584
rect 24748 18544 24788 18584
rect 26956 18544 26987 18584
rect 26987 18544 26996 18584
rect 28108 18544 28115 18584
rect 28115 18544 28148 18584
rect 28876 18544 28916 18584
rect 30892 18544 30923 18584
rect 30923 18544 30932 18584
rect 18316 18460 18356 18500
rect 19276 18460 19316 18500
rect 16972 18376 17012 18416
rect 18220 18376 18260 18416
rect 19948 18460 19988 18500
rect 20908 18460 20948 18500
rect 21100 18460 21140 18500
rect 21868 18460 21908 18500
rect 25324 18460 25364 18500
rect 26284 18460 26324 18500
rect 28204 18460 28244 18500
rect 30988 18460 31028 18500
rect 19852 18376 19892 18416
rect 20140 18376 20180 18416
rect 22732 18376 22772 18416
rect 25036 18376 25076 18416
rect 17260 18292 17300 18332
rect 19372 18292 19412 18332
rect 26092 18292 26132 18332
rect 3340 17956 3380 17996
rect 3724 17956 3764 17996
rect 4684 17956 4724 17996
rect 5068 17956 5108 17996
rect 6796 17956 6836 17996
rect 9004 17956 9044 17996
rect 11500 17956 11540 17996
rect 1324 17872 1364 17912
rect 3916 17872 3956 17912
rect 8812 17872 8852 17912
rect 2572 17788 2612 17828
rect 4300 17788 4340 17828
rect 5164 17788 5204 17828
rect 6796 17788 6836 17828
rect 18660 18124 19028 18164
rect 18220 17956 18260 17996
rect 19756 17956 19796 17996
rect 11212 17788 11252 17828
rect 13036 17788 13076 17828
rect 13708 17788 13748 17828
rect 13900 17788 13940 17828
rect 1708 17704 1748 17744
rect 2284 17704 2324 17744
rect 3532 17704 3572 17744
rect 4780 17704 4820 17744
rect 5260 17704 5300 17744
rect 5740 17704 5780 17744
rect 6028 17704 6068 17744
rect 6508 17704 6548 17744
rect 7660 17704 7700 17744
rect 8428 17704 8468 17744
rect 10060 17704 10100 17744
rect 10348 17704 10388 17744
rect 11308 17704 11348 17744
rect 13420 17704 13460 17744
rect 15436 17704 15476 17744
rect 15628 17704 15668 17744
rect 16204 17704 16244 17744
rect 16492 17704 16532 17744
rect 16684 17704 16724 17744
rect 17548 17704 17588 17744
rect 18220 17704 18231 17744
rect 18231 17704 18260 17744
rect 19852 17704 19892 17744
rect 1612 17620 1652 17660
rect 2572 17620 2612 17660
rect 3340 17620 3369 17660
rect 3369 17620 3380 17660
rect 4012 17620 4052 17660
rect 4876 17620 4916 17660
rect 5068 17620 5108 17660
rect 6700 17620 6740 17660
rect 7276 17620 7316 17660
rect 8716 17620 8756 17660
rect 9484 17620 9524 17660
rect 2476 17536 2516 17576
rect 2956 17536 2996 17576
rect 3628 17536 3668 17576
rect 1036 17452 1076 17492
rect 1324 17452 1364 17492
rect 10636 17620 10676 17660
rect 11020 17620 11060 17660
rect 26188 18208 26228 18248
rect 26434 18124 26802 18164
rect 22636 17956 22676 17996
rect 26860 17956 26900 17996
rect 27532 17956 27572 17996
rect 25324 17872 25364 17912
rect 27148 17788 27188 17828
rect 29836 17872 29876 17912
rect 30988 17872 31028 17912
rect 28396 17788 28436 17828
rect 22348 17704 22388 17744
rect 22924 17704 22939 17744
rect 22939 17704 22964 17744
rect 24460 17704 24500 17744
rect 24844 17704 24884 17744
rect 25036 17704 25076 17744
rect 26092 17704 26132 17744
rect 27340 17704 27380 17744
rect 28588 17704 28619 17744
rect 28619 17704 28628 17744
rect 11404 17620 11435 17660
rect 11435 17620 11444 17660
rect 13900 17620 13940 17660
rect 17260 17620 17300 17660
rect 17836 17620 17876 17660
rect 18124 17620 18164 17660
rect 24364 17620 24404 17660
rect 24652 17620 24683 17660
rect 24683 17620 24692 17660
rect 4780 17536 4820 17576
rect 9292 17536 9332 17576
rect 10732 17536 10772 17576
rect 14476 17536 14516 17576
rect 14860 17536 14900 17576
rect 15436 17536 15476 17576
rect 18028 17536 18059 17576
rect 18059 17536 18068 17576
rect 8908 17452 8948 17492
rect 9964 17452 10004 17492
rect 12556 17452 12596 17492
rect 13516 17452 13556 17492
rect 19276 17452 19316 17492
rect 4352 17368 4720 17408
rect 28108 17620 28148 17660
rect 28300 17620 28340 17660
rect 23596 17536 23636 17576
rect 24268 17536 24308 17576
rect 24460 17536 24500 17576
rect 31276 17536 31316 17576
rect 8428 17368 8468 17408
rect 12126 17368 12494 17408
rect 19900 17368 20268 17408
rect 27674 17368 28042 17408
rect 4972 17284 5012 17324
rect 12940 17284 12980 17324
rect 13228 17284 13268 17324
rect 1612 17200 1652 17240
rect 2284 17200 2324 17240
rect 2188 17116 2228 17156
rect 1324 17032 1355 17072
rect 1355 17032 1364 17072
rect 2092 17032 2132 17072
rect 2476 17116 2516 17156
rect 5164 17200 5204 17240
rect 6220 17200 6260 17240
rect 9100 17200 9140 17240
rect 11020 17200 11060 17240
rect 11404 17200 11444 17240
rect 13708 17200 13748 17240
rect 16876 17200 16907 17240
rect 16907 17200 16916 17240
rect 4972 17116 5012 17156
rect 8236 17116 8276 17156
rect 9196 17147 9236 17156
rect 9196 17116 9227 17147
rect 9227 17116 9236 17147
rect 10636 17116 10676 17156
rect 11884 17116 11924 17156
rect 3628 17032 3668 17072
rect 13612 17116 13652 17156
rect 17932 17200 17972 17240
rect 20428 17200 20468 17240
rect 17836 17116 17876 17156
rect 18028 17116 18068 17156
rect 18220 17116 18260 17156
rect 20620 17116 20660 17156
rect 24556 17200 24596 17240
rect 23980 17116 24020 17156
rect 24268 17116 24308 17156
rect 25036 17116 25076 17156
rect 30892 17116 30932 17156
rect 4492 17032 4532 17072
rect 5548 17032 5588 17072
rect 8908 17032 8939 17072
rect 8939 17032 8948 17072
rect 1612 16948 1652 16988
rect 652 16780 683 16820
rect 683 16780 692 16820
rect 2860 16948 2900 16988
rect 3724 16948 3764 16988
rect 4780 16948 4820 16988
rect 5068 16948 5108 16988
rect 6700 16948 6740 16988
rect 1996 16864 2036 16904
rect 2284 16864 2324 16904
rect 3916 16864 3947 16904
rect 3947 16864 3956 16904
rect 2380 16780 2420 16820
rect 1228 16696 1268 16736
rect 3112 16612 3480 16652
rect 9484 17032 9500 17072
rect 9500 17032 9524 17072
rect 10828 17032 10868 17072
rect 11020 17032 11060 17072
rect 11692 17032 11732 17072
rect 13420 17032 13460 17072
rect 13804 17032 13844 17072
rect 14764 17032 14804 17072
rect 8236 16948 8276 16988
rect 9004 16948 9044 16988
rect 9292 16948 9332 16988
rect 10636 16948 10667 16988
rect 10667 16948 10676 16988
rect 11212 16948 11252 16988
rect 15628 17032 15668 17072
rect 19276 17032 19316 17072
rect 19756 17032 19796 17072
rect 21388 17032 21428 17072
rect 21580 17032 21620 17072
rect 22540 17032 22580 17072
rect 12460 16948 12500 16988
rect 14572 16948 14612 16988
rect 16108 16948 16148 16988
rect 16876 16948 16916 16988
rect 17740 16948 17780 16988
rect 8908 16864 8948 16904
rect 14284 16864 14324 16904
rect 14764 16864 14804 16904
rect 16396 16864 16436 16904
rect 16684 16864 16724 16904
rect 17356 16864 17396 16904
rect 17932 16864 17972 16904
rect 12652 16780 12692 16820
rect 13324 16780 13364 16820
rect 13804 16780 13844 16820
rect 15244 16780 15284 16820
rect 17548 16780 17588 16820
rect 18028 16780 18068 16820
rect 8812 16696 8852 16736
rect 12556 16696 12596 16736
rect 15148 16696 15188 16736
rect 19564 16948 19604 16988
rect 20524 16948 20564 16988
rect 19276 16864 19316 16904
rect 19756 16864 19796 16904
rect 24844 17032 24884 17072
rect 27148 17032 27188 17072
rect 23020 16948 23060 16988
rect 24652 16948 24692 16988
rect 28396 16948 28436 16988
rect 23308 16864 23348 16904
rect 20140 16780 20180 16820
rect 22156 16780 22187 16820
rect 22187 16780 22196 16820
rect 24268 16780 24308 16820
rect 24460 16780 24500 16820
rect 24844 16780 24884 16820
rect 10886 16612 11254 16652
rect 12844 16612 12884 16652
rect 18660 16612 19028 16652
rect 19276 16612 19316 16652
rect 19948 16612 19988 16652
rect 21868 16612 21908 16652
rect 8236 16528 8276 16568
rect 9484 16528 9524 16568
rect 9772 16528 9812 16568
rect 24844 16528 24884 16568
rect 2284 16444 2324 16484
rect 6700 16444 6731 16484
rect 6731 16444 6740 16484
rect 7372 16444 7403 16484
rect 7403 16444 7412 16484
rect 9004 16444 9044 16484
rect 10444 16444 10484 16484
rect 11788 16444 11828 16484
rect 14188 16444 14228 16484
rect 14380 16444 14420 16484
rect 16588 16444 16628 16484
rect 17740 16444 17780 16484
rect 18028 16444 18068 16484
rect 18796 16444 18836 16484
rect 27052 16780 27092 16820
rect 26434 16612 26802 16652
rect 30412 16864 30452 16904
rect 30604 16864 30644 16904
rect 5068 16360 5108 16400
rect 7276 16360 7316 16400
rect 9196 16360 9236 16400
rect 9964 16360 10004 16400
rect 12844 16360 12884 16400
rect 19756 16444 19796 16484
rect 21580 16444 21620 16484
rect 23500 16444 23540 16484
rect 1708 16276 1748 16316
rect 2764 16276 2804 16316
rect 6892 16276 6932 16316
rect 9004 16276 9044 16316
rect 10732 16276 10772 16316
rect 12268 16276 12308 16316
rect 18508 16276 18548 16316
rect 19276 16276 19315 16316
rect 19315 16276 19316 16316
rect 27148 16444 27188 16484
rect 20140 16360 20180 16400
rect 28396 16360 28436 16400
rect 19660 16276 19700 16316
rect 21484 16276 21524 16316
rect 21868 16276 21908 16316
rect 23596 16276 23627 16316
rect 23627 16276 23636 16316
rect 24268 16276 24308 16316
rect 26092 16276 26132 16316
rect 26860 16276 26900 16316
rect 27052 16276 27092 16316
rect 30604 16276 30644 16316
rect 31276 16276 31307 16316
rect 31307 16276 31316 16316
rect 1036 16192 1076 16232
rect 2188 16192 2228 16232
rect 2668 16192 2708 16232
rect 3628 16192 3668 16232
rect 4012 16192 4043 16232
rect 4043 16192 4052 16232
rect 4876 16192 4916 16232
rect 5452 16192 5492 16232
rect 6796 16192 6836 16232
rect 7180 16192 7220 16232
rect 7948 16192 7964 16232
rect 7964 16192 7988 16232
rect 8812 16192 8852 16232
rect 9676 16192 9707 16232
rect 9707 16192 9716 16232
rect 9964 16192 10004 16232
rect 11212 16192 11252 16232
rect 12460 16192 12500 16232
rect 13324 16192 13364 16232
rect 13804 16192 13844 16232
rect 14956 16192 14996 16232
rect 15820 16192 15860 16232
rect 16108 16192 16137 16232
rect 16137 16192 16148 16232
rect 16492 16192 16532 16232
rect 16876 16192 16916 16232
rect 17548 16192 17588 16232
rect 18124 16192 18164 16232
rect 20908 16192 20948 16232
rect 21100 16192 21140 16232
rect 22444 16192 22484 16232
rect 1228 16108 1268 16148
rect 1804 16108 1844 16148
rect 2380 16108 2420 16148
rect 4300 16108 4340 16148
rect 5836 16108 5876 16148
rect 2092 16024 2132 16064
rect 2476 16024 2516 16064
rect 4684 16024 4724 16064
rect 5740 16024 5780 16064
rect 6508 16108 6548 16148
rect 6700 16108 6740 16148
rect 7276 16108 7316 16148
rect 7564 16108 7604 16148
rect 8524 16024 8563 16064
rect 8563 16024 8564 16064
rect 8812 16024 8852 16064
rect 9772 16108 9812 16148
rect 10636 16108 10676 16148
rect 11692 16108 11732 16148
rect 12556 16108 12596 16148
rect 14380 16108 14420 16148
rect 14572 16108 14612 16148
rect 21196 16108 21236 16148
rect 21580 16108 21620 16148
rect 9484 16024 9524 16064
rect 10060 16024 10100 16064
rect 11404 16024 11444 16064
rect 11980 16024 12020 16064
rect 13324 16024 13364 16064
rect 13516 16024 13555 16064
rect 13555 16024 13556 16064
rect 14092 16024 14132 16064
rect 14476 16024 14516 16064
rect 12844 15940 12884 15980
rect 4352 15856 4720 15896
rect 9964 15856 10004 15896
rect 11404 15856 11444 15896
rect 12126 15856 12494 15896
rect 23116 16192 23156 16232
rect 23500 16192 23540 16232
rect 23692 16192 23732 16232
rect 24172 16192 24212 16232
rect 24556 16192 24596 16232
rect 26380 16192 26420 16232
rect 27340 16192 27380 16232
rect 30892 16192 30923 16232
rect 30923 16192 30932 16232
rect 23212 16108 23252 16148
rect 16108 16024 16148 16064
rect 16780 16024 16820 16064
rect 20428 16024 20468 16064
rect 21388 16024 21428 16064
rect 3724 15772 3764 15812
rect 23308 15940 23348 15980
rect 3820 15688 3860 15728
rect 1420 15604 1460 15644
rect 26476 16024 26516 16064
rect 14188 15856 14228 15896
rect 18796 15856 18836 15896
rect 19276 15856 19316 15896
rect 19900 15856 20268 15896
rect 26284 15856 26324 15896
rect 27340 15856 27380 15896
rect 27674 15856 28042 15896
rect 13132 15772 13172 15812
rect 19660 15772 19700 15812
rect 5836 15688 5876 15728
rect 7180 15688 7220 15728
rect 9292 15688 9323 15728
rect 9323 15688 9332 15728
rect 11116 15688 11156 15728
rect 11692 15688 11723 15728
rect 11723 15688 11732 15728
rect 13228 15688 13268 15728
rect 14764 15688 14804 15728
rect 16492 15688 16532 15728
rect 16876 15688 16916 15728
rect 17356 15688 17396 15728
rect 1804 15520 1844 15560
rect 2380 15520 2420 15560
rect 1228 15352 1268 15392
rect 3532 15520 3544 15560
rect 3544 15520 3572 15560
rect 4492 15520 4532 15560
rect 5452 15520 5492 15560
rect 5740 15520 5749 15560
rect 5749 15520 5780 15560
rect 6220 15520 6260 15560
rect 6796 15520 6836 15560
rect 4108 15436 4148 15476
rect 6028 15436 6068 15476
rect 7276 15520 7316 15560
rect 2764 15268 2795 15308
rect 2795 15268 2804 15308
rect 9100 15604 9140 15644
rect 9484 15604 9524 15644
rect 9964 15604 10004 15644
rect 11500 15604 11540 15644
rect 7948 15436 7988 15476
rect 6796 15352 6836 15392
rect 7180 15352 7220 15392
rect 7564 15352 7604 15392
rect 8044 15352 8084 15392
rect 8908 15436 8948 15476
rect 9196 15436 9236 15476
rect 9388 15352 9428 15392
rect 7084 15268 7124 15308
rect 7372 15268 7412 15308
rect 8236 15268 8276 15308
rect 5452 15184 5492 15224
rect 5740 15184 5780 15224
rect 3112 15100 3480 15140
rect 5356 15100 5396 15140
rect 9580 15100 9620 15140
rect 1708 15016 1748 15056
rect 6124 15016 6164 15056
rect 7756 15016 7796 15056
rect 4108 14932 4148 14972
rect 4300 14932 4340 14972
rect 5740 14932 5780 14972
rect 10540 15520 10580 15560
rect 10732 15520 10772 15560
rect 10156 15436 10196 15476
rect 11500 15436 11531 15476
rect 11531 15436 11540 15476
rect 9964 15352 10004 15392
rect 11212 15352 11252 15392
rect 13804 15604 13844 15644
rect 14188 15604 14228 15644
rect 16588 15635 16628 15644
rect 16588 15604 16619 15635
rect 16619 15604 16628 15635
rect 17164 15604 17193 15644
rect 17193 15604 17204 15644
rect 18028 15688 18068 15728
rect 20908 15688 20948 15728
rect 23692 15688 23732 15728
rect 28684 15772 28724 15812
rect 18220 15604 18260 15644
rect 19852 15604 19892 15644
rect 25228 15688 25268 15728
rect 25996 15688 26036 15728
rect 26380 15604 26420 15644
rect 11788 15520 11828 15560
rect 12844 15520 12884 15560
rect 13516 15520 13527 15560
rect 13527 15520 13556 15560
rect 14092 15520 14132 15560
rect 14572 15520 14612 15560
rect 12460 15436 12500 15476
rect 15916 15520 15956 15560
rect 17356 15520 17396 15560
rect 13036 15436 13076 15476
rect 13228 15436 13268 15476
rect 13612 15436 13652 15476
rect 14380 15436 14420 15476
rect 15244 15436 15284 15476
rect 16396 15436 16436 15476
rect 14668 15352 14708 15392
rect 15820 15352 15860 15392
rect 16588 15352 16628 15392
rect 17740 15520 17780 15560
rect 18028 15520 18059 15560
rect 18059 15520 18068 15560
rect 19084 15520 19124 15560
rect 20620 15520 20660 15560
rect 21484 15520 21524 15560
rect 24172 15520 24212 15560
rect 25036 15520 25076 15560
rect 25228 15520 25268 15560
rect 18316 15436 18356 15476
rect 25900 15520 25940 15560
rect 26476 15520 26501 15560
rect 26501 15520 26516 15560
rect 26860 15520 26900 15560
rect 27052 15520 27092 15560
rect 27436 15520 27447 15560
rect 27447 15520 27476 15560
rect 19660 15436 19700 15476
rect 23692 15436 23732 15476
rect 26956 15436 26996 15476
rect 18700 15352 18740 15392
rect 20428 15352 20468 15392
rect 14956 15268 14996 15308
rect 16684 15268 16724 15308
rect 17644 15268 17675 15308
rect 17675 15268 17684 15308
rect 20812 15268 20852 15308
rect 21292 15268 21332 15308
rect 19564 15184 19604 15224
rect 21580 15184 21620 15224
rect 10886 15100 11254 15140
rect 15820 15100 15860 15140
rect 16300 15100 16340 15140
rect 18660 15100 19028 15140
rect 22156 15100 22196 15140
rect 11788 15016 11828 15056
rect 17356 15016 17396 15056
rect 7084 14932 7124 14972
rect 7948 14932 7988 14972
rect 1228 14848 1268 14888
rect 1708 14848 1748 14888
rect 2956 14764 2996 14804
rect 8236 14848 8276 14888
rect 9100 14848 9140 14888
rect 10156 14932 10196 14972
rect 4108 14764 4148 14804
rect 1228 14680 1268 14720
rect 1804 14680 1844 14720
rect 2380 14680 2420 14720
rect 2860 14680 2900 14720
rect 3532 14680 3572 14720
rect 1036 14596 1067 14636
rect 1067 14596 1076 14636
rect 1324 14596 1364 14636
rect 3436 14596 3476 14636
rect 3724 14596 3764 14636
rect 1900 14512 1940 14552
rect 1228 14428 1268 14468
rect 4108 14428 4148 14468
rect 940 14344 980 14384
rect 2188 14344 2228 14384
rect 2764 14344 2804 14384
rect 1804 14260 1844 14300
rect 5740 14680 5764 14720
rect 5764 14680 5780 14720
rect 6796 14680 6836 14720
rect 7084 14680 7124 14720
rect 7756 14764 7796 14804
rect 8140 14764 8180 14804
rect 8524 14764 8564 14804
rect 10348 14848 10388 14888
rect 10252 14764 10292 14804
rect 21484 15016 21524 15056
rect 11596 14932 11636 14972
rect 11884 14932 11924 14972
rect 13228 14932 13268 14972
rect 17836 14932 17876 14972
rect 18700 14932 18740 14972
rect 12940 14764 12980 14804
rect 14764 14764 14787 14804
rect 14787 14764 14804 14804
rect 16492 14764 16532 14804
rect 17164 14764 17204 14804
rect 17452 14764 17492 14804
rect 17644 14764 17684 14804
rect 18604 14764 18644 14804
rect 26284 15352 26324 15392
rect 30892 15520 30923 15560
rect 30923 15520 30932 15560
rect 25324 15268 25364 15308
rect 26434 15100 26802 15140
rect 25036 15016 25076 15056
rect 26188 14932 26228 14972
rect 19756 14848 19796 14888
rect 21196 14848 21236 14888
rect 20908 14764 20948 14804
rect 21100 14764 21140 14804
rect 21484 14764 21524 14804
rect 8332 14680 8372 14720
rect 9196 14680 9227 14720
rect 9227 14680 9236 14720
rect 9484 14680 9524 14720
rect 9964 14680 10004 14720
rect 10444 14680 10463 14720
rect 10463 14680 10484 14720
rect 10732 14680 10772 14720
rect 11212 14680 11224 14720
rect 11224 14680 11252 14720
rect 11404 14680 11444 14720
rect 12556 14680 12596 14720
rect 13132 14680 13163 14720
rect 13163 14680 13172 14720
rect 13708 14680 13724 14720
rect 13724 14680 13748 14720
rect 13996 14680 14036 14720
rect 14668 14680 14708 14720
rect 15340 14680 15380 14720
rect 15820 14680 15860 14720
rect 16396 14680 16436 14720
rect 4492 14596 4532 14636
rect 5452 14596 5492 14636
rect 6124 14596 6164 14636
rect 6412 14596 6452 14636
rect 6892 14596 6932 14636
rect 17836 14680 17852 14720
rect 17852 14680 17876 14720
rect 18700 14680 18740 14720
rect 18892 14680 18932 14720
rect 19564 14680 19604 14720
rect 21580 14680 21620 14720
rect 22444 14680 22484 14720
rect 22924 14680 22964 14720
rect 23980 14680 24020 14720
rect 24652 14764 24692 14804
rect 25228 14764 25268 14804
rect 26860 14764 26900 14804
rect 27148 14764 27188 14804
rect 30412 15436 30452 15476
rect 28876 15268 28916 15308
rect 29356 15268 29396 15308
rect 28588 14848 28628 14888
rect 31084 14848 31124 14888
rect 24748 14680 24777 14720
rect 24777 14680 24788 14720
rect 24940 14680 24980 14720
rect 25420 14680 25460 14720
rect 26668 14680 26708 14720
rect 7660 14596 7700 14636
rect 9004 14596 9044 14636
rect 14188 14596 14228 14636
rect 15916 14596 15956 14636
rect 16108 14596 16148 14636
rect 16876 14596 16916 14636
rect 17644 14596 17684 14636
rect 19084 14596 19124 14636
rect 19660 14596 19700 14636
rect 20428 14596 20468 14636
rect 27244 14680 27284 14720
rect 27532 14680 27572 14720
rect 27820 14680 27860 14720
rect 28492 14680 28532 14720
rect 28972 14680 29012 14720
rect 30508 14680 30548 14720
rect 24268 14596 24308 14636
rect 26764 14596 26804 14636
rect 29356 14596 29396 14636
rect 5836 14512 5867 14552
rect 5867 14512 5876 14552
rect 13516 14512 13547 14552
rect 13547 14512 13556 14552
rect 13804 14512 13844 14552
rect 16012 14512 16051 14552
rect 16051 14512 16052 14552
rect 16588 14512 16628 14552
rect 17740 14512 17771 14552
rect 17771 14512 17780 14552
rect 17932 14512 17972 14552
rect 18604 14512 18644 14552
rect 23308 14512 23348 14552
rect 5932 14428 5972 14468
rect 11692 14428 11732 14468
rect 24364 14428 24404 14468
rect 4352 14344 4720 14384
rect 5068 14344 5108 14384
rect 6892 14344 6932 14384
rect 7564 14344 7604 14384
rect 12126 14344 12494 14384
rect 19660 14344 19700 14384
rect 19900 14344 20268 14384
rect 27674 14344 28042 14384
rect 7468 14260 7508 14300
rect 10348 14260 10388 14300
rect 10540 14260 10580 14300
rect 14092 14260 14132 14300
rect 14572 14260 14612 14300
rect 15244 14260 15284 14300
rect 18220 14260 18260 14300
rect 1612 14176 1652 14216
rect 2380 14176 2420 14216
rect 5452 14176 5492 14216
rect 5644 14176 5675 14216
rect 5675 14176 5684 14216
rect 7276 14176 7316 14216
rect 10444 14176 10484 14216
rect 10636 14176 10676 14216
rect 2764 14092 2804 14132
rect 5836 14092 5876 14132
rect 652 13504 692 13544
rect 27148 14260 27188 14300
rect 14764 14176 14795 14216
rect 14795 14176 14804 14216
rect 15340 14176 15380 14216
rect 16204 14176 16244 14216
rect 18892 14176 18932 14216
rect 20428 14176 20468 14216
rect 21292 14176 21332 14216
rect 24940 14176 24980 14216
rect 25228 14176 25268 14216
rect 26092 14176 26132 14216
rect 27052 14176 27092 14216
rect 27244 14176 27284 14216
rect 9004 14092 9044 14132
rect 9388 14092 9428 14132
rect 10540 14092 10580 14132
rect 11212 14092 11252 14132
rect 15148 14092 15188 14132
rect 1324 14008 1364 14048
rect 1708 14008 1739 14048
rect 1739 14008 1748 14048
rect 2188 14008 2228 14048
rect 3724 14008 3764 14048
rect 5932 14008 5972 14048
rect 7756 14008 7796 14048
rect 10348 14008 10388 14048
rect 10732 14008 10772 14048
rect 11308 14008 11348 14048
rect 172 13252 212 13292
rect 1228 13924 1268 13964
rect 1612 13756 1652 13796
rect 2764 13756 2804 13796
rect 3532 13924 3572 13964
rect 3112 13588 3480 13628
rect 3724 13420 3764 13460
rect 17644 14092 17684 14132
rect 21580 14092 21620 14132
rect 22252 14092 22292 14132
rect 23692 14092 23732 14132
rect 24172 14092 24212 14132
rect 24460 14092 24500 14132
rect 12460 14008 12500 14048
rect 14188 14008 14228 14048
rect 14668 14008 14697 14048
rect 14697 14008 14708 14048
rect 5452 13924 5492 13964
rect 6028 13924 6051 13964
rect 6051 13924 6068 13964
rect 6316 13924 6356 13964
rect 6892 13924 6932 13964
rect 8332 13924 8372 13964
rect 8908 13924 8948 13964
rect 10156 13924 10179 13964
rect 10179 13924 10196 13964
rect 12652 13924 12692 13964
rect 12940 13924 12980 13964
rect 5164 13756 5204 13796
rect 6412 13840 6452 13880
rect 7852 13840 7892 13880
rect 8140 13840 8180 13880
rect 9964 13840 10004 13880
rect 11404 13840 11444 13880
rect 15244 14008 15284 14048
rect 15052 13924 15092 13964
rect 15340 13924 15380 13964
rect 17740 14008 17780 14048
rect 18796 14008 18836 14048
rect 20236 14008 20249 14048
rect 20249 14008 20276 14048
rect 20812 14008 20852 14048
rect 21484 14008 21524 14048
rect 22444 14008 22484 14048
rect 23308 14008 23317 14048
rect 23317 14008 23348 14048
rect 24652 14008 24692 14048
rect 24940 14008 24980 14048
rect 16780 13924 16820 13964
rect 17548 13924 17588 13964
rect 20620 13924 20660 13964
rect 16300 13840 16340 13880
rect 17932 13840 17972 13880
rect 11596 13756 11636 13796
rect 13804 13756 13844 13796
rect 14572 13756 14612 13796
rect 14764 13756 14804 13796
rect 17164 13756 17204 13796
rect 21484 13756 21524 13796
rect 9004 13672 9044 13712
rect 12748 13672 12788 13712
rect 16876 13672 16916 13712
rect 6124 13588 6164 13628
rect 10886 13588 11254 13628
rect 18660 13588 19028 13628
rect 7948 13504 7988 13544
rect 9196 13504 9236 13544
rect 9676 13504 9716 13544
rect 12460 13504 12500 13544
rect 15724 13504 15764 13544
rect 17260 13504 17300 13544
rect 5740 13420 5780 13460
rect 5548 13336 5588 13376
rect 6604 13420 6644 13460
rect 7468 13420 7508 13460
rect 6124 13336 6164 13376
rect 6700 13336 6740 13376
rect 7852 13336 7892 13376
rect 8908 13336 8948 13376
rect 10636 13420 10676 13460
rect 11308 13420 11348 13460
rect 4780 13252 4811 13292
rect 4811 13252 4820 13292
rect 5644 13252 5684 13292
rect 6412 13252 6452 13292
rect 6892 13252 6932 13292
rect 7564 13252 7604 13292
rect 1420 13168 1460 13208
rect 7948 13252 7988 13292
rect 8524 13252 8564 13292
rect 3340 13168 3380 13208
rect 3724 13168 3764 13208
rect 4876 13168 4916 13208
rect 6124 13168 6164 13208
rect 6700 13168 6721 13208
rect 6721 13168 6740 13208
rect 7084 13168 7124 13208
rect 7468 13168 7479 13208
rect 7479 13168 7508 13208
rect 10348 13252 10371 13292
rect 10371 13252 10388 13292
rect 10636 13252 10676 13292
rect 14380 13420 14420 13460
rect 15532 13420 15572 13460
rect 16300 13420 16340 13460
rect 17452 13420 17492 13460
rect 13324 13336 13364 13376
rect 13804 13336 13844 13376
rect 14764 13336 14804 13376
rect 11404 13252 11444 13292
rect 12748 13252 12788 13292
rect 12940 13252 12980 13292
rect 15244 13336 15284 13376
rect 17740 13336 17780 13376
rect 15628 13252 15668 13292
rect 16972 13252 17012 13292
rect 17164 13252 17204 13292
rect 17356 13252 17396 13292
rect 18220 13252 18260 13292
rect 22636 13504 22676 13544
rect 20140 13420 20180 13460
rect 23980 13924 24020 13964
rect 24268 13924 24308 13964
rect 25516 14008 25556 14048
rect 27340 14092 27380 14132
rect 25804 14008 25844 14048
rect 26188 14008 26228 14048
rect 27052 14008 27092 14048
rect 27628 14008 27632 14048
rect 27632 14008 27668 14048
rect 28588 14008 28628 14048
rect 30604 14008 30644 14048
rect 30892 14008 30923 14048
rect 30923 14008 30932 14048
rect 26860 13924 26890 13964
rect 26890 13924 26900 13964
rect 27148 13924 27188 13964
rect 28972 13924 29012 13964
rect 31084 13924 31124 13964
rect 23500 13840 23540 13880
rect 25324 13840 25364 13880
rect 26284 13840 26324 13880
rect 26668 13840 26708 13880
rect 28780 13840 28820 13880
rect 27340 13756 27380 13796
rect 27628 13756 27668 13796
rect 30508 13756 30548 13796
rect 26434 13588 26802 13628
rect 24268 13420 24308 13460
rect 25900 13420 25940 13460
rect 26956 13420 26996 13460
rect 19660 13336 19700 13376
rect 25228 13336 25268 13376
rect 26764 13336 26804 13376
rect 29932 13336 29972 13376
rect 8332 13168 8372 13208
rect 9100 13168 9140 13208
rect 11020 13168 11043 13208
rect 11043 13168 11060 13208
rect 13132 13168 13172 13208
rect 14380 13168 14420 13208
rect 14764 13168 14771 13208
rect 14771 13168 14804 13208
rect 15532 13168 15572 13208
rect 15724 13168 15749 13208
rect 15749 13168 15764 13208
rect 16012 13168 16052 13208
rect 16588 13168 16628 13208
rect 17836 13168 17867 13208
rect 17867 13168 17876 13208
rect 18316 13168 18345 13208
rect 18345 13168 18356 13208
rect 20236 13252 20276 13292
rect 21292 13252 21332 13292
rect 21484 13252 21524 13292
rect 23308 13252 23348 13292
rect 24652 13252 24692 13292
rect 5164 13084 5204 13124
rect 5548 13084 5588 13124
rect 6028 13084 6068 13124
rect 7948 13084 7988 13124
rect 6508 13000 6548 13040
rect 7564 13000 7604 13040
rect 8620 13000 8660 13040
rect 8908 13000 8948 13040
rect 10156 13084 10196 13124
rect 10444 13084 10484 13124
rect 10924 13084 10964 13124
rect 12556 13084 12596 13124
rect 12748 13084 12788 13124
rect 13420 13084 13460 13124
rect 14092 13084 14132 13124
rect 13228 13000 13268 13040
rect 14764 13000 14804 13040
rect 3628 12916 3668 12956
rect 7372 12916 7412 12956
rect 8428 12916 8468 12956
rect 10156 12916 10196 12956
rect 11404 12916 11444 12956
rect 17452 13084 17492 13124
rect 17740 13084 17780 13124
rect 18892 13084 18932 13124
rect 15244 13000 15284 13040
rect 19756 13168 19796 13208
rect 20812 13168 20852 13208
rect 18124 13000 18155 13040
rect 18155 13000 18164 13040
rect 18508 13000 18548 13040
rect 26860 13252 26900 13292
rect 28108 13252 28148 13292
rect 28396 13252 28436 13292
rect 30700 13252 30740 13292
rect 21388 13168 21428 13208
rect 22252 13168 22292 13208
rect 22540 13168 22580 13208
rect 24460 13168 24461 13208
rect 24461 13168 24500 13208
rect 25228 13168 25268 13208
rect 25900 13168 25940 13208
rect 27052 13168 27057 13208
rect 27057 13168 27092 13208
rect 27340 13168 27380 13208
rect 28780 13168 28820 13208
rect 28972 13168 29012 13208
rect 30604 13168 30644 13208
rect 23692 13084 23732 13124
rect 24172 13084 24212 13124
rect 25804 13084 25844 13124
rect 20812 13000 20852 13040
rect 21484 13000 21524 13040
rect 23884 13000 23924 13040
rect 24268 13000 24308 13040
rect 15436 12916 15476 12956
rect 23788 12916 23828 12956
rect 24556 12916 24596 12956
rect 25228 12916 25268 12956
rect 4352 12832 4720 12872
rect 12126 12832 12494 12872
rect 15340 12832 15380 12872
rect 16972 12832 17012 12872
rect 17164 12832 17204 12872
rect 19900 12832 20268 12872
rect 23116 12832 23156 12872
rect 23692 12832 23732 12872
rect 27674 12832 28042 12872
rect 3724 12748 3764 12788
rect 5356 12748 5396 12788
rect 940 12664 980 12704
rect 3340 12664 3380 12704
rect 4204 12664 4244 12704
rect 7948 12748 7988 12788
rect 9388 12748 9428 12788
rect 13516 12748 13556 12788
rect 14380 12748 14420 12788
rect 16204 12748 16244 12788
rect 18124 12748 18164 12788
rect 6028 12664 6068 12704
rect 6700 12664 6740 12704
rect 8524 12664 8564 12704
rect 8908 12664 8948 12704
rect 4492 12580 4532 12620
rect 4972 12580 5012 12620
rect 7372 12580 7412 12620
rect 1324 12496 1364 12536
rect 2284 12496 2324 12536
rect 2764 12496 2804 12536
rect 2668 12412 2708 12452
rect 1900 12328 1940 12368
rect 8140 12580 8180 12620
rect 11308 12664 11348 12704
rect 13036 12664 13067 12704
rect 13067 12664 13076 12704
rect 14572 12664 14603 12704
rect 14603 12664 14612 12704
rect 17836 12664 17876 12704
rect 18412 12664 18452 12704
rect 9484 12580 9524 12620
rect 5836 12496 5876 12536
rect 5644 12412 5684 12452
rect 1324 12244 1364 12284
rect 1228 12160 1268 12200
rect 2668 12160 2708 12200
rect 3112 12076 3480 12116
rect 1804 11908 1844 11948
rect 2764 11908 2804 11948
rect 4492 11908 4523 11948
rect 4523 11908 4532 11948
rect 1900 11740 1940 11780
rect 2860 11740 2900 11780
rect 6316 12412 6356 12452
rect 7084 12412 7107 12452
rect 7107 12412 7124 12452
rect 7276 12328 7316 12368
rect 7468 12244 7508 12284
rect 8332 12496 8372 12536
rect 8524 12496 8547 12536
rect 8547 12496 8564 12536
rect 9100 12496 9140 12536
rect 12556 12580 12596 12620
rect 13996 12580 14036 12620
rect 14476 12580 14516 12620
rect 16876 12580 16916 12620
rect 10636 12496 10657 12536
rect 10657 12496 10676 12536
rect 11116 12496 11156 12536
rect 12748 12496 12755 12536
rect 12755 12496 12788 12536
rect 18604 12580 18644 12620
rect 26380 12748 26420 12788
rect 27244 12748 27284 12788
rect 19180 12664 19220 12704
rect 22540 12664 22580 12704
rect 23884 12664 23924 12704
rect 24460 12664 24500 12704
rect 25708 12664 25748 12704
rect 26284 12664 26324 12704
rect 26956 12664 26987 12704
rect 26987 12664 26996 12704
rect 27532 12664 27572 12704
rect 28588 12664 28628 12704
rect 21196 12580 21236 12620
rect 25420 12580 25460 12620
rect 26860 12580 26900 12620
rect 27052 12580 27092 12620
rect 27244 12580 27284 12620
rect 28108 12580 28148 12620
rect 28396 12580 28436 12620
rect 13324 12496 13364 12536
rect 13612 12496 13652 12536
rect 15340 12496 15380 12536
rect 16492 12496 16532 12536
rect 17164 12496 17204 12536
rect 20716 12496 20756 12536
rect 21484 12496 21524 12536
rect 23212 12496 23252 12536
rect 23692 12496 23732 12536
rect 24460 12496 24500 12536
rect 24652 12496 24692 12536
rect 8620 12412 8660 12452
rect 9676 12412 9716 12452
rect 10828 12412 10868 12452
rect 11788 12412 11828 12452
rect 12940 12412 12980 12452
rect 7948 12328 7988 12368
rect 8908 12328 8948 12368
rect 10732 12328 10772 12368
rect 8140 12244 8180 12284
rect 8332 12244 8372 12284
rect 8716 12244 8756 12284
rect 13036 12328 13076 12368
rect 13612 12244 13652 12284
rect 16588 12244 16628 12284
rect 6988 12160 7028 12200
rect 10348 12160 10388 12200
rect 13516 12160 13556 12200
rect 15724 12160 15764 12200
rect 5164 12076 5204 12116
rect 10886 12076 11254 12116
rect 13132 12076 13172 12116
rect 16492 12076 16532 12116
rect 7372 11992 7412 12032
rect 7564 11992 7604 12032
rect 8236 11992 8276 12032
rect 5740 11824 5780 11864
rect 4972 11740 5012 11780
rect 5836 11740 5876 11780
rect 1420 11656 1460 11696
rect 4108 11656 4148 11696
rect 4876 11656 4916 11696
rect 5260 11656 5300 11696
rect 18508 12244 18548 12284
rect 22060 12412 22100 12452
rect 20812 12328 20852 12368
rect 20140 12244 20180 12284
rect 22636 12244 22676 12284
rect 10636 11992 10676 12032
rect 12556 11992 12596 12032
rect 14476 11992 14516 12032
rect 16108 11992 16148 12032
rect 6988 11824 7028 11864
rect 6700 11740 6740 11780
rect 10444 11908 10484 11948
rect 7372 11824 7412 11864
rect 7660 11740 7700 11780
rect 7084 11656 7124 11696
rect 7276 11656 7316 11696
rect 7564 11656 7604 11696
rect 1132 11572 1172 11612
rect 2860 11572 2900 11612
rect 8225 11824 8265 11864
rect 10348 11824 10388 11864
rect 10540 11824 10580 11864
rect 10924 11824 10964 11864
rect 11500 11908 11540 11948
rect 12652 11908 12692 11948
rect 13036 11908 13067 11948
rect 13067 11908 13076 11948
rect 11596 11824 11636 11864
rect 13132 11824 13172 11864
rect 9004 11740 9044 11780
rect 9676 11740 9716 11780
rect 9964 11740 10004 11780
rect 11500 11740 11540 11780
rect 12748 11740 12788 11780
rect 13804 11908 13844 11948
rect 16204 11908 16244 11948
rect 16492 11908 16532 11948
rect 13996 11824 14036 11864
rect 14764 11824 14804 11864
rect 15244 11824 15284 11864
rect 12940 11740 12980 11780
rect 13900 11740 13940 11780
rect 14572 11740 14612 11780
rect 16108 11824 16148 11864
rect 16396 11824 16436 11864
rect 15340 11740 15380 11780
rect 15724 11740 15764 11780
rect 18660 12076 19028 12116
rect 18604 11908 18644 11948
rect 16588 11824 16628 11864
rect 21292 11824 21332 11864
rect 17740 11740 17780 11780
rect 20620 11740 20660 11780
rect 21964 11740 22004 11780
rect 22636 11740 22676 11780
rect 22828 11740 22868 11780
rect 23884 12412 23924 12452
rect 24556 12412 24596 12452
rect 25708 12412 25748 12452
rect 26476 12496 26516 12536
rect 26764 12496 26804 12536
rect 27436 12496 27476 12536
rect 26188 12412 26228 12452
rect 27820 12412 27860 12452
rect 28204 12412 28244 12452
rect 30604 12496 30635 12536
rect 30635 12496 30644 12536
rect 29932 12412 29972 12452
rect 25804 12328 25844 12368
rect 28492 12328 28532 12368
rect 23980 12244 24020 12284
rect 23500 12160 23540 12200
rect 23692 12160 23732 12200
rect 24268 12160 24308 12200
rect 30700 12160 30740 12200
rect 26434 12076 26802 12116
rect 26188 11992 26228 12032
rect 25708 11908 25748 11948
rect 26092 11908 26132 11948
rect 31276 11824 31316 11864
rect 23596 11740 23636 11780
rect 24940 11740 24980 11780
rect 25420 11740 25460 11780
rect 26188 11740 26228 11780
rect 28204 11740 28244 11780
rect 28972 11740 29012 11780
rect 8908 11656 8948 11696
rect 9196 11656 9236 11696
rect 9772 11656 9812 11696
rect 10156 11656 10196 11696
rect 10540 11656 10580 11696
rect 11020 11656 11060 11696
rect 11212 11656 11252 11696
rect 13516 11656 13545 11696
rect 13545 11656 13556 11696
rect 14092 11656 14111 11696
rect 14111 11656 14132 11696
rect 14284 11656 14324 11696
rect 14764 11656 14804 11696
rect 15436 11656 15465 11696
rect 15465 11656 15476 11696
rect 15820 11656 15860 11696
rect 6988 11572 7028 11612
rect 8524 11572 8564 11612
rect 11596 11572 11636 11612
rect 11788 11572 11828 11612
rect 13228 11572 13268 11612
rect 16588 11656 16613 11696
rect 16613 11656 16628 11696
rect 17452 11656 17492 11696
rect 18124 11656 18155 11696
rect 18155 11656 18164 11696
rect 15532 11572 15572 11612
rect 3436 11488 3476 11528
rect 3820 11488 3860 11528
rect 5260 11488 5300 11528
rect 5740 11488 5771 11528
rect 5771 11488 5780 11528
rect 16396 11572 16436 11612
rect 20428 11656 20468 11696
rect 20716 11656 20756 11696
rect 21388 11656 21428 11696
rect 21868 11656 21908 11696
rect 22540 11656 22580 11696
rect 23980 11656 24020 11696
rect 25324 11656 25364 11696
rect 26860 11656 26900 11696
rect 27532 11656 27572 11696
rect 27820 11656 27860 11696
rect 28300 11656 28340 11696
rect 28492 11656 28517 11696
rect 28517 11656 28532 11696
rect 28780 11656 28820 11696
rect 30700 11656 30731 11696
rect 30731 11656 30740 11696
rect 21580 11572 21620 11612
rect 23212 11572 23252 11612
rect 23500 11572 23540 11612
rect 24172 11572 24212 11612
rect 25516 11572 25556 11612
rect 28684 11572 28724 11612
rect 31180 11572 31220 11612
rect 8620 11488 8660 11528
rect 14476 11488 14507 11528
rect 14507 11488 14516 11528
rect 15436 11488 15467 11528
rect 15467 11488 15476 11528
rect 16012 11488 16052 11528
rect 19180 11488 19220 11528
rect 21484 11488 21524 11528
rect 23884 11488 23924 11528
rect 27340 11488 27380 11528
rect 28588 11488 28628 11528
rect 4012 11404 4052 11444
rect 6604 11404 6644 11444
rect 8236 11404 8276 11444
rect 9964 11404 10004 11444
rect 4352 11320 4720 11360
rect 5548 11320 5588 11360
rect 8332 11320 8372 11360
rect 8716 11320 8756 11360
rect 12126 11320 12494 11360
rect 12748 11320 12788 11360
rect 13036 11320 13076 11360
rect 16396 11320 16436 11360
rect 6508 11236 6548 11276
rect 16108 11236 16148 11276
rect 4204 11152 4235 11192
rect 4235 11152 4244 11192
rect 4780 11152 4811 11192
rect 4811 11152 4820 11192
rect 6988 11152 7028 11192
rect 7180 11152 7220 11192
rect 8044 11152 8084 11192
rect 8428 11152 8468 11192
rect 9100 11152 9140 11192
rect 10540 11152 10555 11192
rect 10555 11152 10580 11192
rect 11500 11152 11540 11192
rect 11788 11152 11828 11192
rect 12940 11152 12980 11192
rect 13900 11152 13940 11192
rect 15820 11152 15860 11192
rect 16684 11152 16724 11192
rect 16876 11152 16916 11192
rect 1324 11068 1364 11108
rect 1612 11068 1652 11108
rect 4300 11068 4340 11108
rect 6220 11068 6260 11108
rect 10156 11068 10196 11108
rect 11596 11068 11636 11108
rect 12172 11068 12212 11108
rect 15148 11068 15188 11108
rect 2092 10984 2132 11024
rect 2860 10984 2900 11024
rect 3436 10984 3448 11024
rect 3448 10984 3476 11024
rect 4396 10984 4420 11024
rect 4420 10984 4436 11024
rect 5260 10984 5300 11024
rect 5548 10984 5588 11024
rect 6124 10984 6164 11024
rect 7372 10984 7412 11024
rect 7660 10984 7700 11024
rect 8140 10984 8180 11024
rect 8332 10984 8357 11024
rect 8357 10984 8372 11024
rect 8908 10984 8909 11024
rect 8909 10984 8948 11024
rect 1324 10900 1364 10940
rect 2668 10900 2708 10940
rect 1132 10816 1172 10856
rect 1516 10732 1556 10772
rect 4588 10900 4628 10940
rect 4684 10816 4724 10856
rect 5740 10900 5780 10940
rect 6316 10900 6356 10940
rect 7276 10900 7316 10940
rect 7852 10900 7892 10940
rect 8236 10900 8259 10940
rect 8259 10900 8276 10940
rect 4876 10816 4916 10856
rect 4204 10732 4244 10772
rect 9964 10984 10004 11024
rect 10252 10984 10292 11024
rect 10444 10984 10475 11024
rect 10475 10984 10484 11024
rect 11020 10984 11060 11024
rect 11884 10984 11924 11024
rect 16108 11068 16148 11108
rect 17644 11068 17684 11108
rect 13804 10984 13829 11024
rect 13829 10984 13844 11024
rect 9772 10900 9812 10940
rect 10156 10900 10196 10940
rect 11500 10900 11540 10940
rect 11788 10900 11828 10940
rect 9580 10816 9620 10856
rect 10348 10816 10388 10856
rect 6604 10732 6635 10772
rect 6635 10732 6644 10772
rect 8908 10732 8948 10772
rect 11692 10732 11732 10772
rect 13612 10942 13652 10982
rect 13324 10900 13364 10940
rect 13996 10900 14036 10940
rect 14284 10900 14324 10940
rect 14956 10984 14996 11024
rect 15244 10984 15284 11024
rect 13516 10816 13556 10856
rect 19900 11320 20268 11360
rect 24556 11320 24596 11360
rect 27674 11320 28042 11360
rect 19756 11236 19796 11276
rect 23980 11152 24020 11192
rect 16300 10984 16340 11024
rect 17164 10984 17204 11024
rect 17932 10984 17972 11024
rect 19084 10984 19124 11024
rect 20620 11068 20660 11108
rect 21196 11068 21236 11108
rect 21484 11068 21524 11108
rect 22252 11068 22292 11108
rect 24172 11068 24212 11108
rect 25036 11068 25076 11108
rect 15340 10900 15380 10940
rect 16972 10900 17012 10940
rect 15436 10816 15439 10856
rect 15439 10816 15476 10856
rect 16012 10816 16052 10856
rect 16396 10816 16436 10856
rect 17644 10900 17684 10940
rect 17836 10900 17876 10940
rect 21100 10984 21140 11024
rect 21388 10984 21428 11024
rect 21964 10984 21995 11024
rect 21995 10984 22004 11024
rect 22828 10984 22868 11024
rect 23212 10984 23252 11024
rect 23500 10984 23531 11024
rect 23531 10984 23540 11024
rect 23884 10984 23924 11024
rect 24460 10984 24500 11024
rect 25996 10984 26036 11024
rect 26860 11152 26900 11192
rect 28780 11152 28820 11192
rect 26956 11068 26996 11108
rect 28588 11068 28628 11108
rect 31276 11068 31307 11108
rect 31307 11068 31316 11108
rect 27340 10984 27380 11024
rect 28108 10984 28148 11024
rect 29356 10984 29396 11024
rect 30892 10984 30923 11024
rect 30923 10984 30932 11024
rect 18892 10900 18923 10940
rect 18923 10900 18932 10940
rect 19180 10900 19220 10940
rect 20716 10900 20756 10940
rect 25420 10900 25460 10940
rect 29548 10900 29588 10940
rect 30988 10900 31028 10940
rect 13996 10732 14036 10772
rect 16108 10732 16148 10772
rect 17932 10732 17972 10772
rect 19948 10816 19988 10856
rect 6796 10648 6836 10688
rect 3112 10564 3480 10604
rect 10886 10564 11254 10604
rect 8140 10480 8180 10520
rect 8620 10480 8660 10520
rect 3724 10396 3764 10436
rect 4972 10396 5012 10436
rect 7276 10396 7316 10436
rect 9292 10396 9332 10436
rect 12748 10396 12788 10436
rect 6604 10312 6644 10352
rect 2284 10228 2324 10268
rect 4492 10228 4532 10268
rect 4684 10228 4724 10268
rect 6220 10228 6260 10268
rect 1036 10144 1076 10184
rect 1324 10144 1364 10184
rect 1996 10144 2036 10184
rect 2188 10144 2228 10184
rect 2956 10144 2996 10184
rect 3916 10144 3956 10184
rect 7180 10312 7220 10352
rect 7084 10228 7124 10268
rect 7948 10312 7988 10352
rect 8524 10312 8564 10352
rect 9004 10312 9044 10352
rect 10732 10312 10772 10352
rect 7372 10228 7412 10268
rect 7756 10228 7796 10268
rect 8236 10228 8276 10268
rect 8620 10228 8660 10268
rect 10540 10228 10580 10268
rect 11116 10312 11156 10352
rect 11788 10312 11828 10352
rect 13228 10312 13268 10352
rect 11404 10228 11444 10268
rect 11980 10228 12020 10268
rect 12364 10228 12404 10268
rect 28492 10816 28532 10856
rect 23500 10732 23540 10772
rect 24844 10732 24884 10772
rect 29068 10732 29108 10772
rect 29356 10732 29396 10772
rect 30412 10732 30452 10772
rect 13612 10564 13652 10604
rect 13900 10564 13940 10604
rect 18660 10564 19028 10604
rect 20428 10564 20468 10604
rect 21292 10564 21332 10604
rect 26434 10564 26802 10604
rect 20620 10480 20660 10520
rect 21388 10480 21428 10520
rect 25132 10480 25172 10520
rect 14956 10396 14987 10436
rect 14987 10396 14996 10436
rect 17260 10396 17300 10436
rect 14668 10312 14708 10352
rect 14092 10228 14132 10268
rect 14572 10228 14612 10268
rect 14860 10228 14900 10268
rect 16876 10312 16916 10352
rect 17548 10312 17588 10352
rect 15340 10228 15380 10268
rect 15820 10228 15860 10268
rect 16396 10228 16436 10268
rect 17452 10228 17492 10268
rect 19084 10312 19124 10352
rect 19564 10396 19604 10436
rect 23212 10396 23252 10436
rect 24460 10396 24500 10436
rect 24652 10396 24692 10436
rect 25804 10396 25844 10436
rect 29548 10396 29588 10436
rect 20716 10312 20756 10352
rect 20908 10312 20948 10352
rect 21100 10312 21140 10352
rect 23692 10312 23732 10352
rect 24076 10312 24116 10352
rect 25420 10312 25460 10352
rect 27532 10312 27572 10352
rect 21580 10228 21620 10268
rect 21964 10228 22004 10268
rect 24556 10228 24596 10268
rect 28300 10228 28340 10268
rect 30604 10228 30644 10268
rect 4972 10144 5012 10184
rect 5356 10144 5396 10184
rect 5548 10144 5588 10184
rect 6796 10144 6836 10184
rect 7852 10144 7892 10184
rect 8908 10144 8948 10184
rect 9868 10144 9908 10184
rect 10636 10144 10676 10184
rect 11788 10144 11828 10184
rect 12172 10144 12193 10184
rect 12193 10144 12212 10184
rect 13324 10144 13364 10184
rect 13900 10144 13940 10184
rect 2764 10060 2804 10100
rect 4588 10060 4628 10100
rect 6508 10060 6548 10100
rect 7564 10060 7604 10100
rect 3052 9976 3092 10016
rect 5068 9976 5108 10016
rect 5836 9976 5876 10016
rect 6604 9976 6644 10016
rect 7948 9976 7988 10016
rect 2572 9808 2612 9848
rect 9196 10060 9236 10100
rect 14956 10144 14996 10184
rect 15532 10144 15572 10184
rect 16108 10144 16148 10184
rect 16588 10144 16628 10184
rect 17644 10144 17675 10184
rect 17675 10144 17684 10184
rect 18604 10144 18644 10184
rect 19003 10144 19043 10184
rect 19948 10144 19988 10184
rect 20332 10144 20360 10184
rect 20360 10144 20372 10184
rect 21388 10144 21428 10184
rect 22636 10144 22676 10184
rect 23500 10144 23540 10184
rect 24940 10144 24980 10184
rect 25324 10144 25364 10184
rect 27436 10144 27476 10184
rect 28108 10144 28148 10184
rect 29068 10144 29108 10184
rect 30508 10144 30548 10184
rect 11980 10060 12020 10100
rect 14380 10060 14420 10100
rect 16876 10060 16916 10100
rect 17164 10060 17204 10100
rect 17836 10060 17876 10100
rect 19660 10060 19700 10100
rect 20428 10060 20468 10100
rect 30412 10060 30452 10100
rect 15820 9976 15860 10016
rect 17548 9976 17588 10016
rect 19852 9976 19883 10016
rect 19883 9976 19892 10016
rect 23788 9976 23828 10016
rect 24844 9976 24884 10016
rect 27052 9976 27092 10016
rect 27340 9976 27380 10016
rect 8044 9892 8084 9932
rect 10444 9892 10484 9932
rect 14284 9892 14324 9932
rect 17260 9892 17300 9932
rect 20428 9892 20468 9932
rect 20716 9892 20756 9932
rect 23308 9892 23348 9932
rect 29356 9892 29396 9932
rect 4352 9808 4720 9848
rect 9388 9808 9428 9848
rect 11596 9808 11636 9848
rect 12126 9808 12494 9848
rect 17452 9808 17492 9848
rect 19900 9808 20268 9848
rect 20620 9808 20660 9848
rect 24460 9808 24500 9848
rect 25612 9808 25652 9848
rect 27674 9808 28042 9848
rect 3628 9724 3668 9764
rect 1036 9472 1076 9512
rect 1516 9472 1556 9512
rect 7564 9724 7604 9764
rect 2188 9640 2228 9680
rect 3052 9640 3092 9680
rect 4300 9640 4340 9680
rect 5932 9640 5972 9680
rect 2956 9556 2996 9596
rect 7468 9640 7499 9680
rect 7499 9640 7508 9680
rect 7852 9640 7892 9680
rect 8908 9640 8948 9680
rect 6618 9556 6658 9596
rect 8332 9556 8361 9596
rect 8361 9556 8372 9596
rect 16012 9724 16052 9764
rect 21676 9724 21716 9764
rect 9196 9640 9236 9680
rect 10348 9640 10388 9680
rect 10828 9640 10868 9680
rect 11404 9640 11444 9680
rect 11596 9640 11636 9680
rect 11884 9640 11924 9680
rect 12364 9640 12404 9680
rect 14956 9640 14996 9680
rect 17164 9640 17204 9680
rect 18316 9640 18356 9680
rect 18508 9640 18548 9680
rect 19372 9640 19412 9680
rect 19852 9640 19892 9680
rect 22636 9640 22676 9680
rect 10540 9556 10580 9596
rect 11212 9556 11252 9596
rect 13516 9556 13556 9596
rect 18700 9556 18740 9596
rect 19564 9556 19604 9596
rect 20140 9556 20171 9596
rect 20171 9556 20180 9596
rect 2188 9472 2228 9512
rect 2668 9472 2708 9512
rect 5644 9472 5684 9512
rect 5932 9472 5972 9512
rect 7372 9472 7412 9512
rect 7948 9472 7988 9512
rect 8140 9472 8180 9512
rect 1804 9388 1844 9428
rect 1996 9388 2036 9428
rect 2572 9388 2612 9428
rect 2860 9388 2900 9428
rect 5836 9388 5876 9428
rect 6220 9388 6260 9428
rect 10444 9472 10484 9512
rect 10636 9472 10648 9512
rect 10648 9472 10676 9512
rect 10924 9472 10964 9512
rect 7084 9388 7124 9428
rect 7756 9388 7796 9428
rect 8716 9388 8756 9428
rect 5260 9304 5300 9344
rect 11404 9472 11444 9512
rect 11692 9472 11732 9512
rect 12076 9472 12116 9512
rect 12940 9472 12980 9512
rect 13228 9472 13268 9512
rect 13612 9472 13652 9512
rect 13900 9472 13940 9512
rect 14284 9503 14324 9512
rect 14284 9472 14315 9503
rect 14315 9472 14324 9503
rect 11884 9388 11924 9428
rect 13036 9388 13076 9428
rect 14860 9472 14900 9512
rect 15436 9472 15476 9512
rect 14956 9388 14996 9428
rect 13228 9304 13268 9344
rect 15820 9503 15860 9512
rect 15820 9472 15851 9503
rect 15851 9472 15860 9503
rect 16108 9472 16148 9512
rect 17452 9472 17492 9512
rect 17836 9472 17876 9512
rect 19276 9472 19316 9512
rect 17260 9388 17300 9428
rect 17644 9388 17684 9428
rect 18316 9388 18356 9428
rect 19180 9388 19220 9428
rect 19468 9388 19508 9428
rect 18700 9304 18740 9344
rect 1324 9220 1364 9260
rect 3628 9220 3668 9260
rect 5932 9220 5972 9260
rect 8332 9220 8372 9260
rect 13612 9220 13652 9260
rect 14380 9220 14420 9260
rect 6028 9136 6068 9176
rect 13228 9136 13268 9176
rect 268 9052 308 9092
rect 3112 9052 3480 9092
rect 9772 9052 9812 9092
rect 10886 9052 11254 9092
rect 18660 9052 19028 9092
rect 9196 8968 9236 9008
rect 11404 8968 11444 9008
rect 1228 8884 1259 8924
rect 1259 8884 1268 8924
rect 1996 8884 2036 8924
rect 2572 8884 2612 8924
rect 3916 8884 3947 8924
rect 3947 8884 3956 8924
rect 8332 8884 8363 8924
rect 8363 8884 8372 8924
rect 2380 8800 2420 8840
rect 2764 8800 2804 8840
rect 2284 8716 2324 8756
rect 3916 8632 3956 8672
rect 4300 8632 4340 8672
rect 1804 8548 1844 8588
rect 2380 8548 2420 8588
rect 5164 8716 5204 8756
rect 19948 9304 19988 9344
rect 20140 9304 20180 9344
rect 24844 9556 24884 9596
rect 25804 9556 25844 9596
rect 27052 9724 27092 9764
rect 27436 9640 27476 9680
rect 28108 9640 28148 9680
rect 28684 9640 28724 9680
rect 26860 9556 26900 9596
rect 28300 9556 28340 9596
rect 30220 9556 30260 9596
rect 30508 9556 30548 9596
rect 31180 9556 31220 9596
rect 23308 9472 23348 9512
rect 23788 9472 23819 9512
rect 23819 9472 23828 9512
rect 24364 9472 24376 9512
rect 24376 9472 24404 9512
rect 20428 9388 20468 9428
rect 20908 9388 20939 9428
rect 20939 9388 20948 9428
rect 21772 9388 21812 9428
rect 23500 9388 23540 9428
rect 25036 9472 25076 9512
rect 25900 9472 25940 9512
rect 27244 9472 27284 9512
rect 27532 9472 27563 9512
rect 27563 9472 27572 9512
rect 28108 9472 28148 9512
rect 30412 9472 30452 9512
rect 30892 9472 30923 9512
rect 30923 9472 30932 9512
rect 24652 9388 24692 9428
rect 26284 9388 26324 9428
rect 27052 9388 27092 9428
rect 29356 9388 29387 9428
rect 29387 9388 29396 9428
rect 31084 9388 31124 9428
rect 23308 9304 23348 9344
rect 24460 9304 24500 9344
rect 26956 9304 26996 9344
rect 28300 9304 28340 9344
rect 28972 9304 29012 9344
rect 23788 9220 23819 9260
rect 23819 9220 23828 9260
rect 26860 9220 26900 9260
rect 20428 9136 20468 9176
rect 21964 9136 22004 9176
rect 23692 9052 23732 9092
rect 19948 8968 19988 9008
rect 21292 8968 21332 9008
rect 21580 8968 21620 9008
rect 12844 8884 12884 8924
rect 13708 8884 13748 8924
rect 14572 8884 14612 8924
rect 16684 8884 16724 8924
rect 12076 8800 12116 8840
rect 9100 8716 9140 8756
rect 11212 8716 11252 8756
rect 11404 8716 11444 8756
rect 13612 8716 13652 8756
rect 14572 8716 14612 8756
rect 15052 8716 15092 8756
rect 6028 8632 6068 8672
rect 7084 8632 7124 8672
rect 9004 8632 9044 8672
rect 9292 8632 9332 8672
rect 9772 8632 9812 8672
rect 10348 8632 10388 8672
rect 11500 8632 11507 8672
rect 11507 8632 11540 8672
rect 11692 8632 11732 8672
rect 12268 8632 12299 8672
rect 12299 8632 12308 8672
rect 17548 8800 17588 8840
rect 18124 8800 18164 8840
rect 15724 8716 15747 8756
rect 15747 8716 15764 8756
rect 16108 8716 16148 8756
rect 16876 8716 16916 8756
rect 12460 8632 12500 8672
rect 14764 8632 14804 8672
rect 15436 8632 15476 8672
rect 18028 8716 18068 8756
rect 18508 8716 18548 8756
rect 18316 8672 18356 8693
rect 16684 8632 16713 8672
rect 16713 8632 16724 8672
rect 18316 8653 18355 8672
rect 18355 8653 18356 8672
rect 20524 8800 20564 8840
rect 21772 8800 21812 8840
rect 24556 8800 24596 8840
rect 23308 8716 23348 8756
rect 24460 8716 24500 8756
rect 19564 8632 19604 8672
rect 23404 8632 23444 8672
rect 23980 8632 24020 8672
rect 26434 9052 26802 9092
rect 27532 8884 27572 8924
rect 28972 8884 29012 8924
rect 24844 8800 24884 8840
rect 25996 8800 26036 8840
rect 26572 8800 26612 8840
rect 30988 8800 31028 8840
rect 24940 8716 24980 8756
rect 28876 8716 28916 8756
rect 30124 8716 30164 8756
rect 26956 8632 26996 8672
rect 28108 8632 28148 8672
rect 29356 8632 29396 8672
rect 29836 8632 29876 8672
rect 30508 8632 30547 8672
rect 30547 8632 30548 8672
rect 5740 8548 5771 8588
rect 5771 8548 5780 8588
rect 6988 8548 7028 8588
rect 8812 8548 8852 8588
rect 13996 8548 14036 8588
rect 16300 8548 16340 8588
rect 16876 8548 16916 8588
rect 17164 8548 17204 8588
rect 18316 8548 18356 8588
rect 19084 8548 19124 8588
rect 19756 8548 19796 8588
rect 23884 8548 23924 8588
rect 748 8464 788 8504
rect 7276 8464 7316 8504
rect 10444 8464 10484 8504
rect 11500 8464 11540 8504
rect 1804 8380 1844 8420
rect 4352 8296 4720 8336
rect 3820 8212 3860 8252
rect 14380 8464 14420 8504
rect 16780 8464 16820 8504
rect 17836 8464 17876 8504
rect 17068 8380 17108 8420
rect 12126 8296 12494 8336
rect 17932 8296 17972 8336
rect 19276 8296 19316 8336
rect 14956 8212 14996 8252
rect 18412 8212 18452 8252
rect 28780 8464 28820 8504
rect 30412 8464 30452 8504
rect 19900 8296 20268 8336
rect 27674 8296 28042 8336
rect 25036 8212 25076 8252
rect 2764 8128 2804 8168
rect 3532 8128 3572 8168
rect 4108 8128 4148 8168
rect 5164 8128 5204 8168
rect 6988 8128 7028 8168
rect 16684 8128 16724 8168
rect 16876 8128 16916 8168
rect 17356 8128 17396 8168
rect 18124 8128 18164 8168
rect 19084 8128 19124 8168
rect 19468 8128 19508 8168
rect 19852 8128 19892 8168
rect 23116 8128 23156 8168
rect 28108 8128 28148 8168
rect 28876 8128 28916 8168
rect 29836 8128 29876 8168
rect 30124 8128 30164 8168
rect 2476 8044 2516 8084
rect 2380 7960 2420 8000
rect 1516 7876 1556 7916
rect 3052 7960 3092 8000
rect 5548 7960 5579 8000
rect 5579 7960 5588 8000
rect 6892 8044 6932 8084
rect 7276 8044 7316 8084
rect 12364 8044 12404 8084
rect 12556 8044 12596 8084
rect 17932 8044 17961 8084
rect 17961 8044 17972 8084
rect 1708 7792 1748 7832
rect 6700 7960 6740 8000
rect 7084 7960 7124 8000
rect 7852 7960 7892 8000
rect 8908 7960 8948 8000
rect 9676 7960 9716 8000
rect 3532 7792 3572 7832
rect 7372 7876 7412 7916
rect 14092 7960 14132 8000
rect 15628 7960 15668 8000
rect 16108 7960 16148 8000
rect 17068 7960 17108 8000
rect 18412 7960 18452 8000
rect 19276 7960 19305 8000
rect 19305 7960 19316 8000
rect 20428 7960 20468 8000
rect 15148 7876 15188 7916
rect 15340 7876 15380 7916
rect 18604 7876 18627 7916
rect 18627 7876 18644 7916
rect 7276 7792 7316 7832
rect 12748 7792 12788 7832
rect 19468 7876 19508 7916
rect 18220 7792 18260 7832
rect 18412 7792 18452 7832
rect 2764 7708 2804 7748
rect 7084 7708 7124 7748
rect 9484 7708 9524 7748
rect 14956 7708 14996 7748
rect 460 7624 500 7664
rect 1804 7624 1844 7664
rect 14284 7624 14324 7664
rect 3112 7540 3480 7580
rect 10886 7540 11254 7580
rect 18660 7540 19028 7580
rect 1612 7456 1652 7496
rect 17068 7456 17108 7496
rect 1516 7372 1547 7412
rect 1547 7372 1556 7412
rect 2956 7372 2996 7412
rect 4108 7372 4148 7412
rect 7276 7372 7316 7412
rect 8908 7372 8948 7412
rect 12364 7372 12404 7412
rect 12748 7372 12779 7412
rect 12779 7372 12788 7412
rect 15724 7372 15764 7412
rect 18412 7372 18452 7412
rect 2764 7204 2804 7244
rect 4492 7204 4532 7244
rect 4780 7204 4820 7244
rect 1516 7120 1556 7160
rect 1708 7120 1748 7160
rect 2188 7120 2228 7160
rect 3532 7120 3572 7160
rect 4108 7120 4148 7160
rect 20428 7372 20459 7412
rect 20459 7372 20468 7412
rect 22828 8044 22868 8084
rect 23788 8044 23828 8084
rect 26860 8044 26900 8084
rect 29932 8044 29972 8084
rect 21676 7991 21716 8000
rect 21676 7960 21716 7991
rect 21964 7960 22004 8000
rect 22636 7960 22676 8000
rect 23980 7960 24020 8000
rect 25996 7960 26027 8000
rect 26027 7960 26036 8000
rect 30028 7960 30068 8000
rect 30316 7960 30356 8000
rect 24652 7876 24692 7916
rect 26572 7876 26612 7916
rect 28396 7876 28436 7916
rect 29836 7876 29876 7916
rect 31084 7792 31124 7832
rect 21484 7708 21524 7748
rect 30604 7708 30644 7748
rect 26434 7540 26802 7580
rect 21484 7372 21524 7412
rect 23500 7372 23540 7412
rect 28396 7372 28436 7412
rect 30028 7372 30068 7412
rect 9484 7288 9524 7328
rect 24652 7288 24692 7328
rect 28876 7288 28916 7328
rect 8236 7204 8276 7244
rect 4972 7120 4983 7160
rect 4983 7120 5012 7160
rect 6700 7120 6740 7160
rect 6892 7120 6923 7160
rect 6923 7120 6932 7160
rect 8140 7120 8180 7160
rect 8620 7120 8660 7160
rect 1228 7036 1268 7076
rect 1516 6952 1556 6992
rect 1996 6952 2036 6992
rect 2188 6952 2228 6992
rect 1900 6784 1940 6824
rect 4012 7036 4052 7076
rect 2860 6952 2900 6992
rect 4352 6784 4720 6824
rect 9388 7036 9428 7076
rect 2764 6700 2804 6740
rect 3532 6700 3572 6740
rect 2188 6616 2228 6656
rect 3628 6532 3668 6572
rect 4972 6700 5012 6740
rect 6220 6616 6251 6656
rect 6251 6616 6260 6656
rect 8716 6952 8747 6992
rect 8747 6952 8756 6992
rect 10156 7193 10196 7202
rect 10156 7162 10196 7193
rect 8620 6616 8660 6656
rect 14284 7204 14324 7244
rect 11788 7120 11828 7160
rect 12556 7120 12587 7160
rect 12587 7120 12596 7160
rect 13036 7120 13076 7160
rect 13420 7036 13460 7076
rect 11788 6952 11828 6992
rect 12556 6952 12596 6992
rect 12126 6784 12494 6824
rect 8140 6532 8180 6572
rect 9004 6532 9044 6572
rect 10060 6532 10100 6572
rect 12940 6532 12980 6572
rect 19084 7204 19124 7244
rect 26764 7204 26804 7244
rect 27532 7204 27571 7244
rect 27571 7204 27572 7244
rect 28780 7204 28820 7244
rect 29740 7288 29780 7328
rect 30316 7204 30356 7244
rect 30604 7204 30610 7244
rect 30610 7204 30644 7244
rect 15148 7120 15188 7160
rect 15628 7120 15668 7160
rect 17932 7120 17972 7160
rect 18604 7120 18644 7160
rect 20044 7120 20084 7160
rect 21292 7120 21332 7160
rect 21484 7120 21524 7160
rect 23116 7120 23156 7160
rect 23500 7120 23540 7160
rect 25036 7120 25064 7160
rect 25064 7120 25076 7160
rect 26284 7120 26324 7160
rect 28108 7120 28148 7160
rect 29644 7120 29684 7160
rect 30028 7120 30068 7160
rect 30700 7120 30740 7160
rect 14860 7036 14900 7076
rect 20524 7036 20564 7076
rect 18412 6952 18452 6992
rect 17932 6868 17972 6908
rect 15148 6616 15188 6656
rect 16204 6616 16244 6656
rect 16972 6616 17012 6656
rect 15340 6532 15380 6572
rect 24364 7036 24404 7076
rect 28204 7036 28235 7076
rect 28235 7036 28244 7076
rect 28780 7036 28820 7076
rect 29260 7036 29300 7076
rect 29548 7036 29588 7076
rect 30124 7036 30164 7076
rect 20620 6952 20660 6992
rect 23212 6952 23252 6992
rect 23404 6952 23444 6992
rect 23596 6952 23636 6992
rect 23980 6952 24020 6992
rect 24268 6952 24308 6992
rect 29164 6952 29204 6992
rect 23884 6868 23924 6908
rect 19900 6784 20268 6824
rect 23596 6784 23636 6824
rect 18220 6700 18260 6740
rect 20524 6700 20564 6740
rect 20620 6616 20660 6656
rect 27674 6784 28042 6824
rect 22540 6616 22580 6656
rect 26764 6616 26795 6656
rect 26795 6616 26804 6656
rect 29548 6616 29579 6656
rect 29579 6616 29588 6656
rect 17932 6532 17972 6572
rect 23404 6532 23444 6572
rect 28396 6532 28436 6572
rect 29164 6532 29204 6572
rect 29452 6532 29492 6572
rect 1612 6448 1652 6488
rect 2188 6448 2228 6488
rect 2476 6448 2516 6488
rect 4204 6448 4244 6488
rect 4396 6448 4436 6488
rect 8236 6479 8276 6488
rect 8236 6448 8276 6479
rect 9196 6448 9236 6488
rect 9484 6448 9524 6488
rect 9676 6448 9716 6488
rect 11980 6448 12020 6488
rect 14284 6448 14324 6488
rect 14956 6448 14996 6488
rect 16396 6448 16436 6488
rect 17548 6448 17588 6488
rect 18124 6448 18125 6488
rect 18125 6448 18164 6488
rect 19180 6448 19220 6488
rect 20332 6448 20363 6488
rect 20363 6448 20372 6488
rect 22060 6448 22100 6488
rect 22348 6448 22388 6488
rect 23500 6448 23540 6488
rect 25228 6448 25259 6488
rect 25259 6448 25268 6488
rect 27820 6448 27860 6488
rect 28300 6448 28340 6488
rect 28780 6448 28820 6488
rect 30604 6448 30644 6488
rect 556 6364 596 6404
rect 2284 6364 2324 6404
rect 2764 6364 2804 6404
rect 3532 6364 3572 6404
rect 3916 6364 3956 6404
rect 6028 6364 6059 6404
rect 6059 6364 6068 6404
rect 7084 6364 7124 6404
rect 11500 6364 11540 6404
rect 13900 6364 13940 6404
rect 14188 6364 14228 6404
rect 14860 6364 14891 6404
rect 14891 6364 14900 6404
rect 16492 6364 16532 6404
rect 17644 6364 17684 6404
rect 22252 6364 22292 6404
rect 24172 6364 24212 6404
rect 24940 6364 24980 6404
rect 25612 6364 25652 6404
rect 27340 6364 27380 6404
rect 28012 6364 28052 6404
rect 29260 6364 29300 6404
rect 30508 6364 30514 6404
rect 30514 6364 30548 6404
rect 2860 6280 2900 6320
rect 5932 6280 5972 6320
rect 6604 6280 6644 6320
rect 12556 6280 12596 6320
rect 13420 6280 13460 6320
rect 16780 6280 16820 6320
rect 20140 6280 20180 6320
rect 22828 6280 22868 6320
rect 25516 6280 25556 6320
rect 4300 6196 4340 6236
rect 16108 6196 16139 6236
rect 16139 6196 16148 6236
rect 18412 6196 18452 6236
rect 20716 6196 20756 6236
rect 25996 6196 26027 6236
rect 26027 6196 26036 6236
rect 76 6112 116 6152
rect 6796 6112 6836 6152
rect 18508 6112 18548 6152
rect 28780 6112 28820 6152
rect 29260 6112 29300 6152
rect 30892 6112 30932 6152
rect 3112 6028 3480 6068
rect 6508 6028 6548 6068
rect 7084 6028 7124 6068
rect 10886 6028 11254 6068
rect 18660 6028 19028 6068
rect 26434 6028 26802 6068
rect 6700 5944 6740 5984
rect 17740 5944 17780 5984
rect 17932 5944 17972 5984
rect 21964 5944 22004 5984
rect 27820 5944 27860 5984
rect 29644 5944 29684 5984
rect 4396 5860 4436 5900
rect 4684 5776 4724 5816
rect 1228 5692 1268 5732
rect 2476 5692 2507 5732
rect 2507 5692 2516 5732
rect 3532 5692 3572 5732
rect 4204 5692 4244 5732
rect 652 5608 692 5648
rect 1708 5608 1748 5648
rect 2188 5608 2228 5648
rect 2860 5608 2900 5648
rect 2668 5440 2708 5480
rect 16492 5860 16523 5900
rect 16523 5860 16532 5900
rect 20428 5860 20468 5900
rect 21484 5860 21515 5900
rect 21515 5860 21524 5900
rect 25228 5860 25268 5900
rect 25612 5860 25652 5900
rect 30028 5860 30068 5900
rect 5740 5776 5780 5816
rect 6892 5776 6932 5816
rect 10060 5776 10100 5816
rect 17644 5776 17684 5816
rect 18412 5776 18452 5816
rect 22348 5776 22388 5816
rect 23116 5776 23156 5816
rect 29164 5776 29204 5816
rect 29836 5776 29876 5816
rect 6412 5692 6452 5732
rect 9100 5692 9140 5732
rect 10252 5692 10292 5732
rect 11308 5692 11348 5732
rect 12556 5692 12596 5732
rect 13036 5692 13076 5732
rect 3724 5608 3764 5648
rect 4300 5608 4340 5648
rect 4876 5608 4899 5648
rect 4899 5608 4916 5648
rect 5740 5608 5780 5648
rect 6124 5608 6164 5648
rect 7084 5608 7124 5648
rect 8716 5608 8756 5648
rect 4684 5524 4724 5564
rect 6316 5524 6356 5564
rect 8908 5524 8948 5564
rect 16396 5692 16436 5732
rect 16780 5692 16820 5732
rect 18028 5692 18068 5732
rect 18316 5692 18356 5732
rect 10060 5608 10100 5648
rect 11212 5608 11243 5648
rect 11243 5608 11252 5648
rect 12460 5608 12489 5648
rect 12489 5608 12500 5648
rect 12748 5608 12788 5648
rect 13228 5608 13268 5648
rect 14572 5608 14612 5648
rect 14860 5608 14900 5648
rect 17548 5608 17588 5648
rect 17836 5608 17876 5648
rect 21964 5608 22004 5648
rect 3724 5440 3764 5480
rect 4876 5440 4916 5480
rect 5932 5440 5972 5480
rect 6700 5440 6740 5480
rect 8140 5440 8180 5480
rect 1228 5188 1268 5228
rect 11884 5524 11924 5564
rect 4352 5272 4720 5312
rect 6892 5272 6932 5312
rect 8716 5272 8756 5312
rect 1708 5020 1748 5060
rect 3532 5104 3572 5144
rect 4108 5104 4148 5144
rect 11404 5440 11444 5480
rect 12940 5440 12980 5480
rect 6028 5104 6068 5144
rect 5356 5020 5396 5060
rect 8620 5020 8660 5060
rect 12126 5272 12494 5312
rect 12748 5356 12788 5396
rect 14572 5356 14612 5396
rect 12748 5188 12788 5228
rect 14476 5188 14516 5228
rect 12076 5020 12116 5060
rect 1516 4936 1556 4976
rect 1804 4936 1844 4976
rect 2380 4936 2420 4976
rect 3532 4936 3572 4976
rect 5452 4936 5492 4976
rect 7372 4936 7379 4976
rect 7379 4936 7412 4976
rect 8812 4936 8852 4976
rect 9004 4936 9044 4976
rect 9484 4936 9524 4976
rect 10252 4936 10292 4976
rect 10924 4936 10964 4976
rect 11980 4936 11986 4976
rect 11986 4936 12020 4976
rect 12556 4936 12596 4976
rect 13420 4936 13460 4976
rect 16108 5524 16148 5564
rect 18124 5524 18164 5564
rect 18124 5356 18164 5396
rect 15628 5272 15668 5312
rect 19900 5272 20268 5312
rect 20716 5440 20747 5480
rect 20747 5440 20756 5480
rect 16492 5188 16532 5228
rect 18412 5188 18452 5228
rect 16588 5020 16628 5060
rect 17356 5020 17396 5060
rect 18316 5020 18356 5060
rect 18796 5020 18836 5060
rect 29740 5692 29771 5732
rect 29771 5692 29780 5732
rect 30604 5860 30635 5900
rect 30635 5860 30644 5900
rect 22540 5608 22580 5648
rect 24076 5608 24116 5648
rect 25996 5608 26036 5648
rect 27148 5608 27188 5648
rect 28108 5608 28148 5648
rect 29452 5608 29492 5648
rect 29644 5608 29684 5648
rect 30124 5608 30164 5648
rect 30892 5608 30932 5648
rect 22252 5440 22292 5480
rect 24940 5440 24980 5480
rect 24556 5356 24596 5396
rect 21580 5104 21611 5144
rect 21611 5104 21620 5144
rect 23212 5188 23252 5228
rect 22924 5104 22955 5144
rect 22955 5104 22964 5144
rect 24172 5104 24212 5144
rect 18988 5020 19028 5060
rect 20716 5020 20756 5060
rect 28876 5524 28916 5564
rect 29548 5524 29588 5564
rect 30316 5524 30356 5564
rect 29452 5356 29492 5396
rect 27674 5272 28042 5312
rect 27532 5188 27572 5228
rect 15820 4936 15860 4976
rect 16012 4936 16052 4976
rect 16780 4936 16820 4976
rect 17164 4936 17193 4976
rect 17193 4936 17204 4976
rect 17644 4936 17684 4976
rect 18124 4936 18164 4976
rect 20524 4936 20564 4976
rect 21676 4936 21716 4976
rect 23116 4936 23156 4976
rect 23500 4936 23540 4976
rect 23884 4936 23924 4976
rect 25708 4936 25748 4976
rect 30508 5104 30539 5144
rect 30539 5104 30548 5144
rect 27244 5020 27284 5060
rect 27532 5020 27572 5060
rect 26092 4936 26132 4976
rect 27148 4936 27188 4976
rect 28012 4936 28052 4976
rect 28300 4936 28329 4976
rect 28329 4936 28340 4976
rect 29068 4936 29080 4976
rect 29080 4936 29108 4976
rect 29356 4936 29396 4976
rect 30508 4936 30548 4976
rect 3628 4852 3668 4892
rect 7468 4852 7499 4892
rect 7499 4852 7508 4892
rect 10636 4852 10676 4892
rect 11212 4852 11252 4892
rect 11884 4852 11924 4892
rect 13036 4852 13076 4892
rect 15916 4852 15956 4892
rect 13228 4768 13268 4808
rect 7756 4684 7796 4724
rect 10060 4684 10100 4724
rect 13132 4684 13172 4724
rect 8812 4600 8852 4640
rect 3112 4516 3480 4556
rect 10886 4516 11254 4556
rect 19084 4852 19124 4892
rect 24844 4852 24884 4892
rect 28588 4852 28628 4892
rect 17260 4768 17300 4808
rect 23500 4768 23540 4808
rect 24076 4768 24116 4808
rect 28492 4768 28532 4808
rect 17068 4684 17108 4724
rect 19084 4684 19124 4724
rect 20524 4684 20564 4724
rect 23116 4684 23156 4724
rect 27244 4684 27284 4724
rect 30316 4684 30356 4724
rect 28204 4600 28244 4640
rect 18660 4516 19028 4556
rect 26434 4516 26802 4556
rect 11884 4432 11924 4472
rect 13036 4432 13076 4472
rect 1804 4348 1844 4388
rect 3532 4348 3572 4388
rect 7372 4348 7412 4388
rect 8524 4348 8564 4388
rect 1612 4264 1652 4304
rect 9484 4348 9524 4388
rect 11596 4348 11636 4388
rect 12748 4348 12788 4388
rect 13420 4348 13460 4388
rect 16396 4348 16436 4388
rect 18316 4348 18356 4388
rect 20716 4348 20756 4388
rect 5356 4180 5396 4220
rect 6892 4180 6932 4220
rect 13900 4264 13940 4304
rect 15052 4264 15092 4304
rect 18028 4264 18068 4304
rect 10252 4180 10292 4220
rect 11500 4180 11540 4220
rect 12556 4180 12596 4220
rect 28012 4432 28052 4472
rect 26092 4348 26132 4388
rect 1132 4096 1172 4136
rect 1612 4096 1652 4136
rect 2188 4096 2228 4136
rect 2380 4096 2420 4136
rect 4972 4096 5012 4136
rect 5452 4096 5492 4136
rect 7276 4096 7316 4136
rect 8524 4096 8555 4136
rect 8555 4096 8564 4136
rect 8812 4096 8852 4136
rect 9964 4096 10004 4136
rect 11308 4096 11348 4136
rect 11596 4096 11636 4136
rect 13228 4096 13268 4136
rect 13420 4096 13460 4136
rect 16012 4096 16043 4136
rect 16043 4096 16052 4136
rect 16492 4096 16532 4136
rect 16684 4096 16724 4136
rect 17548 4096 17555 4136
rect 17555 4096 17588 4136
rect 18028 4096 18068 4136
rect 18316 4096 18356 4136
rect 21100 4096 21140 4136
rect 22924 4096 22964 4136
rect 24172 4096 24212 4136
rect 25420 4096 25460 4136
rect 26380 4180 26420 4220
rect 28300 4264 28340 4304
rect 27148 4180 27188 4220
rect 2860 4012 2900 4052
rect 3916 4012 3956 4052
rect 6604 4012 6644 4052
rect 11884 4012 11924 4052
rect 13900 4012 13940 4052
rect 652 3928 692 3968
rect 1516 3928 1556 3968
rect 4876 3928 4916 3968
rect 5644 3844 5684 3884
rect 4352 3760 4720 3800
rect 2188 3676 2228 3716
rect 3916 3676 3956 3716
rect 8716 3928 8756 3968
rect 10060 3928 10091 3968
rect 10091 3928 10100 3968
rect 11308 3928 11339 3968
rect 11339 3928 11348 3968
rect 12556 3928 12596 3968
rect 15916 3928 15956 3968
rect 16684 3928 16724 3968
rect 19468 3928 19499 3968
rect 19499 3928 19508 3968
rect 5452 3592 5492 3632
rect 5740 3592 5780 3632
rect 6028 3592 6068 3632
rect 6796 3592 6836 3632
rect 1420 3508 1460 3548
rect 3820 3508 3860 3548
rect 8812 3508 8852 3548
rect 10732 3592 10772 3632
rect 1132 3424 1172 3464
rect 1996 3424 2036 3464
rect 4684 3424 4724 3464
rect 4876 3424 4916 3464
rect 6124 3424 6164 3464
rect 6508 3424 6548 3464
rect 8524 3424 8564 3464
rect 10732 3424 10772 3464
rect 2476 3340 2516 3380
rect 10156 3340 10196 3380
rect 4684 3256 4724 3296
rect 4972 3256 5012 3296
rect 6124 3256 6164 3296
rect 6892 3256 6932 3296
rect 3532 3172 3572 3212
rect 7084 3172 7124 3212
rect 12126 3760 12494 3800
rect 13036 3592 13076 3632
rect 13324 3592 13355 3632
rect 13355 3592 13364 3632
rect 11884 3508 11924 3548
rect 26476 4096 26492 4136
rect 26492 4096 26516 4136
rect 28012 4180 28052 4220
rect 29356 4264 29396 4304
rect 30220 4264 30260 4304
rect 30700 4180 30740 4220
rect 27436 4096 27476 4136
rect 29740 4096 29780 4136
rect 30316 4096 30356 4136
rect 25804 4012 25844 4052
rect 23596 3928 23636 3968
rect 19900 3760 20268 3800
rect 17644 3676 17684 3716
rect 16588 3592 16628 3632
rect 17356 3592 17396 3632
rect 17548 3592 17588 3632
rect 20524 3676 20564 3716
rect 18316 3508 18356 3548
rect 11788 3424 11828 3464
rect 12172 3424 12212 3464
rect 12460 3424 12500 3464
rect 13228 3424 13268 3464
rect 13804 3424 13833 3464
rect 13833 3424 13844 3464
rect 14284 3424 14324 3464
rect 14572 3424 14612 3464
rect 15052 3424 15059 3464
rect 15059 3424 15092 3464
rect 15820 3424 15860 3464
rect 16492 3424 16532 3464
rect 18124 3424 18136 3464
rect 18136 3424 18164 3464
rect 18508 3424 18548 3464
rect 16396 3340 16436 3380
rect 22252 3592 22283 3632
rect 22283 3592 22292 3632
rect 22828 3592 22868 3632
rect 19276 3424 19316 3464
rect 19660 3424 19700 3464
rect 20140 3424 20180 3464
rect 20524 3424 20564 3464
rect 21676 3424 21716 3464
rect 21964 3424 22004 3464
rect 22636 3424 22676 3464
rect 24844 3928 24875 3968
rect 24875 3928 24884 3968
rect 26572 4012 26612 4052
rect 27340 4012 27380 4052
rect 28204 4012 28244 4052
rect 30508 4012 30548 4052
rect 28780 3928 28820 3968
rect 25420 3844 25460 3884
rect 27674 3760 28042 3800
rect 25324 3676 25364 3716
rect 26380 3676 26420 3716
rect 27148 3676 27188 3716
rect 28204 3676 28244 3716
rect 29740 3676 29780 3716
rect 25420 3592 25460 3632
rect 25804 3592 25844 3632
rect 26572 3592 26612 3632
rect 29356 3592 29396 3632
rect 28588 3508 28628 3548
rect 28876 3508 28916 3548
rect 24172 3424 24212 3464
rect 24940 3424 24980 3464
rect 27052 3424 27092 3464
rect 27532 3424 27572 3464
rect 28204 3424 28244 3464
rect 28780 3424 28820 3464
rect 30412 3424 30452 3464
rect 23212 3340 23252 3380
rect 13132 3256 13172 3296
rect 14572 3256 14612 3296
rect 17644 3256 17684 3296
rect 30220 3340 30260 3380
rect 25708 3256 25748 3296
rect 14476 3172 14507 3212
rect 14507 3172 14516 3212
rect 19276 3172 19316 3212
rect 20236 3172 20276 3212
rect 23788 3172 23828 3212
rect 28780 3172 28820 3212
rect 29356 3172 29396 3212
rect 8716 3088 8756 3128
rect 12172 3088 12212 3128
rect 14860 3088 14900 3128
rect 18220 3088 18260 3128
rect 21004 3088 21044 3128
rect 22924 3088 22964 3128
rect 24940 3088 24980 3128
rect 3112 3004 3480 3044
rect 10886 3004 11254 3044
rect 18660 3004 19028 3044
rect 26434 3004 26802 3044
rect 3916 2836 3956 2876
rect 7468 2836 7508 2876
rect 10636 2836 10676 2876
rect 13228 2836 13268 2876
rect 13708 2836 13748 2876
rect 17068 2836 17108 2876
rect 18508 2836 18548 2876
rect 21100 2836 21140 2876
rect 22828 2836 22868 2876
rect 28876 2836 28916 2876
rect 2476 2752 2516 2792
rect 4588 2752 4628 2792
rect 4876 2752 4916 2792
rect 1132 2668 1172 2708
rect 1324 2668 1347 2708
rect 1347 2668 1364 2708
rect 3628 2668 3668 2708
rect 6700 2752 6740 2792
rect 6892 2752 6932 2792
rect 7084 2668 7124 2708
rect 3532 2584 3563 2624
rect 3563 2584 3572 2624
rect 4588 2584 4628 2624
rect 5836 2584 5876 2624
rect 15916 2752 15956 2792
rect 16204 2752 16244 2792
rect 17356 2752 17396 2792
rect 19276 2752 19316 2792
rect 22636 2752 22676 2792
rect 9388 2668 9428 2708
rect 12460 2668 12491 2708
rect 12491 2668 12500 2708
rect 14764 2668 14804 2708
rect 16396 2668 16436 2708
rect 17644 2668 17684 2708
rect 19180 2668 19220 2708
rect 8908 2584 8948 2624
rect 11500 2584 11540 2624
rect 12172 2584 12212 2624
rect 12556 2584 12596 2624
rect 13132 2584 13163 2624
rect 13163 2584 13172 2624
rect 13708 2584 13748 2624
rect 14476 2584 14516 2624
rect 14860 2584 14900 2624
rect 17164 2584 17204 2624
rect 18508 2584 18548 2624
rect 19660 2584 19700 2624
rect 20236 2584 20247 2624
rect 20247 2584 20276 2624
rect 1516 2500 1556 2540
rect 2092 2500 2132 2540
rect 2860 2500 2900 2540
rect 4780 2500 4820 2540
rect 13036 2500 13076 2540
rect 14284 2500 14324 2540
rect 5740 2416 5780 2456
rect 4352 2248 4720 2288
rect 2092 2080 2132 2120
rect 1996 1912 2027 1952
rect 2027 1912 2036 1952
rect 4396 1912 4436 1952
rect 4780 1912 4820 1952
rect 6892 2080 6932 2120
rect 6028 1996 6068 2036
rect 6412 1912 6452 1952
rect 11308 2416 11348 2456
rect 16204 2500 16244 2540
rect 16588 2500 16628 2540
rect 17068 2500 17108 2540
rect 16684 2416 16724 2456
rect 17356 2416 17396 2456
rect 10156 2332 10196 2372
rect 11596 2332 11636 2372
rect 23212 2668 23252 2708
rect 23884 2668 23924 2708
rect 24076 2668 24116 2708
rect 26860 2752 26900 2792
rect 20620 2584 20660 2624
rect 21964 2584 22004 2624
rect 22156 2584 22196 2624
rect 22924 2584 22964 2624
rect 23788 2584 23828 2624
rect 20140 2500 20180 2540
rect 21868 2500 21908 2540
rect 21580 2416 21620 2456
rect 22348 2416 22388 2456
rect 22636 2416 22676 2456
rect 19756 2332 19796 2372
rect 22540 2332 22580 2372
rect 12126 2248 12494 2288
rect 13804 2248 13844 2288
rect 19900 2248 20268 2288
rect 18412 2164 18452 2204
rect 22156 2164 22196 2204
rect 10732 2080 10763 2120
rect 10763 2080 10772 2120
rect 13132 2080 13172 2120
rect 13804 2080 13844 2120
rect 10156 1996 10196 2036
rect 10636 1996 10676 2036
rect 8908 1912 8948 1952
rect 10732 1912 10772 1952
rect 11788 1912 11828 1952
rect 12172 1912 12212 1952
rect 12364 1996 12404 2036
rect 14284 2080 14315 2120
rect 14315 2080 14324 2120
rect 15820 2080 15860 2120
rect 18316 2080 18356 2120
rect 12556 1912 12596 1952
rect 13036 1912 13076 1952
rect 13324 1912 13364 1952
rect 13516 1912 13556 1952
rect 30316 2752 30356 2792
rect 29356 2668 29396 2708
rect 25228 2584 25268 2624
rect 25804 2584 25844 2624
rect 28204 2584 28244 2624
rect 23596 2500 23636 2540
rect 25996 2500 26036 2540
rect 28780 2500 28820 2540
rect 24172 2332 24212 2372
rect 24268 2248 24308 2288
rect 27674 2248 28042 2288
rect 21964 2080 22004 2120
rect 23116 2080 23156 2120
rect 27532 2080 27572 2120
rect 23980 1996 24020 2036
rect 16780 1912 16820 1952
rect 21868 1912 21908 1952
rect 22348 1912 22388 1952
rect 24172 1912 24203 1952
rect 24203 1912 24212 1952
rect 24460 1912 24500 1952
rect 25324 1912 25364 1952
rect 2668 1828 2708 1868
rect 3820 1828 3860 1868
rect 11500 1828 11540 1868
rect 17644 1828 17684 1868
rect 19180 1828 19220 1868
rect 20908 1828 20948 1868
rect 22636 1828 22676 1868
rect 22828 1828 22868 1868
rect 23500 1828 23540 1868
rect 24268 1828 24308 1868
rect 26860 1828 26900 1868
rect 28108 1828 28148 1868
rect 5836 1744 5876 1784
rect 6124 1744 6164 1784
rect 7564 1744 7604 1784
rect 16780 1744 16820 1784
rect 21004 1744 21044 1784
rect 23788 1744 23828 1784
rect 29836 1912 29876 1952
rect 30988 1912 31028 1952
rect 30988 1744 31028 1784
rect 4780 1660 4820 1700
rect 5740 1660 5780 1700
rect 13420 1660 13460 1700
rect 14764 1660 14804 1700
rect 18220 1660 18260 1700
rect 19084 1660 19124 1700
rect 23308 1660 23348 1700
rect 30796 1660 30836 1700
rect 2092 1576 2132 1616
rect 5932 1576 5972 1616
rect 6700 1576 6740 1616
rect 10732 1576 10772 1616
rect 3112 1492 3480 1532
rect 10886 1492 11254 1532
rect 18660 1492 19028 1532
rect 26434 1492 26802 1532
rect 4876 1408 4916 1448
rect 5548 1408 5588 1448
rect 13516 1408 13556 1448
rect 19660 1408 19700 1448
rect 8428 1324 8468 1364
rect 12556 1324 12596 1364
rect 12844 1324 12884 1364
rect 16876 1324 16916 1364
rect 23500 1324 23540 1364
rect 24460 1324 24500 1364
rect 29836 1324 29876 1364
rect 2668 1240 2708 1280
rect 4972 1240 5012 1280
rect 5164 1240 5204 1280
rect 11788 1240 11828 1280
rect 13036 1240 13076 1280
rect 13324 1240 13364 1280
rect 15052 1240 15092 1280
rect 19180 1240 19220 1280
rect 7564 1156 7604 1196
rect 16780 1156 16820 1196
rect 19084 1156 19124 1196
rect 5836 1114 5876 1154
rect 3820 1072 3860 1112
rect 4396 1072 4427 1112
rect 4427 1072 4436 1112
rect 4876 1072 4916 1112
rect 8524 1072 8564 1112
rect 10732 1072 10772 1112
rect 11596 1072 11636 1112
rect 12364 1072 12404 1112
rect 12940 1072 12980 1112
rect 13420 1072 13460 1112
rect 14764 1072 14804 1112
rect 15052 1072 15092 1112
rect 20908 1240 20948 1280
rect 21580 1240 21620 1280
rect 25324 1240 25364 1280
rect 23788 1156 23828 1196
rect 25228 1156 25268 1196
rect 30316 1156 30356 1196
rect 30796 1156 30827 1196
rect 30827 1156 30836 1196
rect 23116 1072 23147 1112
rect 23147 1072 23156 1112
rect 24076 1072 24116 1112
rect 25996 1072 26036 1112
rect 27532 1072 27572 1112
rect 30412 1072 30443 1112
rect 30443 1072 30452 1112
rect 5932 988 5972 1028
rect 5548 904 5579 944
rect 5579 904 5588 944
rect 6028 904 6068 944
rect 6412 820 6452 860
rect 4352 736 4720 776
rect 5740 736 5780 776
rect 10636 988 10676 1028
rect 11308 988 11348 1028
rect 12652 988 12692 1028
rect 13516 988 13547 1028
rect 13547 988 13556 1028
rect 12556 820 12596 860
rect 12126 736 12494 776
rect 18220 988 18260 1028
rect 19756 988 19796 1028
rect 23308 988 23348 1028
rect 15052 820 15092 860
rect 19900 736 20268 776
rect 27674 736 28042 776
<< metal3 >>
rect 3128 28600 3208 29000
rect 3896 28600 3976 29000
rect 4664 28600 4744 29000
rect 5432 28600 5512 29000
rect 6200 28600 6280 29000
rect 6968 28600 7048 29000
rect 7736 28600 7816 29000
rect 8504 28600 8584 29000
rect 9272 28600 9352 29000
rect 10040 28600 10120 29000
rect 10808 28600 10888 29000
rect 11576 28600 11656 29000
rect 12344 28600 12424 29000
rect 13112 28600 13192 29000
rect 13880 28600 13960 29000
rect 14648 28600 14728 29000
rect 15416 28600 15496 29000
rect 16184 28600 16264 29000
rect 16396 28664 16436 28673
rect 3148 27488 3188 28600
rect 3628 27656 3668 27665
rect 3148 27439 3188 27448
rect 3532 27572 3572 27581
rect 3112 27236 3480 27245
rect 3112 27187 3480 27196
rect 3532 26984 3572 27532
rect 3532 26935 3572 26944
rect 3628 26144 3668 27616
rect 3724 27404 3764 27413
rect 3724 26984 3764 27364
rect 3916 27068 3956 28600
rect 4684 28160 4724 28600
rect 4684 28120 4820 28160
rect 4352 27992 4720 28001
rect 4352 27943 4720 27952
rect 3916 27019 3956 27028
rect 3724 26228 3764 26944
rect 4780 26732 4820 28120
rect 4780 26683 4820 26692
rect 4876 26816 4916 26825
rect 4780 26564 4820 26573
rect 4352 26480 4720 26489
rect 4352 26431 4720 26440
rect 3724 26179 3764 26188
rect 3628 26095 3668 26104
rect 4204 25808 4244 25817
rect 3112 25724 3480 25733
rect 3112 25675 3480 25684
rect 3052 25388 3092 25397
rect 2572 25304 2612 25313
rect 2188 24632 2228 24641
rect 1900 24464 1940 24473
rect 1900 23876 1940 24424
rect 1900 23827 1940 23836
rect 2188 23708 2228 24592
rect 2188 23372 2228 23668
rect 2188 23323 2228 23332
rect 2572 23792 2612 25264
rect 3052 24464 3092 25348
rect 3052 24415 3092 24424
rect 4204 24632 4244 25768
rect 4780 25220 4820 26524
rect 4352 24968 4720 24977
rect 4352 24919 4720 24928
rect 4780 24884 4820 25180
rect 4780 24835 4820 24844
rect 4876 24716 4916 26776
rect 5452 26732 5492 28600
rect 5740 27572 5780 27581
rect 5452 26683 5492 26692
rect 5548 26984 5588 26993
rect 5068 26144 5108 26153
rect 5068 25472 5108 26104
rect 5068 25423 5108 25432
rect 5164 26060 5204 26069
rect 3532 24380 3572 24389
rect 3112 24212 3480 24221
rect 3112 24163 3480 24172
rect 844 23120 884 23129
rect 844 22532 884 23080
rect 844 22483 884 22492
rect 2092 22952 2132 22961
rect 2092 22364 2132 22912
rect 2092 22315 2132 22324
rect 2572 22280 2612 23752
rect 3532 23792 3572 24340
rect 3532 23743 3572 23752
rect 3628 24296 3668 24305
rect 3628 23624 3668 24256
rect 4204 23792 4244 24592
rect 4396 24632 4436 24641
rect 4396 23876 4436 24592
rect 3628 23120 3668 23584
rect 3628 23060 3668 23080
rect 3532 23020 3668 23060
rect 4108 23752 4204 23792
rect 3112 22700 3480 22709
rect 3112 22651 3480 22660
rect 364 21776 404 21785
rect 172 21736 364 21776
rect 76 18836 116 18845
rect 76 6152 116 18796
rect 172 13292 212 21736
rect 364 21727 404 21736
rect 652 21608 692 21617
rect 652 21020 692 21568
rect 652 20971 692 20980
rect 1996 21272 2036 21281
rect 1228 20684 1268 20693
rect 556 20516 596 20525
rect 460 20432 500 20441
rect 172 13243 212 13252
rect 268 16484 308 16493
rect 268 9092 308 16444
rect 268 9043 308 9052
rect 460 7664 500 20392
rect 460 7615 500 7624
rect 556 6404 596 20476
rect 940 20180 980 20189
rect 748 19760 788 19769
rect 652 16820 692 16829
rect 652 13544 692 16780
rect 652 13495 692 13504
rect 748 8504 788 19720
rect 844 19592 884 19601
rect 844 14216 884 19552
rect 940 14384 980 20140
rect 1228 19928 1268 20644
rect 1228 19879 1268 19888
rect 1324 20348 1364 20357
rect 1324 19844 1364 20308
rect 1324 19795 1364 19804
rect 1420 20264 1460 20273
rect 1324 19424 1364 19433
rect 1132 19340 1172 19349
rect 1036 19088 1076 19097
rect 1036 17492 1076 19048
rect 1132 18752 1172 19300
rect 1132 18703 1172 18712
rect 1036 17443 1076 17452
rect 1228 18500 1268 18509
rect 1228 16736 1268 18460
rect 1324 17912 1364 19384
rect 1420 17996 1460 20224
rect 1804 20096 1844 20105
rect 1708 20012 1748 20021
rect 1708 19340 1748 19972
rect 1804 19424 1844 20056
rect 1804 19375 1844 19384
rect 1708 19256 1748 19300
rect 1420 17947 1460 17956
rect 1516 19172 1556 19181
rect 1708 19176 1748 19216
rect 1324 17863 1364 17872
rect 1324 17492 1364 17501
rect 1324 17072 1364 17452
rect 1324 17023 1364 17032
rect 1228 16687 1268 16696
rect 1036 16232 1076 16241
rect 1036 16097 1076 16192
rect 1228 16148 1268 16157
rect 1228 15392 1268 16108
rect 1228 15343 1268 15352
rect 1420 15644 1460 15653
rect 1228 14888 1268 14897
rect 1228 14720 1268 14848
rect 1228 14671 1268 14680
rect 940 14335 980 14344
rect 1036 14636 1076 14645
rect 844 14176 980 14216
rect 940 12704 980 14176
rect 940 12655 980 12664
rect 1036 10184 1076 14596
rect 1324 14636 1364 14645
rect 1228 14468 1268 14477
rect 1228 13964 1268 14428
rect 1228 13915 1268 13924
rect 1324 14048 1364 14596
rect 1324 12536 1364 14008
rect 1324 12487 1364 12496
rect 1420 13208 1460 15604
rect 1324 12284 1364 12293
rect 1228 12200 1268 12209
rect 1132 11612 1172 11621
rect 1132 10856 1172 11572
rect 1132 10807 1172 10816
rect 1036 9512 1076 10144
rect 1036 9463 1076 9472
rect 748 8455 788 8464
rect 1228 8924 1268 12160
rect 1324 11108 1364 12244
rect 1324 11059 1364 11068
rect 1420 11696 1460 13168
rect 1324 10940 1364 10949
rect 1324 10184 1364 10900
rect 1324 10135 1364 10144
rect 556 6355 596 6364
rect 1228 7076 1268 8884
rect 76 6103 116 6112
rect 1228 5732 1268 7036
rect 652 5648 692 5657
rect 652 3968 692 5608
rect 1228 5228 1268 5692
rect 1132 5188 1228 5228
rect 1132 4136 1172 5188
rect 1228 5179 1268 5188
rect 1324 9260 1364 9269
rect 1132 4087 1172 4096
rect 652 3919 692 3928
rect 1132 3464 1172 3473
rect 1132 2708 1172 3424
rect 1132 2659 1172 2668
rect 1324 2708 1364 9220
rect 1420 3548 1460 11656
rect 1516 10940 1556 19132
rect 1900 19172 1940 19181
rect 1804 19004 1844 19013
rect 1612 18920 1652 18929
rect 1612 17660 1652 18880
rect 1708 18500 1748 18509
rect 1708 17996 1748 18460
rect 1708 17947 1748 17956
rect 1612 17240 1652 17620
rect 1612 16988 1652 17200
rect 1612 16939 1652 16948
rect 1708 17744 1748 17753
rect 1612 16316 1652 16325
rect 1612 14216 1652 16276
rect 1708 16316 1748 17704
rect 1708 16267 1748 16276
rect 1804 16316 1844 18964
rect 1900 18752 1940 19132
rect 1900 18703 1940 18712
rect 1996 18584 2036 21232
rect 2284 20852 2324 20861
rect 2284 20096 2324 20812
rect 2284 20047 2324 20056
rect 2572 20768 2612 22240
rect 2860 21608 2900 21617
rect 2668 21440 2708 21449
rect 2668 20852 2708 21400
rect 2668 20803 2708 20812
rect 2764 21356 2804 21365
rect 2380 19844 2420 19853
rect 2188 19340 2228 19349
rect 2092 19256 2132 19265
rect 2092 19121 2132 19216
rect 2188 19172 2228 19300
rect 2188 19123 2228 19132
rect 2380 19172 2420 19804
rect 2380 19123 2420 19132
rect 2092 18836 2132 18845
rect 2092 18701 2132 18796
rect 1804 16267 1844 16276
rect 1900 18544 2036 18584
rect 2092 18584 2132 18593
rect 1804 16148 1844 16157
rect 1804 15560 1844 16108
rect 1804 15511 1844 15520
rect 1612 14167 1652 14176
rect 1708 15056 1748 15065
rect 1708 14888 1748 15016
rect 1708 14048 1748 14848
rect 1804 14720 1844 14729
rect 1804 14300 1844 14680
rect 1900 14552 1940 18544
rect 2092 18332 2132 18544
rect 2476 18584 2516 18593
rect 2092 18283 2132 18292
rect 2284 18500 2324 18509
rect 2188 18248 2228 18257
rect 2188 17240 2228 18208
rect 2188 17156 2228 17200
rect 2284 17744 2324 18460
rect 2284 17240 2324 17704
rect 2284 17191 2324 17200
rect 2476 17576 2516 18544
rect 2572 17828 2612 20728
rect 2764 20180 2804 21316
rect 2860 20768 2900 21568
rect 3112 21188 3480 21197
rect 3112 21139 3480 21148
rect 2860 20719 2900 20728
rect 3148 20768 3188 20777
rect 2668 20140 2804 20180
rect 2956 20684 2996 20693
rect 2668 20096 2708 20140
rect 2668 20047 2708 20056
rect 2860 20096 2900 20105
rect 2860 19928 2900 20056
rect 2668 19888 2900 19928
rect 2956 19928 2996 20644
rect 3148 20264 3188 20728
rect 3148 20215 3188 20224
rect 3436 20768 3476 20777
rect 3436 20180 3476 20728
rect 3436 20131 3476 20140
rect 3340 20096 3380 20107
rect 3340 20012 3380 20056
rect 3340 19963 3380 19972
rect 2668 19340 2708 19888
rect 2956 19879 2996 19888
rect 2860 19760 2900 19769
rect 2860 19625 2900 19720
rect 3112 19676 3480 19685
rect 3112 19627 3480 19636
rect 2668 19291 2708 19300
rect 2956 19508 2996 19517
rect 2764 19256 2804 19265
rect 2764 18752 2804 19216
rect 2860 19172 2900 19181
rect 2956 19172 2996 19468
rect 3148 19340 3188 19349
rect 3148 19205 3188 19300
rect 2900 19132 2996 19172
rect 3052 19172 3092 19181
rect 2860 19123 2900 19132
rect 3052 19004 3092 19132
rect 3340 19172 3380 19181
rect 3532 19172 3572 23020
rect 3628 22868 3668 22877
rect 3628 22280 3668 22828
rect 3628 22231 3668 22240
rect 4108 21608 4148 23752
rect 4204 23743 4244 23752
rect 4300 23836 4396 23876
rect 4300 23624 4340 23836
rect 4396 23827 4436 23836
rect 4780 23708 4820 23717
rect 4876 23708 4916 24676
rect 4820 23668 4916 23708
rect 4972 24632 5012 24641
rect 4972 23708 5012 24592
rect 5164 24632 5204 26020
rect 5548 26060 5588 26944
rect 5740 26144 5780 27532
rect 6220 26732 6260 28600
rect 6700 27572 6740 27581
rect 6700 26984 6740 27532
rect 6700 26935 6740 26944
rect 6220 26683 6260 26692
rect 6316 26816 6356 26825
rect 5740 26095 5780 26104
rect 5836 26228 5876 26237
rect 5548 26011 5588 26020
rect 5836 25976 5876 26188
rect 5740 25936 5876 25976
rect 6220 26144 6260 26153
rect 5644 25388 5684 25397
rect 5068 24464 5108 24473
rect 5068 24329 5108 24424
rect 5164 24128 5204 24592
rect 5164 24079 5204 24088
rect 5260 25304 5300 25313
rect 5260 24044 5300 25264
rect 5548 25304 5588 25313
rect 5452 24884 5492 24893
rect 5548 24884 5588 25264
rect 5492 24844 5588 24884
rect 5452 24835 5492 24844
rect 5644 24800 5684 25348
rect 5740 25304 5780 25936
rect 5740 25255 5780 25264
rect 5644 24632 5684 24760
rect 5644 24464 5684 24592
rect 5644 24415 5684 24424
rect 5836 25136 5876 25145
rect 5836 24464 5876 25096
rect 5836 24415 5876 24424
rect 6220 24632 6260 26104
rect 6316 25556 6356 26776
rect 6316 25507 6356 25516
rect 5260 23995 5300 24004
rect 5356 24380 5396 24389
rect 4780 23659 4820 23668
rect 4972 23659 5012 23668
rect 5356 23708 5396 24340
rect 5356 23659 5396 23668
rect 5548 23792 5588 23801
rect 4204 23584 4340 23624
rect 5260 23624 5300 23633
rect 4204 23288 4244 23584
rect 4352 23456 4720 23465
rect 4352 23407 4720 23416
rect 5260 23456 5300 23584
rect 4204 23248 4340 23288
rect 4300 23036 4340 23248
rect 4876 23204 4916 23213
rect 5260 23204 5300 23416
rect 4916 23164 5300 23204
rect 4876 23155 4916 23164
rect 4300 22364 4340 22996
rect 4300 22112 4340 22324
rect 4204 22072 4340 22112
rect 4972 22280 5012 22289
rect 4204 21776 4244 22072
rect 4352 21944 4720 21953
rect 4352 21895 4720 21904
rect 4204 21736 4340 21776
rect 4108 21559 4148 21568
rect 4012 21524 4052 21533
rect 3916 20684 3956 20693
rect 3820 20180 3860 20189
rect 3628 20096 3668 20105
rect 3628 19424 3668 20056
rect 3628 19375 3668 19384
rect 3724 20012 3764 20021
rect 3380 19132 3572 19172
rect 3340 19123 3380 19132
rect 2764 18703 2804 18712
rect 2860 18964 3092 19004
rect 2668 18584 2708 18593
rect 2668 18449 2708 18544
rect 2764 18500 2804 18509
rect 2764 18332 2804 18460
rect 2572 17779 2612 17788
rect 2668 18292 2804 18332
rect 2668 17828 2708 18292
rect 2092 17072 2132 17081
rect 1900 14503 1940 14512
rect 1996 16904 2036 16913
rect 1804 14251 1844 14260
rect 1708 13999 1748 14008
rect 1612 13796 1652 13805
rect 1612 11108 1652 13756
rect 1900 12368 1940 12377
rect 1612 11059 1652 11068
rect 1804 11948 1844 11957
rect 1516 10900 1652 10940
rect 1516 10772 1556 10781
rect 1516 9512 1556 10732
rect 1516 9463 1556 9472
rect 1516 7916 1556 7925
rect 1516 7412 1556 7876
rect 1612 7496 1652 10900
rect 1804 9428 1844 11908
rect 1900 11780 1940 12328
rect 1900 11731 1940 11740
rect 1996 10352 2036 16864
rect 2092 16064 2132 17032
rect 2188 16232 2228 17116
rect 2476 17156 2516 17536
rect 2284 16904 2324 16913
rect 2284 16484 2324 16864
rect 2284 16435 2324 16444
rect 2380 16820 2420 16829
rect 2188 16097 2228 16192
rect 2380 16148 2420 16780
rect 2092 16015 2132 16024
rect 2380 15560 2420 16108
rect 2476 16064 2516 17116
rect 2476 16015 2516 16024
rect 2572 17660 2612 17669
rect 2380 15511 2420 15520
rect 2380 14720 2420 14729
rect 2188 14384 2228 14393
rect 2188 14048 2228 14344
rect 2380 14216 2420 14680
rect 2380 14167 2420 14176
rect 2228 14008 2324 14048
rect 2188 13999 2228 14008
rect 2284 12536 2324 14008
rect 2284 12487 2324 12496
rect 2572 11276 2612 17620
rect 2668 16232 2708 17788
rect 2860 16988 2900 18964
rect 3148 18836 3188 18845
rect 3148 18701 3188 18796
rect 3724 18668 3764 19972
rect 3820 19172 3860 20140
rect 3916 20096 3956 20644
rect 3916 19340 3956 20056
rect 3916 19291 3956 19300
rect 3820 19123 3860 19132
rect 2956 18584 2996 18593
rect 2956 18080 2996 18544
rect 3112 18164 3480 18173
rect 3112 18115 3480 18124
rect 2956 18031 2996 18040
rect 3340 17996 3380 18005
rect 3340 17660 3380 17956
rect 3724 17996 3764 18628
rect 4012 18332 4052 21484
rect 4108 21104 4148 21113
rect 4108 20348 4148 21064
rect 4204 20768 4244 20863
rect 4300 20852 4340 21736
rect 4972 21692 5012 22240
rect 4972 21643 5012 21652
rect 4684 21608 4724 21617
rect 4684 21473 4724 21568
rect 4972 21524 5012 21533
rect 4300 20803 4340 20812
rect 4684 21188 4724 21197
rect 4204 20719 4244 20728
rect 4684 20768 4724 21148
rect 4972 21020 5012 21484
rect 4972 20971 5012 20980
rect 5164 21440 5204 21449
rect 4724 20728 4820 20768
rect 4684 20719 4724 20728
rect 4300 20684 4340 20693
rect 4300 20600 4340 20644
rect 4108 20299 4148 20308
rect 4204 20560 4340 20600
rect 4204 20096 4244 20560
rect 4352 20432 4720 20441
rect 4352 20383 4720 20392
rect 4204 20012 4244 20056
rect 4204 19932 4244 19972
rect 4300 20096 4340 20107
rect 4300 20012 4340 20056
rect 4300 19963 4340 19972
rect 4492 20096 4532 20105
rect 4204 19508 4244 19517
rect 4204 18752 4244 19468
rect 4492 19424 4532 20056
rect 4588 19760 4628 19769
rect 4588 19625 4628 19720
rect 4492 19256 4532 19384
rect 4780 19340 4820 20728
rect 5164 20684 5204 21400
rect 5260 20768 5300 23164
rect 5548 23036 5588 23752
rect 5548 22280 5588 22996
rect 5548 22231 5588 22240
rect 5932 23120 5972 23129
rect 5644 22112 5684 22121
rect 5644 21692 5684 22072
rect 5260 20719 5300 20728
rect 5356 21608 5396 21648
rect 5644 21643 5684 21652
rect 5356 21524 5396 21568
rect 5356 21020 5396 21484
rect 5164 20635 5204 20644
rect 5164 20096 5204 20105
rect 4972 20012 5012 20021
rect 4780 19291 4820 19300
rect 4876 19928 4916 19937
rect 4492 19207 4532 19216
rect 4352 18920 4720 18929
rect 4352 18871 4720 18880
rect 4204 18703 4244 18712
rect 4780 18668 4820 18677
rect 4012 18283 4052 18292
rect 4300 18584 4340 18593
rect 3340 17611 3380 17620
rect 3532 17744 3572 17753
rect 2860 16939 2900 16948
rect 2956 17576 2996 17585
rect 2668 16183 2708 16192
rect 2764 16316 2804 16325
rect 2764 15308 2804 16276
rect 2764 15259 2804 15268
rect 2956 14804 2996 17536
rect 3112 16652 3480 16661
rect 3112 16603 3480 16612
rect 3532 15560 3572 17704
rect 3628 17576 3668 17585
rect 3628 17072 3668 17536
rect 3628 17023 3668 17032
rect 3724 16988 3764 17956
rect 3916 17912 3956 17921
rect 3916 17744 3956 17872
rect 4300 17828 4340 18544
rect 4300 17779 4340 17788
rect 4684 18500 4724 18509
rect 4684 17996 4724 18460
rect 3916 17695 3956 17704
rect 4012 17660 4052 17669
rect 4052 17620 4148 17660
rect 4012 17611 4052 17620
rect 4108 17240 4148 17620
rect 4684 17576 4724 17956
rect 4780 17744 4820 18628
rect 4780 17695 4820 17704
rect 4876 17660 4916 19888
rect 4972 18752 5012 19972
rect 5164 19508 5204 20056
rect 5164 19459 5204 19468
rect 4972 18703 5012 18712
rect 5068 18500 5108 18509
rect 4876 17611 4916 17620
rect 4972 18080 5012 18089
rect 4684 17527 4724 17536
rect 4780 17576 4820 17585
rect 4352 17408 4720 17417
rect 4352 17359 4720 17368
rect 4492 17240 4532 17249
rect 4108 17200 4340 17240
rect 3724 16939 3764 16948
rect 3916 16904 3956 16913
rect 3532 15511 3572 15520
rect 3628 16232 3668 16241
rect 3112 15140 3480 15149
rect 3112 15091 3480 15100
rect 2956 14755 2996 14764
rect 2860 14720 2900 14729
rect 2764 14680 2860 14720
rect 2764 14384 2804 14680
rect 2860 14652 2900 14680
rect 3532 14720 3572 14729
rect 3436 14636 3476 14645
rect 3436 14501 3476 14596
rect 2764 14335 2804 14344
rect 2764 14132 2804 14141
rect 2764 13796 2804 14092
rect 3532 13964 3572 14680
rect 3532 13915 3572 13924
rect 2764 13747 2804 13756
rect 3112 13628 3480 13637
rect 3112 13579 3480 13588
rect 3340 13208 3380 13217
rect 3340 12704 3380 13168
rect 3628 12956 3668 16192
rect 3724 15812 3764 15821
rect 3724 15677 3764 15772
rect 3820 15728 3860 15737
rect 3724 14636 3764 14645
rect 3724 14048 3764 14596
rect 3724 13460 3764 14008
rect 3724 13411 3764 13420
rect 3628 12907 3668 12916
rect 3724 13208 3764 13217
rect 3724 12788 3764 13168
rect 3724 12739 3764 12748
rect 3340 12655 3380 12664
rect 2764 12536 2804 12545
rect 2572 11227 2612 11236
rect 2668 12452 2708 12461
rect 2668 12200 2708 12412
rect 1804 8588 1844 9388
rect 1804 8539 1844 8548
rect 1900 10312 2036 10352
rect 2092 11024 2132 11033
rect 1804 8420 1844 8429
rect 1612 7447 1652 7456
rect 1708 7832 1748 7841
rect 1516 7363 1556 7372
rect 1516 7160 1556 7169
rect 1516 6992 1556 7120
rect 1708 7160 1748 7792
rect 1708 7111 1748 7120
rect 1804 7664 1844 8380
rect 1516 4976 1556 6952
rect 1516 4927 1556 4936
rect 1612 6488 1652 6497
rect 1612 4304 1652 6448
rect 1612 4255 1652 4264
rect 1708 5648 1748 5657
rect 1708 5060 1748 5608
rect 1612 4136 1652 4145
rect 1708 4136 1748 5020
rect 1804 4976 1844 7624
rect 1900 6824 1940 10312
rect 1996 10184 2036 10193
rect 1996 9428 2036 10144
rect 1996 9379 2036 9388
rect 1996 8924 2036 8933
rect 1996 6992 2036 8884
rect 1996 6943 2036 6952
rect 1900 6775 1940 6784
rect 1804 4388 1844 4936
rect 1804 4339 1844 4348
rect 1652 4096 1748 4136
rect 1612 4087 1652 4096
rect 1420 3499 1460 3508
rect 1516 3968 1556 3977
rect 1324 2659 1364 2668
rect 1516 2540 1556 3928
rect 1516 2491 1556 2500
rect 1996 3464 2036 3473
rect 1996 1952 2036 3424
rect 1996 1903 2036 1912
rect 2092 2540 2132 10984
rect 2668 10940 2708 12160
rect 2764 11948 2804 12496
rect 3112 12116 3480 12125
rect 3112 12067 3480 12076
rect 2764 11899 2804 11908
rect 2860 11780 2900 11789
rect 2860 11612 2900 11740
rect 2860 11024 2900 11572
rect 2860 10975 2900 10984
rect 3436 11528 3476 11537
rect 3436 11024 3476 11488
rect 3820 11528 3860 15688
rect 3820 11479 3860 11488
rect 3436 10975 3476 10984
rect 2284 10436 2324 10445
rect 2284 10268 2324 10396
rect 2188 10184 2228 10193
rect 2188 9680 2228 10144
rect 2188 9631 2228 9640
rect 2188 9512 2228 9521
rect 2284 9512 2324 10228
rect 2572 9848 2612 9857
rect 2668 9848 2708 10900
rect 3112 10604 3480 10613
rect 3112 10555 3480 10564
rect 3724 10436 3764 10445
rect 2956 10184 2996 10193
rect 2612 9808 2708 9848
rect 2764 10100 2804 10109
rect 2228 9472 2324 9512
rect 2188 9463 2228 9472
rect 2284 8756 2324 9472
rect 2380 9680 2420 9689
rect 2380 8840 2420 9640
rect 2572 9428 2612 9808
rect 2572 8924 2612 9388
rect 2572 8875 2612 8884
rect 2668 9512 2708 9521
rect 2764 9512 2804 10060
rect 2956 9596 2996 10144
rect 3532 10184 3572 10193
rect 3052 10016 3092 10025
rect 3052 9680 3092 9976
rect 3052 9631 3092 9640
rect 2956 9547 2996 9556
rect 2708 9472 2804 9512
rect 2420 8800 2516 8840
rect 2380 8791 2420 8800
rect 2188 7160 2228 7169
rect 2188 6992 2228 7120
rect 2188 6656 2228 6952
rect 2188 6607 2228 6616
rect 2188 6488 2228 6497
rect 2188 5648 2228 6448
rect 2284 6404 2324 8716
rect 2380 8588 2420 8597
rect 2380 8000 2420 8548
rect 2476 8084 2516 8800
rect 2476 8035 2516 8044
rect 2380 7951 2420 7960
rect 2284 6355 2324 6364
rect 2476 6488 2516 6497
rect 2476 5732 2516 6448
rect 2476 5683 2516 5692
rect 2188 5599 2228 5608
rect 2668 5480 2708 9472
rect 2860 9428 2900 9437
rect 2764 8840 2804 8849
rect 2764 8168 2804 8800
rect 2764 8119 2804 8128
rect 2764 7748 2804 7757
rect 2764 7244 2804 7708
rect 2764 7195 2804 7204
rect 2860 7160 2900 9388
rect 3112 9092 3480 9101
rect 3112 9043 3480 9052
rect 3532 8168 3572 10144
rect 3532 8119 3572 8128
rect 3628 9764 3668 9773
rect 3628 9260 3668 9724
rect 3052 8000 3092 8009
rect 2956 7960 3052 8000
rect 2956 7412 2996 7960
rect 3052 7951 3092 7960
rect 3532 7832 3572 7841
rect 3112 7580 3480 7589
rect 3112 7531 3480 7540
rect 2956 7363 2996 7372
rect 2860 6992 2900 7120
rect 3532 7160 3572 7792
rect 3532 7111 3572 7120
rect 2860 6943 2900 6952
rect 2764 6740 2804 6749
rect 2764 6404 2804 6700
rect 2764 6355 2804 6364
rect 3532 6740 3572 6749
rect 3532 6404 3572 6700
rect 3628 6572 3668 9220
rect 3724 8084 3764 10396
rect 3916 10352 3956 16864
rect 4012 16232 4052 16241
rect 4012 11444 4052 16192
rect 4300 16148 4340 17200
rect 4492 17072 4532 17200
rect 4492 17023 4532 17032
rect 4780 16988 4820 17536
rect 4972 17324 5012 18040
rect 5068 17996 5108 18460
rect 5164 18080 5204 18175
rect 5164 18031 5204 18040
rect 5068 17947 5108 17956
rect 5164 17828 5204 17837
rect 4972 17275 5012 17284
rect 5068 17660 5108 17669
rect 4780 16939 4820 16948
rect 4972 17156 5012 17165
rect 4876 16232 4916 16241
rect 4300 16099 4340 16108
rect 4684 16064 4724 16159
rect 4684 16015 4724 16024
rect 4352 15896 4720 15905
rect 4352 15847 4720 15856
rect 4492 15728 4532 15737
rect 4492 15560 4532 15688
rect 4108 15476 4148 15485
rect 4108 14972 4148 15436
rect 4300 14972 4340 14981
rect 4108 14804 4148 14932
rect 4108 14755 4148 14764
rect 4204 14932 4300 14972
rect 4108 14468 4148 14477
rect 4108 14333 4148 14428
rect 4108 14216 4148 14225
rect 4108 12536 4148 14176
rect 4204 12704 4244 14932
rect 4300 14923 4340 14932
rect 4492 14636 4532 15520
rect 4492 14587 4532 14596
rect 4352 14384 4720 14393
rect 4352 14335 4720 14344
rect 4876 13544 4916 16192
rect 4876 13495 4916 13504
rect 4780 13292 4820 13301
rect 4352 12872 4720 12881
rect 4352 12823 4720 12832
rect 4204 12655 4244 12664
rect 4492 12620 4532 12629
rect 4108 12496 4244 12536
rect 4012 11395 4052 11404
rect 4108 11696 4148 11705
rect 3820 10312 3956 10352
rect 3820 8252 3860 10312
rect 3916 10184 3956 10193
rect 3916 8924 3956 10144
rect 3916 8672 3956 8884
rect 3916 8623 3956 8632
rect 3820 8203 3860 8212
rect 4108 8168 4148 11656
rect 4204 11192 4244 12496
rect 4492 11948 4532 12580
rect 4492 11899 4532 11908
rect 4352 11360 4720 11369
rect 4352 11311 4720 11320
rect 4204 11057 4244 11152
rect 4780 11192 4820 13252
rect 4876 13292 4916 13301
rect 4876 13208 4916 13252
rect 4876 13157 4916 13168
rect 4972 12620 5012 17116
rect 5068 16988 5108 17620
rect 5164 17240 5204 17788
rect 5260 17828 5300 17837
rect 5260 17744 5300 17788
rect 5260 17693 5300 17704
rect 5164 17191 5204 17200
rect 5068 16400 5108 16948
rect 5068 16351 5108 16360
rect 5356 15140 5396 20980
rect 5740 20852 5780 20861
rect 5452 20768 5492 20777
rect 5452 20684 5492 20728
rect 5452 20633 5492 20644
rect 5548 20600 5588 20609
rect 5548 20012 5588 20560
rect 5740 20096 5780 20812
rect 5740 20047 5780 20056
rect 5548 19963 5588 19972
rect 5836 19928 5876 19937
rect 5836 19340 5876 19888
rect 5836 19291 5876 19300
rect 5740 19256 5780 19265
rect 5548 19172 5588 19181
rect 5548 18668 5588 19132
rect 5740 18752 5780 19216
rect 5740 18703 5780 18712
rect 5644 18668 5684 18677
rect 5548 18628 5644 18668
rect 5644 18533 5684 18628
rect 5932 18668 5972 23080
rect 6220 23120 6260 24592
rect 6892 25472 6932 25481
rect 6892 24548 6932 25432
rect 6988 25136 7028 28600
rect 7468 27404 7508 27413
rect 7468 26816 7508 27364
rect 7468 26767 7508 26776
rect 7756 26648 7796 28600
rect 8524 27908 8564 28600
rect 9292 27908 9332 28600
rect 10060 28244 10100 28600
rect 10060 28195 10100 28204
rect 8524 27868 8660 27908
rect 8524 27740 8564 27749
rect 7756 26599 7796 26608
rect 8236 27572 8276 27581
rect 8236 26312 8276 27532
rect 8524 26900 8564 27700
rect 8524 26851 8564 26860
rect 8620 26648 8660 27868
rect 9292 27859 9332 27868
rect 9292 27572 9332 27581
rect 8620 26599 8660 26608
rect 8716 27152 8756 27161
rect 8236 26263 8276 26272
rect 8332 26312 8372 26321
rect 8332 26144 8372 26272
rect 8716 26312 8756 27112
rect 9292 26984 9332 27532
rect 9292 26935 9332 26944
rect 9676 27404 9716 27413
rect 9196 26732 9236 26741
rect 8716 26263 8756 26272
rect 8908 26312 8948 26321
rect 8332 26095 8372 26104
rect 8908 26060 8948 26272
rect 6988 25087 7028 25096
rect 8140 25892 8180 25901
rect 8140 25136 8180 25852
rect 8140 25087 8180 25096
rect 8332 25724 8372 25733
rect 8332 24716 8372 25684
rect 8908 25388 8948 26020
rect 9100 26228 9140 26237
rect 9004 25976 9044 26004
rect 9100 25976 9140 26188
rect 9196 26144 9236 26692
rect 9676 26312 9716 27364
rect 10348 27404 10388 27413
rect 10252 26732 10292 26741
rect 9676 26263 9716 26272
rect 10060 26312 10100 26321
rect 10156 26312 10196 26321
rect 10100 26272 10156 26312
rect 10060 26244 10100 26272
rect 10156 26263 10196 26272
rect 9196 26095 9236 26104
rect 9964 26144 10004 26239
rect 9964 26095 10004 26104
rect 10156 26144 10196 26153
rect 9044 25936 9140 25976
rect 9004 25927 9044 25936
rect 9100 25556 9140 25936
rect 6892 24499 6932 24508
rect 8236 24548 8276 24557
rect 6220 23071 6260 23080
rect 7084 23960 7124 23969
rect 7084 23036 7124 23920
rect 7468 23792 7508 23801
rect 7084 22987 7124 22996
rect 7372 23120 7412 23129
rect 6028 22448 6068 22457
rect 6028 22280 6068 22408
rect 6028 22231 6068 22240
rect 6508 22448 6548 22457
rect 6412 22028 6452 22037
rect 6316 20684 6356 20693
rect 6124 19928 6164 19937
rect 5932 18619 5972 18628
rect 6028 19172 6068 19181
rect 6028 18500 6068 19132
rect 5740 17744 5780 17753
rect 5548 17072 5588 17081
rect 5452 16232 5492 16241
rect 5452 16097 5492 16192
rect 5452 15560 5492 15571
rect 5452 15476 5492 15520
rect 5452 15427 5492 15436
rect 5356 15091 5396 15100
rect 5452 15224 5492 15233
rect 5452 14636 5492 15184
rect 5452 14587 5492 14596
rect 4972 12571 5012 12580
rect 5068 14384 5108 14393
rect 4972 11780 5012 11789
rect 4780 11143 4820 11152
rect 4876 11696 4916 11705
rect 4300 11108 4340 11117
rect 4300 10973 4340 11068
rect 4876 11108 4916 11656
rect 4876 11059 4916 11068
rect 4396 11024 4436 11033
rect 4396 10889 4436 10984
rect 4492 10940 4532 10949
rect 4588 10940 4628 10968
rect 4532 10900 4588 10940
rect 4108 8119 4148 8128
rect 4204 10772 4244 10781
rect 3724 8044 3860 8084
rect 3628 6523 3668 6532
rect 2668 5431 2708 5440
rect 2860 6320 2900 6329
rect 2860 5648 2900 6280
rect 3112 6068 3480 6077
rect 3112 6019 3480 6028
rect 3532 5732 3572 6364
rect 3532 5683 3572 5692
rect 2380 4976 2420 4985
rect 2188 4136 2228 4145
rect 2188 3716 2228 4096
rect 2380 4136 2420 4936
rect 2380 4087 2420 4096
rect 2188 3667 2228 3676
rect 2860 4052 2900 5608
rect 3724 5648 3764 5657
rect 3724 5480 3764 5608
rect 3532 5144 3572 5153
rect 3532 4976 3572 5104
rect 3112 4556 3480 4565
rect 3112 4507 3480 4516
rect 3532 4388 3572 4936
rect 3628 4892 3668 4901
rect 3724 4892 3764 5440
rect 3668 4852 3764 4892
rect 3628 4843 3668 4852
rect 3820 4808 3860 8044
rect 4204 7580 4244 10732
rect 4492 10268 4532 10900
rect 4588 10891 4628 10900
rect 4492 10219 4532 10228
rect 4684 10856 4724 10865
rect 4684 10268 4724 10816
rect 4588 10184 4628 10195
rect 4588 10100 4628 10144
rect 4684 10133 4724 10228
rect 4876 10856 4916 10865
rect 4876 10184 4916 10816
rect 4972 10436 5012 11740
rect 4972 10387 5012 10396
rect 4972 10184 5012 10279
rect 4876 10144 4972 10184
rect 4972 10135 5012 10144
rect 4588 10051 4628 10060
rect 5068 10016 5108 14344
rect 5452 14300 5492 14311
rect 5452 14216 5492 14260
rect 5452 14167 5492 14176
rect 5452 13964 5492 13973
rect 5164 13796 5204 13805
rect 5164 13124 5204 13756
rect 5164 13075 5204 13084
rect 5260 13292 5300 13301
rect 5164 12116 5204 12125
rect 5164 11024 5204 12076
rect 5260 11696 5300 13252
rect 5260 11647 5300 11656
rect 5356 12788 5396 12797
rect 5164 10975 5204 10984
rect 5260 11528 5300 11537
rect 5260 11024 5300 11488
rect 5260 10975 5300 10984
rect 5356 10184 5396 12748
rect 5452 11360 5492 13924
rect 5548 13376 5588 17032
rect 5740 16064 5780 17704
rect 6028 17744 6068 18460
rect 6028 17695 6068 17704
rect 5740 16015 5780 16024
rect 5836 16148 5876 16157
rect 5836 15728 5876 16108
rect 5836 15679 5876 15688
rect 5740 15560 5780 15569
rect 5740 15224 5780 15520
rect 5740 14972 5780 15184
rect 5740 14923 5780 14932
rect 6028 15476 6068 15485
rect 6028 15392 6068 15436
rect 5740 14720 5780 14729
rect 5644 14216 5684 14225
rect 5644 14081 5684 14176
rect 5548 13327 5588 13336
rect 5740 13460 5780 14680
rect 5932 14636 5972 14645
rect 5836 14552 5876 14561
rect 5836 14132 5876 14512
rect 5932 14468 5972 14596
rect 5932 14419 5972 14428
rect 6028 14216 6068 15352
rect 6124 15056 6164 19888
rect 6316 19340 6356 20644
rect 6412 19844 6452 21988
rect 6508 21524 6548 22408
rect 6508 21475 6548 21484
rect 7276 21356 7316 21365
rect 7180 21316 7276 21356
rect 7180 20852 7220 21316
rect 7276 21307 7316 21316
rect 7084 20812 7180 20852
rect 6700 20180 6740 20189
rect 6700 20096 6740 20140
rect 6700 20045 6740 20056
rect 6988 20096 7028 20105
rect 6412 19795 6452 19804
rect 6796 20012 6836 20021
rect 6316 19291 6356 19300
rect 6604 19256 6644 19265
rect 6604 18668 6644 19216
rect 6604 18584 6644 18628
rect 6604 18533 6644 18544
rect 6700 19088 6740 19097
rect 6220 18500 6260 18509
rect 6220 17240 6260 18460
rect 6508 18500 6548 18509
rect 6220 17191 6260 17200
rect 6316 18332 6356 18341
rect 6316 16064 6356 18292
rect 6508 17744 6548 18460
rect 6508 17695 6548 17704
rect 6700 17660 6740 19048
rect 6796 18248 6836 19972
rect 6988 19844 7028 20056
rect 6988 19424 7028 19804
rect 6988 19375 7028 19384
rect 6892 19004 6932 19013
rect 6892 18752 6932 18964
rect 6892 18703 6932 18712
rect 6796 18199 6836 18208
rect 6892 18584 6932 18593
rect 6892 18500 6932 18544
rect 6796 17996 6836 18005
rect 6796 17828 6836 17956
rect 6796 17779 6836 17788
rect 6892 17828 6932 18460
rect 6892 17779 6932 17788
rect 6700 17611 6740 17620
rect 6700 16988 6740 16997
rect 6700 16484 6740 16948
rect 6700 16435 6740 16444
rect 6796 16316 6836 16325
rect 6796 16232 6836 16276
rect 6796 16181 6836 16192
rect 6892 16316 6932 16325
rect 6316 16015 6356 16024
rect 6508 16148 6548 16157
rect 6124 15007 6164 15016
rect 6220 15560 6260 15569
rect 6028 14167 6068 14176
rect 6124 14636 6164 14645
rect 5836 14083 5876 14092
rect 5644 13292 5684 13301
rect 5548 13208 5588 13219
rect 5548 13124 5588 13168
rect 5644 13157 5684 13252
rect 5548 13075 5588 13084
rect 5644 12452 5684 12461
rect 5548 11360 5588 11369
rect 5452 11320 5548 11360
rect 5548 11024 5588 11320
rect 5548 10975 5588 10984
rect 5356 10135 5396 10144
rect 5548 10184 5588 10193
rect 5068 9967 5108 9976
rect 4352 9848 4720 9857
rect 4352 9799 4720 9808
rect 4300 9680 4340 9689
rect 4300 8672 4340 9640
rect 5548 9680 5588 10144
rect 5548 9631 5588 9640
rect 5644 9596 5684 12412
rect 5740 11864 5780 13420
rect 5932 14048 5972 14057
rect 5836 13376 5876 13385
rect 5836 12536 5876 13336
rect 5836 12487 5876 12496
rect 5740 11815 5780 11824
rect 5836 11780 5876 11789
rect 5836 11645 5876 11740
rect 5740 11528 5780 11537
rect 5740 10940 5780 11488
rect 5740 10891 5780 10900
rect 5644 9512 5684 9556
rect 5644 9461 5684 9472
rect 5836 10016 5876 10025
rect 5836 9428 5876 9976
rect 5932 9680 5972 14008
rect 6028 13964 6068 13973
rect 6028 13124 6068 13924
rect 6124 13628 6164 14596
rect 6220 14636 6260 15520
rect 6508 15476 6548 16108
rect 6220 14587 6260 14596
rect 6412 14636 6452 14645
rect 6124 13579 6164 13588
rect 6316 13964 6356 13973
rect 6124 13376 6164 13471
rect 6124 13327 6164 13336
rect 6220 13460 6260 13469
rect 6028 12704 6068 13084
rect 6028 12655 6068 12664
rect 6124 13208 6164 13217
rect 6220 13206 6260 13420
rect 6164 13168 6260 13206
rect 6124 13166 6260 13168
rect 5932 9631 5972 9640
rect 6028 11780 6068 11789
rect 5836 9379 5876 9388
rect 5932 9512 5972 9521
rect 5260 9344 5300 9353
rect 4300 8623 4340 8632
rect 5164 8756 5204 8765
rect 4352 8336 4720 8345
rect 4352 8287 4720 8296
rect 5164 8168 5204 8716
rect 5164 8119 5204 8128
rect 4012 7540 4244 7580
rect 4012 7076 4052 7540
rect 4108 7412 4148 7421
rect 4108 7160 4148 7372
rect 4108 7111 4148 7120
rect 4492 7244 4532 7253
rect 4012 7027 4052 7036
rect 4108 6992 4148 7001
rect 3532 4339 3572 4348
rect 3724 4768 3860 4808
rect 3916 6404 3956 6413
rect 2476 3380 2516 3389
rect 2476 2792 2516 3340
rect 2476 2743 2516 2752
rect 2092 2120 2132 2500
rect 2860 2540 2900 4012
rect 3532 3212 3572 3221
rect 3112 3044 3480 3053
rect 3112 2995 3480 3004
rect 3532 2624 3572 3172
rect 3724 2900 3764 4768
rect 3916 4640 3956 6364
rect 4108 5144 4148 6952
rect 4492 6992 4532 7204
rect 4492 6943 4532 6952
rect 4780 7244 4820 7253
rect 4780 6992 4820 7204
rect 4780 6943 4820 6952
rect 4972 7160 5012 7169
rect 4352 6824 4720 6833
rect 4352 6775 4720 6784
rect 4972 6740 5012 7120
rect 4972 6691 5012 6700
rect 4204 6488 4244 6497
rect 4204 5732 4244 6448
rect 4396 6488 4436 6497
rect 4204 5683 4244 5692
rect 4300 6236 4340 6245
rect 4300 5648 4340 6196
rect 4396 5900 4436 6448
rect 4396 5851 4436 5860
rect 4300 5599 4340 5608
rect 4684 5816 4724 5825
rect 4684 5564 4724 5776
rect 4684 5515 4724 5524
rect 4876 5648 4916 5657
rect 4876 5480 4916 5608
rect 4352 5312 4720 5321
rect 4352 5263 4720 5272
rect 4108 5095 4148 5104
rect 4876 4640 4916 5440
rect 3628 2860 3764 2900
rect 3820 4600 3956 4640
rect 4780 4600 4916 4640
rect 3820 3548 3860 4600
rect 3628 2708 3668 2860
rect 3628 2659 3668 2668
rect 3532 2575 3572 2584
rect 2860 2491 2900 2500
rect 2092 1616 2132 2080
rect 2092 1567 2132 1576
rect 2668 1868 2708 1877
rect 2668 1280 2708 1828
rect 3820 1868 3860 3508
rect 3916 4052 3956 4061
rect 3916 3716 3956 4012
rect 4352 3800 4720 3809
rect 4352 3751 4720 3760
rect 3916 2876 3956 3676
rect 4684 3464 4724 3473
rect 4684 3296 4724 3424
rect 4684 3247 4724 3256
rect 3916 2827 3956 2836
rect 4588 2792 4628 2801
rect 4588 2624 4628 2752
rect 4588 2575 4628 2584
rect 4780 2540 4820 4600
rect 4972 4136 5012 4145
rect 4352 2288 4720 2297
rect 4352 2239 4720 2248
rect 3112 1532 3480 1541
rect 3112 1483 3480 1492
rect 2668 1231 2708 1240
rect 3820 1112 3860 1828
rect 3820 1063 3860 1072
rect 4396 1952 4436 1961
rect 4396 1112 4436 1912
rect 4780 1952 4820 2500
rect 4780 1700 4820 1912
rect 4780 1651 4820 1660
rect 4876 3968 4916 3977
rect 4876 3464 4916 3928
rect 4876 2792 4916 3424
rect 4972 3296 5012 4096
rect 5260 4136 5300 9304
rect 5932 9260 5972 9472
rect 5932 9211 5972 9220
rect 6028 9176 6068 11740
rect 6124 11024 6164 13166
rect 6316 12452 6356 13924
rect 6412 13880 6452 14596
rect 6412 13831 6452 13840
rect 6412 13292 6452 13303
rect 6412 13208 6452 13252
rect 6412 13159 6452 13168
rect 6508 13040 6548 15436
rect 6700 16148 6740 16157
rect 6508 12991 6548 13000
rect 6604 13460 6644 13469
rect 6604 12956 6644 13420
rect 6700 13376 6740 16108
rect 6892 15896 6932 16276
rect 6892 15847 6932 15856
rect 6988 16316 7028 16325
rect 6796 15560 6836 15569
rect 6796 15392 6836 15520
rect 6796 15343 6836 15352
rect 6892 15476 6932 15485
rect 6700 13327 6740 13336
rect 6796 14720 6836 14729
rect 6604 12907 6644 12916
rect 6700 13208 6740 13217
rect 6700 12704 6740 13168
rect 6700 12655 6740 12664
rect 6316 12403 6356 12412
rect 6700 11780 6740 11875
rect 6700 11731 6740 11740
rect 6604 11444 6644 11453
rect 6316 11360 6356 11369
rect 6124 10975 6164 10984
rect 6220 11108 6260 11117
rect 6220 10268 6260 11068
rect 6220 10219 6260 10228
rect 6316 10940 6356 11320
rect 6508 11276 6548 11285
rect 6508 11141 6548 11236
rect 6604 11024 6644 11404
rect 6796 11360 6836 14680
rect 6892 14636 6932 15436
rect 6892 14587 6932 14596
rect 6892 14384 6932 14393
rect 6892 13964 6932 14344
rect 6892 13915 6932 13924
rect 6892 13292 6932 13301
rect 6892 13157 6932 13252
rect 6988 12788 7028 16276
rect 7084 15980 7124 20812
rect 7180 20803 7220 20812
rect 7276 20768 7316 20777
rect 7276 20096 7316 20728
rect 7276 20047 7316 20056
rect 7372 20012 7412 23080
rect 7468 23036 7508 23752
rect 8044 23624 8084 23633
rect 7468 22987 7508 22996
rect 7852 23288 7892 23297
rect 7852 22952 7892 23248
rect 8044 23120 8084 23584
rect 8044 23071 8084 23080
rect 7852 22903 7892 22912
rect 7660 22532 7700 22541
rect 7372 19963 7412 19972
rect 7564 20012 7604 20021
rect 7180 19928 7220 19937
rect 7180 18584 7220 19888
rect 7276 19508 7316 19517
rect 7276 19004 7316 19468
rect 7564 19088 7604 19972
rect 7660 19424 7700 22492
rect 8044 22280 8084 22289
rect 7948 21356 7988 21365
rect 7852 20852 7892 20861
rect 7756 20096 7796 20105
rect 7756 19961 7796 20056
rect 7660 19375 7700 19384
rect 7756 19508 7796 19517
rect 7564 19039 7604 19048
rect 7276 18955 7316 18964
rect 7660 18668 7700 18677
rect 7564 18584 7604 18593
rect 7180 18535 7220 18544
rect 7468 18544 7564 18584
rect 7372 18500 7412 18509
rect 7276 17660 7316 17669
rect 7276 16400 7316 17620
rect 7372 16484 7412 18460
rect 7372 16435 7412 16444
rect 7084 15931 7124 15940
rect 7180 16232 7220 16241
rect 7180 15728 7220 16192
rect 7276 16148 7316 16360
rect 7276 16099 7316 16108
rect 7180 15679 7220 15688
rect 7276 15560 7316 15569
rect 7276 15425 7316 15520
rect 7180 15392 7220 15401
rect 7084 15308 7124 15317
rect 7084 14972 7124 15268
rect 7084 14923 7124 14932
rect 7180 15308 7220 15352
rect 7372 15308 7412 15317
rect 7180 15268 7372 15308
rect 7084 14720 7124 14731
rect 7084 14636 7124 14680
rect 7084 14587 7124 14596
rect 6796 11311 6836 11320
rect 6892 12748 7028 12788
rect 7084 13208 7124 13217
rect 6604 10984 6836 11024
rect 6316 10016 6356 10900
rect 6604 10772 6644 10781
rect 6604 10352 6644 10732
rect 6796 10688 6836 10984
rect 6796 10639 6836 10648
rect 6604 10303 6644 10312
rect 6796 10352 6836 10361
rect 6508 10268 6548 10277
rect 6508 10100 6548 10228
rect 6796 10184 6836 10312
rect 6796 10135 6836 10144
rect 6892 10184 6932 12748
rect 7084 12452 7124 13168
rect 7180 13040 7220 15268
rect 7372 15259 7412 15268
rect 7468 14300 7508 18544
rect 7564 18535 7604 18544
rect 7660 18332 7700 18628
rect 7756 18416 7796 19468
rect 7852 19256 7892 20812
rect 7852 19207 7892 19216
rect 7948 19088 7988 21316
rect 8044 20768 8084 22240
rect 8044 20719 8084 20728
rect 8140 20600 8180 20609
rect 8140 20012 8180 20560
rect 7756 18367 7796 18376
rect 7852 19048 7988 19088
rect 8044 19928 8084 19937
rect 7660 17744 7700 18292
rect 7660 17695 7700 17704
rect 7564 16232 7604 16241
rect 7564 16148 7604 16192
rect 7564 16097 7604 16108
rect 7756 15980 7796 15989
rect 7564 15896 7604 15905
rect 7564 15392 7604 15856
rect 7564 15343 7604 15352
rect 7756 15056 7796 15940
rect 7756 14804 7796 15016
rect 7756 14755 7796 14764
rect 7660 14636 7700 14645
rect 7468 14251 7508 14260
rect 7564 14384 7604 14393
rect 7180 12991 7220 13000
rect 7276 14216 7316 14225
rect 7124 12412 7220 12452
rect 7084 12403 7124 12412
rect 6988 12200 7028 12209
rect 6988 11864 7028 12160
rect 6988 11815 7028 11824
rect 7084 11696 7124 11705
rect 6988 11612 7028 11621
rect 6988 11192 7028 11572
rect 7084 11561 7124 11656
rect 6988 11143 7028 11152
rect 7180 11192 7220 12412
rect 7276 12368 7316 14176
rect 7468 13460 7508 13469
rect 7468 13208 7508 13420
rect 7372 12956 7412 12965
rect 7372 12620 7412 12916
rect 7372 12571 7412 12580
rect 7468 12452 7508 13168
rect 7564 13460 7604 14344
rect 7564 13292 7604 13420
rect 7564 13208 7604 13252
rect 7564 13159 7604 13168
rect 7276 12319 7316 12328
rect 7372 12412 7508 12452
rect 7564 13040 7604 13049
rect 7564 12452 7604 13000
rect 7372 12032 7412 12412
rect 7564 12403 7604 12412
rect 7660 12536 7700 14596
rect 7852 14468 7892 19048
rect 7948 16232 7988 16241
rect 7948 15476 7988 16192
rect 8044 15812 8084 19888
rect 8140 19340 8180 19972
rect 8140 19291 8180 19300
rect 8140 18752 8180 18761
rect 8140 18584 8180 18712
rect 8140 18535 8180 18544
rect 8236 17156 8276 24508
rect 8332 23624 8372 24676
rect 8524 25136 8564 25145
rect 8524 24548 8564 25096
rect 8908 24716 8948 25348
rect 8908 24667 8948 24676
rect 9004 25516 9100 25556
rect 9004 25304 9044 25516
rect 9100 25507 9140 25516
rect 9292 26060 9332 26069
rect 8716 24632 8756 24641
rect 8524 24499 8564 24508
rect 8620 24592 8716 24632
rect 8332 23575 8372 23584
rect 8620 24212 8660 24592
rect 8716 24583 8756 24592
rect 9004 24632 9044 25264
rect 9292 25304 9332 26020
rect 10060 25976 10100 25985
rect 9868 25892 9908 25901
rect 9868 25724 9908 25852
rect 10060 25841 10100 25936
rect 9868 25675 9908 25684
rect 10156 25556 10196 26104
rect 10156 25507 10196 25516
rect 9292 24800 9332 25264
rect 9964 25388 10004 25397
rect 9676 25052 9716 25061
rect 9292 24760 9620 24800
rect 8620 23708 8660 24172
rect 9004 23876 9044 24592
rect 9580 24632 9620 24760
rect 9580 24583 9620 24592
rect 9004 23827 9044 23836
rect 9100 23960 9140 23969
rect 8332 22868 8372 22877
rect 8332 22280 8372 22828
rect 8620 22364 8660 23668
rect 8620 22315 8660 22324
rect 8716 23624 8756 23633
rect 8332 22231 8372 22240
rect 8716 22280 8756 23584
rect 8908 23204 8948 23213
rect 8716 22231 8756 22240
rect 8812 23120 8852 23129
rect 8812 21608 8852 23080
rect 8908 22196 8948 23164
rect 9100 23036 9140 23920
rect 9292 23960 9332 23969
rect 9292 23792 9332 23920
rect 9292 23743 9332 23752
rect 9100 22987 9140 22996
rect 9676 22448 9716 25012
rect 9868 24968 9908 24977
rect 9772 24548 9812 24559
rect 9772 24464 9812 24508
rect 9772 24415 9812 24424
rect 9676 22399 9716 22408
rect 8908 22147 8948 22156
rect 8236 17107 8276 17116
rect 8332 21356 8372 21365
rect 8044 15763 8084 15772
rect 8236 16988 8276 16997
rect 8236 16568 8276 16948
rect 7948 14972 7988 15436
rect 8044 15644 8084 15653
rect 8044 15392 8084 15604
rect 8044 15257 8084 15352
rect 8236 15308 8276 16528
rect 8236 15259 8276 15268
rect 7948 14923 7988 14932
rect 8236 14888 8276 14897
rect 7852 14419 7892 14428
rect 8140 14804 8180 14813
rect 7372 11983 7412 11992
rect 7468 12284 7508 12293
rect 7372 11864 7412 11873
rect 7180 11143 7220 11152
rect 7276 11696 7316 11705
rect 7276 11528 7316 11656
rect 7276 10940 7316 11488
rect 7372 11024 7412 11824
rect 7372 10975 7412 10984
rect 7276 10436 7316 10900
rect 7276 10387 7316 10396
rect 7180 10352 7220 10361
rect 6548 10060 6644 10100
rect 6508 10051 6548 10060
rect 6316 9967 6356 9976
rect 6604 10016 6644 10060
rect 6604 9967 6644 9976
rect 6700 9932 6740 9941
rect 6618 9596 6658 9605
rect 6700 9596 6740 9892
rect 6892 9932 6932 10144
rect 6988 10268 7028 10277
rect 7084 10268 7124 10296
rect 7028 10228 7084 10268
rect 6988 10016 7028 10228
rect 7084 10219 7124 10228
rect 6988 9967 7028 9976
rect 6892 9883 6932 9892
rect 6658 9556 6740 9596
rect 6618 9547 6658 9556
rect 6028 8672 6068 9136
rect 6028 8623 6068 8632
rect 6220 9428 6260 9437
rect 5740 8588 5780 8597
rect 5548 8000 5588 8009
rect 5740 8000 5780 8548
rect 5588 7960 5780 8000
rect 5548 7951 5588 7960
rect 5740 5816 5780 7960
rect 6220 6656 6260 9388
rect 7084 9428 7124 9437
rect 7180 9428 7220 10312
rect 7372 10268 7412 10277
rect 7372 10100 7412 10228
rect 7124 9388 7220 9428
rect 7276 10060 7412 10100
rect 7084 9379 7124 9388
rect 7084 8672 7124 8681
rect 6988 8588 7028 8597
rect 6988 8168 7028 8548
rect 6988 8119 7028 8128
rect 6892 8084 6932 8093
rect 6700 8000 6740 8009
rect 6700 7160 6740 7960
rect 6700 7111 6740 7120
rect 6892 7160 6932 8044
rect 7084 8000 7124 8632
rect 7276 8504 7316 10060
rect 7372 9848 7412 9857
rect 7372 9512 7412 9808
rect 7468 9680 7508 12244
rect 7564 12032 7604 12041
rect 7564 11696 7604 11992
rect 7660 11780 7700 12496
rect 7660 11731 7700 11740
rect 7756 14048 7796 14057
rect 7564 11647 7604 11656
rect 7660 11024 7700 11033
rect 7660 10856 7700 10984
rect 7660 10807 7700 10816
rect 7564 10604 7604 10613
rect 7564 10100 7604 10564
rect 7756 10268 7796 14008
rect 7852 13880 7892 13889
rect 7852 13376 7892 13840
rect 8140 13880 8180 14764
rect 8140 13831 8180 13840
rect 7852 10940 7892 13336
rect 7948 13544 7988 13553
rect 7948 13292 7988 13504
rect 7948 13243 7988 13252
rect 8044 13544 8084 13553
rect 7948 13124 7988 13133
rect 7948 12788 7988 13084
rect 7948 12739 7988 12748
rect 7852 10891 7892 10900
rect 7948 12368 7988 12377
rect 7948 10352 7988 12328
rect 8044 11192 8084 13504
rect 8140 13208 8180 13217
rect 8140 12620 8180 13168
rect 8140 12571 8180 12580
rect 8236 12536 8276 14848
rect 8332 14720 8372 21316
rect 8524 20180 8564 20189
rect 8812 20180 8852 21568
rect 9292 22112 9332 22121
rect 9004 21440 9044 21449
rect 9004 21188 9044 21400
rect 9004 20852 9044 21148
rect 9292 20852 9332 22072
rect 9388 21608 9428 21617
rect 9388 21356 9428 21568
rect 9388 21307 9428 21316
rect 9676 21356 9716 21365
rect 9292 20812 9428 20852
rect 9004 20803 9044 20812
rect 8428 19928 8468 19937
rect 8428 17744 8468 19888
rect 8428 17408 8468 17704
rect 8428 17359 8468 17368
rect 8524 16484 8564 20140
rect 8524 16435 8564 16444
rect 8620 20140 8852 20180
rect 9004 20432 9044 20441
rect 8332 13964 8372 14680
rect 8428 16232 8468 16241
rect 8428 14048 8468 16192
rect 8524 16064 8564 16073
rect 8620 16064 8660 20140
rect 9004 20096 9044 20392
rect 9004 20047 9044 20056
rect 8716 20012 8756 20021
rect 8716 19172 8756 19972
rect 8716 19123 8756 19132
rect 8908 19340 8948 19349
rect 8812 19088 8852 19097
rect 8812 18668 8852 19048
rect 8908 18752 8948 19300
rect 9292 19256 9332 19265
rect 9004 19172 9044 19181
rect 9004 18920 9044 19132
rect 9004 18871 9044 18880
rect 9292 19172 9332 19216
rect 8908 18703 8948 18712
rect 9292 18752 9332 19132
rect 9292 18703 9332 18712
rect 8812 18619 8852 18628
rect 9004 18668 9044 18677
rect 8812 18500 8852 18509
rect 8812 17912 8852 18460
rect 9004 17996 9044 18628
rect 9004 17947 9044 17956
rect 9100 18500 9140 18509
rect 8564 16024 8660 16064
rect 8716 17660 8756 17669
rect 8524 15929 8564 16024
rect 8524 14804 8564 14813
rect 8524 14468 8564 14764
rect 8524 14419 8564 14428
rect 8428 14008 8564 14048
rect 8332 13915 8372 13924
rect 8524 13292 8564 14008
rect 8716 13376 8756 17620
rect 8812 16736 8852 17872
rect 8908 17492 8948 17501
rect 8908 17072 8948 17452
rect 9100 17240 9140 18460
rect 9100 17191 9140 17200
rect 9292 17576 9332 17585
rect 8908 17023 8948 17032
rect 9196 17156 9236 17165
rect 9004 16988 9044 16997
rect 8908 16904 8948 16913
rect 8908 16769 8948 16864
rect 8812 16232 8852 16696
rect 9004 16484 9044 16948
rect 9004 16435 9044 16444
rect 9196 16400 9236 17116
rect 8812 16183 8852 16192
rect 9004 16316 9044 16325
rect 8716 13327 8756 13336
rect 8812 16064 8852 16073
rect 8332 13208 8372 13217
rect 8332 13073 8372 13168
rect 8428 12956 8468 12965
rect 8332 12536 8372 12631
rect 8236 12496 8332 12536
rect 8044 11143 8084 11152
rect 8140 12284 8180 12293
rect 8140 11024 8180 12244
rect 8236 12032 8276 12496
rect 8332 12487 8372 12496
rect 8332 12368 8372 12377
rect 8332 12284 8372 12328
rect 8332 12233 8372 12244
rect 8236 11983 8276 11992
rect 8225 11864 8265 11873
rect 8265 11824 8276 11864
rect 8225 11815 8276 11824
rect 8236 11696 8276 11815
rect 8236 11647 8276 11656
rect 8140 10975 8180 10984
rect 8236 11444 8276 11453
rect 8236 10940 8276 11404
rect 7948 10303 7988 10312
rect 8140 10520 8180 10529
rect 7756 10219 7796 10228
rect 7564 9764 7604 10060
rect 7564 9715 7604 9724
rect 7852 10184 7892 10193
rect 8140 10184 8180 10480
rect 8236 10268 8276 10900
rect 8332 11360 8372 11369
rect 8332 11024 8372 11320
rect 8332 10889 8372 10984
rect 8428 11192 8468 12916
rect 8524 12704 8564 13252
rect 8524 12655 8564 12664
rect 8620 13040 8660 13049
rect 8524 12536 8564 12547
rect 8524 12452 8564 12496
rect 8524 11612 8564 12412
rect 8620 12452 8660 13000
rect 8620 12403 8660 12412
rect 8716 12956 8756 12965
rect 8524 11563 8564 11572
rect 8716 12284 8756 12916
rect 8620 11528 8660 11537
rect 8620 11393 8660 11488
rect 8716 11360 8756 12244
rect 8716 11311 8756 11320
rect 8236 10219 8276 10228
rect 7468 9631 7508 9640
rect 7852 9680 7892 10144
rect 7948 10144 8180 10184
rect 7948 10016 7988 10144
rect 7948 9967 7988 9976
rect 8044 9932 8084 9941
rect 8044 9764 8084 9892
rect 8044 9715 8084 9724
rect 7852 9631 7892 9640
rect 7372 9463 7412 9472
rect 7948 9596 7988 9605
rect 7948 9512 7988 9556
rect 7948 9461 7988 9472
rect 8140 9512 8180 10144
rect 8428 10016 8468 11152
rect 8716 11192 8756 11201
rect 8620 10520 8660 10529
rect 8620 10385 8660 10480
rect 8524 10352 8564 10361
rect 8524 10217 8564 10312
rect 8620 10268 8660 10277
rect 8620 10133 8660 10228
rect 8428 9967 8468 9976
rect 8332 9932 8372 9941
rect 8332 9596 8372 9892
rect 8716 9764 8756 11152
rect 8716 9715 8756 9724
rect 8332 9547 8372 9556
rect 8140 9463 8180 9472
rect 7276 8455 7316 8464
rect 7756 9428 7796 9437
rect 7276 8084 7316 8093
rect 7316 8044 7412 8084
rect 7276 8035 7316 8044
rect 7084 7951 7124 7960
rect 7372 7916 7412 8044
rect 7372 7867 7412 7876
rect 7276 7832 7316 7841
rect 6892 7111 6932 7120
rect 7084 7748 7124 7757
rect 6220 6607 6260 6616
rect 6028 6404 6068 6413
rect 5740 5767 5780 5776
rect 5932 6320 5972 6329
rect 5740 5648 5780 5657
rect 5356 5060 5396 5069
rect 5356 4220 5396 5020
rect 5356 4171 5396 4180
rect 5452 4976 5492 4985
rect 5260 4087 5300 4096
rect 5452 4136 5492 4936
rect 5452 3632 5492 4096
rect 5452 3583 5492 3592
rect 5644 3884 5684 3893
rect 4972 3247 5012 3256
rect 5644 2900 5684 3844
rect 5740 3632 5780 5608
rect 5932 5480 5972 6280
rect 5932 5431 5972 5440
rect 6028 5144 6068 6364
rect 7084 6404 7124 7708
rect 7276 7412 7316 7792
rect 7276 7363 7316 7372
rect 6604 6320 6644 6329
rect 6508 6068 6548 6077
rect 6412 5732 6452 5741
rect 6124 5692 6412 5732
rect 6124 5648 6164 5692
rect 6412 5683 6452 5692
rect 6124 5599 6164 5608
rect 6028 5095 6068 5104
rect 6316 5564 6356 5573
rect 6316 4976 6356 5524
rect 6316 4927 6356 4936
rect 5740 3583 5780 3592
rect 6028 3632 6068 3641
rect 5644 2860 5780 2900
rect 4396 1063 4436 1072
rect 4876 1448 4916 2752
rect 5740 2456 5780 2860
rect 5740 2407 5780 2416
rect 5836 2624 5876 2633
rect 5836 1784 5876 2584
rect 5740 1700 5780 1709
rect 4876 1112 4916 1408
rect 5548 1448 5588 1457
rect 4972 1280 5012 1289
rect 5164 1280 5204 1289
rect 5012 1240 5164 1280
rect 4972 1231 5012 1240
rect 5164 1231 5204 1240
rect 4876 1063 4916 1072
rect 5548 944 5588 1408
rect 5548 895 5588 904
rect 4352 776 4720 785
rect 4352 727 4720 736
rect 5740 776 5780 1660
rect 5836 1154 5876 1744
rect 6028 2036 6068 3592
rect 5836 1105 5876 1114
rect 5932 1616 5972 1625
rect 5932 1028 5972 1576
rect 5932 979 5972 988
rect 6028 944 6068 1996
rect 6124 3464 6164 3473
rect 6124 3296 6164 3424
rect 6508 3464 6548 6028
rect 6604 4052 6644 6280
rect 6796 6152 6836 6161
rect 6700 5984 6740 5993
rect 6700 5480 6740 5944
rect 6700 5431 6740 5440
rect 6604 4003 6644 4012
rect 6796 3632 6836 6112
rect 7084 6068 7124 6364
rect 7084 6019 7124 6028
rect 6796 3583 6836 3592
rect 6892 5816 6932 5825
rect 6932 5776 7124 5816
rect 6892 5312 6932 5776
rect 7084 5648 7124 5776
rect 7084 5599 7124 5608
rect 6892 4220 6932 5272
rect 7372 4976 7412 4985
rect 7372 4388 7412 4936
rect 7372 4339 7412 4348
rect 7468 4892 7508 4901
rect 6508 3415 6548 3424
rect 6124 1784 6164 3256
rect 6892 3296 6932 4180
rect 7276 4136 7316 4145
rect 7276 4001 7316 4096
rect 6892 3247 6932 3256
rect 7084 3212 7124 3221
rect 6700 2792 6740 2801
rect 6124 1735 6164 1744
rect 6412 1952 6452 1961
rect 6028 895 6068 904
rect 6412 860 6452 1912
rect 6700 1616 6740 2752
rect 6892 2792 6932 2801
rect 6892 2120 6932 2752
rect 7084 2708 7124 3172
rect 7468 2876 7508 4852
rect 7756 4724 7796 9388
rect 8716 9428 8756 9437
rect 8332 9260 8372 9269
rect 8332 8924 8372 9220
rect 8332 8875 8372 8884
rect 7852 8000 7892 8009
rect 7852 7865 7892 7960
rect 8236 7244 8276 7253
rect 8140 7160 8180 7169
rect 8140 6572 8180 7120
rect 8140 5480 8180 6532
rect 8236 6488 8276 7204
rect 8620 7160 8660 7169
rect 8620 6656 8660 7120
rect 8716 6992 8756 9388
rect 8812 8588 8852 16024
rect 8908 15476 8948 15485
rect 8908 15341 8948 15436
rect 9004 14888 9044 16276
rect 9196 15728 9236 16360
rect 9196 15679 9236 15688
rect 9292 16988 9332 17536
rect 9292 15728 9332 16948
rect 9388 15896 9428 20812
rect 9484 17660 9524 17669
rect 9484 17408 9524 17620
rect 9484 17359 9524 17368
rect 9484 17072 9524 17081
rect 9484 16820 9524 17032
rect 9484 16771 9524 16780
rect 9484 16568 9524 16577
rect 9484 16064 9524 16528
rect 9676 16232 9716 21316
rect 9772 19508 9812 19517
rect 9772 19340 9812 19468
rect 9772 18500 9812 19300
rect 9772 18451 9812 18460
rect 9676 16183 9716 16192
rect 9772 16568 9812 16577
rect 9484 16015 9524 16024
rect 9772 16148 9812 16528
rect 9388 15856 9620 15896
rect 9292 15679 9332 15688
rect 9100 15644 9140 15653
rect 9484 15644 9524 15653
rect 9100 15476 9140 15604
rect 9388 15604 9484 15644
rect 9100 15427 9140 15436
rect 9196 15476 9236 15485
rect 9100 14888 9140 14897
rect 9004 14848 9100 14888
rect 9004 14636 9044 14645
rect 9004 14132 9044 14596
rect 8908 13964 8948 13973
rect 8908 13544 8948 13924
rect 9004 13712 9044 14092
rect 9004 13663 9044 13672
rect 8908 13504 9044 13544
rect 8908 13376 8948 13385
rect 8908 13241 8948 13336
rect 8908 13040 8948 13049
rect 8908 12704 8948 13000
rect 8908 12655 8948 12664
rect 8908 12368 8948 12377
rect 8908 12233 8948 12328
rect 9004 11780 9044 13504
rect 9100 13208 9140 14848
rect 9196 14720 9236 15436
rect 9388 15392 9428 15604
rect 9484 15595 9524 15604
rect 9388 15343 9428 15352
rect 9580 15308 9620 15856
rect 9196 13544 9236 14680
rect 9484 15268 9620 15308
rect 9484 14720 9524 15268
rect 9580 15140 9620 15149
rect 9620 15100 9716 15140
rect 9580 15091 9620 15100
rect 9196 13495 9236 13504
rect 9388 14132 9428 14141
rect 9100 13124 9140 13168
rect 9100 13075 9140 13084
rect 9388 12788 9428 14092
rect 9388 12739 9428 12748
rect 9484 12620 9524 14680
rect 9676 14720 9716 15100
rect 9196 12580 9484 12620
rect 9004 11731 9044 11740
rect 9100 12536 9140 12545
rect 8908 11696 8948 11705
rect 8908 11612 8948 11656
rect 8908 11572 9044 11612
rect 8908 11024 8948 11033
rect 8908 10772 8948 10984
rect 9004 10856 9044 11572
rect 9100 11192 9140 12496
rect 9196 11696 9236 12580
rect 9484 12571 9524 12580
rect 9580 14636 9620 14645
rect 9196 11647 9236 11656
rect 9100 11143 9140 11152
rect 9100 10856 9140 10865
rect 9004 10816 9100 10856
rect 8908 10723 8948 10732
rect 9004 10352 9044 10447
rect 9004 10303 9044 10312
rect 8908 10184 8948 10193
rect 8908 9680 8948 10144
rect 9004 10184 9044 10193
rect 9004 10016 9044 10144
rect 9004 9965 9044 9976
rect 8908 9631 8948 9640
rect 9100 8756 9140 10816
rect 9580 10856 9620 14596
rect 9676 13544 9716 14680
rect 9676 13495 9716 13504
rect 9676 12536 9716 12545
rect 9676 12452 9716 12496
rect 9676 12401 9716 12412
rect 9580 10807 9620 10816
rect 9676 11780 9716 11789
rect 9292 10436 9332 10445
rect 9196 10184 9236 10195
rect 9196 10100 9236 10144
rect 9196 10051 9236 10060
rect 9196 9680 9236 9689
rect 9196 9545 9236 9640
rect 8812 8539 8852 8548
rect 9004 8672 9044 8681
rect 8908 8000 8948 8009
rect 8908 7412 8948 7960
rect 8908 7363 8948 7372
rect 8716 6943 8756 6952
rect 8620 6607 8660 6616
rect 8236 6439 8276 6448
rect 9004 6572 9044 8632
rect 8140 5431 8180 5440
rect 8716 5648 8756 5657
rect 8716 5312 8756 5608
rect 8716 5263 8756 5272
rect 8908 5564 8948 5573
rect 8620 5060 8660 5069
rect 7756 4675 7796 4684
rect 8428 4976 8468 4985
rect 7468 2827 7508 2836
rect 7084 2659 7124 2668
rect 6892 2071 6932 2080
rect 6700 1567 6740 1576
rect 7564 1784 7604 1793
rect 7564 1196 7604 1744
rect 8428 1364 8468 4936
rect 8620 4925 8660 5020
rect 8812 4976 8852 4985
rect 8812 4640 8852 4936
rect 8524 4388 8564 4397
rect 8524 4136 8564 4348
rect 8524 3464 8564 4096
rect 8812 4136 8852 4600
rect 8524 3415 8564 3424
rect 8716 3968 8756 3977
rect 8716 3128 8756 3928
rect 8812 3548 8852 4096
rect 8812 3499 8852 3508
rect 8716 3079 8756 3088
rect 8908 2624 8948 5524
rect 9004 4976 9044 6532
rect 9100 5732 9140 8716
rect 9196 9008 9236 9017
rect 9196 6488 9236 8968
rect 9292 8672 9332 10396
rect 9676 10100 9716 11740
rect 9772 11696 9812 16108
rect 9772 11647 9812 11656
rect 9772 10940 9812 10949
rect 9772 10805 9812 10900
rect 9868 10184 9908 24928
rect 9964 24716 10004 25348
rect 9964 24667 10004 24676
rect 10156 25136 10196 25145
rect 10156 24716 10196 25096
rect 10156 24667 10196 24676
rect 10252 24548 10292 26692
rect 10252 24499 10292 24508
rect 10060 23876 10100 23885
rect 10060 23741 10100 23836
rect 10252 23288 10292 23297
rect 9964 22112 10004 22121
rect 9964 21524 10004 22072
rect 9964 21475 10004 21484
rect 10156 22112 10196 22121
rect 10060 20180 10100 20275
rect 10060 20131 10100 20140
rect 9964 19256 10004 19267
rect 9964 19172 10004 19216
rect 9964 19123 10004 19132
rect 10060 17744 10100 17753
rect 9964 17492 10004 17501
rect 9964 16400 10004 17452
rect 10060 17240 10100 17704
rect 10060 17191 10100 17200
rect 9964 16351 10004 16360
rect 9964 16232 10004 16241
rect 9964 16097 10004 16192
rect 10060 16064 10100 16073
rect 10060 15929 10100 16024
rect 9964 15896 10004 15905
rect 9964 15812 10004 15856
rect 9964 15772 10100 15812
rect 9964 15644 10004 15653
rect 9964 15509 10004 15604
rect 9964 15392 10004 15401
rect 9964 15257 10004 15352
rect 10060 14804 10100 15772
rect 10156 15476 10196 22072
rect 10156 15427 10196 15436
rect 10060 14755 10100 14764
rect 10156 14972 10196 14981
rect 9964 14720 10004 14729
rect 9964 13880 10004 14680
rect 9964 13831 10004 13840
rect 10156 13964 10196 14932
rect 10252 14972 10292 23248
rect 10348 19760 10388 27364
rect 10540 27404 10580 27413
rect 10444 26564 10484 26573
rect 10444 25892 10484 26524
rect 10444 25843 10484 25852
rect 10444 25724 10484 25733
rect 10444 25220 10484 25684
rect 10540 25724 10580 27364
rect 10828 27404 10868 28600
rect 11596 27824 11636 28600
rect 12364 28412 12404 28600
rect 12364 28363 12404 28372
rect 12126 27992 12494 28001
rect 12126 27943 12494 27952
rect 11596 27775 11636 27784
rect 11788 27908 11828 27917
rect 11692 27740 11732 27749
rect 10828 27355 10868 27364
rect 11596 27656 11636 27665
rect 10886 27236 11254 27245
rect 10886 27187 11254 27196
rect 10828 26900 10868 26909
rect 10540 25675 10580 25684
rect 10636 26144 10676 26153
rect 10540 25556 10580 25565
rect 10540 25388 10580 25516
rect 10540 25339 10580 25348
rect 10444 25171 10484 25180
rect 10444 24800 10484 24809
rect 10444 24665 10484 24760
rect 10540 24548 10580 24557
rect 10444 24380 10484 24389
rect 10444 24212 10484 24340
rect 10444 24163 10484 24172
rect 10540 24044 10580 24508
rect 10540 23995 10580 24004
rect 10444 23792 10484 23801
rect 10444 23036 10484 23752
rect 10444 22987 10484 22996
rect 10540 23624 10580 23633
rect 10540 23204 10580 23584
rect 10444 21440 10484 21449
rect 10444 20768 10484 21400
rect 10444 20719 10484 20728
rect 10348 19720 10484 19760
rect 10252 14923 10292 14932
rect 10348 17744 10388 17753
rect 10348 14888 10388 17704
rect 10444 16484 10484 19720
rect 10444 16435 10484 16444
rect 10444 16232 10484 16241
rect 10444 14888 10484 16192
rect 10540 15728 10580 23164
rect 10636 22784 10676 26104
rect 10828 25976 10868 26860
rect 11404 26564 11444 26573
rect 11404 26312 11444 26524
rect 11404 26263 11444 26272
rect 11596 26312 11636 27616
rect 11692 27068 11732 27700
rect 11692 27019 11732 27028
rect 10828 25927 10868 25936
rect 11308 26144 11348 26153
rect 10886 25724 11254 25733
rect 10886 25675 11254 25684
rect 11116 25556 11156 25565
rect 10732 25472 10772 25481
rect 10732 23960 10772 25432
rect 11116 25388 11156 25516
rect 11308 25556 11348 26104
rect 11500 26060 11540 26069
rect 11308 25507 11348 25516
rect 11404 25892 11444 25901
rect 11116 25339 11156 25348
rect 10828 25304 10868 25313
rect 10828 25169 10868 25264
rect 11116 25220 11156 25229
rect 10924 25052 10964 25061
rect 10924 24632 10964 25012
rect 10924 24583 10964 24592
rect 11116 24548 11156 25180
rect 11116 24413 11156 24508
rect 11308 25052 11348 25061
rect 10886 24212 11254 24221
rect 10886 24163 11254 24172
rect 10828 23960 10868 23969
rect 10732 23920 10828 23960
rect 10828 23288 10868 23920
rect 10924 23792 10964 23801
rect 10964 23752 11060 23792
rect 10924 23743 10964 23752
rect 10924 23288 10964 23297
rect 10828 23248 10924 23288
rect 10924 23239 10964 23248
rect 11020 22952 11060 23752
rect 11212 23624 11252 23633
rect 11212 23204 11252 23584
rect 11212 23155 11252 23164
rect 11020 22903 11060 22912
rect 11116 23120 11156 23129
rect 11116 22952 11156 23080
rect 11116 22903 11156 22912
rect 10636 22735 10676 22744
rect 10886 22700 11254 22709
rect 10886 22651 11254 22660
rect 11212 22532 11252 22541
rect 10636 22448 10676 22457
rect 10636 17660 10676 22408
rect 11212 21608 11252 22492
rect 11212 21559 11252 21568
rect 11308 22280 11348 25012
rect 11404 24632 11444 25852
rect 11500 25640 11540 26020
rect 11500 25591 11540 25600
rect 11500 25472 11540 25481
rect 11500 24968 11540 25432
rect 11500 24919 11540 24928
rect 11596 25304 11636 26272
rect 11596 24716 11636 25264
rect 11692 25808 11732 25817
rect 11692 25136 11732 25768
rect 11692 25087 11732 25096
rect 11596 24667 11636 24676
rect 11404 22448 11444 24592
rect 11692 24632 11732 24641
rect 11500 24464 11540 24473
rect 11500 23120 11540 24424
rect 11692 24044 11732 24592
rect 11692 23995 11732 24004
rect 11692 23456 11732 23465
rect 11692 23204 11732 23416
rect 11692 23155 11732 23164
rect 11500 23060 11540 23080
rect 11500 23020 11636 23060
rect 11404 22399 11444 22408
rect 11500 22952 11540 22961
rect 10732 21524 10772 21533
rect 10732 20768 10772 21484
rect 11308 21524 11348 22240
rect 11500 21608 11540 22912
rect 11596 22532 11636 23020
rect 11596 22483 11636 22492
rect 11692 22952 11732 22961
rect 11692 21776 11732 22912
rect 11788 22280 11828 27868
rect 12460 26900 12500 26909
rect 12500 26860 12692 26900
rect 12460 26851 12500 26860
rect 12126 26480 12494 26489
rect 12126 26431 12494 26440
rect 12556 26480 12596 26489
rect 11980 26396 12020 26405
rect 11884 26228 11924 26237
rect 11884 25136 11924 26188
rect 11980 26144 12020 26356
rect 12556 26228 12596 26440
rect 12556 26179 12596 26188
rect 11980 26095 12020 26104
rect 12460 26144 12500 26153
rect 12460 25976 12500 26104
rect 12460 25927 12500 25936
rect 12652 26144 12692 26860
rect 11980 25892 12020 25901
rect 11980 25757 12020 25852
rect 12652 25304 12692 26104
rect 12748 26816 12788 26825
rect 12748 25976 12788 26776
rect 12844 26648 12884 26657
rect 12844 26228 12884 26608
rect 12940 26480 12980 26489
rect 12940 26345 12980 26440
rect 12844 26179 12884 26188
rect 12940 26144 12980 26239
rect 12940 26095 12980 26104
rect 12748 25927 12788 25936
rect 12844 26060 12884 26069
rect 12844 25556 12884 26020
rect 12844 25507 12884 25516
rect 12940 25976 12980 25985
rect 12652 25255 12692 25264
rect 11884 24464 11924 25096
rect 11884 23876 11924 24424
rect 11884 23288 11924 23836
rect 11884 23239 11924 23248
rect 11980 25220 12020 25229
rect 11788 22231 11828 22240
rect 11980 23036 12020 25180
rect 12126 24968 12494 24977
rect 12126 24919 12494 24928
rect 12652 24548 12692 24557
rect 12556 23876 12596 23971
rect 12556 23827 12596 23836
rect 12126 23456 12494 23465
rect 12126 23407 12494 23416
rect 12460 23288 12500 23297
rect 12460 23204 12500 23248
rect 12460 23153 12500 23164
rect 11692 21727 11732 21736
rect 11500 21559 11540 21568
rect 11692 21608 11732 21617
rect 11732 21568 11828 21608
rect 11692 21559 11732 21568
rect 11308 21475 11348 21484
rect 11404 21440 11444 21449
rect 10886 21188 11254 21197
rect 10886 21139 11254 21148
rect 11404 21188 11444 21400
rect 11404 21139 11444 21148
rect 10732 20096 10772 20728
rect 11212 21020 11252 21029
rect 11020 20684 11060 20693
rect 10924 20600 10964 20609
rect 10924 20264 10964 20560
rect 10924 20215 10964 20224
rect 10732 20047 10772 20056
rect 11020 20096 11060 20644
rect 11020 20047 11060 20056
rect 11212 20096 11252 20980
rect 11500 21020 11540 21029
rect 11212 20047 11252 20056
rect 11404 20936 11444 20945
rect 11404 20012 11444 20896
rect 11500 20885 11540 20980
rect 11692 20852 11732 20861
rect 11404 19963 11444 19972
rect 11596 20768 11636 20777
rect 10732 19928 10772 19937
rect 10732 19340 10772 19888
rect 11500 19844 11540 19853
rect 10886 19676 11254 19685
rect 10886 19627 11254 19636
rect 10732 19291 10772 19300
rect 10924 19424 10964 19433
rect 10924 19088 10964 19384
rect 10924 19039 10964 19048
rect 11308 19340 11348 19349
rect 10828 19004 10868 19013
rect 10828 18668 10868 18964
rect 11308 18752 11348 19300
rect 11500 19340 11540 19804
rect 11596 19676 11636 20728
rect 11596 19627 11636 19636
rect 11404 19256 11444 19265
rect 11404 19004 11444 19216
rect 11404 18955 11444 18964
rect 11308 18703 11348 18712
rect 10828 18619 10868 18628
rect 11212 18584 11252 18593
rect 11212 18449 11252 18544
rect 11500 18584 11540 19300
rect 11692 18920 11732 20812
rect 11692 18871 11732 18880
rect 11788 18752 11828 21568
rect 11980 21440 12020 22996
rect 12556 23120 12596 23129
rect 12556 22985 12596 23080
rect 12460 22952 12500 22961
rect 12076 22616 12116 22625
rect 12076 22364 12116 22576
rect 12076 22315 12116 22324
rect 12460 22364 12500 22912
rect 12460 22315 12500 22324
rect 12364 22280 12404 22289
rect 12364 22145 12404 22240
rect 12652 22196 12692 24508
rect 12844 23624 12884 23633
rect 12652 22147 12692 22156
rect 12748 22532 12788 22541
rect 12126 21944 12494 21953
rect 12126 21895 12494 21904
rect 12748 21776 12788 22492
rect 12844 22448 12884 23584
rect 12940 23204 12980 25936
rect 13036 25472 13076 25481
rect 13036 24548 13076 25432
rect 13036 24499 13076 24508
rect 12940 23155 12980 23164
rect 12844 22399 12884 22408
rect 12844 22196 12884 22205
rect 12844 22061 12884 22156
rect 13036 22196 13076 22205
rect 11980 21391 12020 21400
rect 12364 21440 12404 21449
rect 12364 21104 12404 21400
rect 12364 21055 12404 21064
rect 11980 20936 12020 20945
rect 11884 20768 11924 20777
rect 11884 20516 11924 20728
rect 11884 20467 11924 20476
rect 11980 20348 12020 20896
rect 12748 20684 12788 21736
rect 13036 21608 13076 22156
rect 13132 21776 13172 28600
rect 13900 28580 13940 28600
rect 13900 28531 13940 28540
rect 14668 28160 14708 28600
rect 14668 28111 14708 28120
rect 15436 28076 15476 28600
rect 15436 28027 15476 28036
rect 16204 27908 16244 28600
rect 16204 27859 16244 27868
rect 15148 27656 15188 27665
rect 13324 27404 13364 27413
rect 13324 26984 13364 27364
rect 13804 27404 13844 27413
rect 13324 25304 13364 26944
rect 13708 26984 13748 26993
rect 13708 26060 13748 26944
rect 13804 26480 13844 27364
rect 14476 27404 14516 27413
rect 13804 26431 13844 26440
rect 14380 26816 14420 26825
rect 13708 26011 13748 26020
rect 14380 26144 14420 26776
rect 13324 23060 13364 25264
rect 14380 24632 14420 26104
rect 14476 26144 14516 27364
rect 14668 27404 14708 27413
rect 14668 26648 14708 27364
rect 14668 26599 14708 26608
rect 15148 26312 15188 27616
rect 15724 27572 15764 27581
rect 15724 26984 15764 27532
rect 15724 26935 15764 26944
rect 16204 26816 16244 26825
rect 15148 26263 15188 26272
rect 16108 26480 16148 26489
rect 14476 26095 14516 26104
rect 15820 26144 15860 26153
rect 16108 26144 16148 26440
rect 15860 26104 16108 26144
rect 15820 26095 15860 26104
rect 16108 26095 16148 26104
rect 16204 26060 16244 26776
rect 16204 26011 16244 26020
rect 15148 25724 15188 25733
rect 14668 25472 14708 25481
rect 14188 24464 14228 24473
rect 13900 24380 13940 24389
rect 13228 23020 13364 23060
rect 13420 24128 13460 24137
rect 13228 22028 13268 23020
rect 13324 22280 13364 22289
rect 13324 22145 13364 22240
rect 13228 21979 13268 21988
rect 13132 21727 13172 21736
rect 12126 20432 12494 20441
rect 12126 20383 12494 20392
rect 11980 20299 12020 20308
rect 11980 19676 12020 19685
rect 11884 19508 11924 19517
rect 11884 19256 11924 19468
rect 11980 19424 12020 19636
rect 11980 19375 12020 19384
rect 11884 19207 11924 19216
rect 12460 19340 12500 19349
rect 12460 19256 12500 19300
rect 12460 19205 12500 19216
rect 11500 18535 11540 18544
rect 11596 18712 11828 18752
rect 11980 19172 12020 19181
rect 11404 18500 11444 18509
rect 11020 18332 11060 18341
rect 10732 18292 11020 18332
rect 10732 17744 10772 18292
rect 11020 18283 11060 18292
rect 10886 18164 11254 18173
rect 10886 18115 11254 18124
rect 11212 17828 11252 17837
rect 11212 17744 11252 17788
rect 11308 17744 11348 17753
rect 10732 17704 10868 17744
rect 11212 17704 11308 17744
rect 10636 17611 10676 17620
rect 10732 17576 10772 17585
rect 10636 17408 10676 17417
rect 10636 17156 10676 17368
rect 10636 17107 10676 17116
rect 10540 15679 10580 15688
rect 10636 16988 10676 16997
rect 10636 16148 10676 16948
rect 10732 16316 10772 17536
rect 10828 17408 10868 17704
rect 11308 17695 11348 17704
rect 10828 17359 10868 17368
rect 11020 17660 11060 17669
rect 11020 17240 11060 17620
rect 11404 17660 11444 18460
rect 11404 17611 11444 17620
rect 11500 17996 11540 18005
rect 11020 17191 11060 17200
rect 11404 17240 11444 17249
rect 11404 17105 11444 17200
rect 10828 17072 10868 17081
rect 10828 16937 10868 17032
rect 11020 17072 11060 17081
rect 11020 16904 11060 17032
rect 11020 16855 11060 16864
rect 11212 16988 11252 16997
rect 11212 16853 11252 16948
rect 10886 16652 11254 16661
rect 10886 16603 11254 16612
rect 10732 16267 10772 16276
rect 10540 15560 10580 15569
rect 10540 15425 10580 15520
rect 10444 14848 10580 14888
rect 10348 14839 10388 14848
rect 10252 14804 10292 14813
rect 10252 14669 10292 14764
rect 10444 14720 10484 14729
rect 10348 14300 10388 14309
rect 10348 14048 10388 14260
rect 10444 14216 10484 14680
rect 10540 14300 10580 14848
rect 10540 14251 10580 14260
rect 10444 14167 10484 14176
rect 10636 14216 10676 16108
rect 11212 16232 11252 16241
rect 11116 15728 11156 15737
rect 10732 15560 10772 15569
rect 10732 15392 10772 15520
rect 10732 15343 10772 15352
rect 11116 15308 11156 15688
rect 11212 15392 11252 16192
rect 11404 16064 11444 16073
rect 11404 15896 11444 16024
rect 11404 15847 11444 15856
rect 11500 15644 11540 17956
rect 11500 15595 11540 15604
rect 11212 15343 11252 15352
rect 11500 15476 11540 15485
rect 11116 15259 11156 15268
rect 10886 15140 11254 15149
rect 10886 15091 11254 15100
rect 10732 14972 10772 14981
rect 10732 14720 10772 14932
rect 10732 14671 10772 14680
rect 11212 14720 11252 14729
rect 11404 14720 11444 14729
rect 10636 14167 10676 14176
rect 10348 13999 10388 14008
rect 10540 14132 10580 14141
rect 10156 13124 10196 13924
rect 10156 13075 10196 13084
rect 10348 13292 10388 13301
rect 10156 12956 10196 12965
rect 9964 11780 10004 11789
rect 9964 11645 10004 11740
rect 10156 11696 10196 12916
rect 9964 11444 10004 11453
rect 9964 11024 10004 11404
rect 10156 11108 10196 11656
rect 10156 11059 10196 11068
rect 10348 12200 10388 13252
rect 10444 13124 10484 13152
rect 10540 13124 10580 14092
rect 11212 14132 11252 14680
rect 11212 14083 11252 14092
rect 11308 14680 11404 14720
rect 10732 14048 10772 14057
rect 10636 13460 10676 13469
rect 10636 13292 10676 13420
rect 10636 13243 10676 13252
rect 10484 13084 10580 13124
rect 10444 13075 10484 13084
rect 10348 11864 10388 12160
rect 9964 10975 10004 10984
rect 10252 11024 10292 11033
rect 10156 10940 10196 10951
rect 10156 10856 10196 10900
rect 10156 10807 10196 10816
rect 9868 10135 9908 10144
rect 10060 10100 10100 10109
rect 9676 10060 9812 10100
rect 9388 9848 9428 9857
rect 9388 9713 9428 9808
rect 9292 8623 9332 8632
rect 9772 9092 9812 10060
rect 10060 9092 10100 10060
rect 10252 9512 10292 10984
rect 10348 10856 10388 11824
rect 10444 11948 10484 11957
rect 10444 11024 10484 11908
rect 10540 11864 10580 13084
rect 10636 12536 10676 12545
rect 10636 12032 10676 12496
rect 10732 12368 10772 14008
rect 11308 14048 11348 14680
rect 11404 14671 11444 14680
rect 10886 13628 11254 13637
rect 10886 13579 11254 13588
rect 11116 13460 11156 13469
rect 11116 13376 11156 13420
rect 11308 13460 11348 14008
rect 11308 13411 11348 13420
rect 11404 13880 11444 13889
rect 10924 13336 11156 13376
rect 10924 13124 10964 13336
rect 10924 13075 10964 13084
rect 11020 13208 11060 13217
rect 10732 12319 10772 12328
rect 10828 12452 10868 12461
rect 10828 12317 10868 12412
rect 11020 12452 11060 13168
rect 11020 12403 11060 12412
rect 11116 12536 11156 13336
rect 11404 13292 11444 13840
rect 11404 12956 11444 13252
rect 11404 12907 11444 12916
rect 11116 12284 11156 12496
rect 11116 12235 11156 12244
rect 11308 12704 11348 12713
rect 10636 11983 10676 11992
rect 10732 12200 10772 12209
rect 10540 11815 10580 11824
rect 10540 11696 10580 11705
rect 10540 11561 10580 11656
rect 10444 10975 10484 10984
rect 10540 11192 10580 11201
rect 10540 10856 10580 11152
rect 10348 10807 10388 10816
rect 10444 10816 10580 10856
rect 10444 10100 10484 10816
rect 10540 10688 10580 10697
rect 10540 10268 10580 10648
rect 10732 10352 10772 12160
rect 10886 12116 11254 12125
rect 10886 12067 11254 12076
rect 10924 11864 10964 11873
rect 10924 11696 10964 11824
rect 11020 11696 11060 11705
rect 10924 11656 11020 11696
rect 11020 11647 11060 11656
rect 11212 11696 11252 11705
rect 11020 11024 11060 11033
rect 11020 10889 11060 10984
rect 11212 10772 11252 11656
rect 11308 10940 11348 12664
rect 11500 11948 11540 15436
rect 11596 14972 11636 18712
rect 11980 18668 12020 19132
rect 12556 19172 12596 19181
rect 12126 18920 12494 18929
rect 12126 18871 12494 18880
rect 11980 18619 12020 18628
rect 11788 18584 11828 18593
rect 11692 18500 11732 18509
rect 11692 17072 11732 18460
rect 11692 16820 11732 17032
rect 11692 16771 11732 16780
rect 11788 16484 11828 18544
rect 12556 17492 12596 19132
rect 12556 17443 12596 17452
rect 12126 17408 12494 17417
rect 12126 17359 12494 17368
rect 11884 17156 11924 17165
rect 11884 17072 11924 17116
rect 11884 17021 11924 17032
rect 11788 16435 11828 16444
rect 12460 16988 12500 16997
rect 12268 16316 12308 16325
rect 12268 16232 12308 16276
rect 12460 16232 12500 16948
rect 12652 16820 12692 16829
rect 12556 16736 12596 16745
rect 12556 16601 12596 16696
rect 12652 16685 12692 16780
rect 12748 16400 12788 20644
rect 12940 20684 12980 20693
rect 12940 20549 12980 20644
rect 13036 19844 13076 21568
rect 13324 21608 13364 21617
rect 13324 20684 13364 21568
rect 13324 20635 13364 20644
rect 13420 20264 13460 24088
rect 13900 23792 13940 24340
rect 13900 23743 13940 23752
rect 14188 23792 14228 24424
rect 14380 23876 14420 24592
rect 14380 23827 14420 23836
rect 14476 25304 14516 25313
rect 14476 24968 14516 25264
rect 14188 23743 14228 23752
rect 13612 23708 13652 23717
rect 13612 23120 13652 23668
rect 13612 23071 13652 23080
rect 14476 22616 14516 24928
rect 14668 23036 14708 25432
rect 14860 24632 14900 24641
rect 14860 23792 14900 24592
rect 15148 24548 15188 25684
rect 15340 25304 15380 25313
rect 15340 24800 15380 25264
rect 15340 24751 15380 24760
rect 16012 25136 16052 25145
rect 15148 23876 15188 24508
rect 15148 23827 15188 23836
rect 15244 24380 15284 24389
rect 14860 23743 14900 23752
rect 15244 23792 15284 24340
rect 16012 24044 16052 25096
rect 16012 23995 16052 24004
rect 16108 24632 16148 24641
rect 15244 23743 15284 23752
rect 15820 23540 15860 23549
rect 15820 23120 15860 23500
rect 16108 23204 16148 24592
rect 16108 23155 16148 23164
rect 15820 23071 15860 23080
rect 16012 23120 16052 23129
rect 14668 22987 14708 22996
rect 14476 22567 14516 22576
rect 15244 22280 15284 22291
rect 15244 22196 15284 22240
rect 15244 22147 15284 22156
rect 13612 21608 13652 21617
rect 13612 21020 13652 21568
rect 13612 20971 13652 20980
rect 14476 21440 14516 21449
rect 14476 20852 14516 21400
rect 14476 20803 14516 20812
rect 15052 21020 15092 21029
rect 14380 20684 14420 20693
rect 14092 20600 14132 20609
rect 14092 20516 14132 20560
rect 14092 20465 14132 20476
rect 12844 18080 12884 18089
rect 12844 17324 12884 18040
rect 13036 17828 13076 19804
rect 13228 20096 13268 20105
rect 13420 20096 13460 20224
rect 13268 20056 13460 20096
rect 13516 20180 13556 20189
rect 13228 19340 13268 20056
rect 13228 19291 13268 19300
rect 13516 19256 13556 20140
rect 14380 20180 14420 20644
rect 14380 20131 14420 20140
rect 14476 20264 14516 20273
rect 13516 19207 13556 19216
rect 13708 20012 13748 20021
rect 13132 19172 13172 19181
rect 13132 18584 13172 19132
rect 13132 18535 13172 18544
rect 13420 18752 13460 18761
rect 13036 17779 13076 17788
rect 13420 17744 13460 18712
rect 13708 18584 13748 19972
rect 13612 18332 13652 18341
rect 12940 17324 12980 17333
rect 12844 17284 12940 17324
rect 12940 17275 12980 17284
rect 13228 17324 13268 17333
rect 12844 17072 12884 17081
rect 12844 16652 12884 17032
rect 12844 16603 12884 16612
rect 12268 16192 12460 16232
rect 12460 16183 12500 16192
rect 12652 16360 12788 16400
rect 12844 16400 12884 16409
rect 11692 16148 11732 16157
rect 11692 15728 11732 16108
rect 12556 16148 12596 16157
rect 11692 15679 11732 15688
rect 11980 16064 12020 16073
rect 11788 15560 11828 15569
rect 11596 14923 11636 14932
rect 11692 15056 11732 15065
rect 11692 14468 11732 15016
rect 11788 15056 11828 15520
rect 11788 15007 11828 15016
rect 11692 14419 11732 14428
rect 11884 14972 11924 14981
rect 11500 11899 11540 11908
rect 11596 13796 11636 13805
rect 11596 11864 11636 13756
rect 11788 13292 11828 13301
rect 11788 12452 11828 13252
rect 11788 12403 11828 12412
rect 11596 11815 11636 11824
rect 11500 11780 11540 11789
rect 11500 11192 11540 11740
rect 11884 11696 11924 14932
rect 11500 11143 11540 11152
rect 11596 11612 11636 11621
rect 11596 11108 11636 11572
rect 11596 11059 11636 11068
rect 11788 11612 11828 11621
rect 11788 11192 11828 11572
rect 11308 10891 11348 10900
rect 11500 10940 11540 10949
rect 11500 10805 11540 10900
rect 11788 10940 11828 11152
rect 11884 11024 11924 11656
rect 11884 10975 11924 10984
rect 11788 10891 11828 10900
rect 11884 10856 11924 10865
rect 11692 10772 11732 10781
rect 11212 10732 11348 10772
rect 10886 10604 11254 10613
rect 10886 10555 11254 10564
rect 10732 10303 10772 10312
rect 11116 10352 11156 10361
rect 10540 10219 10580 10228
rect 10636 10184 10676 10193
rect 10444 10060 10580 10100
rect 10444 9932 10484 9941
rect 10252 9463 10292 9472
rect 10348 9680 10388 9689
rect 10060 9052 10292 9092
rect 9772 8672 9812 9052
rect 9772 8623 9812 8632
rect 9676 8000 9716 8009
rect 9484 7748 9524 7757
rect 9484 7328 9524 7708
rect 9196 6439 9236 6448
rect 9388 7076 9428 7085
rect 9100 5683 9140 5692
rect 9004 4927 9044 4936
rect 9388 2708 9428 7036
rect 9484 6488 9524 7288
rect 9484 6439 9524 6448
rect 9676 6488 9716 7960
rect 10156 7202 10196 7211
rect 10156 7160 10196 7162
rect 9676 6439 9716 6448
rect 10060 7120 10196 7160
rect 10060 6572 10100 7120
rect 10252 7076 10292 9052
rect 10348 8672 10388 9640
rect 10444 9512 10484 9892
rect 10540 9596 10580 10060
rect 10636 9680 10676 10144
rect 11116 9848 11156 10312
rect 10636 9631 10676 9640
rect 10732 9808 11156 9848
rect 10540 9547 10580 9556
rect 10444 9463 10484 9472
rect 10636 9512 10676 9521
rect 10636 9176 10676 9472
rect 10636 9127 10676 9136
rect 10348 8623 10388 8632
rect 10444 8504 10484 8513
rect 10444 8369 10484 8464
rect 10060 5816 10100 6532
rect 9964 5776 10060 5816
rect 9484 4976 9524 4985
rect 9484 4388 9524 4936
rect 9484 4339 9524 4348
rect 9964 4136 10004 5776
rect 10060 5767 10100 5776
rect 10156 7036 10292 7076
rect 9964 4087 10004 4096
rect 10060 5648 10100 5657
rect 10060 4724 10100 5608
rect 10060 3968 10100 4684
rect 10060 3919 10100 3928
rect 10156 3380 10196 7036
rect 10252 5732 10292 5741
rect 10252 4976 10292 5692
rect 10252 4220 10292 4936
rect 10252 4171 10292 4180
rect 10636 4892 10676 4901
rect 10156 3331 10196 3340
rect 10636 2876 10676 4852
rect 10732 3632 10772 9808
rect 10828 9680 10868 9689
rect 10828 9545 10868 9640
rect 11212 9596 11252 9605
rect 10924 9512 10964 9521
rect 10924 9377 10964 9472
rect 11212 9461 11252 9556
rect 10886 9092 11254 9101
rect 10886 9043 11254 9052
rect 11212 8756 11252 8765
rect 11308 8756 11348 10732
rect 11404 10268 11444 10277
rect 11404 10133 11444 10228
rect 11596 9848 11636 9857
rect 11404 9680 11444 9689
rect 11404 9512 11444 9640
rect 11596 9680 11636 9808
rect 11596 9631 11636 9640
rect 11692 9512 11732 10732
rect 11788 10352 11828 10361
rect 11788 10184 11828 10312
rect 11788 10135 11828 10144
rect 11884 9680 11924 10816
rect 11980 10268 12020 16024
rect 12126 15896 12494 15905
rect 12126 15847 12494 15856
rect 12460 15476 12500 15485
rect 12556 15476 12596 16108
rect 12500 15436 12596 15476
rect 12460 15427 12500 15436
rect 12556 14720 12596 14729
rect 12126 14384 12494 14393
rect 12126 14335 12494 14344
rect 12460 14048 12500 14057
rect 12460 13544 12500 14008
rect 12460 13495 12500 13504
rect 12556 13124 12596 14680
rect 12652 14300 12692 16360
rect 12844 15980 12884 16360
rect 12844 15931 12884 15940
rect 13132 15812 13172 15823
rect 13132 15728 13172 15772
rect 13132 15679 13172 15688
rect 13228 15728 13268 17284
rect 13420 17072 13460 17704
rect 13420 17023 13460 17032
rect 13516 18248 13556 18257
rect 13516 17492 13556 18208
rect 13324 16820 13364 16829
rect 13324 16232 13364 16780
rect 13324 16064 13364 16192
rect 13324 16015 13364 16024
rect 13516 16064 13556 17452
rect 13612 17156 13652 18292
rect 13708 17828 13748 18544
rect 13708 17240 13748 17788
rect 13708 17191 13748 17200
rect 13804 19928 13844 19937
rect 13804 19256 13844 19888
rect 13804 17828 13844 19216
rect 14476 19256 14516 20224
rect 15052 20096 15092 20980
rect 14956 19424 14996 19433
rect 14476 19088 14516 19216
rect 14476 18752 14516 19048
rect 14860 19340 14900 19349
rect 14476 18584 14516 18712
rect 14476 18535 14516 18544
rect 14572 19004 14612 19013
rect 13900 17828 13940 17856
rect 13804 17788 13900 17828
rect 13612 16400 13652 17116
rect 13804 17072 13844 17788
rect 13900 17779 13940 17788
rect 13804 17023 13844 17032
rect 13900 17660 13940 17669
rect 13612 16351 13652 16360
rect 13804 16820 13844 16829
rect 13516 16015 13556 16024
rect 13804 16232 13844 16780
rect 13228 15679 13268 15688
rect 13804 15644 13844 16192
rect 13804 15595 13844 15604
rect 12652 14251 12692 14260
rect 12844 15560 12884 15569
rect 12556 13075 12596 13084
rect 12652 13964 12692 13973
rect 12126 12872 12494 12881
rect 12126 12823 12494 12832
rect 12556 12620 12596 12629
rect 12556 12032 12596 12580
rect 12556 11983 12596 11992
rect 12652 12452 12692 13924
rect 12748 13712 12788 13721
rect 12748 13292 12788 13672
rect 12748 13243 12788 13252
rect 12652 11948 12692 12412
rect 12652 11899 12692 11908
rect 12748 13124 12788 13133
rect 12748 12536 12788 13084
rect 12748 11780 12788 12496
rect 12126 11360 12494 11369
rect 12126 11311 12494 11320
rect 12748 11360 12788 11740
rect 12748 11311 12788 11320
rect 11980 10219 12020 10228
rect 12172 11108 12212 11117
rect 12172 10184 12212 11068
rect 12748 10436 12788 10445
rect 12172 10135 12212 10144
rect 12364 10268 12404 10277
rect 11884 9631 11924 9640
rect 11980 10100 12020 10109
rect 11444 9472 11540 9512
rect 11404 9463 11444 9472
rect 11404 9008 11444 9103
rect 11404 8959 11444 8968
rect 11252 8716 11348 8756
rect 11212 8707 11252 8716
rect 10886 7580 11254 7589
rect 10886 7531 11254 7540
rect 10886 6068 11254 6077
rect 10886 6019 11254 6028
rect 11308 5732 11348 8716
rect 11308 5683 11348 5692
rect 11404 8756 11444 8765
rect 11212 5648 11252 5657
rect 10924 5060 10964 5069
rect 10924 4976 10964 5020
rect 10924 4925 10964 4936
rect 11212 4892 11252 5608
rect 11404 5480 11444 8716
rect 11500 8672 11540 9472
rect 11500 8623 11540 8632
rect 11980 9512 12020 10060
rect 12364 10016 12404 10228
rect 12364 9967 12404 9976
rect 12126 9848 12494 9857
rect 12126 9799 12494 9808
rect 12364 9680 12404 9689
rect 12076 9512 12116 9521
rect 11980 9472 12076 9512
rect 11692 9344 11732 9472
rect 11692 8672 11732 9304
rect 11692 8623 11732 8632
rect 11884 9428 11924 9437
rect 11404 5431 11444 5440
rect 11500 8504 11540 8513
rect 11500 6404 11540 8464
rect 11788 7160 11828 7169
rect 11788 6992 11828 7120
rect 11788 6943 11828 6952
rect 11212 4843 11252 4852
rect 10886 4556 11254 4565
rect 10886 4507 11254 4516
rect 11500 4220 11540 6364
rect 11884 5564 11924 9388
rect 12076 8840 12116 9472
rect 12076 8791 12116 8800
rect 12268 8672 12308 8681
rect 12364 8672 12404 9640
rect 12748 9512 12788 10396
rect 12748 9463 12788 9472
rect 12844 8924 12884 15520
rect 12940 15560 12980 15569
rect 12940 14804 12980 15520
rect 13516 15560 13556 15569
rect 12940 14755 12980 14764
rect 13036 15476 13076 15485
rect 12940 13964 12980 13973
rect 12940 13292 12980 13924
rect 12940 13157 12980 13252
rect 13036 12704 13076 15436
rect 13228 15476 13268 15485
rect 13228 14972 13268 15436
rect 13228 14923 13268 14932
rect 13132 14720 13172 14729
rect 13132 14552 13172 14680
rect 13132 14503 13172 14512
rect 13516 14552 13556 15520
rect 13516 14503 13556 14512
rect 13612 15476 13652 15485
rect 13324 13376 13364 13385
rect 13132 13208 13172 13217
rect 13132 12872 13172 13168
rect 13228 13124 13268 13133
rect 13228 13040 13268 13084
rect 13228 12989 13268 13000
rect 13132 12832 13268 12872
rect 13036 12655 13076 12664
rect 12940 12452 12980 12461
rect 12940 12317 12980 12412
rect 13036 12368 13076 12377
rect 13036 11948 13076 12328
rect 12940 11864 12980 11904
rect 13036 11899 13076 11908
rect 13132 12116 13172 12125
rect 12940 11780 12980 11824
rect 13132 11864 13172 12076
rect 13228 12032 13268 12832
rect 13324 12536 13364 13336
rect 13324 12487 13364 12496
rect 13420 13124 13460 13133
rect 13420 12368 13460 13084
rect 13612 13040 13652 15436
rect 13612 12991 13652 13000
rect 13708 14720 13748 14729
rect 13228 11983 13268 11992
rect 13324 12328 13460 12368
rect 13516 12788 13556 12797
rect 13324 11864 13364 12328
rect 13516 12200 13556 12748
rect 13612 12620 13652 12629
rect 13612 12536 13652 12580
rect 13612 12452 13652 12496
rect 13612 12403 13652 12412
rect 13516 12151 13556 12160
rect 13612 12284 13652 12293
rect 13132 11815 13172 11824
rect 13228 11824 13364 11864
rect 13516 12032 13556 12041
rect 12940 11192 12980 11740
rect 13228 11612 13268 11824
rect 13132 11572 13228 11612
rect 12940 11143 12980 11152
rect 13036 11360 13076 11369
rect 13036 10016 13076 11320
rect 13036 9967 13076 9976
rect 12844 8875 12884 8884
rect 12940 9680 12980 9689
rect 12940 9512 12980 9640
rect 12460 8672 12500 8681
rect 12308 8632 12460 8672
rect 12268 8623 12308 8632
rect 12460 8623 12500 8632
rect 12126 8336 12494 8345
rect 12126 8287 12494 8296
rect 12364 8084 12404 8093
rect 12556 8084 12596 8093
rect 12404 8044 12556 8084
rect 12364 7412 12404 8044
rect 12556 8035 12596 8044
rect 12364 7363 12404 7372
rect 12748 7832 12788 7841
rect 12748 7412 12788 7792
rect 12748 7363 12788 7372
rect 12556 7160 12596 7169
rect 12556 6992 12596 7120
rect 12126 6824 12494 6833
rect 12126 6775 12494 6784
rect 11980 6488 12020 6497
rect 11980 6353 12020 6448
rect 12556 6320 12596 6952
rect 12940 7160 12980 9472
rect 13036 9428 13076 9437
rect 13036 9293 13076 9388
rect 13036 7160 13076 7188
rect 12940 7120 13036 7160
rect 12940 6572 12980 7120
rect 13036 7111 13076 7120
rect 12940 6404 12980 6532
rect 12940 6355 12980 6364
rect 12556 6271 12596 6280
rect 12556 5732 12596 5741
rect 11884 5515 11924 5524
rect 12460 5648 12500 5657
rect 12460 5513 12500 5608
rect 12556 5480 12596 5692
rect 13036 5732 13076 5741
rect 12748 5648 12788 5657
rect 13036 5648 13076 5692
rect 12788 5608 12980 5648
rect 12748 5599 12788 5608
rect 12940 5480 12980 5608
rect 13036 5597 13076 5608
rect 12556 5440 12788 5480
rect 12748 5396 12788 5440
rect 12940 5431 12980 5440
rect 12748 5347 12788 5356
rect 12126 5312 12494 5321
rect 12126 5263 12494 5272
rect 12748 5228 12788 5237
rect 12076 5060 12116 5069
rect 11980 5020 12076 5060
rect 11980 4976 12020 5020
rect 12076 5011 12116 5020
rect 11980 4927 12020 4936
rect 12556 4976 12596 4985
rect 11884 4892 11924 4901
rect 11884 4472 11924 4852
rect 11884 4423 11924 4432
rect 11308 4136 11348 4145
rect 11308 3968 11348 4096
rect 11308 3919 11348 3928
rect 10732 3583 10772 3592
rect 10636 2827 10676 2836
rect 10732 3464 10772 3473
rect 9388 2659 9428 2668
rect 8908 1952 8948 2584
rect 10156 2372 10196 2381
rect 10156 2036 10196 2332
rect 10732 2120 10772 3424
rect 10886 3044 11254 3053
rect 10886 2995 11254 3004
rect 11500 2624 11540 4180
rect 11596 4388 11636 4397
rect 11596 4136 11636 4348
rect 12556 4220 12596 4936
rect 12748 4388 12788 5188
rect 13036 4892 13076 4901
rect 13036 4472 13076 4852
rect 13132 4724 13172 11572
rect 13228 11477 13268 11572
rect 13516 11696 13556 11992
rect 13516 11528 13556 11656
rect 13324 10940 13364 10949
rect 13324 10688 13364 10900
rect 13516 10856 13556 11488
rect 13612 10982 13652 12244
rect 13612 10933 13652 10942
rect 13516 10807 13556 10816
rect 13324 10639 13364 10648
rect 13612 10604 13652 10613
rect 13228 10352 13268 10361
rect 13268 10312 13460 10352
rect 13228 10303 13268 10312
rect 13324 10184 13364 10193
rect 13228 10016 13268 10025
rect 13228 9512 13268 9976
rect 13228 9463 13268 9472
rect 13228 9344 13268 9353
rect 13228 9176 13268 9304
rect 13228 9127 13268 9136
rect 13228 8924 13268 8933
rect 13228 5648 13268 8884
rect 13228 5060 13268 5608
rect 13228 5011 13268 5020
rect 13132 4675 13172 4684
rect 13228 4808 13268 4817
rect 13036 4423 13076 4432
rect 12748 4339 12788 4348
rect 12556 4171 12596 4180
rect 11596 4087 11636 4096
rect 13228 4136 13268 4768
rect 13228 4087 13268 4096
rect 11884 4052 11924 4061
rect 11884 3548 11924 4012
rect 12556 3968 12596 3977
rect 12126 3800 12494 3809
rect 12126 3751 12494 3760
rect 11884 3499 11924 3508
rect 10732 2071 10772 2080
rect 11308 2456 11348 2465
rect 10156 1987 10196 1996
rect 10636 2036 10676 2045
rect 8908 1903 8948 1912
rect 8428 1315 8468 1324
rect 7564 1147 7604 1156
rect 8524 1112 8564 1121
rect 8524 977 8564 1072
rect 10636 1028 10676 1996
rect 10732 1952 10772 1961
rect 10732 1616 10772 1912
rect 10732 1112 10772 1576
rect 10886 1532 11254 1541
rect 10886 1483 11254 1492
rect 10732 1063 10772 1072
rect 10636 979 10676 988
rect 11308 1028 11348 2416
rect 11500 1868 11540 2584
rect 11788 3464 11828 3473
rect 11500 1819 11540 1828
rect 11596 2372 11636 2381
rect 11596 1112 11636 2332
rect 11788 1952 11828 3424
rect 12172 3464 12212 3473
rect 12172 3128 12212 3424
rect 12172 2624 12212 3088
rect 12460 3464 12500 3473
rect 12460 2708 12500 3424
rect 12460 2659 12500 2668
rect 12172 2575 12212 2584
rect 12556 2624 12596 3928
rect 12556 2575 12596 2584
rect 13036 3632 13076 3641
rect 13036 2540 13076 3592
rect 13324 3632 13364 10144
rect 13420 9260 13460 10312
rect 13516 9596 13556 9605
rect 13516 9260 13556 9556
rect 13612 9596 13652 10564
rect 13612 9512 13652 9556
rect 13612 9461 13652 9472
rect 13612 9260 13652 9269
rect 13516 9220 13612 9260
rect 13420 9211 13460 9220
rect 13612 8756 13652 9220
rect 13708 8924 13748 14680
rect 13804 14552 13844 14561
rect 13804 14417 13844 14512
rect 13804 13796 13844 13805
rect 13804 13376 13844 13756
rect 13804 13327 13844 13336
rect 13804 13040 13844 13049
rect 13804 11948 13844 13000
rect 13804 11024 13844 11908
rect 13900 11948 13940 17620
rect 14476 17576 14516 17585
rect 14476 17441 14516 17536
rect 14380 16988 14420 16997
rect 14284 16904 14324 16913
rect 14188 16484 14228 16493
rect 14092 16064 14132 16073
rect 14092 15560 14132 16024
rect 14188 15896 14228 16444
rect 14188 15847 14228 15856
rect 14092 15511 14132 15520
rect 14188 15644 14228 15653
rect 14092 14804 14132 14813
rect 13996 14720 14036 14729
rect 13996 14585 14036 14680
rect 14092 14300 14132 14764
rect 14188 14636 14228 15604
rect 14188 14587 14228 14596
rect 14092 14251 14132 14260
rect 14188 14048 14228 14057
rect 14092 13292 14132 13301
rect 14092 13124 14132 13252
rect 14092 13075 14132 13084
rect 13996 12620 14036 12629
rect 13996 12485 14036 12580
rect 13900 11899 13940 11908
rect 13996 11864 14036 11873
rect 13900 11780 13940 11789
rect 13900 11192 13940 11740
rect 13900 11143 13940 11152
rect 13804 10975 13844 10984
rect 13900 11024 13940 11033
rect 13900 10604 13940 10984
rect 13996 10940 14036 11824
rect 13996 10891 14036 10900
rect 14092 11696 14132 11705
rect 14188 11696 14228 14008
rect 14284 12452 14324 16864
rect 14380 16484 14420 16948
rect 14572 16988 14612 18964
rect 14860 18584 14900 19300
rect 14860 18535 14900 18544
rect 14764 18332 14804 18341
rect 14764 17072 14804 18292
rect 14572 16939 14612 16948
rect 14668 17032 14764 17072
rect 14380 16435 14420 16444
rect 14380 16148 14420 16157
rect 14380 15476 14420 16108
rect 14572 16148 14612 16157
rect 14476 16064 14516 16073
rect 14476 15929 14516 16024
rect 14380 13460 14420 15436
rect 14572 15560 14612 16108
rect 14572 14720 14612 15520
rect 14572 14671 14612 14680
rect 14668 15392 14708 17032
rect 14764 17023 14804 17032
rect 14860 17576 14900 17585
rect 14764 16904 14804 16913
rect 14764 15728 14804 16864
rect 14764 15560 14804 15688
rect 14764 15511 14804 15520
rect 14668 14720 14708 15352
rect 14668 14671 14708 14680
rect 14764 14804 14804 14813
rect 14380 13411 14420 13420
rect 14572 14300 14612 14309
rect 14572 13796 14612 14260
rect 14764 14216 14804 14764
rect 14764 14167 14804 14176
rect 14380 13208 14420 13217
rect 14380 12788 14420 13168
rect 14380 12739 14420 12748
rect 14476 13124 14516 13133
rect 14476 12620 14516 13084
rect 14572 12704 14612 13756
rect 14668 14048 14708 14057
rect 14668 13040 14708 14008
rect 14764 13796 14804 13805
rect 14764 13376 14804 13756
rect 14764 13327 14804 13336
rect 14668 12991 14708 13000
rect 14764 13208 14804 13217
rect 14764 13040 14804 13168
rect 14572 12655 14612 12664
rect 14476 12571 14516 12580
rect 14572 12536 14612 12545
rect 14284 12412 14420 12452
rect 14284 11696 14324 11791
rect 14188 11656 14284 11696
rect 13900 10555 13940 10564
rect 13996 10772 14036 10781
rect 13900 10184 13940 10193
rect 13900 9512 13940 10144
rect 13900 9463 13940 9472
rect 13708 8875 13748 8884
rect 13612 8707 13652 8716
rect 13996 8588 14036 10732
rect 14092 10268 14132 11656
rect 14284 11647 14324 11656
rect 14380 11528 14420 12412
rect 14284 11488 14420 11528
rect 14476 12032 14516 12041
rect 14476 11528 14516 11992
rect 14284 11192 14324 11488
rect 14476 11479 14516 11488
rect 14572 11780 14612 12496
rect 14764 12116 14804 13000
rect 14764 12067 14804 12076
rect 14572 11192 14612 11740
rect 14284 11143 14324 11152
rect 14476 11152 14612 11192
rect 14668 11948 14708 11957
rect 14284 10940 14324 10949
rect 14284 10352 14324 10900
rect 14092 10219 14132 10228
rect 14188 10312 14324 10352
rect 14188 10016 14228 10312
rect 14188 9967 14228 9976
rect 14380 10100 14420 10109
rect 14284 9932 14324 9941
rect 14284 9512 14324 9892
rect 14284 9463 14324 9472
rect 13996 8539 14036 8548
rect 14380 9260 14420 10060
rect 14380 8504 14420 9220
rect 14380 8455 14420 8464
rect 14092 8000 14132 8009
rect 14092 7865 14132 7960
rect 14284 7664 14324 7673
rect 14284 7244 14324 7624
rect 13420 7076 13460 7085
rect 13420 6320 13460 7036
rect 13900 6488 13940 6528
rect 13420 6271 13460 6280
rect 13516 6404 13556 6413
rect 13420 4976 13460 4985
rect 13420 4388 13460 4936
rect 13420 4339 13460 4348
rect 13324 3583 13364 3592
rect 13420 4136 13460 4145
rect 13228 3464 13268 3473
rect 13036 2491 13076 2500
rect 13132 3296 13172 3305
rect 13132 2624 13172 3256
rect 13228 2876 13268 3424
rect 13420 2900 13460 4096
rect 13228 2827 13268 2836
rect 13324 2860 13460 2900
rect 12126 2288 12494 2297
rect 12126 2239 12494 2248
rect 13132 2120 13172 2584
rect 13132 2071 13172 2080
rect 12364 2036 12404 2045
rect 11788 1280 11828 1912
rect 12172 1952 12212 1961
rect 12172 1817 12212 1912
rect 11788 1231 11828 1240
rect 11596 1063 11636 1072
rect 12364 1112 12404 1996
rect 12364 1063 12404 1072
rect 12556 1952 12596 1961
rect 12556 1364 12596 1912
rect 11308 979 11348 988
rect 6412 811 6452 820
rect 12556 860 12596 1324
rect 12652 1952 12692 1961
rect 13036 1952 13076 1961
rect 12652 1028 12692 1912
rect 12844 1912 13036 1952
rect 12844 1364 12884 1912
rect 13036 1903 13076 1912
rect 13324 1952 13364 2860
rect 12844 1315 12884 1324
rect 13036 1280 13076 1289
rect 12940 1112 12980 1121
rect 13036 1112 13076 1240
rect 13324 1280 13364 1912
rect 13516 1952 13556 6364
rect 13900 6404 13940 6448
rect 14284 6488 14324 7204
rect 14284 6439 14324 6448
rect 13900 4304 13940 6364
rect 14188 6404 14228 6413
rect 14188 6269 14228 6364
rect 14476 5228 14516 11152
rect 14572 10940 14612 10949
rect 14572 10268 14612 10900
rect 14668 10520 14708 11908
rect 14764 11864 14804 11873
rect 14764 11696 14804 11824
rect 14764 11647 14804 11656
rect 14668 10352 14708 10480
rect 14668 10303 14708 10312
rect 14572 10219 14612 10228
rect 14860 10268 14900 17536
rect 14956 16232 14996 19384
rect 15052 19172 15092 20056
rect 15052 19123 15092 19132
rect 15148 20852 15188 20861
rect 15148 19088 15188 20812
rect 15916 20684 15956 20693
rect 15916 20549 15956 20644
rect 15820 20096 15860 20105
rect 15820 19256 15860 20056
rect 15820 19207 15860 19216
rect 15916 20096 15956 20105
rect 15148 16736 15188 19048
rect 15436 19088 15476 19097
rect 15436 17744 15476 19048
rect 15724 19088 15764 19097
rect 15436 17576 15476 17704
rect 15436 17527 15476 17536
rect 15628 17744 15668 17753
rect 15628 17240 15668 17704
rect 15628 17191 15668 17200
rect 15628 17072 15668 17081
rect 15148 16687 15188 16696
rect 15244 16820 15284 16829
rect 14956 15476 14996 16192
rect 15244 15476 15284 16780
rect 14956 15436 15092 15476
rect 14956 15308 14996 15317
rect 14956 11024 14996 15268
rect 15052 14132 15092 15436
rect 15244 15427 15284 15436
rect 15340 14720 15380 14729
rect 15244 14300 15284 14309
rect 15052 14083 15092 14092
rect 15148 14132 15188 14141
rect 14956 10975 14996 10984
rect 15052 13964 15092 13973
rect 14956 10688 14996 10697
rect 14956 10436 14996 10648
rect 14956 10387 14996 10396
rect 14860 9512 14900 10228
rect 14956 10184 14996 10193
rect 14956 9932 14996 10144
rect 14956 9680 14996 9892
rect 14956 9631 14996 9640
rect 14860 9463 14900 9472
rect 14956 9428 14996 9437
rect 14572 8924 14612 8933
rect 14572 8756 14612 8884
rect 14572 8707 14612 8716
rect 14956 8924 14996 9388
rect 14764 8672 14804 8681
rect 14572 5648 14612 5657
rect 14572 5396 14612 5608
rect 14572 5347 14612 5356
rect 14476 5179 14516 5188
rect 13900 4052 13940 4264
rect 13900 4003 13940 4012
rect 13804 3464 13844 3473
rect 13804 2900 13844 3424
rect 13708 2876 13844 2900
rect 13748 2860 13844 2876
rect 14284 3464 14324 3473
rect 13708 2624 13748 2836
rect 13708 2575 13748 2584
rect 14284 2540 14324 3424
rect 14572 3464 14612 3473
rect 14572 3296 14612 3424
rect 14572 3247 14612 3256
rect 14476 3212 14516 3221
rect 14476 2624 14516 3172
rect 14764 2708 14804 8632
rect 14956 8252 14996 8884
rect 15052 8756 15092 13924
rect 15148 12452 15188 14092
rect 15244 14048 15284 14260
rect 15340 14216 15380 14680
rect 15628 14384 15668 17032
rect 15724 14552 15764 19048
rect 15916 18416 15956 20056
rect 15916 18367 15956 18376
rect 16012 16736 16052 23080
rect 16396 23060 16436 28624
rect 23096 28600 23176 29000
rect 23864 28600 23944 29000
rect 24632 28600 24712 29000
rect 25400 28600 25480 29000
rect 26168 28600 26248 29000
rect 26936 28600 27016 29000
rect 27704 28600 27784 29000
rect 28472 28600 28552 29000
rect 29240 28600 29320 29000
rect 30008 28600 30088 29000
rect 30776 28600 30856 29000
rect 17644 28412 17684 28421
rect 17068 27656 17108 27665
rect 16780 27572 16820 27581
rect 16780 26900 16820 27532
rect 17068 27068 17108 27616
rect 17068 27019 17108 27028
rect 17644 26900 17684 28372
rect 20428 28244 20468 28253
rect 19900 27992 20268 28001
rect 19900 27943 20268 27952
rect 17836 27824 17876 27833
rect 17740 27572 17780 27581
rect 17740 27068 17780 27532
rect 17740 27019 17780 27028
rect 17644 26860 17780 26900
rect 16780 26851 16820 26860
rect 17068 26816 17108 26825
rect 16972 26396 17012 26405
rect 16588 26144 16628 26153
rect 16492 25976 16532 25985
rect 16492 25304 16532 25936
rect 16492 25255 16532 25264
rect 16588 25220 16628 26104
rect 16588 25171 16628 25180
rect 16972 24632 17012 26356
rect 17068 26396 17108 26776
rect 17164 26396 17204 26424
rect 17068 26356 17164 26396
rect 17068 25724 17108 26356
rect 17164 26347 17204 26356
rect 17452 26312 17492 26321
rect 17068 25675 17108 25684
rect 17356 26228 17396 26237
rect 17356 25640 17396 26188
rect 17356 25591 17396 25600
rect 17452 25388 17492 26272
rect 17356 25304 17396 25313
rect 17452 25304 17492 25348
rect 17396 25264 17492 25304
rect 17356 25255 17396 25264
rect 16972 24296 17012 24592
rect 17356 25052 17396 25061
rect 16300 23020 16436 23060
rect 16588 23288 16628 23297
rect 16108 22280 16148 22289
rect 16108 21608 16148 22240
rect 16108 21559 16148 21568
rect 16108 21020 16148 21029
rect 16108 20684 16148 20980
rect 16108 19088 16148 20644
rect 16108 19039 16148 19048
rect 16108 18500 16148 18509
rect 16108 18365 16148 18460
rect 16204 17744 16244 17753
rect 15820 16232 15860 16241
rect 15820 16097 15860 16192
rect 15916 15560 15956 15569
rect 15820 15520 15916 15560
rect 15820 15392 15860 15520
rect 15916 15511 15956 15520
rect 15820 15343 15860 15352
rect 15820 15140 15860 15149
rect 15820 14720 15860 15100
rect 15820 14671 15860 14680
rect 15724 14503 15764 14512
rect 15916 14636 15956 14645
rect 15628 14344 15860 14384
rect 15340 14167 15380 14176
rect 15244 13999 15284 14008
rect 15340 13964 15380 13973
rect 15244 13376 15284 13385
rect 15244 13292 15284 13336
rect 15244 13241 15284 13252
rect 15244 13040 15284 13049
rect 15244 12536 15284 13000
rect 15340 12872 15380 13924
rect 15724 13544 15764 13553
rect 15532 13460 15572 13469
rect 15532 13292 15572 13420
rect 15532 13208 15572 13252
rect 15340 12823 15380 12832
rect 15436 12956 15476 12965
rect 15244 12487 15284 12496
rect 15340 12536 15380 12545
rect 15148 11780 15188 12412
rect 15148 11108 15188 11740
rect 15244 11864 15284 11873
rect 15244 11612 15284 11824
rect 15244 11563 15284 11572
rect 15340 11780 15380 12496
rect 15340 11276 15380 11740
rect 15436 12116 15476 12916
rect 15436 11696 15476 12076
rect 15436 11647 15476 11656
rect 15532 11612 15572 13168
rect 15628 13292 15668 13303
rect 15628 13208 15668 13252
rect 15628 13159 15668 13168
rect 15724 13208 15764 13504
rect 15724 13159 15764 13168
rect 15820 13040 15860 14344
rect 15532 11563 15572 11572
rect 15628 13000 15860 13040
rect 15340 11227 15380 11236
rect 15436 11528 15476 11537
rect 15148 11059 15188 11068
rect 15244 11024 15284 11033
rect 15244 10889 15284 10984
rect 15340 10940 15380 10949
rect 15340 10268 15380 10900
rect 15436 10856 15476 11488
rect 15436 10807 15476 10816
rect 15340 10219 15380 10228
rect 15532 10184 15572 10279
rect 15532 10135 15572 10144
rect 15052 8707 15092 8716
rect 15436 9512 15476 9521
rect 15628 9512 15668 13000
rect 15724 12200 15764 12209
rect 15724 11780 15764 12160
rect 15724 11731 15764 11740
rect 15820 11696 15860 11705
rect 15820 11192 15860 11656
rect 15916 11444 15956 14596
rect 16012 14552 16052 16696
rect 16108 16988 16148 16997
rect 16108 16232 16148 16948
rect 16108 16183 16148 16192
rect 16108 16064 16148 16073
rect 16108 14804 16148 16024
rect 16108 14755 16148 14764
rect 16012 14503 16052 14512
rect 16108 14636 16148 14645
rect 16012 13208 16052 13217
rect 16108 13208 16148 14596
rect 16204 14216 16244 17704
rect 16300 15140 16340 23020
rect 16492 21524 16532 21533
rect 16396 21356 16436 21365
rect 16396 21188 16436 21316
rect 16396 20768 16436 21148
rect 16492 20852 16532 21484
rect 16588 20936 16628 23248
rect 16972 23120 17012 24256
rect 17164 24464 17204 24473
rect 17164 23876 17204 24424
rect 17164 23827 17204 23836
rect 16972 23071 17012 23080
rect 17356 23120 17396 25012
rect 17452 24632 17492 25264
rect 17548 25976 17588 25985
rect 17548 25304 17588 25936
rect 17548 24800 17588 25264
rect 17548 24751 17588 24760
rect 17644 25136 17684 25145
rect 17452 24583 17492 24592
rect 17356 23071 17396 23080
rect 17644 23120 17684 25096
rect 17644 23071 17684 23080
rect 16588 20887 16628 20896
rect 16780 22868 16820 22877
rect 16492 20803 16532 20812
rect 16396 20719 16436 20728
rect 16396 20096 16436 20105
rect 16396 19508 16436 20056
rect 16396 19459 16436 19468
rect 16588 20096 16628 20105
rect 16492 18500 16532 18509
rect 16492 17744 16532 18460
rect 16492 17695 16532 17704
rect 16396 16904 16436 16913
rect 16396 15476 16436 16864
rect 16588 16484 16628 20056
rect 16684 19088 16724 19097
rect 16684 18752 16724 19048
rect 16684 18703 16724 18712
rect 16684 18584 16724 18593
rect 16684 18449 16724 18544
rect 16684 17744 16724 17753
rect 16684 16904 16724 17704
rect 16684 16855 16724 16864
rect 16588 16435 16628 16444
rect 16492 16232 16532 16241
rect 16492 15728 16532 16192
rect 16780 16064 16820 22828
rect 17644 22196 17684 22205
rect 17644 21608 17684 22156
rect 17740 21776 17780 26860
rect 17740 21727 17780 21736
rect 17836 21692 17876 27784
rect 19084 27656 19124 27665
rect 18660 27236 19028 27245
rect 18660 27187 19028 27196
rect 18124 27152 18164 27161
rect 18124 26312 18164 27112
rect 18028 26144 18068 26153
rect 18124 26144 18164 26272
rect 18068 26104 18164 26144
rect 18892 26396 18932 26405
rect 18892 26144 18932 26356
rect 18028 26095 18068 26104
rect 18892 26095 18932 26104
rect 18028 25976 18068 25985
rect 17932 25808 17972 25817
rect 17932 25220 17972 25768
rect 17932 25171 17972 25180
rect 18028 24716 18068 25936
rect 18660 25724 19028 25733
rect 18660 25675 19028 25684
rect 18700 25388 18740 25397
rect 18700 25304 18740 25348
rect 18700 25253 18740 25264
rect 18892 25304 18932 25399
rect 18892 25255 18932 25264
rect 18124 25220 18164 25229
rect 18124 24800 18164 25180
rect 18892 25136 18932 25145
rect 18124 24751 18164 24760
rect 18220 25052 18260 25061
rect 18028 24667 18068 24676
rect 18220 24716 18260 25012
rect 18892 24800 18932 25096
rect 18892 24751 18932 24760
rect 18220 24667 18260 24676
rect 18988 24716 19028 24725
rect 19084 24716 19124 27616
rect 20140 27656 20180 27665
rect 19660 27404 19700 27413
rect 19660 26900 19700 27364
rect 19276 26396 19316 26405
rect 19180 25808 19220 25817
rect 19180 25673 19220 25768
rect 19276 25220 19316 26356
rect 19564 26312 19604 26321
rect 19468 26144 19508 26153
rect 19276 25171 19316 25180
rect 19372 25892 19412 25901
rect 19028 24676 19124 24716
rect 18988 24667 19028 24676
rect 18412 24632 18452 24641
rect 18412 24044 18452 24592
rect 19084 24592 19316 24632
rect 19084 24548 19124 24592
rect 19084 24499 19124 24508
rect 19180 24464 19220 24473
rect 19084 24380 19124 24389
rect 18660 24212 19028 24221
rect 18660 24163 19028 24172
rect 18412 23995 18452 24004
rect 18892 23960 18932 23969
rect 17932 23792 17972 23801
rect 17932 23624 17972 23752
rect 17932 23288 17972 23584
rect 17932 23239 17972 23248
rect 18412 23792 18452 23801
rect 17932 23120 17972 23129
rect 17932 22952 17972 23080
rect 18412 23120 18452 23752
rect 18892 23204 18932 23920
rect 19084 23960 19124 24340
rect 19084 23911 19124 23920
rect 18892 23155 18932 23164
rect 18988 23792 19028 23801
rect 18988 23120 19028 23752
rect 18452 23080 18548 23120
rect 18412 23071 18452 23080
rect 17932 22912 18452 22952
rect 17836 21652 17972 21692
rect 17068 21524 17108 21533
rect 17068 20264 17108 21484
rect 17548 21524 17588 21533
rect 17068 20215 17108 20224
rect 17260 20852 17300 20861
rect 17260 20264 17300 20812
rect 17548 20852 17588 21484
rect 17548 20803 17588 20812
rect 17644 20684 17684 21568
rect 17644 20635 17684 20644
rect 17836 21524 17876 21533
rect 17260 20215 17300 20224
rect 17836 20264 17876 21484
rect 17932 20768 17972 21652
rect 17932 20719 17972 20728
rect 17836 20215 17876 20224
rect 17107 20105 17147 20152
rect 17068 20096 17147 20105
rect 17068 20047 17147 20056
rect 17452 20096 17492 20105
rect 17356 20012 17396 20021
rect 17260 19928 17300 19937
rect 16972 19676 17012 19685
rect 16876 19172 16916 19181
rect 16876 19037 16916 19132
rect 16876 18668 16916 18677
rect 16972 18668 17012 19636
rect 17260 19340 17300 19888
rect 17356 19508 17396 19972
rect 17356 19459 17396 19468
rect 17452 19760 17492 20056
rect 18124 20096 18164 20105
rect 18124 19961 18164 20056
rect 17260 19291 17300 19300
rect 17164 19172 17204 19181
rect 17164 18668 17204 19132
rect 17356 19172 17396 19181
rect 17356 19037 17396 19132
rect 17452 19088 17492 19720
rect 17644 19844 17684 19853
rect 17644 19508 17684 19804
rect 17644 19459 17684 19468
rect 17548 19256 17588 19265
rect 17548 19121 17588 19216
rect 18220 19256 18260 19265
rect 17452 19039 17492 19048
rect 17644 19088 17684 19097
rect 16972 18628 17108 18668
rect 17164 18628 17300 18668
rect 16876 18500 16916 18628
rect 16876 18451 16916 18460
rect 17068 18500 17108 18628
rect 17068 18451 17108 18460
rect 17164 18500 17204 18509
rect 16972 18416 17012 18425
rect 16876 17240 16916 17249
rect 16876 16988 16916 17200
rect 16876 16939 16916 16948
rect 16780 16015 16820 16024
rect 16876 16232 16916 16241
rect 16492 15679 16532 15688
rect 16876 15728 16916 16192
rect 16876 15679 16916 15688
rect 16396 15427 16436 15436
rect 16588 15644 16628 15653
rect 16300 15091 16340 15100
rect 16588 15392 16628 15604
rect 16492 14804 16532 14813
rect 16204 14167 16244 14176
rect 16396 14720 16436 14729
rect 16300 13880 16340 13889
rect 16300 13460 16340 13840
rect 16300 13411 16340 13420
rect 16052 13168 16148 13208
rect 16300 13208 16340 13217
rect 16012 11696 16052 13168
rect 16204 12788 16244 12797
rect 16108 12032 16148 12041
rect 16108 11864 16148 11992
rect 16204 11948 16244 12748
rect 16204 11899 16244 11908
rect 16108 11815 16148 11824
rect 16300 11696 16340 13168
rect 16396 11864 16436 14680
rect 16492 12536 16532 14764
rect 16588 14552 16628 15352
rect 16588 14503 16628 14512
rect 16684 15308 16724 15317
rect 16588 13208 16628 13217
rect 16588 12620 16628 13168
rect 16588 12571 16628 12580
rect 16492 12116 16532 12496
rect 16492 12067 16532 12076
rect 16588 12284 16628 12293
rect 16396 11815 16436 11824
rect 16492 11948 16532 11957
rect 16012 11656 16244 11696
rect 15916 11395 15956 11404
rect 16012 11528 16052 11537
rect 15820 11143 15860 11152
rect 16012 10856 16052 11488
rect 16108 11276 16148 11285
rect 16108 11108 16148 11236
rect 16108 11059 16148 11068
rect 16012 10807 16052 10816
rect 16108 10772 16148 10781
rect 15820 10436 15860 10445
rect 15820 10268 15860 10396
rect 16108 10352 16148 10732
rect 16108 10303 16148 10312
rect 15820 10219 15860 10228
rect 15476 9472 15668 9512
rect 15724 10184 15764 10193
rect 15436 8672 15476 9472
rect 15724 9344 15764 10144
rect 16108 10184 16148 10193
rect 15820 10016 15860 10025
rect 15820 9512 15860 9976
rect 16108 9932 16148 10144
rect 15820 9377 15860 9472
rect 16012 9764 16052 9773
rect 15724 9295 15764 9304
rect 15436 8623 15476 8632
rect 15724 8756 15764 8765
rect 14956 8203 14996 8212
rect 15628 8000 15668 8009
rect 15148 7916 15188 7925
rect 14956 7748 14996 7757
rect 14860 7076 14900 7085
rect 14860 6404 14900 7036
rect 14956 6488 14996 7708
rect 15148 7160 15188 7876
rect 15148 6656 15188 7120
rect 15148 6607 15188 6616
rect 15340 7916 15380 7925
rect 15340 6572 15380 7876
rect 15340 6523 15380 6532
rect 15628 7160 15668 7960
rect 15724 7412 15764 8716
rect 16012 8504 16052 9724
rect 16012 8455 16052 8464
rect 16108 9512 16148 9892
rect 16108 8756 16148 9472
rect 16108 8000 16148 8716
rect 16108 7951 16148 7960
rect 15724 7363 15764 7372
rect 14956 6439 14996 6448
rect 14860 6355 14900 6364
rect 14860 5648 14900 5657
rect 14860 5513 14900 5608
rect 15628 5312 15668 7120
rect 16204 6656 16244 11656
rect 16300 11024 16340 11656
rect 16396 11612 16436 11621
rect 16396 11477 16436 11572
rect 16396 11360 16436 11369
rect 16396 11225 16436 11320
rect 16300 10975 16340 10984
rect 16396 10856 16436 10865
rect 16396 10268 16436 10816
rect 16396 10219 16436 10228
rect 16204 6607 16244 6616
rect 16300 8588 16340 8597
rect 16108 6236 16148 6245
rect 16108 5564 16148 6196
rect 16108 5515 16148 5524
rect 15628 5263 15668 5272
rect 15820 4976 15860 4985
rect 15052 4304 15092 4313
rect 15052 3464 15092 4264
rect 15052 3415 15092 3424
rect 15820 3464 15860 4936
rect 16012 4976 16052 4985
rect 14764 2659 14804 2668
rect 14860 3128 14900 3137
rect 14476 2575 14516 2584
rect 14860 2624 14900 3088
rect 14860 2575 14900 2584
rect 13804 2288 13844 2297
rect 13804 2120 13844 2248
rect 13804 2071 13844 2080
rect 14284 2120 14324 2500
rect 14284 2071 14324 2080
rect 15820 2120 15860 3424
rect 15916 4892 15956 4901
rect 15916 3968 15956 4852
rect 16012 4136 16052 4936
rect 16012 4087 16052 4096
rect 15916 2792 15956 3928
rect 16300 2900 16340 8548
rect 16492 6572 16532 11908
rect 16588 11864 16628 12244
rect 16588 11815 16628 11824
rect 16588 11696 16628 11705
rect 16588 11561 16628 11656
rect 16684 11192 16724 15268
rect 16876 14636 16916 14645
rect 16780 13964 16820 13973
rect 16780 11948 16820 13924
rect 16876 13712 16916 14596
rect 16876 12620 16916 13672
rect 16972 13544 17012 18376
rect 17164 15644 17204 18460
rect 17260 18332 17300 18628
rect 17548 18584 17588 18595
rect 17356 18500 17396 18509
rect 17356 18365 17396 18460
rect 17548 18500 17588 18544
rect 17548 18451 17588 18460
rect 17260 18283 17300 18292
rect 17548 17744 17588 17753
rect 17164 15595 17204 15604
rect 17260 17660 17300 17669
rect 17164 14804 17204 14813
rect 17164 14720 17204 14764
rect 17164 14669 17204 14680
rect 17164 13796 17204 13805
rect 16972 13504 17108 13544
rect 16972 13292 17012 13301
rect 16972 12872 17012 13252
rect 16972 12823 17012 12832
rect 16876 12571 16916 12580
rect 16780 11899 16820 11908
rect 16684 11143 16724 11152
rect 16780 11444 16820 11453
rect 16492 6523 16532 6532
rect 16588 10184 16628 10193
rect 16396 6488 16436 6497
rect 16396 6320 16436 6448
rect 16396 6271 16436 6280
rect 16492 6404 16532 6413
rect 16492 5900 16532 6364
rect 16492 5851 16532 5860
rect 16396 5732 16436 5741
rect 16396 4388 16436 5692
rect 16396 4339 16436 4348
rect 16492 5228 16532 5237
rect 16492 4136 16532 5188
rect 16588 5060 16628 10144
rect 16684 8924 16724 8933
rect 16684 8789 16724 8884
rect 16684 8672 16724 8681
rect 16684 8168 16724 8632
rect 16780 8504 16820 11404
rect 16876 11192 16916 11201
rect 16876 10352 16916 11152
rect 16876 10303 16916 10312
rect 16972 10940 17012 10949
rect 16876 10100 16916 10109
rect 16876 8756 16916 10060
rect 16876 8707 16916 8716
rect 16780 8455 16820 8464
rect 16876 8588 16916 8597
rect 16684 8119 16724 8128
rect 16876 8168 16916 8548
rect 16876 8119 16916 8128
rect 16972 6656 17012 10900
rect 17068 8420 17108 13504
rect 17164 13292 17204 13756
rect 17260 13544 17300 17620
rect 17356 16904 17396 16913
rect 17356 15812 17396 16864
rect 17548 16820 17588 17704
rect 17548 16232 17588 16780
rect 17548 16097 17588 16192
rect 17356 15728 17396 15772
rect 17356 15677 17396 15688
rect 17356 15560 17396 15569
rect 17356 15056 17396 15520
rect 17644 15308 17684 19048
rect 17932 18752 17972 18761
rect 17836 18584 17876 18593
rect 17836 17660 17876 18544
rect 17932 18500 17972 18712
rect 18220 18752 18260 19216
rect 18220 18703 18260 18712
rect 18124 18584 18164 18593
rect 17932 18451 17972 18460
rect 18028 18500 18068 18509
rect 17876 17620 17972 17660
rect 17836 17611 17876 17620
rect 17932 17240 17972 17620
rect 18028 17576 18068 18460
rect 18124 17828 18164 18544
rect 18316 18500 18356 18509
rect 18220 18416 18260 18425
rect 18220 17996 18260 18376
rect 18220 17947 18260 17956
rect 18124 17788 18260 17828
rect 18220 17744 18260 17788
rect 18220 17695 18260 17704
rect 18028 17441 18068 17536
rect 18124 17660 18164 17669
rect 17932 17191 17972 17200
rect 17836 17156 17876 17165
rect 17740 16988 17780 16997
rect 17740 16853 17780 16948
rect 17836 16736 17876 17116
rect 18028 17156 18068 17165
rect 18124 17156 18164 17620
rect 18068 17116 18164 17156
rect 18028 17107 18068 17116
rect 17932 16904 17972 16913
rect 17932 16769 17972 16864
rect 18028 16820 18068 16829
rect 17740 16696 17876 16736
rect 17740 16484 17780 16696
rect 17740 16435 17780 16444
rect 18028 16484 18068 16780
rect 18028 16435 18068 16444
rect 18124 16232 18164 17116
rect 18220 17240 18260 17249
rect 18220 17156 18260 17200
rect 18220 17105 18260 17116
rect 17836 15772 18068 15812
rect 17644 15259 17684 15268
rect 17740 15560 17780 15569
rect 17356 15007 17396 15016
rect 17260 13495 17300 13504
rect 17452 14804 17492 14813
rect 17644 14804 17684 14813
rect 17452 13460 17492 14764
rect 17548 14764 17644 14804
rect 17548 13964 17588 14764
rect 17644 14755 17684 14764
rect 17548 13915 17588 13924
rect 17644 14636 17684 14645
rect 17644 14132 17684 14596
rect 17740 14552 17780 15520
rect 17836 14972 17876 15772
rect 18028 15728 18068 15772
rect 18028 15679 18068 15688
rect 17836 14923 17876 14932
rect 18028 15560 18068 15569
rect 17740 14503 17780 14512
rect 17836 14720 17876 14729
rect 17452 13411 17492 13420
rect 17164 13243 17204 13252
rect 17356 13292 17396 13301
rect 17164 12872 17204 12881
rect 17164 12536 17204 12832
rect 17164 12487 17204 12496
rect 17356 11612 17396 13252
rect 17356 11563 17396 11572
rect 17452 13124 17492 13133
rect 17452 11696 17492 13084
rect 17260 11276 17300 11285
rect 17164 11024 17204 11033
rect 17164 10100 17204 10984
rect 17260 10436 17300 11236
rect 17260 10387 17300 10396
rect 17356 11024 17396 11033
rect 17164 10051 17204 10060
rect 17260 9932 17300 9941
rect 17068 8371 17108 8380
rect 17164 9680 17204 9689
rect 17164 8588 17204 9640
rect 17260 9428 17300 9892
rect 17260 9379 17300 9388
rect 17068 8000 17108 8009
rect 17068 7496 17108 7960
rect 17068 7447 17108 7456
rect 16972 6607 17012 6616
rect 16588 5011 16628 5020
rect 16684 6572 16724 6581
rect 16684 5648 16724 6532
rect 16780 6320 16820 6329
rect 16780 5732 16820 6280
rect 16780 5683 16820 5692
rect 16492 3464 16532 4096
rect 16684 4136 16724 5608
rect 16780 4976 16820 4985
rect 17164 4976 17204 8548
rect 16780 4841 16820 4936
rect 17068 4936 17164 4976
rect 17068 4724 17108 4936
rect 17164 4927 17204 4936
rect 17260 9260 17300 9269
rect 17260 4808 17300 9220
rect 17356 8168 17396 10984
rect 17452 10268 17492 11656
rect 17644 11696 17684 14092
rect 17740 14048 17780 14057
rect 17740 13376 17780 14008
rect 17836 13544 17876 14680
rect 17932 14552 17972 14561
rect 17932 14417 17972 14512
rect 17836 13495 17876 13504
rect 17932 13880 17972 13889
rect 17740 13327 17780 13336
rect 17932 13292 17972 13840
rect 17836 13208 17876 13217
rect 17644 11108 17684 11656
rect 17644 11059 17684 11068
rect 17740 13124 17780 13133
rect 17740 11780 17780 13084
rect 17836 12704 17876 13168
rect 17836 12655 17876 12664
rect 17644 10940 17684 10949
rect 17644 10688 17684 10900
rect 17548 10436 17588 10445
rect 17548 10352 17588 10396
rect 17548 10301 17588 10312
rect 17452 10219 17492 10228
rect 17644 10184 17684 10648
rect 17644 10135 17684 10144
rect 17548 10016 17588 10025
rect 17452 9848 17492 9857
rect 17452 9512 17492 9808
rect 17452 9463 17492 9472
rect 17548 8840 17588 9976
rect 17644 9428 17684 9437
rect 17644 9293 17684 9388
rect 17548 8791 17588 8800
rect 17356 8119 17396 8128
rect 17740 6572 17780 11740
rect 17932 11024 17972 13252
rect 17932 10975 17972 10984
rect 17836 10940 17876 10949
rect 17836 10805 17876 10900
rect 17932 10772 17972 10781
rect 17836 10352 17876 10361
rect 17836 10100 17876 10312
rect 17836 10051 17876 10060
rect 17836 9512 17876 9521
rect 17836 8504 17876 9472
rect 17836 8455 17876 8464
rect 17932 8336 17972 10732
rect 18028 8756 18068 15520
rect 18124 13040 18164 16192
rect 18220 16232 18260 16241
rect 18220 15644 18260 16192
rect 18220 15595 18260 15604
rect 18316 15560 18356 18460
rect 18316 15476 18356 15520
rect 18316 15425 18356 15436
rect 18220 14300 18260 14309
rect 18220 13292 18260 14260
rect 18220 13124 18260 13252
rect 18316 13544 18356 13553
rect 18316 13208 18356 13504
rect 18316 13159 18356 13168
rect 18220 13075 18260 13084
rect 18124 12991 18164 13000
rect 18412 12980 18452 22912
rect 18508 22532 18548 23080
rect 18988 23071 19028 23080
rect 19084 23624 19124 23633
rect 18660 22700 19028 22709
rect 18660 22651 19028 22660
rect 18604 22532 18644 22541
rect 18508 22492 18604 22532
rect 18604 22112 18644 22492
rect 19084 22364 19124 23584
rect 19084 22315 19124 22324
rect 19180 23120 19220 24424
rect 19276 24044 19316 24592
rect 19372 24548 19412 25852
rect 19468 25304 19508 26104
rect 19564 25556 19604 26272
rect 19564 25507 19604 25516
rect 19468 25255 19508 25264
rect 19372 24499 19412 24508
rect 19660 24464 19700 26860
rect 20140 26816 20180 27616
rect 20140 26767 20180 26776
rect 19900 26480 20268 26489
rect 19900 26431 20268 26440
rect 19948 26312 19988 26321
rect 19948 26144 19988 26272
rect 19948 26095 19988 26104
rect 19852 25976 19892 25985
rect 19756 25556 19796 25565
rect 19756 24632 19796 25516
rect 19852 25472 19892 25936
rect 19852 25304 19892 25432
rect 19852 25255 19892 25264
rect 20140 25892 20180 25901
rect 20140 25304 20180 25852
rect 20140 25255 20180 25264
rect 20332 25556 20372 25565
rect 19900 24968 20268 24977
rect 19900 24919 20268 24928
rect 20332 24884 20372 25516
rect 20332 24835 20372 24844
rect 19756 24583 19796 24592
rect 20236 24800 20276 24809
rect 20236 24632 20276 24760
rect 20236 24583 20276 24592
rect 19660 24424 19796 24464
rect 19276 23995 19316 24004
rect 19468 23960 19508 23969
rect 19180 22280 19220 23080
rect 19276 23204 19316 23213
rect 19276 22448 19316 23164
rect 19372 23036 19412 23045
rect 19372 22532 19412 22996
rect 19372 22483 19412 22492
rect 19276 22399 19316 22408
rect 19180 22231 19220 22240
rect 18604 22063 18644 22072
rect 18988 22196 19028 22205
rect 18988 21608 19028 22156
rect 19468 21776 19508 23920
rect 19660 23792 19700 23801
rect 18988 21559 19028 21568
rect 19084 21736 19508 21776
rect 19564 22868 19604 22877
rect 18660 21188 19028 21197
rect 18660 21139 19028 21148
rect 18988 20684 19028 20693
rect 18988 20180 19028 20644
rect 18988 20131 19028 20140
rect 18508 20096 18548 20105
rect 18508 19340 18548 20056
rect 18660 19676 19028 19685
rect 18660 19627 19028 19636
rect 18508 18416 18548 19300
rect 18988 19172 19028 19181
rect 18988 18584 19028 19132
rect 18988 18449 19028 18544
rect 18508 18367 18548 18376
rect 18660 18164 19028 18173
rect 18660 18115 19028 18124
rect 18660 16652 19028 16661
rect 18660 16603 19028 16612
rect 18796 16484 18836 16493
rect 18508 16316 18548 16325
rect 18508 13208 18548 16276
rect 18796 15896 18836 16444
rect 18796 15847 18836 15856
rect 19084 15560 19124 21736
rect 19276 21608 19316 21617
rect 19180 21356 19220 21365
rect 19180 20348 19220 21316
rect 19276 20852 19316 21568
rect 19276 20803 19316 20812
rect 19180 20299 19220 20308
rect 19276 20096 19316 20105
rect 19084 15511 19124 15520
rect 19180 19256 19220 19265
rect 18700 15392 18740 15403
rect 18700 15308 18740 15352
rect 18700 15259 18740 15268
rect 18660 15140 19028 15149
rect 18660 15091 19028 15100
rect 18700 14972 18740 14981
rect 18604 14804 18644 14899
rect 18604 14755 18644 14764
rect 18700 14720 18740 14932
rect 18604 14636 18644 14647
rect 18604 14552 18644 14596
rect 18700 14585 18740 14680
rect 18892 14720 18932 14729
rect 18604 14503 18644 14512
rect 18892 14216 18932 14680
rect 18892 14167 18932 14176
rect 19084 14636 19124 14645
rect 18796 14132 18836 14141
rect 18796 14048 18836 14092
rect 18796 13997 18836 14008
rect 18660 13628 19028 13637
rect 18660 13579 19028 13588
rect 18548 13168 18644 13208
rect 18508 13159 18548 13168
rect 18316 12940 18452 12980
rect 18508 13040 18548 13049
rect 18124 12788 18164 12797
rect 18124 12653 18164 12748
rect 18124 11780 18164 11789
rect 18124 11696 18164 11740
rect 18124 11645 18164 11656
rect 18220 11612 18260 11621
rect 18124 10100 18164 10109
rect 18124 8924 18164 10060
rect 18124 8840 18164 8884
rect 18124 8789 18164 8800
rect 18028 8707 18068 8716
rect 17932 8084 17972 8296
rect 17932 8035 17972 8044
rect 18124 8168 18164 8177
rect 17932 7160 17972 7171
rect 17932 7076 17972 7120
rect 18124 7160 18164 8128
rect 18220 8000 18260 11572
rect 18316 9680 18356 12940
rect 18316 9631 18356 9640
rect 18412 12704 18452 12713
rect 18316 9428 18356 9437
rect 18316 8693 18356 9388
rect 18316 8644 18356 8653
rect 18316 8588 18356 8597
rect 18316 8084 18356 8548
rect 18412 8252 18452 12664
rect 18508 12284 18548 13000
rect 18604 12620 18644 13168
rect 18892 13124 18932 13133
rect 19084 13124 19124 14596
rect 18932 13084 19124 13124
rect 18892 13075 18932 13084
rect 18604 12571 18644 12580
rect 18508 12235 18548 12244
rect 18660 12116 19028 12125
rect 18660 12067 19028 12076
rect 18604 11948 18644 11957
rect 18604 10772 18644 11908
rect 19084 11276 19124 13084
rect 19180 12704 19220 19216
rect 19276 19088 19316 20056
rect 19468 19844 19508 19853
rect 19468 19256 19508 19804
rect 19276 19039 19316 19048
rect 19372 19172 19412 19181
rect 19372 18752 19412 19132
rect 19372 18703 19412 18712
rect 19468 18668 19508 19216
rect 19468 18584 19508 18628
rect 19276 18500 19316 18511
rect 19468 18504 19508 18544
rect 19276 18416 19316 18460
rect 19564 18416 19604 22828
rect 19660 22196 19700 23752
rect 19756 22448 19796 24424
rect 20332 23708 20372 23717
rect 19900 23456 20268 23465
rect 19900 23407 20268 23416
rect 20332 23288 20372 23668
rect 20332 23120 20372 23248
rect 20332 23071 20372 23080
rect 20428 23456 20468 28204
rect 21388 28160 21428 28169
rect 20524 28076 20564 28085
rect 20524 25136 20564 28036
rect 21100 27908 21140 27917
rect 20812 27488 20852 27497
rect 20716 27068 20756 27077
rect 20716 26144 20756 27028
rect 20812 26900 20852 27448
rect 20812 26851 20852 26860
rect 20908 27320 20948 27329
rect 20716 26095 20756 26104
rect 20620 26060 20660 26069
rect 20620 25304 20660 26020
rect 20620 25255 20660 25264
rect 20812 26060 20852 26069
rect 20908 26060 20948 27280
rect 20852 26020 20948 26060
rect 21004 26144 21044 26153
rect 20524 25096 20756 25136
rect 20428 23060 20468 23416
rect 20428 23020 20564 23060
rect 19756 22399 19796 22408
rect 20332 22868 20372 22877
rect 19660 22147 19700 22156
rect 19900 21944 20268 21953
rect 19900 21895 20268 21904
rect 19852 21692 19892 21701
rect 19756 21440 19796 21449
rect 19756 20096 19796 21400
rect 19852 20768 19892 21652
rect 20140 21692 20180 21701
rect 19852 20719 19892 20728
rect 19948 21608 19988 21617
rect 19948 20684 19988 21568
rect 20140 20852 20180 21652
rect 20140 20803 20180 20812
rect 19948 20635 19988 20644
rect 19900 20432 20268 20441
rect 19900 20383 20268 20392
rect 19852 20096 19892 20105
rect 19756 20056 19852 20096
rect 19852 20047 19892 20056
rect 20236 20012 20276 20021
rect 19660 19928 19700 19937
rect 19660 19424 19700 19888
rect 20236 19844 20276 19972
rect 20236 19795 20276 19804
rect 19660 18500 19700 19384
rect 19660 18451 19700 18460
rect 19756 19340 19796 19349
rect 19276 18367 19316 18376
rect 19468 18376 19604 18416
rect 19372 18332 19412 18341
rect 19276 17492 19316 17501
rect 19276 17072 19316 17452
rect 19276 17023 19316 17032
rect 19276 16904 19316 16913
rect 19276 16769 19316 16864
rect 19276 16652 19316 16661
rect 19276 16316 19316 16612
rect 19276 16267 19316 16276
rect 19180 12655 19220 12664
rect 19276 15896 19316 15905
rect 19180 11528 19220 11537
rect 19180 11393 19220 11488
rect 19084 11236 19220 11276
rect 19084 11024 19124 11033
rect 18892 10940 18932 10949
rect 18892 10805 18932 10900
rect 18508 10732 18644 10772
rect 18508 10016 18548 10732
rect 18660 10604 19028 10613
rect 18660 10555 19028 10564
rect 19084 10352 19124 10984
rect 19180 10940 19220 11236
rect 19180 10772 19220 10900
rect 19180 10723 19220 10732
rect 19084 10303 19124 10312
rect 18604 10184 18644 10193
rect 19003 10184 19043 10193
rect 18644 10144 19003 10184
rect 18604 10135 18644 10144
rect 18508 9680 18548 9976
rect 18508 9631 18548 9640
rect 18700 9596 18740 10144
rect 19003 10135 19043 10144
rect 18700 9344 18740 9556
rect 19276 9512 19316 15856
rect 19372 9680 19412 18292
rect 19372 9631 19412 9640
rect 19276 9463 19316 9472
rect 18700 9295 18740 9304
rect 19180 9428 19220 9437
rect 18660 9092 19028 9101
rect 18660 9043 19028 9052
rect 18412 8203 18452 8212
rect 18508 8756 18548 8765
rect 18316 8044 18452 8084
rect 18412 8000 18452 8044
rect 18220 7960 18356 8000
rect 18124 7111 18164 7120
rect 18220 7832 18260 7841
rect 17932 7027 17972 7036
rect 17548 6532 17780 6572
rect 17932 6908 17972 6917
rect 17932 6572 17972 6868
rect 18220 6740 18260 7792
rect 18220 6691 18260 6700
rect 17548 6488 17588 6532
rect 17932 6523 17972 6532
rect 17548 5648 17588 6448
rect 18124 6488 18164 6497
rect 17644 6404 17684 6413
rect 17644 5816 17684 6364
rect 17740 5984 17780 5993
rect 17932 5984 17972 5993
rect 17780 5944 17932 5984
rect 17740 5935 17780 5944
rect 17932 5935 17972 5944
rect 17644 5767 17684 5776
rect 18028 5732 18068 5741
rect 17836 5648 17876 5657
rect 17588 5608 17836 5648
rect 17356 5060 17396 5069
rect 17356 4976 17396 5020
rect 17356 4925 17396 4936
rect 17260 4759 17300 4768
rect 16724 4096 16820 4136
rect 16684 4087 16724 4096
rect 16684 3968 16724 3977
rect 16492 3415 16532 3424
rect 16588 3632 16628 3641
rect 15916 2743 15956 2752
rect 16204 2860 16340 2900
rect 16396 3380 16436 3389
rect 16204 2792 16244 2860
rect 16204 2743 16244 2752
rect 16396 2708 16436 3340
rect 16396 2659 16436 2668
rect 16204 2624 16244 2633
rect 16204 2540 16244 2584
rect 16204 2489 16244 2500
rect 16588 2540 16628 3592
rect 16588 2491 16628 2500
rect 16684 2456 16724 3928
rect 16684 2407 16724 2416
rect 15820 2071 15860 2080
rect 13516 1817 13556 1912
rect 16780 1952 16820 4096
rect 17068 2876 17108 4684
rect 17548 4136 17588 5608
rect 17836 5599 17876 5608
rect 17068 2540 17108 2836
rect 17356 3632 17396 3641
rect 17356 2792 17396 3592
rect 17548 3632 17588 4096
rect 17644 4976 17684 4985
rect 17644 3716 17684 4936
rect 18028 4304 18068 5692
rect 18124 5564 18164 6448
rect 18316 5900 18356 7960
rect 18412 7951 18452 7960
rect 18412 7832 18452 7841
rect 18412 7412 18452 7792
rect 18412 7363 18452 7372
rect 18412 7076 18452 7087
rect 18412 6992 18452 7036
rect 18412 6943 18452 6952
rect 18124 5515 18164 5524
rect 18220 5860 18356 5900
rect 18412 6236 18452 6245
rect 18124 5396 18164 5405
rect 18124 4976 18164 5356
rect 18124 4927 18164 4936
rect 18028 4136 18068 4264
rect 18028 4087 18068 4096
rect 17644 3667 17684 3676
rect 17548 3583 17588 3592
rect 18124 3464 18164 3473
rect 18220 3464 18260 5860
rect 18412 5816 18452 6196
rect 18508 6152 18548 8716
rect 19084 8588 19124 8597
rect 19084 8168 19124 8548
rect 19084 8119 19124 8128
rect 18604 7916 18644 7925
rect 18604 7781 18644 7876
rect 19084 7916 19124 7925
rect 18660 7580 19028 7589
rect 18660 7531 19028 7540
rect 19084 7244 19124 7876
rect 19084 7195 19124 7204
rect 18604 7160 18644 7169
rect 18604 7025 18644 7120
rect 19180 6488 19220 9388
rect 19468 9428 19508 18376
rect 19756 17996 19796 19300
rect 19900 18920 20268 18929
rect 19900 18871 20268 18880
rect 20236 18752 20276 18761
rect 19756 17947 19796 17956
rect 19852 18584 19892 18593
rect 19852 18416 19892 18544
rect 20236 18584 20276 18712
rect 20236 18535 20276 18544
rect 19852 17744 19892 18376
rect 19948 18500 19988 18509
rect 19948 18365 19988 18460
rect 20140 18416 20180 18425
rect 20140 18281 20180 18376
rect 19852 17695 19892 17704
rect 19900 17408 20268 17417
rect 19900 17359 20268 17368
rect 19756 17072 19796 17081
rect 19564 16988 19604 16997
rect 19564 16853 19604 16948
rect 19756 16904 19796 17032
rect 19756 16484 19796 16864
rect 19948 17072 19988 17081
rect 19948 16652 19988 17032
rect 20140 16820 20180 16829
rect 20140 16685 20180 16780
rect 19948 16603 19988 16612
rect 19756 16435 19796 16444
rect 20140 16400 20180 16409
rect 19660 16316 19700 16325
rect 19660 16181 19700 16276
rect 20140 16265 20180 16360
rect 19900 15896 20268 15905
rect 19900 15847 20268 15856
rect 19660 15812 19700 15821
rect 19564 15476 19604 15485
rect 19564 15224 19604 15436
rect 19564 15175 19604 15184
rect 19660 15476 19700 15772
rect 19564 14720 19604 14815
rect 19564 14671 19604 14680
rect 19660 14636 19700 15436
rect 19852 15644 19892 15653
rect 19852 15056 19892 15604
rect 19852 15007 19892 15016
rect 19660 14587 19700 14596
rect 19756 14888 19796 14897
rect 19660 14384 19700 14393
rect 19660 13376 19700 14344
rect 19660 13327 19700 13336
rect 19660 13208 19700 13217
rect 19660 11360 19700 13168
rect 19756 13208 19796 14848
rect 19900 14384 20268 14393
rect 19900 14335 20268 14344
rect 20236 14048 20276 14057
rect 20140 13460 20180 13469
rect 20140 13325 20180 13420
rect 20236 13292 20276 14008
rect 20236 13243 20276 13252
rect 19756 13159 19796 13168
rect 19900 12872 20268 12881
rect 19900 12823 20268 12832
rect 20140 12284 20180 12293
rect 20140 12149 20180 12244
rect 19660 11276 19700 11320
rect 19900 11360 20268 11369
rect 19900 11311 20268 11320
rect 19756 11276 19796 11285
rect 19660 11236 19756 11276
rect 19756 11227 19796 11236
rect 19948 10856 19988 10865
rect 19564 10436 19604 10445
rect 19564 10301 19604 10396
rect 19948 10184 19988 10816
rect 19948 10135 19988 10144
rect 20332 10184 20372 22828
rect 20524 20852 20564 23020
rect 20524 20803 20564 20812
rect 20620 22112 20660 22121
rect 20428 20768 20468 20777
rect 20428 20096 20468 20728
rect 20620 20684 20660 22072
rect 20620 20549 20660 20644
rect 20428 20047 20468 20056
rect 20524 20012 20564 20021
rect 20524 19424 20564 19972
rect 20716 19928 20756 25096
rect 20812 24128 20852 26020
rect 20812 23876 20852 24088
rect 20812 23827 20852 23836
rect 20908 23120 20948 23129
rect 20908 22196 20948 23080
rect 20908 22147 20948 22156
rect 21004 21524 21044 26104
rect 21100 24548 21140 27868
rect 21196 25472 21236 25481
rect 21196 24716 21236 25432
rect 21196 24667 21236 24676
rect 21100 24508 21236 24548
rect 21100 23036 21140 23045
rect 21100 22280 21140 22996
rect 21100 22231 21140 22240
rect 20908 21484 21044 21524
rect 20908 20684 20948 21484
rect 21004 21356 21044 21365
rect 21004 20852 21044 21316
rect 21004 20803 21044 20812
rect 20908 20264 20948 20644
rect 20908 20215 20948 20224
rect 20716 19879 20756 19888
rect 20908 20012 20948 20021
rect 20524 19375 20564 19384
rect 20812 19340 20852 19349
rect 20812 18668 20852 19300
rect 20908 19256 20948 19972
rect 21100 19844 21140 19853
rect 21100 19340 21140 19804
rect 21196 19424 21236 24508
rect 21196 19375 21236 19384
rect 20948 19216 21044 19256
rect 20908 19207 20948 19216
rect 20812 18619 20852 18628
rect 20908 19088 20948 19097
rect 20908 18500 20948 19048
rect 21004 18584 21044 19216
rect 21004 18535 21044 18544
rect 20908 18451 20948 18460
rect 21100 18500 21140 19300
rect 21388 19256 21428 28120
rect 22732 27656 22772 27665
rect 22252 25976 22292 25985
rect 22252 25388 22292 25936
rect 22252 25339 22292 25348
rect 22732 25304 22772 27616
rect 23116 26900 23156 28600
rect 23116 26851 23156 26860
rect 23308 28580 23348 28589
rect 22732 25255 22772 25264
rect 23116 26648 23156 26657
rect 22828 25136 22868 25145
rect 22828 24632 22868 25096
rect 21580 24380 21620 24389
rect 21484 22196 21524 22205
rect 21580 22196 21620 24340
rect 22348 24296 22388 24305
rect 22252 23624 22292 23633
rect 22252 23120 22292 23584
rect 22348 23540 22388 24256
rect 22732 24044 22772 24053
rect 22732 23792 22772 24004
rect 22732 23743 22772 23752
rect 22348 23491 22388 23500
rect 22252 23071 22292 23080
rect 21772 22868 21812 22877
rect 21772 22364 21812 22828
rect 21772 22315 21812 22324
rect 21524 22156 21620 22196
rect 21484 22147 21524 22156
rect 21580 21608 21620 22156
rect 21964 22280 22004 22289
rect 21964 21776 22004 22240
rect 22252 22280 22292 22289
rect 21964 21727 22004 21736
rect 22060 22196 22100 22205
rect 21580 21559 21620 21568
rect 22060 21608 22100 22156
rect 22252 21776 22292 22240
rect 22252 21727 22292 21736
rect 22540 22112 22580 22121
rect 22060 21559 22100 21568
rect 22348 21524 22388 21533
rect 21388 18668 21428 19216
rect 21388 18619 21428 18628
rect 21868 19424 21908 19433
rect 21100 18451 21140 18460
rect 21868 18500 21908 19384
rect 21868 18451 21908 18460
rect 22348 17744 22388 21484
rect 22444 21440 22484 21449
rect 22444 20852 22484 21400
rect 22444 20803 22484 20812
rect 22348 17695 22388 17704
rect 20428 17240 20468 17249
rect 20468 17200 20660 17240
rect 20428 17191 20468 17200
rect 20620 17156 20660 17200
rect 20620 17107 20660 17116
rect 21388 17072 21428 17081
rect 20524 16988 20564 16997
rect 20428 16064 20468 16073
rect 20428 15392 20468 16024
rect 20428 15343 20468 15352
rect 20428 14636 20468 14645
rect 20428 14216 20468 14596
rect 20428 11696 20468 14176
rect 20428 11561 20468 11656
rect 19660 10100 19700 10109
rect 19564 9596 19604 9605
rect 19564 9461 19604 9556
rect 19468 9379 19508 9388
rect 19564 8672 19604 8681
rect 19660 8672 19700 10060
rect 19852 10016 19892 10025
rect 19468 8632 19564 8672
rect 19604 8632 19700 8672
rect 19756 9976 19852 10016
rect 19276 8336 19316 8345
rect 19276 8000 19316 8296
rect 19468 8168 19508 8632
rect 19564 8623 19604 8632
rect 19756 8588 19796 9976
rect 19852 9967 19892 9976
rect 19900 9848 20268 9857
rect 19900 9799 20268 9808
rect 19852 9680 19892 9689
rect 19852 9008 19892 9640
rect 20140 9596 20180 9605
rect 20140 9461 20180 9556
rect 19852 8959 19892 8968
rect 19948 9428 19988 9437
rect 19948 9344 19988 9388
rect 19948 9008 19988 9304
rect 20140 9344 20180 9353
rect 20140 9209 20180 9304
rect 19948 8959 19988 8968
rect 19756 8539 19796 8548
rect 19900 8336 20268 8345
rect 19900 8287 20268 8296
rect 19468 8033 19508 8128
rect 19852 8168 19892 8177
rect 19276 7951 19316 7960
rect 19852 8000 19892 8128
rect 19852 7951 19892 7960
rect 19180 6439 19220 6448
rect 19468 7916 19508 7925
rect 18508 6103 18548 6112
rect 18660 6068 19028 6077
rect 18660 6019 19028 6028
rect 18412 5767 18452 5776
rect 18316 5732 18356 5741
rect 18316 5060 18356 5692
rect 18316 4388 18356 5020
rect 18316 4339 18356 4348
rect 18412 5228 18452 5237
rect 18164 3424 18260 3464
rect 18124 3415 18164 3424
rect 17068 2491 17108 2500
rect 17164 2624 17204 2633
rect 17164 2489 17204 2584
rect 17356 2456 17396 2752
rect 17356 2407 17396 2416
rect 17644 3296 17684 3305
rect 17644 2708 17684 3256
rect 18220 3128 18260 3424
rect 18220 3079 18260 3088
rect 18316 4136 18356 4145
rect 18316 3548 18356 4096
rect 16820 1912 16916 1952
rect 16780 1903 16820 1912
rect 16780 1784 16820 1793
rect 13324 1231 13364 1240
rect 13420 1700 13460 1709
rect 12980 1072 13076 1112
rect 13420 1112 13460 1660
rect 14764 1700 14804 1709
rect 12940 1044 12980 1072
rect 13420 1063 13460 1072
rect 13516 1448 13556 1457
rect 12652 979 12692 988
rect 13516 1028 13556 1408
rect 14764 1112 14804 1660
rect 14764 1063 14804 1072
rect 15052 1280 15092 1289
rect 15052 1112 15092 1240
rect 16780 1196 16820 1744
rect 16876 1364 16916 1912
rect 17644 1868 17684 2668
rect 18316 2120 18356 3508
rect 18412 2204 18452 5188
rect 18796 5060 18836 5069
rect 18988 5060 19028 5069
rect 18836 5020 18988 5060
rect 18796 5011 18836 5020
rect 18988 5011 19028 5020
rect 19084 4892 19124 4901
rect 19084 4724 19124 4852
rect 19084 4675 19124 4684
rect 18660 4556 19028 4565
rect 18660 4507 19028 4516
rect 19468 3968 19508 7876
rect 20044 7160 20084 7169
rect 20140 7160 20180 7169
rect 20084 7120 20140 7160
rect 20044 7111 20084 7120
rect 20140 7111 20180 7120
rect 19900 6824 20268 6833
rect 19900 6775 20268 6784
rect 20332 6488 20372 10144
rect 20428 10604 20468 10613
rect 20428 10100 20468 10564
rect 20428 10051 20468 10060
rect 20428 9932 20468 9941
rect 20428 9428 20468 9892
rect 20428 9379 20468 9388
rect 20428 9176 20468 9185
rect 20428 9041 20468 9136
rect 20524 8840 20564 16948
rect 20908 16232 20948 16241
rect 20908 15728 20948 16192
rect 20908 15679 20948 15688
rect 21100 16232 21140 16241
rect 20620 15560 20660 15569
rect 20620 13964 20660 15520
rect 20620 13915 20660 13924
rect 20812 15308 20852 15317
rect 20812 14048 20852 15268
rect 20812 13208 20852 14008
rect 20812 13159 20852 13168
rect 20908 14804 20948 14813
rect 20812 13040 20852 13049
rect 20716 12536 20756 12545
rect 20620 11780 20660 11789
rect 20620 11108 20660 11740
rect 20620 10520 20660 11068
rect 20620 10471 20660 10480
rect 20716 11696 20756 12496
rect 20812 12368 20852 13000
rect 20812 12319 20852 12328
rect 20716 10940 20756 11656
rect 20908 11024 20948 14764
rect 21100 14804 21140 16192
rect 21100 14755 21140 14764
rect 21196 16148 21236 16157
rect 21196 14888 21236 16108
rect 21388 16064 21428 17032
rect 21580 17072 21620 17081
rect 21580 16484 21620 17032
rect 22540 17072 22580 22072
rect 22636 20600 22676 20609
rect 22636 17996 22676 20560
rect 22828 19340 22868 24592
rect 22924 24464 22964 24473
rect 22924 23876 22964 24424
rect 22924 23827 22964 23836
rect 22924 22112 22964 22121
rect 22924 21608 22964 22072
rect 22924 21559 22964 21568
rect 23116 20180 23156 26608
rect 23212 24464 23252 24473
rect 23212 24296 23252 24424
rect 23212 24247 23252 24256
rect 23308 23624 23348 28540
rect 23884 26900 23924 28600
rect 23884 26851 23924 26860
rect 23980 27740 24020 27749
rect 23788 26732 23828 26741
rect 23596 26648 23636 26657
rect 23308 23575 23348 23584
rect 23404 26480 23444 26489
rect 23404 21020 23444 26440
rect 23596 25472 23636 26608
rect 23788 25556 23828 26692
rect 23980 26312 24020 27700
rect 24460 27572 24500 27581
rect 24460 26984 24500 27532
rect 24460 26935 24500 26944
rect 24172 26816 24212 26825
rect 23980 26263 24020 26272
rect 24076 26648 24116 26657
rect 24076 26228 24116 26608
rect 24076 26179 24116 26188
rect 23788 25507 23828 25516
rect 23884 26144 23924 26153
rect 23596 25423 23636 25432
rect 23884 25388 23924 26104
rect 24172 26144 24212 26776
rect 24172 26095 24212 26104
rect 24652 26144 24692 28600
rect 24940 27152 24980 27161
rect 24652 26095 24692 26104
rect 24748 26228 24788 26237
rect 24556 25388 24596 25397
rect 23884 25339 23924 25348
rect 24460 25348 24556 25388
rect 23980 25220 24020 25229
rect 23596 23708 23636 23717
rect 23596 23288 23636 23668
rect 23980 23708 24020 25180
rect 24364 25136 24404 25145
rect 24364 24632 24404 25096
rect 24364 24583 24404 24592
rect 24460 24464 24500 25348
rect 24556 25339 24596 25348
rect 24748 25388 24788 26188
rect 24748 25339 24788 25348
rect 24844 26060 24884 26069
rect 24556 24632 24596 24641
rect 24748 24632 24788 24641
rect 24596 24592 24692 24632
rect 24556 24583 24596 24592
rect 24364 24424 24500 24464
rect 24556 24464 24596 24473
rect 23596 23239 23636 23248
rect 23692 23624 23732 23633
rect 23692 23120 23732 23584
rect 23692 23071 23732 23080
rect 23692 22280 23732 22375
rect 23692 22231 23732 22240
rect 23980 22196 24020 23668
rect 24076 23792 24116 23801
rect 24076 23372 24116 23752
rect 24076 23323 24116 23332
rect 24364 23204 24404 24424
rect 24460 24296 24500 24305
rect 24460 23792 24500 24256
rect 24556 23960 24596 24424
rect 24652 24380 24692 24592
rect 24652 24331 24692 24340
rect 24556 23911 24596 23920
rect 24460 23540 24500 23752
rect 24556 23708 24596 23717
rect 24556 23573 24596 23668
rect 24652 23624 24692 23633
rect 24460 23491 24500 23500
rect 24364 23036 24404 23164
rect 24460 23372 24500 23381
rect 24460 23120 24500 23332
rect 24460 23071 24500 23080
rect 24556 23288 24596 23297
rect 24364 22987 24404 22996
rect 24556 23036 24596 23248
rect 24652 23120 24692 23584
rect 24652 23071 24692 23080
rect 24556 22987 24596 22996
rect 24748 22952 24788 24592
rect 24844 24212 24884 26020
rect 24940 25976 24980 27112
rect 25420 26144 25460 28600
rect 25612 27656 25652 27665
rect 25900 27656 25940 27665
rect 25652 27616 25748 27656
rect 25612 27607 25652 27616
rect 25516 27404 25556 27413
rect 25516 26816 25556 27364
rect 25516 26767 25556 26776
rect 25708 26816 25748 27616
rect 25708 26732 25748 26776
rect 25708 26681 25748 26692
rect 25420 26095 25460 26104
rect 25612 26564 25652 26573
rect 24940 25388 24980 25936
rect 25612 25556 25652 26524
rect 25612 25507 25652 25516
rect 25708 26060 25748 26069
rect 25516 25472 25556 25481
rect 24940 25339 24980 25348
rect 25118 25313 25158 25385
rect 25118 25304 25172 25313
rect 25036 25264 25118 25304
rect 24940 25220 24980 25229
rect 24940 24716 24980 25180
rect 25036 24800 25076 25264
rect 25118 25255 25172 25264
rect 25036 24751 25076 24760
rect 25132 25136 25172 25145
rect 24940 24667 24980 24676
rect 24844 24163 24884 24172
rect 25036 24632 25076 24641
rect 24940 23876 24980 23885
rect 24844 23792 24884 23801
rect 24844 23288 24884 23752
rect 24940 23741 24980 23836
rect 24844 23239 24884 23248
rect 24940 23372 24980 23381
rect 24748 22903 24788 22912
rect 24844 23120 24884 23129
rect 24844 22364 24884 23080
rect 24844 22315 24884 22324
rect 24940 23120 24980 23332
rect 23692 22112 23732 22121
rect 23404 20971 23444 20980
rect 23500 22028 23540 22037
rect 23116 20131 23156 20140
rect 22828 19088 22868 19300
rect 23500 19340 23540 21988
rect 22828 19039 22868 19048
rect 23404 19088 23444 19097
rect 22636 17947 22676 17956
rect 22732 18416 22772 18425
rect 22540 17023 22580 17032
rect 22156 16820 22196 16829
rect 21388 16015 21428 16024
rect 21484 16316 21524 16325
rect 21484 15560 21524 16276
rect 21196 12620 21236 14848
rect 21292 15308 21332 15317
rect 21292 14216 21332 15268
rect 21484 15056 21524 15520
rect 21580 16148 21620 16444
rect 21580 15224 21620 16108
rect 21580 15175 21620 15184
rect 21868 16652 21908 16661
rect 21868 16316 21908 16612
rect 21484 15007 21524 15016
rect 21292 13292 21332 14176
rect 21484 14804 21524 14813
rect 21292 13243 21332 13252
rect 21388 14048 21428 14057
rect 21196 11108 21236 12580
rect 21388 13208 21428 14008
rect 21484 14048 21524 14764
rect 21580 14804 21620 14813
rect 21580 14720 21620 14764
rect 21580 14132 21620 14680
rect 21580 14083 21620 14092
rect 21484 13796 21524 14008
rect 21524 13756 21620 13796
rect 21484 13747 21524 13756
rect 21196 11059 21236 11068
rect 21292 11864 21332 11873
rect 21100 11024 21140 11033
rect 20908 10984 21100 11024
rect 20716 10352 20756 10900
rect 20716 9932 20756 10312
rect 20716 9883 20756 9892
rect 20908 10352 20948 10361
rect 20620 9848 20660 9857
rect 20620 9680 20660 9808
rect 20620 9631 20660 9640
rect 20908 9428 20948 10312
rect 21100 10352 21140 10984
rect 21292 10604 21332 11824
rect 21388 11696 21428 13168
rect 21388 11024 21428 11656
rect 21484 13292 21524 13301
rect 21484 13040 21524 13252
rect 21484 12536 21524 13000
rect 21484 11528 21524 12496
rect 21580 13040 21620 13756
rect 21580 11612 21620 13000
rect 21868 11696 21908 16276
rect 22156 15140 22196 16780
rect 22156 15091 22196 15100
rect 22444 16232 22484 16241
rect 22444 14720 22484 16192
rect 22252 14132 22292 14141
rect 22252 13208 22292 14092
rect 22444 14048 22484 14680
rect 22444 13913 22484 14008
rect 22636 13544 22676 13553
rect 22636 13409 22676 13504
rect 22252 13159 22292 13168
rect 22540 13208 22580 13217
rect 22540 12704 22580 13168
rect 22540 12655 22580 12664
rect 22636 12620 22676 12629
rect 22060 12452 22100 12461
rect 21868 11647 21908 11656
rect 21964 11780 22004 11789
rect 21580 11563 21620 11572
rect 21484 11479 21524 11488
rect 21388 10975 21428 10984
rect 21484 11108 21524 11117
rect 21292 10555 21332 10564
rect 21100 10303 21140 10312
rect 21388 10520 21428 10529
rect 21388 10184 21428 10480
rect 21388 10135 21428 10144
rect 20908 9379 20948 9388
rect 20524 8791 20564 8800
rect 21292 9008 21332 9017
rect 20428 8000 20468 8009
rect 20428 7412 20468 7960
rect 20428 7363 20468 7372
rect 21292 7412 21332 8968
rect 21484 7748 21524 11068
rect 21964 11024 22004 11740
rect 21580 10268 21620 10277
rect 21580 9008 21620 10228
rect 21964 10268 22004 10984
rect 22060 11696 22100 12412
rect 22636 12284 22676 12580
rect 22732 12536 22772 18376
rect 22924 17744 22964 17753
rect 22924 14720 22964 17704
rect 22924 14671 22964 14680
rect 23020 16988 23060 16997
rect 22828 13040 22868 13049
rect 22828 12980 22868 13000
rect 23020 13040 23060 16948
rect 23308 16904 23348 16913
rect 23020 12991 23060 13000
rect 23116 16232 23156 16241
rect 22828 12956 22964 12980
rect 22828 12940 22924 12956
rect 22924 12907 22964 12916
rect 23116 12872 23156 16192
rect 23116 12823 23156 12832
rect 23212 16148 23252 16157
rect 23212 12704 23252 16108
rect 23308 15980 23348 16864
rect 23308 15931 23348 15940
rect 23308 14552 23348 14561
rect 23308 14048 23348 14512
rect 23308 13999 23348 14008
rect 23308 13292 23348 13301
rect 23308 12788 23348 13252
rect 23308 12739 23348 12748
rect 23116 12664 23252 12704
rect 22732 12496 23060 12536
rect 22636 12235 22676 12244
rect 22636 11864 22676 11873
rect 22636 11780 22676 11824
rect 22636 11729 22676 11740
rect 22828 11780 22868 11789
rect 22060 11024 22100 11656
rect 22540 11696 22580 11705
rect 22060 10975 22100 10984
rect 22252 11108 22292 11117
rect 22252 10973 22292 11068
rect 21580 8959 21620 8968
rect 21676 9764 21716 9773
rect 21676 8000 21716 9724
rect 21772 9428 21812 9437
rect 21772 8840 21812 9388
rect 21964 9176 22004 10228
rect 21964 9127 22004 9136
rect 21772 8791 21812 8800
rect 21676 7951 21716 7960
rect 21964 8000 22004 8009
rect 21484 7699 21524 7708
rect 21484 7412 21524 7421
rect 21292 7372 21484 7412
rect 20332 6439 20372 6448
rect 20428 7160 20468 7169
rect 20140 6320 20180 6329
rect 20140 6185 20180 6280
rect 20428 5900 20468 7120
rect 21292 7160 21332 7372
rect 21484 7363 21524 7372
rect 21292 7111 21332 7120
rect 21484 7160 21524 7169
rect 20524 7076 20564 7085
rect 20524 6740 20564 7036
rect 20524 6691 20564 6700
rect 20620 6992 20660 7001
rect 20620 6656 20660 6952
rect 20620 6607 20660 6616
rect 20428 5851 20468 5860
rect 20716 6236 20756 6245
rect 20716 5480 20756 6196
rect 21484 5900 21524 7120
rect 21964 5984 22004 7960
rect 22540 6656 22580 11656
rect 22732 11696 22772 11705
rect 22732 11024 22772 11656
rect 22828 11192 22868 11740
rect 22828 11143 22868 11152
rect 22828 11024 22868 11033
rect 22732 10984 22828 11024
rect 22636 10184 22676 10193
rect 22636 9680 22676 10144
rect 22636 8000 22676 9640
rect 22828 8084 22868 10984
rect 22828 8035 22868 8044
rect 22636 7951 22676 7960
rect 23020 7160 23060 12496
rect 23116 8168 23156 12664
rect 23212 12536 23252 12545
rect 23212 11612 23252 12496
rect 23404 11948 23444 19048
rect 23500 18584 23540 19300
rect 23692 19256 23732 22072
rect 23980 21692 24020 22156
rect 23980 21643 24020 21652
rect 24460 22280 24500 22289
rect 23692 18668 23732 19216
rect 24172 20852 24212 20861
rect 24172 19256 24212 20812
rect 24172 19207 24212 19216
rect 24076 19088 24116 19097
rect 24076 18953 24116 19048
rect 23692 18619 23732 18628
rect 24460 18668 24500 22240
rect 24652 21608 24692 21617
rect 24652 21104 24692 21568
rect 24556 20684 24596 20693
rect 24556 20348 24596 20644
rect 24556 20299 24596 20308
rect 24652 19340 24692 21064
rect 24748 21272 24788 21281
rect 24748 20348 24788 21232
rect 24748 20299 24788 20308
rect 24940 20936 24980 23080
rect 24652 19291 24692 19300
rect 24748 19844 24788 19853
rect 24460 18619 24500 18628
rect 24748 19088 24788 19804
rect 23500 18535 23540 18544
rect 24748 18584 24788 19048
rect 24748 18535 24788 18544
rect 24844 19424 24884 19433
rect 24460 17744 24500 17753
rect 24364 17660 24404 17669
rect 23596 17576 23636 17585
rect 23500 16484 23540 16493
rect 23500 16232 23540 16444
rect 23500 16183 23540 16192
rect 23596 16316 23636 17536
rect 24268 17576 24308 17585
rect 23980 17156 24020 17165
rect 23980 16820 24020 17116
rect 24268 17156 24308 17536
rect 24268 17107 24308 17116
rect 23980 16771 24020 16780
rect 24268 16820 24308 16829
rect 23500 13880 23540 13889
rect 23500 13745 23540 13840
rect 23500 13544 23540 13553
rect 23500 12368 23540 13504
rect 23596 12536 23636 16276
rect 24268 16316 24308 16780
rect 24268 16267 24308 16276
rect 23692 16232 23732 16241
rect 24172 16232 24212 16241
rect 23692 15728 23732 16192
rect 23692 15679 23732 15688
rect 23884 16192 24172 16232
rect 23692 15476 23732 15485
rect 23692 14132 23732 15436
rect 23692 14083 23732 14092
rect 23788 14636 23828 14645
rect 23692 13124 23732 13219
rect 23692 13075 23732 13084
rect 23692 12956 23732 12965
rect 23692 12872 23732 12916
rect 23692 12821 23732 12832
rect 23788 12956 23828 14596
rect 23884 13040 23924 16192
rect 24172 16183 24212 16192
rect 24172 15560 24212 15569
rect 24076 15520 24172 15560
rect 23980 14720 24020 14729
rect 23980 14585 24020 14680
rect 23980 13964 24020 13973
rect 23980 13829 24020 13924
rect 23884 12991 23924 13000
rect 24076 13040 24116 15520
rect 24172 15511 24212 15520
rect 24364 14888 24404 17620
rect 24460 17576 24500 17704
rect 24844 17744 24884 19384
rect 24460 17527 24500 17536
rect 24652 17660 24692 17669
rect 24556 17240 24596 17249
rect 24460 16820 24500 16829
rect 24460 16685 24500 16780
rect 24364 14839 24404 14848
rect 24556 16232 24596 17200
rect 24652 16988 24692 17620
rect 24844 17072 24884 17704
rect 24940 17744 24980 20896
rect 25036 20600 25076 24592
rect 25132 23204 25172 25096
rect 25420 25136 25460 25145
rect 25420 24716 25460 25096
rect 25420 24667 25460 24676
rect 25516 23960 25556 25432
rect 25612 25220 25652 25229
rect 25612 24632 25652 25180
rect 25612 24583 25652 24592
rect 25420 23920 25516 23960
rect 25132 23155 25172 23164
rect 25324 23204 25364 23213
rect 25228 22868 25268 22877
rect 25228 22532 25268 22828
rect 25228 22483 25268 22492
rect 25324 22448 25364 23164
rect 25132 22280 25172 22289
rect 25132 22145 25172 22240
rect 25036 20551 25076 20560
rect 25228 21776 25268 21785
rect 25228 20348 25268 21736
rect 25228 20299 25268 20308
rect 24940 17695 24980 17704
rect 25036 20096 25076 20105
rect 25036 19928 25076 20056
rect 25324 20096 25364 22408
rect 25420 20768 25460 23920
rect 25516 23911 25556 23920
rect 25612 23960 25652 23969
rect 25516 23456 25556 23465
rect 25516 23120 25556 23416
rect 25516 23071 25556 23080
rect 25612 21944 25652 23920
rect 25612 21895 25652 21904
rect 25516 21608 25556 21617
rect 25516 21020 25556 21568
rect 25708 21524 25748 26020
rect 25804 25640 25844 25649
rect 25804 25505 25844 25600
rect 25900 25304 25940 27616
rect 26188 26984 26228 28600
rect 26956 27740 26996 28600
rect 27724 28160 27764 28600
rect 27724 28111 27764 28120
rect 27674 27992 28042 28001
rect 27674 27943 28042 27952
rect 26956 27691 26996 27700
rect 28492 27740 28532 28600
rect 29260 27824 29300 28600
rect 30028 28580 30068 28600
rect 30028 28531 30068 28540
rect 29260 27775 29300 27784
rect 29356 28160 29396 28169
rect 28492 27691 28532 27700
rect 29356 27656 29396 28120
rect 29356 27607 29396 27616
rect 27820 27572 27860 27581
rect 27148 27404 27188 27413
rect 26434 27236 26802 27245
rect 26434 27187 26802 27196
rect 26188 26935 26228 26944
rect 26956 27068 26996 27077
rect 26284 26900 26324 26909
rect 26284 26816 26324 26860
rect 26284 26765 26324 26776
rect 25996 26732 26036 26741
rect 25996 26228 26036 26692
rect 25996 26179 26036 26188
rect 26188 26312 26228 26321
rect 26092 26060 26132 26069
rect 25804 24716 25844 24725
rect 25804 24581 25844 24676
rect 25804 24380 25844 24389
rect 25804 23792 25844 24340
rect 25900 23876 25940 25264
rect 25996 25976 26036 25985
rect 25996 23960 26036 25936
rect 25996 23911 26036 23920
rect 26092 25388 26132 26020
rect 25900 23827 25940 23836
rect 25804 23743 25844 23752
rect 25900 23708 25940 23717
rect 25900 23204 25940 23668
rect 26092 23624 26132 25348
rect 26188 24716 26228 26272
rect 26284 26228 26324 26237
rect 26284 25388 26324 26188
rect 26956 26060 26996 27028
rect 27052 26816 27092 26825
rect 27052 26228 27092 26776
rect 27052 26179 27092 26188
rect 26956 26011 26996 26020
rect 27148 26060 27188 27364
rect 27820 26984 27860 27532
rect 28972 27572 29012 27581
rect 27820 26935 27860 26944
rect 28684 27404 28724 27413
rect 27436 26900 27476 26909
rect 27148 26011 27188 26020
rect 27340 26648 27380 26657
rect 27244 25976 27284 25985
rect 26860 25892 26900 25901
rect 26434 25724 26802 25733
rect 26434 25675 26802 25684
rect 26284 25339 26324 25348
rect 26476 25556 26516 25565
rect 26188 24667 26228 24676
rect 26284 25220 26324 25229
rect 26188 23624 26228 23633
rect 26092 23584 26188 23624
rect 26092 23456 26132 23465
rect 25996 23204 26036 23232
rect 25900 23164 25996 23204
rect 25804 22868 25844 22877
rect 25804 22112 25844 22828
rect 25900 22196 25940 23164
rect 25996 23155 26036 23164
rect 25900 22147 25940 22156
rect 25996 23036 26036 23045
rect 25804 22063 25844 22072
rect 25996 21776 26036 22996
rect 26092 22280 26132 23416
rect 26188 22364 26228 23584
rect 26188 22315 26228 22324
rect 26092 22231 26132 22240
rect 26188 22196 26228 22205
rect 26092 21776 26132 21785
rect 25996 21736 26092 21776
rect 25516 20971 25556 20980
rect 25612 21484 25748 21524
rect 25804 21524 25844 21564
rect 25420 20719 25460 20728
rect 25516 20768 25556 20777
rect 25516 20600 25556 20728
rect 25516 20551 25556 20560
rect 25612 20600 25652 21484
rect 25804 21440 25844 21484
rect 25612 20551 25652 20560
rect 25708 21356 25748 21365
rect 25324 20047 25364 20056
rect 25708 20096 25748 21316
rect 25804 20852 25844 21400
rect 25804 20600 25844 20812
rect 25996 21356 26036 21365
rect 25900 20768 25940 20777
rect 25900 20633 25940 20728
rect 25804 20551 25844 20560
rect 25996 20180 26036 21316
rect 26092 20936 26132 21736
rect 26092 20887 26132 20896
rect 25996 20131 26036 20140
rect 25708 20047 25748 20056
rect 25036 19172 25076 19888
rect 25036 18416 25076 19132
rect 25036 17744 25076 18376
rect 25036 17156 25076 17704
rect 25036 17107 25076 17116
rect 25324 19256 25364 19265
rect 25324 18500 25364 19216
rect 25324 17912 25364 18460
rect 24844 17023 24884 17032
rect 24652 16939 24692 16948
rect 24172 14720 24212 14729
rect 24172 14132 24212 14680
rect 24268 14636 24308 14645
rect 24268 14501 24308 14596
rect 24172 13292 24212 14092
rect 24364 14468 24404 14477
rect 24268 13964 24308 13973
rect 24268 13460 24308 13924
rect 24268 13411 24308 13420
rect 24172 13243 24212 13252
rect 24076 12991 24116 13000
rect 24172 13124 24212 13133
rect 23596 12487 23636 12496
rect 23692 12536 23732 12545
rect 23500 12328 23636 12368
rect 23212 11563 23252 11572
rect 23308 11908 23444 11948
rect 23500 12200 23540 12209
rect 23212 11024 23252 11033
rect 23212 10436 23252 10984
rect 23212 10387 23252 10396
rect 23308 10100 23348 11908
rect 23500 11612 23540 12160
rect 23500 11563 23540 11572
rect 23596 11780 23636 12328
rect 23692 12200 23732 12496
rect 23788 12536 23828 12916
rect 24076 12872 24116 12881
rect 23884 12788 23924 12797
rect 23884 12704 23924 12748
rect 23884 12653 23924 12664
rect 23788 12487 23828 12496
rect 23692 12151 23732 12160
rect 23884 12452 23924 12461
rect 23500 11108 23540 11117
rect 23500 11024 23540 11068
rect 23500 10973 23540 10984
rect 23500 10772 23540 10781
rect 23500 10184 23540 10732
rect 23500 10135 23540 10144
rect 23308 10060 23444 10100
rect 23308 9932 23348 9941
rect 23308 9512 23348 9892
rect 23308 9463 23348 9472
rect 23308 9344 23348 9353
rect 23308 8756 23348 9304
rect 23404 8840 23444 10060
rect 23500 9512 23540 9523
rect 23500 9428 23540 9472
rect 23500 9379 23540 9388
rect 23404 8800 23540 8840
rect 23308 8707 23348 8716
rect 23404 8672 23444 8681
rect 23404 8537 23444 8632
rect 23116 8119 23156 8128
rect 23500 7412 23540 8800
rect 23116 7160 23156 7169
rect 23020 7120 23116 7160
rect 23116 7076 23156 7120
rect 23500 7160 23540 7372
rect 23500 7111 23540 7120
rect 23116 6996 23156 7036
rect 22060 6488 22100 6497
rect 22060 6404 22100 6448
rect 22348 6488 22388 6497
rect 22060 6353 22100 6364
rect 22252 6404 22292 6413
rect 21964 5935 22004 5944
rect 21484 5851 21524 5860
rect 19900 5312 20268 5321
rect 19900 5263 20268 5272
rect 20716 5060 20756 5440
rect 21964 5648 22004 5657
rect 19468 3919 19508 3928
rect 20524 4976 20564 4985
rect 20524 4724 20564 4936
rect 19900 3800 20268 3809
rect 19900 3751 20268 3760
rect 20524 3716 20564 4684
rect 20716 4388 20756 5020
rect 20716 4339 20756 4348
rect 21580 5144 21620 5153
rect 18508 3464 18548 3473
rect 19276 3464 19316 3473
rect 18508 2876 18548 3424
rect 19180 3424 19276 3464
rect 18660 3044 19028 3053
rect 18660 2995 19028 3004
rect 18508 2624 18548 2836
rect 19180 2708 19220 3424
rect 19276 3415 19316 3424
rect 19660 3464 19700 3473
rect 19276 3212 19316 3221
rect 19276 2792 19316 3172
rect 19276 2743 19316 2752
rect 19180 2659 19220 2668
rect 18508 2575 18548 2584
rect 19660 2624 19700 3424
rect 18412 2155 18452 2164
rect 18316 2071 18356 2080
rect 17644 1819 17684 1828
rect 19180 1868 19220 1877
rect 16876 1315 16916 1324
rect 18220 1700 18260 1709
rect 16780 1147 16820 1156
rect 13516 979 13556 988
rect 12556 811 12596 820
rect 15052 860 15092 1072
rect 18220 1028 18260 1660
rect 19084 1700 19124 1709
rect 18660 1532 19028 1541
rect 18660 1483 19028 1492
rect 19084 1196 19124 1660
rect 19180 1280 19220 1828
rect 19660 1448 19700 2584
rect 20140 3464 20180 3473
rect 20140 2540 20180 3424
rect 20524 3464 20564 3676
rect 20236 3212 20276 3221
rect 20236 2624 20276 3172
rect 20524 2900 20564 3424
rect 21100 4136 21140 4145
rect 21004 3128 21044 3137
rect 20524 2860 20660 2900
rect 20236 2575 20276 2584
rect 20620 2624 20660 2860
rect 20620 2575 20660 2584
rect 20140 2491 20180 2500
rect 19660 1399 19700 1408
rect 19756 2372 19796 2381
rect 19180 1231 19220 1240
rect 19084 1147 19124 1156
rect 18220 979 18260 988
rect 19756 1028 19796 2332
rect 19900 2288 20268 2297
rect 19900 2239 20268 2248
rect 20908 1868 20948 1877
rect 20908 1280 20948 1828
rect 21004 1784 21044 3088
rect 21100 2876 21140 4096
rect 21100 2827 21140 2836
rect 21004 1735 21044 1744
rect 21580 2456 21620 5104
rect 21676 4976 21716 4985
rect 21676 3464 21716 4936
rect 21676 3415 21716 3424
rect 21964 3464 22004 5608
rect 22252 5480 22292 6364
rect 22348 5816 22388 6448
rect 22348 5767 22388 5776
rect 22540 5648 22580 6616
rect 23212 6992 23252 7001
rect 22540 5599 22580 5608
rect 22828 6320 22868 6329
rect 22252 3632 22292 5440
rect 22252 3583 22292 3592
rect 22828 3632 22868 6280
rect 23116 5816 23156 5825
rect 22924 5144 22964 5153
rect 22924 4136 22964 5104
rect 23116 4976 23156 5776
rect 23212 5228 23252 6952
rect 23404 6992 23444 7001
rect 23404 6572 23444 6952
rect 23596 6992 23636 11740
rect 23692 12032 23732 12041
rect 23692 10772 23732 11992
rect 23884 11780 23924 12412
rect 23980 12284 24020 12293
rect 23980 11864 24020 12244
rect 23980 11815 24020 11824
rect 23884 11731 23924 11740
rect 23980 11696 24020 11705
rect 23884 11528 23924 11537
rect 23884 11024 23924 11488
rect 23980 11192 24020 11656
rect 23980 11143 24020 11152
rect 23884 10975 23924 10984
rect 23692 10732 23924 10772
rect 23692 10352 23732 10361
rect 23692 9092 23732 10312
rect 23788 10016 23828 10025
rect 23788 9512 23828 9976
rect 23788 9463 23828 9472
rect 23692 9043 23732 9052
rect 23788 9260 23828 9269
rect 23788 8084 23828 9220
rect 23884 8588 23924 10732
rect 24076 10352 24116 12832
rect 24172 11612 24212 13084
rect 24172 11563 24212 11572
rect 24268 13040 24308 13049
rect 24268 12200 24308 13000
rect 24076 10303 24116 10312
rect 24172 11108 24212 11117
rect 23980 10100 24020 10109
rect 23980 8672 24020 10060
rect 23980 8623 24020 8632
rect 23884 8539 23924 8548
rect 23788 8035 23828 8044
rect 23596 6943 23636 6952
rect 23980 8000 24020 8009
rect 23980 6992 24020 7960
rect 23884 6908 23924 6917
rect 23596 6824 23636 6833
rect 23884 6824 23924 6868
rect 23636 6784 23924 6824
rect 23596 6775 23636 6784
rect 23404 6523 23444 6532
rect 23212 5179 23252 5188
rect 23500 6488 23540 6497
rect 23116 4724 23156 4936
rect 23500 4976 23540 6448
rect 23500 4808 23540 4936
rect 23500 4759 23540 4768
rect 23884 4976 23924 4985
rect 23116 4675 23156 4684
rect 22924 4087 22964 4096
rect 22828 3583 22868 3592
rect 23596 3968 23636 3977
rect 21964 2624 22004 3424
rect 22636 3464 22676 3473
rect 22636 2792 22676 3424
rect 23212 3380 23252 3389
rect 22924 3128 22964 3137
rect 20908 1231 20948 1240
rect 21580 1280 21620 2416
rect 21868 2540 21908 2549
rect 21868 1952 21908 2500
rect 21964 2120 22004 2584
rect 22156 2624 22196 2633
rect 22636 2624 22676 2752
rect 22156 2204 22196 2584
rect 22540 2584 22676 2624
rect 22828 2876 22868 2885
rect 22156 2155 22196 2164
rect 22348 2456 22388 2465
rect 21964 2071 22004 2080
rect 21868 1903 21908 1912
rect 22348 1952 22388 2416
rect 22540 2372 22580 2584
rect 22540 2323 22580 2332
rect 22636 2456 22676 2465
rect 22348 1903 22388 1912
rect 22636 1868 22676 2416
rect 22636 1819 22676 1828
rect 22828 1868 22868 2836
rect 22924 2624 22964 3088
rect 23212 2708 23252 3340
rect 23212 2659 23252 2668
rect 22924 2575 22964 2584
rect 23596 2540 23636 3928
rect 23788 3212 23828 3221
rect 23788 2624 23828 3172
rect 23884 2708 23924 4936
rect 23884 2659 23924 2668
rect 23788 2575 23828 2584
rect 23596 2491 23636 2500
rect 22828 1819 22868 1828
rect 23116 2120 23156 2129
rect 21580 1231 21620 1240
rect 23116 1112 23156 2080
rect 23980 2036 24020 6952
rect 24172 6824 24212 11068
rect 24268 6992 24308 12160
rect 24364 9596 24404 14428
rect 24460 14132 24500 14141
rect 24460 13964 24500 14092
rect 24460 13915 24500 13924
rect 24460 13208 24500 13217
rect 24460 12704 24500 13168
rect 24460 12655 24500 12664
rect 24556 12956 24596 16192
rect 24844 16820 24884 16829
rect 24844 16568 24884 16780
rect 24652 14804 24692 14813
rect 24652 14669 24692 14764
rect 24748 14720 24788 14729
rect 24652 14048 24692 14057
rect 24652 13913 24692 14008
rect 24460 12536 24500 12545
rect 24460 11360 24500 12496
rect 24556 12452 24596 12916
rect 24652 13292 24692 13301
rect 24652 12536 24692 13252
rect 24652 12487 24692 12496
rect 24556 12403 24596 12412
rect 24556 11360 24596 11369
rect 24460 11320 24556 11360
rect 24460 11024 24500 11033
rect 24460 10436 24500 10984
rect 24460 10387 24500 10396
rect 24556 10268 24596 11320
rect 24748 11108 24788 14680
rect 24748 11059 24788 11068
rect 24844 10772 24884 16528
rect 25228 15728 25268 15737
rect 25036 15560 25076 15569
rect 25036 15056 25076 15520
rect 25036 15007 25076 15016
rect 25228 15560 25268 15688
rect 25228 14804 25268 15520
rect 25324 15308 25364 17872
rect 26092 19172 26132 19181
rect 26188 19172 26228 22156
rect 26284 21524 26324 25180
rect 26476 25136 26516 25516
rect 26668 25388 26708 25397
rect 26476 25087 26516 25096
rect 26572 25304 26612 25313
rect 26380 25052 26420 25061
rect 26380 24800 26420 25012
rect 26380 24751 26420 24760
rect 26572 24800 26612 25264
rect 26572 24751 26612 24760
rect 26668 24548 26708 25348
rect 26764 25388 26804 25397
rect 26764 24716 26804 25348
rect 26764 24667 26804 24676
rect 26860 25304 26900 25852
rect 26956 25724 26996 25733
rect 26956 25640 26996 25684
rect 26956 25589 26996 25600
rect 27244 25556 27284 25936
rect 27340 25808 27380 26608
rect 27340 25759 27380 25768
rect 27244 25507 27284 25516
rect 26956 25388 26996 25483
rect 26956 25339 26996 25348
rect 26860 24884 26900 25264
rect 26668 24499 26708 24508
rect 26434 24212 26802 24221
rect 26434 24163 26802 24172
rect 26572 23960 26612 23969
rect 26380 23792 26420 23801
rect 26380 23036 26420 23752
rect 26572 23624 26612 23920
rect 26860 23792 26900 24844
rect 26956 25220 26996 25229
rect 26956 24632 26996 25180
rect 27436 24716 27476 26860
rect 27628 26816 27668 26825
rect 27436 24667 27476 24676
rect 27532 26732 27572 26741
rect 26956 24497 26996 24592
rect 27340 24632 27380 24641
rect 27532 24632 27572 26692
rect 27628 26681 27668 26776
rect 28492 26816 28532 26825
rect 27674 26480 28042 26489
rect 27674 26431 28042 26440
rect 27628 26144 27668 26153
rect 27628 25388 27668 26104
rect 28492 26144 28532 26776
rect 28684 26228 28724 27364
rect 28684 26179 28724 26188
rect 28780 26900 28820 26909
rect 28012 26060 28052 26069
rect 27628 25339 27668 25348
rect 27820 25976 27860 25985
rect 27820 25388 27860 25936
rect 27820 25339 27860 25348
rect 28012 25388 28052 26020
rect 28492 26009 28532 26104
rect 28780 25976 28820 26860
rect 28780 25927 28820 25936
rect 28012 25304 28052 25348
rect 28396 25892 28436 25901
rect 28012 25224 28052 25264
rect 28204 25304 28244 25313
rect 27674 24968 28042 24977
rect 27674 24919 28042 24928
rect 27724 24632 27764 24641
rect 27532 24592 27724 24632
rect 27764 24592 27860 24632
rect 27148 24380 27188 24389
rect 26860 23743 26900 23752
rect 26956 24044 26996 24053
rect 26572 23575 26612 23584
rect 26860 23624 26900 23633
rect 26860 23120 26900 23584
rect 26860 23071 26900 23080
rect 26956 23288 26996 24004
rect 27148 23960 27188 24340
rect 27340 24128 27380 24592
rect 27724 24583 27764 24592
rect 27340 24079 27380 24088
rect 27532 24464 27572 24473
rect 27148 23911 27188 23920
rect 27532 23624 27572 24424
rect 27820 23792 27860 24592
rect 27820 23657 27860 23752
rect 28108 24548 28148 24557
rect 26380 22868 26420 22996
rect 26668 23036 26708 23045
rect 26668 22901 26708 22996
rect 26380 22819 26420 22828
rect 26860 22868 26900 22877
rect 26434 22700 26802 22709
rect 26434 22651 26802 22660
rect 26380 21776 26420 21785
rect 26380 21692 26420 21736
rect 26380 21641 26420 21652
rect 26860 21692 26900 22828
rect 26860 21557 26900 21652
rect 26284 20936 26324 21484
rect 26572 21524 26612 21533
rect 26572 21389 26612 21484
rect 26434 21188 26802 21197
rect 26434 21139 26802 21148
rect 26572 21020 26612 21029
rect 26476 20936 26516 20945
rect 26284 20896 26476 20936
rect 26476 20887 26516 20896
rect 26476 20768 26516 20777
rect 26476 20600 26516 20728
rect 26476 20551 26516 20560
rect 26572 20012 26612 20980
rect 26764 21020 26804 21029
rect 26764 20885 26804 20980
rect 26764 20348 26804 20357
rect 26572 19963 26612 19972
rect 26668 20264 26708 20273
rect 26132 19132 26228 19172
rect 26284 19928 26324 19937
rect 26092 18332 26132 19132
rect 26284 18500 26324 19888
rect 26668 19844 26708 20224
rect 26764 20213 26804 20308
rect 26668 19795 26708 19804
rect 26434 19676 26802 19685
rect 26434 19627 26802 19636
rect 26956 18584 26996 23248
rect 27436 23540 27476 23549
rect 27148 23204 27188 23213
rect 27052 23036 27092 23045
rect 27052 22448 27092 22996
rect 27052 22399 27092 22408
rect 27052 21692 27092 21701
rect 27052 20768 27092 21652
rect 27148 21440 27188 23164
rect 27436 23204 27476 23500
rect 27436 23155 27476 23164
rect 27340 23036 27380 23045
rect 27244 22868 27284 22877
rect 27244 21524 27284 22828
rect 27340 22028 27380 22996
rect 27532 22364 27572 23584
rect 27674 23456 28042 23465
rect 27674 23407 28042 23416
rect 27724 22868 27764 22877
rect 27340 21776 27380 21988
rect 27340 21727 27380 21736
rect 27436 22280 27476 22320
rect 27532 22315 27572 22324
rect 27628 22616 27668 22625
rect 27436 22196 27476 22240
rect 27436 21608 27476 22156
rect 27628 22112 27668 22576
rect 27724 22280 27764 22828
rect 28108 22448 28148 24508
rect 28204 22616 28244 25264
rect 28396 24716 28436 25852
rect 28972 25640 29012 27532
rect 28972 25591 29012 25600
rect 29452 27572 29492 27581
rect 28684 25304 28724 25313
rect 28684 24800 28724 25264
rect 28684 24751 28724 24760
rect 28300 24676 28396 24716
rect 28300 23792 28340 24676
rect 28396 24667 28436 24676
rect 28300 23743 28340 23752
rect 28396 24548 28436 24557
rect 28204 22567 28244 22576
rect 28108 22408 28244 22448
rect 27724 22231 27764 22240
rect 28108 22280 28148 22289
rect 27436 21559 27476 21568
rect 27532 22072 27668 22112
rect 27340 21524 27380 21533
rect 27244 21484 27340 21524
rect 27148 21391 27188 21400
rect 27052 20600 27092 20728
rect 27244 20852 27284 20861
rect 27244 20717 27284 20812
rect 27340 20768 27380 21484
rect 27436 21272 27476 21281
rect 27436 21020 27476 21232
rect 27436 20971 27476 20980
rect 27340 20728 27476 20768
rect 27436 20684 27476 20728
rect 27436 20635 27476 20644
rect 27052 20348 27092 20560
rect 27052 20299 27092 20308
rect 27148 20600 27188 20609
rect 27148 20264 27188 20560
rect 27052 20012 27092 20021
rect 27052 19004 27092 19972
rect 27052 18955 27092 18964
rect 26956 18535 26996 18544
rect 27148 18752 27188 20224
rect 27340 20600 27380 20609
rect 27340 20180 27380 20560
rect 27436 20348 27476 20357
rect 27436 20264 27476 20308
rect 27532 20264 27572 22072
rect 27674 21944 28042 21953
rect 27674 21895 28042 21904
rect 28108 21692 28148 22240
rect 28204 22196 28244 22408
rect 28396 22364 28436 24508
rect 28780 24380 28820 24389
rect 28396 22315 28436 22324
rect 28492 24044 28532 24053
rect 28492 23876 28532 24004
rect 28204 22156 28436 22196
rect 28108 21643 28148 21652
rect 28396 21944 28436 22156
rect 27628 21608 27668 21617
rect 27628 21473 27668 21568
rect 28300 21524 28340 21533
rect 28012 21356 28052 21365
rect 28012 20852 28052 21316
rect 28204 21020 28244 21029
rect 28052 20812 28148 20852
rect 28012 20803 28052 20812
rect 27820 20768 27860 20777
rect 27820 20633 27860 20728
rect 27674 20432 28042 20441
rect 27674 20383 28042 20392
rect 27532 20224 27668 20264
rect 27436 20213 27476 20224
rect 27340 20131 27380 20140
rect 27628 20180 27668 20224
rect 27628 20131 27668 20140
rect 27532 20096 27572 20105
rect 26284 18451 26324 18460
rect 26092 17744 26132 18292
rect 26092 17695 26132 17704
rect 26188 18248 26228 18257
rect 26092 16316 26132 16325
rect 25996 15728 26036 15737
rect 25324 15259 25364 15268
rect 25900 15560 25940 15569
rect 25228 14755 25268 14764
rect 25612 14888 25652 14897
rect 24940 14720 24980 14729
rect 24940 14216 24980 14680
rect 25420 14720 25460 14729
rect 24940 14167 24980 14176
rect 25228 14216 25268 14225
rect 24940 14048 24980 14057
rect 24980 14008 25172 14048
rect 24940 13999 24980 14008
rect 25132 13964 25172 14008
rect 25036 12872 25076 12881
rect 24556 10219 24596 10228
rect 24652 10436 24692 10445
rect 24364 9512 24404 9556
rect 24364 7076 24404 9472
rect 24460 9848 24500 9857
rect 24460 9344 24500 9808
rect 24652 9428 24692 10396
rect 24844 10016 24884 10732
rect 24940 11780 24980 11789
rect 24940 10184 24980 11740
rect 25036 11108 25076 12832
rect 25036 11059 25076 11068
rect 25132 10520 25172 13924
rect 25228 13376 25268 14176
rect 25228 13327 25268 13336
rect 25324 13880 25364 13889
rect 25228 13208 25268 13217
rect 25228 12956 25268 13168
rect 25228 12907 25268 12916
rect 25132 10471 25172 10480
rect 25324 11696 25364 13840
rect 25420 12620 25460 14680
rect 25516 14048 25556 14057
rect 25516 13913 25556 14008
rect 25420 11780 25460 12580
rect 25420 11731 25460 11740
rect 25324 10184 25364 11656
rect 25516 11696 25556 11705
rect 25516 11612 25556 11656
rect 25516 11561 25556 11572
rect 25420 10940 25460 10949
rect 25420 10352 25460 10900
rect 25420 10303 25460 10312
rect 24980 10144 25076 10184
rect 24940 10135 24980 10144
rect 24844 9967 24884 9976
rect 24652 9379 24692 9388
rect 24844 9596 24884 9605
rect 24460 8756 24500 9304
rect 24460 8707 24500 8716
rect 24556 8840 24596 8849
rect 24364 7027 24404 7036
rect 24268 6943 24308 6952
rect 24172 6784 24308 6824
rect 24172 6404 24212 6413
rect 23980 1987 24020 1996
rect 24076 5648 24116 5657
rect 24076 4808 24116 5608
rect 24172 5144 24212 6364
rect 24172 5095 24212 5104
rect 24076 2708 24116 4768
rect 24172 4136 24212 4145
rect 24172 3464 24212 4096
rect 24172 3415 24212 3424
rect 23500 1868 23540 1877
rect 23116 1063 23156 1072
rect 23308 1700 23348 1709
rect 19756 979 19796 988
rect 23308 1028 23348 1660
rect 23500 1364 23540 1828
rect 23500 1315 23540 1324
rect 23788 1784 23828 1793
rect 23788 1196 23828 1744
rect 23788 1147 23828 1156
rect 24076 1112 24116 2668
rect 24172 2372 24212 2381
rect 24172 1952 24212 2332
rect 24172 1903 24212 1912
rect 24268 2288 24308 6784
rect 24556 5396 24596 8800
rect 24844 8840 24884 9556
rect 25036 9512 25076 10144
rect 25324 10135 25364 10144
rect 25612 9848 25652 14848
rect 25804 14048 25844 14059
rect 25804 13964 25844 14008
rect 25804 13915 25844 13924
rect 25900 13460 25940 15520
rect 25996 14048 26036 15688
rect 26092 14216 26132 16276
rect 26188 14972 26228 18208
rect 26434 18164 26802 18173
rect 26434 18115 26802 18124
rect 26860 17996 26900 18005
rect 26434 16652 26802 16661
rect 26434 16603 26802 16612
rect 26860 16316 26900 17956
rect 27148 17828 27188 18712
rect 27148 17779 27188 17788
rect 27244 19844 27284 19853
rect 27148 17072 27188 17081
rect 26860 16267 26900 16276
rect 27052 16820 27092 16829
rect 27052 16316 27092 16780
rect 27148 16484 27188 17032
rect 27148 16435 27188 16444
rect 27052 16267 27092 16276
rect 26380 16232 26420 16241
rect 26284 15896 26324 15905
rect 26284 15392 26324 15856
rect 26380 15644 26420 16192
rect 26380 15595 26420 15604
rect 26476 16064 26516 16073
rect 26476 15560 26516 16024
rect 26476 15511 26516 15520
rect 26860 15560 26900 15569
rect 26284 15343 26324 15352
rect 26434 15140 26802 15149
rect 26434 15091 26802 15100
rect 26860 14972 26900 15520
rect 27052 15560 27092 15569
rect 27244 15560 27284 19804
rect 27340 19172 27380 19181
rect 27340 17744 27380 19132
rect 27436 19088 27476 19097
rect 27436 18668 27476 19048
rect 27436 18619 27476 18628
rect 27532 17996 27572 20056
rect 28108 19340 28148 20812
rect 28204 20180 28244 20980
rect 28300 20852 28340 21484
rect 28300 20803 28340 20812
rect 28204 20131 28244 20140
rect 28300 20600 28340 20609
rect 28108 19291 28148 19300
rect 28300 19172 28340 20560
rect 27674 18920 28042 18929
rect 27674 18871 28042 18880
rect 27532 17947 27572 17956
rect 28108 18584 28148 18593
rect 27340 17695 27380 17704
rect 28108 17660 28148 18544
rect 28204 18500 28244 18509
rect 28300 18500 28340 19132
rect 28244 18460 28340 18500
rect 28204 18451 28244 18460
rect 28396 17828 28436 21904
rect 28492 21692 28532 23836
rect 28492 20768 28532 21652
rect 28684 23792 28724 23801
rect 28684 23624 28724 23752
rect 28780 23792 28820 24340
rect 29452 24296 29492 27532
rect 29932 27572 29972 27581
rect 29932 25724 29972 27532
rect 30316 27488 30356 27497
rect 29932 25675 29972 25684
rect 30028 25976 30068 25985
rect 29548 24632 29588 24641
rect 29548 24497 29588 24592
rect 29452 24247 29492 24256
rect 29932 24464 29972 24473
rect 28780 23743 28820 23752
rect 29356 23792 29396 23801
rect 28588 21608 28628 21617
rect 28588 21020 28628 21568
rect 28588 20971 28628 20980
rect 28492 20719 28532 20728
rect 28588 20852 28628 20861
rect 28588 19844 28628 20812
rect 28588 19795 28628 19804
rect 28492 19172 28532 19181
rect 28492 18752 28532 19132
rect 28492 18703 28532 18712
rect 28588 19088 28628 19097
rect 28108 17611 28148 17620
rect 28300 17788 28396 17828
rect 28300 17660 28340 17788
rect 28396 17779 28436 17788
rect 28588 17744 28628 19048
rect 28588 17695 28628 17704
rect 27674 17408 28042 17417
rect 27674 17359 28042 17368
rect 27340 16232 27380 16241
rect 27340 15896 27380 16192
rect 27340 15847 27380 15856
rect 27674 15896 28042 15905
rect 27674 15847 28042 15856
rect 27436 15560 27476 15569
rect 27244 15520 27436 15560
rect 26188 14923 26228 14932
rect 26764 14932 26900 14972
rect 26956 15476 26996 15485
rect 26092 14167 26132 14176
rect 26668 14720 26708 14729
rect 26188 14048 26228 14057
rect 25996 14008 26132 14048
rect 25900 13411 25940 13420
rect 25900 13208 25940 13217
rect 25804 13124 25844 13133
rect 25804 12989 25844 13084
rect 25708 12704 25748 12713
rect 25708 12569 25748 12664
rect 25900 12704 25940 13168
rect 25900 12655 25940 12664
rect 25708 12452 25748 12461
rect 25708 11948 25748 12412
rect 25708 11899 25748 11908
rect 25804 12368 25844 12377
rect 25804 11276 25844 12328
rect 26092 11948 26132 14008
rect 26188 12704 26228 14008
rect 26284 13880 26324 13889
rect 26284 13292 26324 13840
rect 26668 13880 26708 14680
rect 26764 14636 26804 14932
rect 26764 14587 26804 14596
rect 26860 14804 26900 14813
rect 26668 13831 26708 13840
rect 26860 13964 26900 14764
rect 26434 13628 26802 13637
rect 26434 13579 26802 13588
rect 26764 13376 26804 13385
rect 26284 13252 26420 13292
rect 26380 12788 26420 13252
rect 26284 12704 26324 12713
rect 26188 12664 26284 12704
rect 26284 12655 26324 12664
rect 26380 12536 26420 12748
rect 26476 12536 26516 12545
rect 26380 12496 26476 12536
rect 26476 12487 26516 12496
rect 26764 12536 26804 13336
rect 26860 13292 26900 13924
rect 26956 13460 26996 15436
rect 27052 14216 27092 15520
rect 27052 14167 27092 14176
rect 27148 14804 27188 14813
rect 27148 14720 27188 14764
rect 27148 14300 27188 14680
rect 26956 13411 26996 13420
rect 27052 14048 27092 14057
rect 26860 13243 26900 13252
rect 27052 13208 27092 14008
rect 27148 13964 27188 14260
rect 27244 14720 27284 14729
rect 27244 14216 27284 14680
rect 27244 14167 27284 14176
rect 27148 13915 27188 13924
rect 27340 14132 27380 14141
rect 27340 13796 27380 14092
rect 27340 13747 27380 13756
rect 27052 13159 27092 13168
rect 27340 13208 27380 13217
rect 27052 12956 27092 12965
rect 26188 12452 26228 12461
rect 26188 12032 26228 12412
rect 26764 12401 26804 12496
rect 26860 12704 26900 12715
rect 26860 12620 26900 12664
rect 26434 12116 26802 12125
rect 26434 12067 26802 12076
rect 26188 11983 26228 11992
rect 26092 11899 26132 11908
rect 26860 11864 26900 12580
rect 26956 12704 26996 12713
rect 26956 12620 26996 12664
rect 26956 12569 26996 12580
rect 27052 12620 27092 12916
rect 27244 12788 27284 12797
rect 27244 12620 27284 12748
rect 27092 12580 27188 12620
rect 27052 12571 27092 12580
rect 26860 11824 26996 11864
rect 26188 11780 26228 11791
rect 26188 11696 26228 11740
rect 26860 11696 26900 11705
rect 26228 11656 26324 11696
rect 26188 11647 26228 11656
rect 25804 11236 25940 11276
rect 25612 9799 25652 9808
rect 25804 10436 25844 10445
rect 25804 9596 25844 10396
rect 25804 9547 25844 9556
rect 25036 9377 25076 9472
rect 25900 9512 25940 11236
rect 25900 9377 25940 9472
rect 25996 11024 26036 11033
rect 24844 8791 24884 8800
rect 25996 8840 26036 10984
rect 24940 8756 24980 8765
rect 24940 8672 24980 8716
rect 24940 8621 24980 8632
rect 25036 8252 25076 8261
rect 24652 7916 24692 7925
rect 24652 7328 24692 7876
rect 24652 7279 24692 7288
rect 25036 7160 25076 8212
rect 25996 8000 26036 8800
rect 25996 7951 26036 7960
rect 26284 9428 26324 11656
rect 26860 11192 26900 11656
rect 26860 11143 26900 11152
rect 26956 11108 26996 11824
rect 26956 11059 26996 11068
rect 26434 10604 26802 10613
rect 26434 10555 26802 10564
rect 27052 10016 27092 10025
rect 27052 9764 27092 9976
rect 26860 9596 26900 9605
rect 26860 9512 26900 9556
rect 26860 9461 26900 9472
rect 25036 7111 25076 7120
rect 26284 7160 26324 9388
rect 27052 9428 27092 9724
rect 26956 9344 26996 9353
rect 26860 9260 26900 9269
rect 26434 9092 26802 9101
rect 26434 9043 26802 9052
rect 26572 8840 26612 8849
rect 26572 7916 26612 8800
rect 26860 8084 26900 9220
rect 26956 8672 26996 9304
rect 26956 8623 26996 8632
rect 26860 8035 26900 8044
rect 26572 7867 26612 7876
rect 26434 7580 26802 7589
rect 26434 7531 26802 7540
rect 26284 7111 26324 7120
rect 26764 7244 26804 7253
rect 26764 6656 26804 7204
rect 26764 6607 26804 6616
rect 25228 6488 25268 6497
rect 24940 6404 24980 6413
rect 24940 5480 24980 6364
rect 25228 5900 25268 6448
rect 25612 6404 25652 6413
rect 25228 5851 25268 5860
rect 25516 6320 25556 6329
rect 25516 5648 25556 6280
rect 25612 5900 25652 6364
rect 25612 5851 25652 5860
rect 25996 6236 26036 6245
rect 25516 5599 25556 5608
rect 25996 5648 26036 6196
rect 26434 6068 26802 6077
rect 26434 6019 26802 6028
rect 25996 5599 26036 5608
rect 24940 5431 24980 5440
rect 24556 5347 24596 5356
rect 25708 4976 25748 4985
rect 24844 4892 24884 4901
rect 24844 3968 24884 4852
rect 24844 3919 24884 3928
rect 25420 4136 25460 4145
rect 25420 3884 25460 4096
rect 25324 3716 25364 3725
rect 24940 3464 24980 3473
rect 24940 3128 24980 3424
rect 24940 3079 24980 3088
rect 24268 1868 24308 2248
rect 25228 2624 25268 2633
rect 24268 1819 24308 1828
rect 24460 1952 24500 1961
rect 24460 1364 24500 1912
rect 24460 1315 24500 1324
rect 25228 1196 25268 2584
rect 25324 1952 25364 3676
rect 25420 3632 25460 3844
rect 25420 3583 25460 3592
rect 25708 3296 25748 4936
rect 26092 4976 26132 4985
rect 26092 4388 26132 4936
rect 26434 4556 26802 4565
rect 26434 4507 26802 4516
rect 26092 4339 26132 4348
rect 26380 4220 26420 4229
rect 25804 4052 25844 4061
rect 25804 3632 25844 4012
rect 26380 3716 26420 4180
rect 26476 4136 26516 4145
rect 26476 4001 26516 4096
rect 26572 4052 26612 4061
rect 26380 3667 26420 3676
rect 25804 3583 25844 3592
rect 26572 3632 26612 4012
rect 26572 3583 26612 3592
rect 27052 3464 27092 9388
rect 27148 5648 27188 12580
rect 27244 12571 27284 12580
rect 27340 11696 27380 13168
rect 27436 12872 27476 15520
rect 27820 14888 27860 14897
rect 27436 12823 27476 12832
rect 27532 14720 27572 14729
rect 27532 12704 27572 14680
rect 27820 14720 27860 14848
rect 27820 14671 27860 14680
rect 27674 14384 28042 14393
rect 27674 14335 28042 14344
rect 27628 14048 27668 14057
rect 27628 13796 27668 14008
rect 27628 13747 27668 13756
rect 28108 13292 28148 13301
rect 27674 12872 28042 12881
rect 27674 12823 28042 12832
rect 27532 12655 27572 12664
rect 28108 12620 28148 13252
rect 28108 12571 28148 12580
rect 27340 11647 27380 11656
rect 27436 12536 27476 12545
rect 27340 11528 27380 11537
rect 27340 11024 27380 11488
rect 27340 10975 27380 10984
rect 27436 10184 27476 12496
rect 27820 12452 27860 12461
rect 27340 10016 27380 10025
rect 27244 9512 27284 9521
rect 27340 9512 27380 9976
rect 27436 9848 27476 10144
rect 27436 9799 27476 9808
rect 27532 11696 27572 11705
rect 27532 10352 27572 11656
rect 27820 11696 27860 12412
rect 28204 12452 28244 12461
rect 28204 11780 28244 12412
rect 28204 11731 28244 11740
rect 27820 11647 27860 11656
rect 28300 11696 28340 17620
rect 28396 16988 28436 16997
rect 28396 16400 28436 16948
rect 28396 16351 28436 16360
rect 28684 15812 28724 23584
rect 29356 23288 29396 23752
rect 29356 23120 29396 23248
rect 29356 23071 29396 23080
rect 29932 23036 29972 24424
rect 30028 23876 30068 25936
rect 30316 25388 30356 27448
rect 30316 25339 30356 25348
rect 30412 27404 30452 27413
rect 30028 23827 30068 23836
rect 29932 22987 29972 22996
rect 28972 22784 29012 22793
rect 28780 22112 28820 22121
rect 28780 21524 28820 22072
rect 28972 21776 29012 22744
rect 30124 22700 30164 22709
rect 28972 21727 29012 21736
rect 29452 22280 29492 22289
rect 29452 21776 29492 22240
rect 30124 22280 30164 22660
rect 30220 22616 30260 22625
rect 30220 22364 30260 22576
rect 30220 22315 30260 22324
rect 29452 21727 29492 21736
rect 30028 21776 30068 21787
rect 30028 21692 30068 21736
rect 30028 21643 30068 21652
rect 28780 21475 28820 21484
rect 29644 21608 29684 21617
rect 28780 21356 28820 21365
rect 28780 20852 28820 21316
rect 29644 21020 29684 21568
rect 30124 21272 30164 22240
rect 30412 21860 30452 27364
rect 30796 27068 30836 28600
rect 30796 27019 30836 27028
rect 31084 27488 31124 27497
rect 31084 26900 31124 27448
rect 31084 26851 31124 26860
rect 30892 26816 30932 26825
rect 30892 25304 30932 26776
rect 31180 26144 31220 26153
rect 30604 24464 30644 24473
rect 30412 21811 30452 21820
rect 30508 23204 30548 23213
rect 30124 21223 30164 21232
rect 30220 21776 30260 21785
rect 30220 21440 30260 21736
rect 29644 20971 29684 20980
rect 28780 20803 28820 20812
rect 30220 20768 30260 21400
rect 30220 20719 30260 20728
rect 30508 21608 30548 23164
rect 29452 20096 29492 20105
rect 28876 20012 28916 20021
rect 28780 19844 28820 19853
rect 28780 18668 28820 19804
rect 28780 18619 28820 18628
rect 28876 18584 28916 19972
rect 29452 18752 29492 20056
rect 30316 20096 30356 20105
rect 30316 19508 30356 20056
rect 30508 20096 30548 21568
rect 30604 20852 30644 24424
rect 30796 22784 30836 22793
rect 30796 22364 30836 22744
rect 30796 22315 30836 22324
rect 30892 21776 30932 25264
rect 30892 21727 30932 21736
rect 30988 26060 31028 26069
rect 30988 23288 31028 26020
rect 30988 21608 31028 23248
rect 31084 25976 31124 25985
rect 31084 22280 31124 25936
rect 31084 22028 31124 22240
rect 31084 21979 31124 21988
rect 30988 21559 31028 21568
rect 30604 20803 30644 20812
rect 31180 20264 31220 26104
rect 31276 24548 31316 24557
rect 31276 24044 31316 24508
rect 31276 23995 31316 24004
rect 31180 20215 31220 20224
rect 30508 20047 30548 20056
rect 30316 19459 30356 19468
rect 30892 20012 30932 20021
rect 29452 18703 29492 18712
rect 29836 19340 29876 19349
rect 28876 18535 28916 18544
rect 29836 17912 29876 19300
rect 29836 17863 29876 17872
rect 30892 19256 30932 19972
rect 30892 18584 30932 19216
rect 30892 17156 30932 18544
rect 30988 18500 31028 18509
rect 30988 17912 31028 18460
rect 30988 17863 31028 17872
rect 28684 15763 28724 15772
rect 30412 16904 30452 16913
rect 30412 15476 30452 16864
rect 30604 16904 30644 16913
rect 30604 16316 30644 16864
rect 30604 16267 30644 16276
rect 30892 16232 30932 17116
rect 31276 17576 31316 17585
rect 31276 16316 31316 17536
rect 31276 16267 31316 16276
rect 30892 16183 30932 16192
rect 30412 15427 30452 15436
rect 30892 15560 30932 15569
rect 28876 15308 28916 15317
rect 28396 14888 28436 14897
rect 28396 13292 28436 14848
rect 28588 14888 28628 14897
rect 28492 14720 28532 14729
rect 28492 14585 28532 14680
rect 28396 13243 28436 13252
rect 28588 14048 28628 14848
rect 28876 14720 28916 15268
rect 29356 15308 29396 15317
rect 28876 14671 28916 14680
rect 28972 14804 29012 14844
rect 28972 14720 29012 14764
rect 28396 12704 28436 12713
rect 28396 12620 28436 12664
rect 28588 12704 28628 14008
rect 28972 13964 29012 14680
rect 29356 14636 29396 15268
rect 29356 14587 29396 14596
rect 30508 14720 30548 14729
rect 28972 13915 29012 13924
rect 28780 13880 28820 13889
rect 28780 13208 28820 13840
rect 30508 13796 30548 14680
rect 29932 13376 29972 13385
rect 28780 13159 28820 13168
rect 28972 13208 29012 13217
rect 28588 12655 28628 12664
rect 28396 12569 28436 12580
rect 28300 11647 28340 11656
rect 28396 12452 28436 12461
rect 28204 11612 28244 11621
rect 27674 11360 28042 11369
rect 27674 11311 28042 11320
rect 28108 11024 28148 11033
rect 28108 10889 28148 10984
rect 27436 9680 27476 9689
rect 27532 9680 27572 10312
rect 28108 10184 28148 10193
rect 27674 9848 28042 9857
rect 27674 9799 28042 9808
rect 27476 9640 27572 9680
rect 27628 9680 27668 9689
rect 27436 9631 27476 9640
rect 27284 9472 27380 9512
rect 27532 9512 27572 9521
rect 27244 9463 27284 9472
rect 27532 8924 27572 9472
rect 27532 8875 27572 8884
rect 27628 8660 27668 9640
rect 28108 9680 28148 10144
rect 28108 9631 28148 9640
rect 28108 9512 28148 9521
rect 28204 9512 28244 11572
rect 28148 9472 28244 9512
rect 28108 9463 28148 9472
rect 27532 8620 27668 8660
rect 28108 8672 28148 8681
rect 27532 7244 27572 8620
rect 27674 8336 28042 8345
rect 27674 8287 28042 8296
rect 27340 6404 27380 6413
rect 27188 5608 27284 5648
rect 27148 5599 27188 5608
rect 27244 5060 27284 5608
rect 27148 4976 27188 4985
rect 27148 4220 27188 4936
rect 27244 4724 27284 5020
rect 27244 4675 27284 4684
rect 27148 3716 27188 4180
rect 27340 4052 27380 6364
rect 27532 5228 27572 7204
rect 28108 8168 28148 8632
rect 28108 7160 28148 8128
rect 28108 7111 28148 7120
rect 28204 7076 28244 9472
rect 28300 10268 28340 10277
rect 28300 9596 28340 10228
rect 28300 9344 28340 9556
rect 28300 9295 28340 9304
rect 28396 7916 28436 12412
rect 28492 12368 28532 12377
rect 28492 11696 28532 12328
rect 28972 11780 29012 13168
rect 29932 12452 29972 13336
rect 30508 12980 30548 13756
rect 29932 12403 29972 12412
rect 30316 12940 30548 12980
rect 30604 14048 30644 14057
rect 30604 13208 30644 14008
rect 30892 14048 30932 15520
rect 30892 13999 30932 14008
rect 31084 14888 31124 14897
rect 31084 13964 31124 14848
rect 31084 13915 31124 13924
rect 28972 11731 29012 11740
rect 28492 10856 28532 11656
rect 28780 11696 28820 11705
rect 28684 11612 28724 11621
rect 28492 10807 28532 10816
rect 28588 11528 28628 11537
rect 28588 11108 28628 11488
rect 28588 10100 28628 11068
rect 28396 7867 28436 7876
rect 28492 10060 28628 10100
rect 28396 7412 28436 7421
rect 27674 6824 28042 6833
rect 27674 6775 28042 6784
rect 27820 6488 27860 6497
rect 27820 5984 27860 6448
rect 27820 5935 27860 5944
rect 28012 6404 28052 6413
rect 28012 5648 28052 6364
rect 28012 5599 28052 5608
rect 28108 5648 28148 5657
rect 27674 5312 28042 5321
rect 27674 5263 28042 5272
rect 27340 4003 27380 4012
rect 27436 5188 27532 5228
rect 27436 4136 27476 5188
rect 27532 5179 27572 5188
rect 27436 4001 27476 4096
rect 27532 5060 27572 5069
rect 27148 3667 27188 3676
rect 27052 3415 27092 3424
rect 27532 3464 27572 5020
rect 28012 4976 28052 5004
rect 28108 4976 28148 5608
rect 28052 4936 28148 4976
rect 28012 4927 28052 4936
rect 28012 4472 28052 4481
rect 28012 4220 28052 4432
rect 28012 4171 28052 4180
rect 27674 3800 28042 3809
rect 27674 3751 28042 3760
rect 25708 2624 25748 3256
rect 26434 3044 26802 3053
rect 26434 2995 26802 3004
rect 26860 2792 26900 2801
rect 25804 2624 25844 2633
rect 25708 2584 25804 2624
rect 25804 2575 25844 2584
rect 25324 1280 25364 1912
rect 25324 1231 25364 1240
rect 25996 2540 26036 2549
rect 25228 1147 25268 1156
rect 24076 1063 24116 1072
rect 25996 1112 26036 2500
rect 26860 1868 26900 2752
rect 26860 1819 26900 1828
rect 27532 2120 27572 3424
rect 27674 2288 28042 2297
rect 27674 2239 28042 2248
rect 26434 1532 26802 1541
rect 26434 1483 26802 1492
rect 25996 1063 26036 1072
rect 27532 1112 27572 2080
rect 28108 1868 28148 4936
rect 28204 4640 28244 7036
rect 28300 7076 28340 7085
rect 28300 6488 28340 7036
rect 28396 6572 28436 7372
rect 28396 6523 28436 6532
rect 28300 6439 28340 6448
rect 28204 4591 28244 4600
rect 28300 4976 28340 4985
rect 28300 4304 28340 4936
rect 28492 4808 28532 10060
rect 28684 9680 28724 11572
rect 28780 11192 28820 11656
rect 28780 11143 28820 11152
rect 29356 11024 29396 11033
rect 28684 9631 28724 9640
rect 29068 10772 29108 10781
rect 29068 10184 29108 10732
rect 29356 10772 29396 10984
rect 29356 10723 29396 10732
rect 29548 10940 29588 10949
rect 29548 10436 29588 10900
rect 29548 10387 29588 10396
rect 28972 9344 29012 9353
rect 28972 8924 29012 9304
rect 28972 8875 29012 8884
rect 28876 8756 28916 8765
rect 28780 8504 28820 8513
rect 28780 7244 28820 8464
rect 28876 8168 28916 8716
rect 28876 8119 28916 8128
rect 28780 7195 28820 7204
rect 28876 7328 28916 7337
rect 28780 7076 28820 7085
rect 28780 6941 28820 7036
rect 28780 6488 28820 6497
rect 28780 6152 28820 6448
rect 28780 6103 28820 6112
rect 28876 5564 28916 7288
rect 28876 5515 28916 5524
rect 29068 4976 29108 10144
rect 29356 9932 29396 9941
rect 29356 9428 29396 9892
rect 30220 9596 30260 9605
rect 30220 9461 30260 9556
rect 29356 8672 29396 9388
rect 30124 8756 30164 8765
rect 29356 8623 29396 8632
rect 29836 8672 29876 8681
rect 29836 8168 29876 8632
rect 29836 8119 29876 8128
rect 30124 8168 30164 8716
rect 30124 8119 30164 8128
rect 29932 8084 29972 8093
rect 29836 7916 29876 7925
rect 29740 7328 29780 7337
rect 29644 7160 29684 7169
rect 29260 7076 29300 7085
rect 29164 6992 29204 7001
rect 29164 6572 29204 6952
rect 29164 5816 29204 6532
rect 29164 5767 29204 5776
rect 29260 6404 29300 7036
rect 29548 7076 29588 7085
rect 29548 6656 29588 7036
rect 29260 6152 29300 6364
rect 29068 4927 29108 4936
rect 28492 4759 28532 4768
rect 28588 4892 28628 4901
rect 28300 4255 28340 4264
rect 28204 4052 28244 4061
rect 28204 3716 28244 4012
rect 28204 3667 28244 3676
rect 28588 3548 28628 4852
rect 28588 3499 28628 3508
rect 28780 3968 28820 3977
rect 28204 3464 28244 3473
rect 28204 2624 28244 3424
rect 28780 3464 28820 3928
rect 28780 3415 28820 3424
rect 28876 3548 28916 3557
rect 28204 2575 28244 2584
rect 28780 3212 28820 3221
rect 28780 2540 28820 3172
rect 28876 2876 28916 3508
rect 29260 3212 29300 6112
rect 29452 6572 29492 6581
rect 29452 5648 29492 6532
rect 29452 5396 29492 5608
rect 29548 5564 29588 6616
rect 29644 5984 29684 7120
rect 29644 5935 29684 5944
rect 29740 5732 29780 7288
rect 29836 5816 29876 7876
rect 29836 5767 29876 5776
rect 29740 5683 29780 5692
rect 29548 5515 29588 5524
rect 29644 5648 29684 5657
rect 29644 5513 29684 5608
rect 29452 5347 29492 5356
rect 29356 4976 29396 4985
rect 29356 4304 29396 4936
rect 29356 3632 29396 4264
rect 29740 4136 29780 4145
rect 29740 3716 29780 4096
rect 29740 3667 29780 3676
rect 29356 3583 29396 3592
rect 29356 3212 29396 3221
rect 29260 3172 29356 3212
rect 28876 2827 28916 2836
rect 29356 2708 29396 3172
rect 29932 2900 29972 8044
rect 30028 8000 30068 8009
rect 30028 7412 30068 7960
rect 30316 8000 30356 12940
rect 30604 12536 30644 13168
rect 30412 10772 30452 10781
rect 30412 10100 30452 10732
rect 30604 10268 30644 12496
rect 30700 13292 30740 13301
rect 30700 12200 30740 13252
rect 30700 11696 30740 12160
rect 30700 11647 30740 11656
rect 31276 11864 31316 11873
rect 31180 11612 31220 11621
rect 30604 10219 30644 10228
rect 30892 11024 30932 11033
rect 30412 10051 30452 10060
rect 30508 10184 30548 10193
rect 30508 9596 30548 10144
rect 30316 7951 30356 7960
rect 30412 9512 30452 9521
rect 30412 8504 30452 9472
rect 30508 8672 30548 9556
rect 30892 9512 30932 10984
rect 30892 9463 30932 9472
rect 30988 10940 31028 10949
rect 30988 8840 31028 10900
rect 31180 9596 31220 11572
rect 31276 11108 31316 11824
rect 31276 11059 31316 11068
rect 31180 9547 31220 9556
rect 30988 8791 31028 8800
rect 31084 9428 31124 9437
rect 30508 8623 30548 8632
rect 30028 7363 30068 7372
rect 30316 7244 30356 7253
rect 30028 7160 30068 7169
rect 30028 5900 30068 7120
rect 30028 5851 30068 5860
rect 30124 7076 30164 7085
rect 30124 5648 30164 7036
rect 30124 5513 30164 5608
rect 30316 5564 30356 7204
rect 30316 5515 30356 5524
rect 30316 4724 30356 4733
rect 30220 4304 30260 4313
rect 30220 3380 30260 4264
rect 30316 4136 30356 4684
rect 30316 4087 30356 4096
rect 30220 3331 30260 3340
rect 30412 3464 30452 8464
rect 31084 7832 31124 9388
rect 31084 7783 31124 7792
rect 30604 7748 30644 7757
rect 30604 7244 30644 7708
rect 30604 7195 30644 7204
rect 30700 7160 30740 7169
rect 30604 6488 30644 6497
rect 30508 6404 30548 6413
rect 30508 5144 30548 6364
rect 30604 5900 30644 6448
rect 30604 5851 30644 5860
rect 30508 5095 30548 5104
rect 30508 4976 30548 4985
rect 30508 4052 30548 4936
rect 30700 4220 30740 7120
rect 30892 6152 30932 6161
rect 30892 5648 30932 6112
rect 30892 5599 30932 5608
rect 30700 4171 30740 4180
rect 30508 4003 30548 4012
rect 29356 2659 29396 2668
rect 29836 2860 29972 2900
rect 28780 2491 28820 2500
rect 28108 1819 28148 1828
rect 29836 1952 29876 2860
rect 29836 1364 29876 1912
rect 29836 1315 29876 1324
rect 30316 2792 30356 2801
rect 30316 1196 30356 2752
rect 30316 1147 30356 1156
rect 27532 1063 27572 1072
rect 30412 1112 30452 3424
rect 30988 1952 31028 1961
rect 30988 1784 31028 1912
rect 30988 1735 31028 1744
rect 30796 1700 30836 1709
rect 30796 1196 30836 1660
rect 30796 1147 30836 1156
rect 30412 1063 30452 1072
rect 23308 979 23348 988
rect 15052 811 15092 820
rect 5740 727 5780 736
rect 12126 776 12494 785
rect 12126 727 12494 736
rect 19900 776 20268 785
rect 19900 727 20268 736
rect 27674 776 28042 785
rect 27674 727 28042 736
<< via3 >>
rect 3112 27196 3480 27236
rect 4352 27952 4720 27992
rect 4352 26440 4720 26480
rect 3112 25684 3480 25724
rect 4352 24928 4720 24968
rect 3112 24172 3480 24212
rect 3112 22660 3480 22700
rect 556 20476 596 20516
rect 268 16444 308 16484
rect 1708 19216 1748 19256
rect 1036 16192 1076 16232
rect 1612 16276 1652 16316
rect 2284 20812 2324 20852
rect 2188 19300 2228 19340
rect 2092 19216 2132 19256
rect 2092 18796 2132 18836
rect 1804 16276 1844 16316
rect 2476 18544 2516 18584
rect 2188 17200 2228 17240
rect 3112 21148 3480 21188
rect 3148 20224 3188 20264
rect 3340 20056 3380 20096
rect 2860 19720 2900 19760
rect 3112 19636 3480 19676
rect 2668 19300 2708 19340
rect 3148 19300 3188 19340
rect 5068 24424 5108 24464
rect 5644 24760 5684 24800
rect 4352 23416 4720 23456
rect 4352 21904 4720 21944
rect 3916 20644 3956 20684
rect 2668 18544 2708 18584
rect 2668 17788 2708 17828
rect 2188 16192 2228 16232
rect 3148 18796 3188 18836
rect 3112 18124 3480 18164
rect 2956 18040 2996 18080
rect 4684 21568 4724 21608
rect 4300 20812 4340 20852
rect 4204 20728 4244 20768
rect 4352 20392 4720 20432
rect 4204 20056 4244 20096
rect 4300 19972 4340 20012
rect 4588 19720 4628 19760
rect 5356 21568 5396 21608
rect 5356 20980 5396 21020
rect 4352 18880 4720 18920
rect 3532 17704 3572 17744
rect 3112 16612 3480 16652
rect 3916 17704 3956 17744
rect 4684 17536 4724 17576
rect 4352 17368 4720 17408
rect 3112 15100 3480 15140
rect 3436 14596 3476 14636
rect 3112 13588 3480 13628
rect 3724 15772 3764 15812
rect 2572 11236 2612 11276
rect 3112 12076 3480 12116
rect 2284 10396 2324 10436
rect 3112 10564 3480 10604
rect 2380 9640 2420 9680
rect 3532 10144 3572 10184
rect 3112 9052 3480 9092
rect 3112 7540 3480 7580
rect 2860 7120 2900 7160
rect 4492 17200 4532 17240
rect 5164 18040 5204 18080
rect 4684 16024 4724 16064
rect 4352 15856 4720 15896
rect 4492 15688 4532 15728
rect 4108 14428 4148 14468
rect 4108 14176 4148 14216
rect 4352 14344 4720 14384
rect 4876 13504 4916 13544
rect 4352 12832 4720 12872
rect 4352 11320 4720 11360
rect 4204 11152 4244 11192
rect 4876 13252 4916 13292
rect 5260 17788 5300 17828
rect 5452 20644 5492 20684
rect 5740 20056 5780 20096
rect 5644 18628 5684 18668
rect 8332 26272 8372 26312
rect 8908 26272 8948 26312
rect 10348 27364 10388 27404
rect 10060 26272 10100 26312
rect 9964 26104 10004 26144
rect 10156 26104 10196 26144
rect 5452 16192 5492 16232
rect 5452 15436 5492 15476
rect 4300 11068 4340 11108
rect 4876 11068 4916 11108
rect 4396 10984 4436 11024
rect 4492 10900 4532 10940
rect 3112 6028 3480 6068
rect 3112 4516 3480 4556
rect 4684 10228 4724 10268
rect 4588 10144 4628 10184
rect 4972 10144 5012 10184
rect 5452 14260 5492 14300
rect 5260 13252 5300 13292
rect 5164 10984 5204 11024
rect 6028 15352 6068 15392
rect 5740 14680 5780 14720
rect 5644 14176 5684 14216
rect 5932 14596 5972 14636
rect 6700 20056 6740 20096
rect 6604 18628 6644 18668
rect 6892 18460 6932 18500
rect 6892 17788 6932 17828
rect 6796 16276 6836 16316
rect 6316 16024 6356 16064
rect 6028 14176 6068 14216
rect 5644 13252 5684 13292
rect 5548 13168 5588 13208
rect 4352 9808 4720 9848
rect 5548 9640 5588 9680
rect 5836 13336 5876 13376
rect 5836 11740 5876 11780
rect 5644 9556 5684 9596
rect 6508 15436 6548 15476
rect 6220 14596 6260 14636
rect 6124 13336 6164 13376
rect 6220 13420 6260 13460
rect 6028 11740 6068 11780
rect 4352 8296 4720 8336
rect 4108 6952 4148 6992
rect 3112 3004 3480 3044
rect 4492 6952 4532 6992
rect 4780 6952 4820 6992
rect 4972 7120 5012 7160
rect 4352 6784 4720 6824
rect 4352 5272 4720 5312
rect 4352 3760 4720 3800
rect 4352 2248 4720 2288
rect 3112 1492 3480 1532
rect 6412 13168 6452 13208
rect 6892 15856 6932 15896
rect 6988 16276 7028 16316
rect 6892 15436 6932 15476
rect 6604 12916 6644 12956
rect 6700 11740 6740 11780
rect 6316 11320 6356 11360
rect 6508 11236 6548 11276
rect 6892 13252 6932 13292
rect 7372 19972 7412 20012
rect 7756 20056 7796 20096
rect 7084 15940 7124 15980
rect 7276 15520 7316 15560
rect 7084 14596 7124 14636
rect 6796 11320 6836 11360
rect 6796 10312 6836 10352
rect 6508 10228 6548 10268
rect 7564 16192 7604 16232
rect 7756 15940 7796 15980
rect 7564 15856 7604 15896
rect 7180 13000 7220 13040
rect 7084 11656 7124 11696
rect 7564 13420 7604 13460
rect 7564 13168 7604 13208
rect 7564 12412 7604 12452
rect 9100 25516 9140 25556
rect 10060 25936 10100 25976
rect 9868 25852 9908 25892
rect 9772 24424 9812 24464
rect 8044 15772 8084 15812
rect 8044 15604 8084 15644
rect 8044 15352 8084 15392
rect 7852 14428 7892 14468
rect 7660 12496 7700 12536
rect 7276 11488 7316 11528
rect 6892 10144 6932 10184
rect 6316 9976 6356 10016
rect 6700 9892 6740 9932
rect 6988 10228 7028 10268
rect 6988 9976 7028 10016
rect 6892 9892 6932 9932
rect 6700 7960 6740 8000
rect 7372 9808 7412 9848
rect 7660 10816 7700 10856
rect 7564 10564 7604 10604
rect 8044 13504 8084 13544
rect 8140 13168 8180 13208
rect 8524 16444 8564 16484
rect 8428 16192 8468 16232
rect 9292 19132 9332 19172
rect 8524 16024 8564 16064
rect 8524 14428 8564 14468
rect 8908 16864 8948 16904
rect 8716 13336 8756 13376
rect 8524 13252 8564 13292
rect 8332 13168 8372 13208
rect 8332 12496 8372 12536
rect 8332 12328 8372 12368
rect 8236 11656 8276 11696
rect 8332 10984 8372 11024
rect 8524 12412 8564 12452
rect 8716 12916 8756 12956
rect 8620 11488 8660 11528
rect 8044 9724 8084 9764
rect 7948 9556 7988 9596
rect 8716 11152 8756 11192
rect 8620 10480 8660 10520
rect 8524 10312 8564 10352
rect 8620 10228 8660 10268
rect 8428 9976 8468 10016
rect 8332 9892 8372 9932
rect 8716 9724 8756 9764
rect 5260 4096 5300 4136
rect 6316 4936 6356 4976
rect 4352 736 4720 776
rect 7276 4096 7316 4136
rect 7852 7960 7892 8000
rect 8908 15436 8948 15476
rect 9196 15688 9236 15728
rect 9484 17368 9524 17408
rect 9484 16780 9524 16820
rect 9772 18460 9812 18500
rect 9100 15436 9140 15476
rect 8908 13336 8948 13376
rect 8908 12328 8948 12368
rect 9100 13084 9140 13124
rect 9676 14680 9716 14720
rect 9580 14596 9620 14636
rect 9100 10816 9140 10856
rect 9004 10312 9044 10352
rect 9004 10144 9044 10184
rect 9004 9976 9044 10016
rect 9676 12496 9716 12536
rect 9292 10396 9332 10436
rect 9196 10144 9236 10184
rect 9196 9640 9236 9680
rect 8620 5020 8660 5060
rect 8428 4936 8468 4976
rect 9772 10900 9812 10940
rect 10060 23836 10100 23876
rect 10060 20140 10100 20180
rect 9964 19132 10004 19172
rect 10060 17200 10100 17240
rect 9964 16192 10004 16232
rect 10060 16024 10100 16064
rect 9964 15604 10004 15644
rect 9964 15352 10004 15392
rect 10060 14764 10100 14804
rect 12126 27952 12494 27992
rect 10828 27364 10868 27404
rect 10886 27196 11254 27236
rect 10540 25684 10580 25724
rect 10540 25516 10580 25556
rect 10444 25180 10484 25220
rect 10444 24760 10484 24800
rect 10252 14932 10292 14972
rect 10444 16192 10484 16232
rect 10886 25684 11254 25724
rect 11116 25516 11156 25556
rect 10828 25264 10868 25304
rect 11116 25180 11156 25220
rect 11116 24508 11156 24548
rect 10886 24172 11254 24212
rect 11116 22912 11156 22952
rect 10886 22660 11254 22700
rect 11212 22492 11252 22532
rect 11500 25600 11540 25640
rect 11692 23164 11732 23204
rect 11500 22912 11540 22952
rect 11596 22492 11636 22532
rect 12126 26440 12494 26480
rect 12556 26440 12596 26480
rect 12460 25936 12500 25976
rect 11980 25852 12020 25892
rect 12940 26440 12980 26480
rect 12940 26104 12980 26144
rect 12940 25936 12980 25976
rect 11884 23248 11924 23288
rect 12126 24928 12494 24968
rect 12652 24508 12692 24548
rect 12556 23836 12596 23876
rect 12126 23416 12494 23456
rect 12460 23248 12500 23288
rect 10886 21148 11254 21188
rect 11500 20980 11540 21020
rect 10886 19636 11254 19676
rect 11500 19300 11540 19340
rect 11212 18544 11252 18584
rect 12556 23080 12596 23120
rect 12364 22240 12404 22280
rect 12126 21904 12494 21944
rect 12844 22156 12884 22196
rect 11884 20728 11924 20768
rect 14380 26104 14420 26144
rect 13324 22240 13364 22280
rect 12126 20392 12494 20432
rect 11884 19216 11924 19256
rect 12460 19300 12500 19340
rect 11500 18544 11540 18584
rect 10886 18124 11254 18164
rect 10636 17368 10676 17408
rect 10540 15688 10580 15728
rect 10828 17368 10868 17408
rect 11404 17200 11444 17240
rect 10828 17032 10868 17072
rect 11020 16864 11060 16904
rect 11212 16948 11252 16988
rect 10886 16612 11254 16652
rect 10540 15520 10580 15560
rect 10252 14764 10292 14804
rect 10732 15352 10772 15392
rect 11116 15268 11156 15308
rect 10886 15100 11254 15140
rect 10732 14932 10772 14972
rect 9964 11740 10004 11780
rect 10156 10816 10196 10856
rect 9388 9808 9428 9848
rect 10060 10060 10100 10100
rect 10886 13588 11254 13628
rect 11116 13420 11156 13460
rect 10828 12412 10868 12452
rect 11020 12412 11060 12452
rect 11116 12244 11156 12284
rect 10732 12160 10772 12200
rect 10540 11656 10580 11696
rect 10540 10648 10580 10688
rect 10886 12076 11254 12116
rect 11020 10984 11060 11024
rect 12126 18880 12494 18920
rect 11692 16780 11732 16820
rect 12126 17368 12494 17408
rect 11884 17032 11924 17072
rect 12652 16780 12692 16820
rect 12556 16696 12596 16736
rect 12940 20644 12980 20684
rect 13324 20644 13364 20684
rect 15820 23080 15860 23120
rect 15244 22156 15284 22196
rect 14092 20476 14132 20516
rect 12844 17032 12884 17072
rect 11692 15016 11732 15056
rect 11788 13252 11828 13292
rect 11884 11656 11924 11696
rect 11308 10900 11348 10940
rect 11500 10900 11540 10940
rect 11884 10816 11924 10856
rect 10886 10564 11254 10604
rect 10252 9472 10292 9512
rect 10636 9640 10676 9680
rect 10636 9136 10676 9176
rect 10444 8464 10484 8504
rect 9484 4936 9524 4976
rect 10828 9640 10868 9680
rect 11212 9556 11252 9596
rect 10924 9472 10964 9512
rect 10886 9052 11254 9092
rect 11404 10228 11444 10268
rect 12126 15856 12494 15896
rect 12126 14344 12494 14384
rect 13132 15688 13172 15728
rect 13612 16360 13652 16400
rect 12652 14260 12692 14300
rect 12126 12832 12494 12872
rect 12652 12412 12692 12452
rect 12126 11320 12494 11360
rect 11404 8968 11444 9008
rect 10886 7540 11254 7580
rect 10886 6028 11254 6068
rect 10924 5020 10964 5060
rect 12364 9976 12404 10016
rect 12126 9808 12494 9848
rect 11692 9304 11732 9344
rect 10886 4516 11254 4556
rect 12748 9472 12788 9512
rect 12940 15520 12980 15560
rect 12940 13252 12980 13292
rect 13132 14512 13172 14552
rect 13228 13084 13268 13124
rect 12940 12412 12980 12452
rect 12940 11824 12980 11864
rect 13612 13000 13652 13040
rect 13228 11992 13268 12032
rect 13612 12580 13652 12620
rect 13612 12412 13652 12452
rect 13516 11992 13556 12032
rect 13036 9976 13076 10016
rect 12940 9640 12980 9680
rect 12126 8296 12494 8336
rect 12126 6784 12494 6824
rect 11980 6448 12020 6488
rect 13036 9388 13076 9428
rect 12940 6364 12980 6404
rect 12460 5608 12500 5648
rect 13036 5608 13076 5648
rect 12126 5272 12494 5312
rect 10886 3004 11254 3044
rect 13516 11488 13556 11528
rect 13324 10648 13364 10688
rect 13228 9976 13268 10016
rect 13228 8884 13268 8924
rect 13228 5020 13268 5060
rect 12126 3760 12494 3800
rect 8524 1072 8564 1112
rect 10886 1492 11254 1532
rect 13420 9220 13460 9260
rect 13612 9556 13652 9596
rect 13804 14512 13844 14552
rect 13804 13000 13844 13040
rect 14476 17536 14516 17576
rect 14380 16948 14420 16988
rect 14092 14764 14132 14804
rect 13996 14680 14036 14720
rect 14092 13252 14132 13292
rect 13996 12580 14036 12620
rect 13900 11908 13940 11948
rect 13900 10984 13940 11024
rect 14476 16024 14516 16064
rect 14572 14680 14612 14720
rect 14764 15520 14804 15560
rect 14476 13084 14516 13124
rect 14668 13000 14708 13040
rect 14572 12496 14612 12536
rect 14284 11656 14324 11696
rect 13996 10732 14036 10772
rect 14764 12076 14804 12116
rect 14284 11152 14324 11192
rect 14668 11908 14708 11948
rect 14188 9976 14228 10016
rect 14092 7960 14132 8000
rect 13900 6448 13940 6488
rect 13516 6364 13556 6404
rect 12126 2248 12494 2288
rect 12172 1912 12212 1952
rect 12652 1912 12692 1952
rect 14188 6364 14228 6404
rect 14572 10900 14612 10940
rect 14668 10480 14708 10520
rect 15916 20644 15956 20684
rect 15916 20056 15956 20096
rect 15628 17200 15668 17240
rect 15052 14092 15092 14132
rect 14956 10648 14996 10688
rect 14956 9892 14996 9932
rect 14956 8884 14996 8924
rect 19900 27952 20268 27992
rect 17452 25348 17492 25388
rect 16108 20644 16148 20684
rect 16108 18460 16148 18500
rect 16012 16696 16052 16736
rect 15820 16192 15860 16232
rect 15724 14512 15764 14552
rect 15244 13252 15284 13292
rect 15724 13504 15764 13544
rect 15532 13252 15572 13292
rect 15244 12496 15284 12536
rect 15148 12412 15188 12452
rect 15148 11740 15188 11780
rect 15244 11824 15284 11864
rect 15244 11572 15284 11612
rect 15436 12076 15476 12116
rect 15628 13168 15668 13208
rect 15340 11236 15380 11276
rect 15244 10984 15284 11024
rect 15532 10144 15572 10184
rect 16108 14764 16148 14804
rect 17548 25264 17588 25304
rect 16684 18544 16724 18584
rect 18660 27196 19028 27236
rect 17932 25768 17972 25808
rect 18660 25684 19028 25724
rect 18700 25348 18740 25388
rect 18892 25264 18932 25304
rect 19180 25768 19220 25808
rect 18660 24172 19028 24212
rect 17068 20056 17107 20096
rect 17107 20056 17108 20096
rect 16876 19132 16916 19172
rect 18124 20056 18164 20096
rect 17356 19132 17396 19172
rect 17548 19216 17588 19256
rect 16876 18460 16916 18500
rect 17164 18460 17204 18500
rect 16300 13168 16340 13208
rect 16588 12580 16628 12620
rect 16492 11908 16532 11948
rect 15916 11404 15956 11444
rect 15820 10396 15860 10436
rect 16108 10312 16148 10352
rect 15724 10144 15764 10184
rect 16108 9892 16148 9932
rect 15820 9472 15860 9512
rect 15724 9304 15764 9344
rect 16012 8464 16052 8504
rect 14860 5608 14900 5648
rect 16300 11656 16340 11696
rect 16396 11572 16436 11612
rect 16396 11320 16436 11360
rect 16588 11656 16628 11696
rect 17548 18544 17588 18584
rect 17356 18460 17396 18500
rect 17164 14680 17204 14720
rect 16780 11908 16820 11948
rect 16780 11404 16820 11444
rect 16492 6532 16532 6572
rect 16396 6280 16436 6320
rect 16684 8884 16724 8924
rect 17548 16192 17588 16232
rect 17356 15772 17396 15812
rect 17932 18460 17972 18500
rect 18028 17536 18068 17576
rect 17740 16948 17780 16988
rect 17932 16864 17972 16904
rect 18220 17200 18260 17240
rect 17740 15520 17780 15560
rect 17644 14596 17684 14636
rect 17356 11572 17396 11612
rect 17452 13084 17492 13124
rect 17260 11236 17300 11276
rect 17356 10984 17396 11024
rect 16684 6532 16724 6572
rect 16684 5608 16724 5648
rect 16780 4936 16820 4976
rect 17260 9220 17300 9260
rect 17932 14512 17972 14552
rect 17836 13504 17876 13544
rect 17932 13252 17972 13292
rect 17644 11656 17684 11696
rect 17644 10648 17684 10688
rect 17548 10396 17588 10436
rect 17644 9388 17684 9428
rect 17836 10900 17876 10940
rect 17836 10312 17876 10352
rect 18220 16192 18260 16232
rect 18316 15520 18356 15560
rect 18316 13504 18356 13544
rect 18220 13084 18260 13124
rect 18660 22660 19028 22700
rect 19900 26440 20268 26480
rect 19900 24928 20268 24968
rect 18988 22156 19028 22196
rect 18660 21148 19028 21188
rect 18660 19636 19028 19676
rect 18988 18544 19028 18584
rect 18508 18376 18548 18416
rect 18660 18124 19028 18164
rect 18660 16612 19028 16652
rect 18700 15268 18740 15308
rect 18660 15100 19028 15140
rect 18604 14764 18644 14804
rect 18700 14680 18740 14720
rect 18604 14596 18644 14636
rect 18796 14092 18836 14132
rect 18660 13588 19028 13628
rect 18508 13168 18548 13208
rect 18124 12748 18164 12788
rect 18124 11740 18164 11780
rect 18220 11572 18260 11612
rect 18124 10060 18164 10100
rect 18124 8884 18164 8924
rect 18124 8128 18164 8168
rect 18660 12076 19028 12116
rect 19468 18544 19508 18584
rect 19900 23416 20268 23456
rect 19660 22156 19700 22196
rect 19900 21904 20268 21944
rect 19900 20392 20268 20432
rect 19660 18460 19700 18500
rect 19276 18376 19316 18416
rect 19276 16864 19316 16904
rect 19180 11488 19220 11528
rect 18892 10900 18932 10940
rect 18660 10564 19028 10604
rect 19180 10732 19220 10772
rect 18508 9976 18548 10016
rect 18660 9052 19028 9092
rect 18124 7120 18164 7160
rect 17932 7036 17972 7076
rect 17644 6364 17684 6404
rect 17356 4936 17396 4976
rect 16204 2584 16244 2624
rect 13516 1912 13556 1952
rect 18412 7036 18452 7076
rect 18604 7876 18644 7916
rect 19084 7876 19124 7916
rect 18660 7540 19028 7580
rect 18604 7120 18644 7160
rect 19900 18880 20268 18920
rect 19852 18544 19892 18584
rect 19948 18460 19988 18500
rect 20140 18376 20180 18416
rect 19900 17368 20268 17408
rect 19564 16948 19604 16988
rect 19948 17032 19988 17072
rect 20140 16780 20180 16820
rect 20140 16360 20180 16400
rect 19660 16276 19700 16316
rect 19900 15856 20268 15896
rect 19564 15436 19604 15476
rect 19564 14680 19604 14720
rect 19852 15016 19892 15056
rect 19660 13168 19700 13208
rect 19900 14344 20268 14384
rect 20140 13420 20180 13460
rect 19900 12832 20268 12872
rect 20140 12244 20180 12284
rect 19660 11320 19700 11360
rect 19900 11320 20268 11360
rect 19564 10396 19604 10436
rect 20620 20644 20660 20684
rect 20428 11656 20468 11696
rect 19564 9556 19604 9596
rect 19900 9808 20268 9848
rect 20140 9556 20180 9596
rect 19852 8968 19892 9008
rect 19948 9388 19988 9428
rect 20140 9304 20180 9344
rect 19900 8296 20268 8336
rect 19468 8128 19508 8168
rect 19852 7960 19892 8000
rect 18660 6028 19028 6068
rect 17164 2584 17204 2624
rect 18660 4516 19028 4556
rect 20140 7120 20180 7160
rect 19900 6784 20268 6824
rect 20428 9136 20468 9176
rect 20812 14008 20852 14048
rect 20620 11740 20660 11780
rect 23884 26860 23924 26900
rect 23980 23668 24020 23708
rect 23692 22240 23732 22280
rect 24556 23668 24596 23708
rect 24460 23500 24500 23540
rect 24556 23248 24596 23288
rect 24364 22996 24404 23036
rect 25708 26776 25748 26816
rect 24940 25348 24980 25388
rect 25132 25264 25158 25304
rect 25158 25264 25172 25304
rect 24940 23836 24980 23876
rect 24844 23248 24884 23288
rect 24844 23080 24884 23120
rect 22828 19048 22868 19088
rect 21388 14008 21428 14048
rect 21580 14764 21620 14804
rect 20620 9640 20660 9680
rect 21580 13000 21620 13040
rect 22444 14008 22484 14048
rect 22636 13504 22676 13544
rect 22636 12580 22676 12620
rect 22924 17704 22964 17744
rect 22828 13000 22868 13040
rect 23020 13000 23060 13040
rect 22924 12916 22964 12956
rect 23308 12748 23348 12788
rect 22636 11824 22676 11864
rect 22060 11656 22100 11696
rect 22060 10984 22100 11024
rect 22252 11068 22292 11108
rect 20428 7120 20468 7160
rect 20140 6280 20180 6320
rect 22732 11656 22772 11696
rect 22828 11152 22868 11192
rect 24076 19048 24116 19088
rect 23980 16780 24020 16820
rect 23500 13840 23540 13880
rect 23500 13504 23540 13544
rect 23788 14596 23828 14636
rect 23692 13084 23732 13124
rect 23692 12916 23732 12956
rect 23980 14680 24020 14720
rect 23980 13924 24020 13964
rect 24460 16780 24500 16820
rect 24364 14848 24404 14888
rect 25132 23164 25172 23204
rect 25132 22240 25172 22280
rect 24940 17704 24980 17744
rect 25612 23920 25652 23960
rect 25804 25600 25844 25640
rect 27724 28120 27764 28160
rect 27674 27952 28042 27992
rect 29356 28120 29396 28160
rect 26434 27196 26802 27236
rect 26284 26860 26324 26900
rect 25804 24676 25844 24716
rect 25996 23920 26036 23960
rect 25900 23836 25940 23876
rect 26434 25684 26802 25724
rect 25804 22828 25844 22868
rect 25516 20980 25556 21020
rect 25804 21484 25844 21524
rect 25420 20728 25460 20768
rect 25516 20560 25556 20600
rect 25900 20728 25940 20768
rect 24172 14680 24212 14720
rect 24268 14596 24308 14636
rect 24172 13252 24212 13292
rect 24076 13000 24116 13040
rect 23596 12496 23636 12536
rect 24076 12832 24116 12872
rect 23884 12748 23924 12788
rect 23788 12496 23828 12536
rect 23884 12412 23924 12452
rect 23500 11068 23540 11108
rect 23500 9472 23540 9512
rect 23404 8632 23444 8672
rect 23116 7036 23156 7076
rect 22060 6364 22100 6404
rect 19900 5272 20268 5312
rect 19900 3760 20268 3800
rect 18660 3004 19028 3044
rect 18660 1492 19028 1532
rect 19900 2248 20268 2288
rect 23692 11992 23732 12032
rect 23980 11824 24020 11864
rect 23884 11740 23924 11780
rect 23980 10060 24020 10100
rect 24460 13924 24500 13964
rect 24652 14764 24692 14804
rect 24652 14008 24692 14048
rect 24748 11068 24788 11108
rect 26764 25348 26804 25388
rect 26956 25600 26996 25640
rect 26956 25348 26996 25388
rect 26434 24172 26802 24212
rect 27628 26776 27668 26816
rect 26956 24592 26996 24632
rect 27674 26440 28042 26480
rect 27628 26104 27668 26144
rect 28492 26104 28532 26144
rect 27628 25348 27668 25388
rect 28012 25264 28052 25304
rect 27674 24928 28042 24968
rect 27820 23752 27860 23792
rect 26668 22996 26708 23036
rect 26380 22828 26420 22868
rect 26860 22828 26900 22868
rect 26434 22660 26802 22700
rect 26380 21736 26420 21776
rect 26860 21652 26900 21692
rect 26572 21484 26612 21524
rect 26434 21148 26802 21188
rect 26476 20560 26516 20600
rect 26764 20980 26804 21020
rect 26764 20308 26804 20348
rect 26668 19804 26708 19844
rect 26434 19636 26802 19676
rect 27436 23500 27476 23540
rect 27052 22996 27092 23036
rect 27052 21652 27092 21692
rect 27674 23416 28042 23456
rect 27724 22828 27764 22868
rect 27436 22240 27476 22280
rect 27052 20728 27092 20768
rect 27244 20812 27284 20852
rect 27148 20560 27188 20600
rect 27436 20308 27476 20348
rect 27674 21904 28042 21944
rect 27628 21568 27668 21608
rect 27820 20728 27860 20768
rect 27674 20392 28042 20432
rect 25612 14848 25652 14888
rect 25132 13924 25172 13964
rect 25036 12832 25076 12872
rect 24364 9556 24404 9596
rect 25516 14008 25556 14048
rect 25516 11656 25556 11696
rect 25804 13924 25844 13964
rect 26434 18124 26802 18164
rect 26434 16612 26802 16652
rect 27244 19804 27284 19844
rect 26434 15100 26802 15140
rect 27674 18880 28042 18920
rect 28684 23752 28724 23792
rect 29548 24592 29588 24632
rect 28588 19804 28628 19844
rect 27674 17368 28042 17408
rect 27674 15856 28042 15896
rect 25804 13084 25844 13124
rect 25708 12664 25748 12704
rect 25900 12664 25940 12704
rect 26434 13588 26802 13628
rect 27148 14680 27188 14720
rect 27052 12916 27092 12956
rect 26764 12496 26804 12536
rect 26860 12664 26900 12704
rect 26434 12076 26802 12116
rect 26956 12580 26996 12620
rect 26188 11656 26228 11696
rect 25036 9472 25076 9512
rect 25900 9472 25940 9512
rect 24940 8632 24980 8672
rect 26434 10564 26802 10604
rect 26860 9472 26900 9512
rect 26434 9052 26802 9092
rect 26434 7540 26802 7580
rect 25516 5608 25556 5648
rect 26434 6028 26802 6068
rect 26434 4516 26802 4556
rect 26476 4096 26516 4136
rect 27820 14848 27860 14888
rect 27436 12832 27476 12872
rect 27674 14344 28042 14384
rect 27628 14008 27668 14048
rect 27674 12832 28042 12872
rect 27340 11656 27380 11696
rect 27436 9808 27476 9848
rect 30028 21736 30068 21776
rect 29644 21568 29684 21608
rect 28396 14848 28436 14888
rect 28492 14680 28532 14720
rect 28876 14680 28916 14720
rect 28972 14764 29012 14804
rect 28396 12664 28436 12704
rect 28396 12412 28436 12452
rect 28204 11572 28244 11612
rect 27674 11320 28042 11360
rect 28108 10984 28148 11024
rect 27674 9808 28042 9848
rect 27628 9640 27668 9680
rect 27674 8296 28042 8336
rect 27674 6784 28042 6824
rect 28012 5608 28052 5648
rect 27674 5272 28042 5312
rect 27436 4096 27476 4136
rect 27674 3760 28042 3800
rect 26434 3004 26802 3044
rect 27674 2248 28042 2288
rect 26434 1492 26802 1532
rect 28300 7036 28340 7076
rect 28780 7036 28820 7076
rect 30220 9556 30260 9596
rect 29644 5608 29684 5648
rect 30124 5608 30164 5648
rect 12126 736 12494 776
rect 19900 736 20268 776
rect 27674 736 28042 776
<< metal4 >>
rect 27715 28120 27724 28160
rect 27764 28120 29356 28160
rect 29396 28120 29405 28160
rect 4343 27952 4352 27992
rect 4720 27952 4729 27992
rect 12117 27952 12126 27992
rect 12494 27952 12503 27992
rect 19891 27952 19900 27992
rect 20268 27952 20277 27992
rect 27665 27952 27674 27992
rect 28042 27952 28051 27992
rect 10339 27364 10348 27404
rect 10388 27364 10828 27404
rect 10868 27364 10877 27404
rect 3103 27196 3112 27236
rect 3480 27196 3489 27236
rect 10877 27196 10886 27236
rect 11254 27196 11263 27236
rect 18651 27196 18660 27236
rect 19028 27196 19037 27236
rect 26425 27196 26434 27236
rect 26802 27196 26811 27236
rect 23875 26860 23884 26900
rect 23924 26860 26284 26900
rect 26324 26860 26333 26900
rect 25699 26776 25708 26816
rect 25748 26776 27628 26816
rect 27668 26776 27677 26816
rect 4343 26440 4352 26480
rect 4720 26440 4729 26480
rect 12117 26440 12126 26480
rect 12494 26440 12503 26480
rect 12547 26440 12556 26480
rect 12596 26440 12940 26480
rect 12980 26440 12989 26480
rect 19891 26440 19900 26480
rect 20268 26440 20277 26480
rect 27665 26440 27674 26480
rect 28042 26440 28051 26480
rect 8323 26272 8332 26312
rect 8372 26272 8908 26312
rect 8948 26272 10060 26312
rect 10100 26272 10109 26312
rect 9955 26104 9964 26144
rect 10004 26104 10156 26144
rect 10196 26104 10205 26144
rect 12931 26104 12940 26144
rect 12980 26104 14380 26144
rect 14420 26104 14429 26144
rect 27619 26104 27628 26144
rect 27668 26104 28492 26144
rect 28532 26104 28541 26144
rect 10051 25936 10060 25976
rect 10100 25936 12460 25976
rect 12500 25936 12940 25976
rect 12980 25936 12989 25976
rect 9859 25852 9868 25892
rect 9908 25852 11980 25892
rect 12020 25852 12029 25892
rect 17923 25768 17932 25808
rect 17972 25768 19180 25808
rect 19220 25768 19229 25808
rect 3103 25684 3112 25724
rect 3480 25684 3489 25724
rect 10445 25684 10540 25724
rect 10580 25684 10589 25724
rect 10877 25684 10886 25724
rect 11254 25684 11263 25724
rect 18651 25684 18660 25724
rect 19028 25684 19037 25724
rect 26425 25684 26434 25724
rect 26802 25684 26811 25724
rect 11491 25600 11500 25640
rect 11540 25600 11549 25640
rect 25795 25600 25804 25640
rect 25844 25600 26956 25640
rect 26996 25600 27005 25640
rect 11500 25556 11540 25600
rect 9091 25516 9100 25556
rect 9140 25516 10540 25556
rect 10580 25516 11116 25556
rect 11156 25516 11540 25556
rect 17443 25348 17452 25388
rect 17492 25348 18700 25388
rect 18740 25348 18749 25388
rect 24931 25348 24940 25388
rect 24980 25348 26764 25388
rect 26804 25348 26956 25388
rect 26996 25348 27628 25388
rect 27668 25348 27677 25388
rect 10531 25264 10540 25304
rect 10580 25264 10828 25304
rect 10868 25264 10877 25304
rect 17539 25264 17548 25304
rect 17588 25264 18892 25304
rect 18932 25264 18941 25304
rect 25123 25264 25132 25304
rect 25172 25264 28012 25304
rect 28052 25264 28061 25304
rect 10435 25180 10444 25220
rect 10484 25180 11116 25220
rect 11156 25180 11165 25220
rect 4343 24928 4352 24968
rect 4720 24928 4729 24968
rect 12117 24928 12126 24968
rect 12494 24928 12503 24968
rect 19891 24928 19900 24968
rect 20268 24928 20277 24968
rect 27665 24928 27674 24968
rect 28042 24928 28051 24968
rect 5635 24760 5644 24800
rect 5684 24760 10444 24800
rect 10484 24760 10493 24800
rect 25709 24676 25804 24716
rect 25844 24676 25853 24716
rect 26947 24592 26956 24632
rect 26996 24592 29548 24632
rect 29588 24592 29597 24632
rect 11107 24508 11116 24548
rect 11156 24508 12652 24548
rect 12692 24508 12701 24548
rect 5059 24424 5068 24464
rect 5108 24424 9772 24464
rect 9812 24424 9821 24464
rect 3103 24172 3112 24212
rect 3480 24172 3489 24212
rect 10877 24172 10886 24212
rect 11254 24172 11263 24212
rect 18651 24172 18660 24212
rect 19028 24172 19037 24212
rect 26425 24172 26434 24212
rect 26802 24172 26811 24212
rect 25603 23920 25612 23960
rect 25652 23920 25996 23960
rect 26036 23920 26045 23960
rect 10051 23836 10060 23876
rect 10100 23836 12556 23876
rect 12596 23836 12605 23876
rect 24931 23836 24940 23876
rect 24980 23836 25900 23876
rect 25940 23836 25949 23876
rect 27811 23752 27820 23792
rect 27860 23752 28684 23792
rect 28724 23752 28733 23792
rect 23971 23668 23980 23708
rect 24020 23668 24556 23708
rect 24596 23668 24605 23708
rect 24451 23500 24460 23540
rect 24500 23500 27436 23540
rect 27476 23500 27485 23540
rect 4343 23416 4352 23456
rect 4720 23416 4729 23456
rect 12117 23416 12126 23456
rect 12494 23416 12503 23456
rect 19891 23416 19900 23456
rect 20268 23416 20277 23456
rect 27665 23416 27674 23456
rect 28042 23416 28051 23456
rect 11875 23248 11884 23288
rect 11924 23248 12460 23288
rect 12500 23248 12509 23288
rect 24547 23248 24556 23288
rect 24596 23248 24844 23288
rect 24884 23248 24893 23288
rect 11683 23164 11692 23204
rect 11732 23164 12596 23204
rect 12556 23120 12596 23164
rect 24844 23164 25132 23204
rect 25172 23164 25181 23204
rect 24844 23120 24884 23164
rect 12547 23080 12556 23120
rect 12596 23080 15820 23120
rect 15860 23080 15869 23120
rect 24835 23080 24844 23120
rect 24884 23080 24893 23120
rect 24355 22996 24364 23036
rect 24404 22996 26668 23036
rect 26708 22996 27052 23036
rect 27092 22996 27101 23036
rect 11107 22912 11116 22952
rect 11156 22912 11500 22952
rect 11540 22912 11549 22952
rect 25709 22828 25804 22868
rect 25844 22828 25853 22868
rect 26371 22828 26380 22868
rect 26420 22828 26860 22868
rect 26900 22828 27724 22868
rect 27764 22828 27773 22868
rect 3103 22660 3112 22700
rect 3480 22660 3489 22700
rect 10877 22660 10886 22700
rect 11254 22660 11263 22700
rect 18651 22660 18660 22700
rect 19028 22660 19037 22700
rect 26425 22660 26434 22700
rect 26802 22660 26811 22700
rect 11203 22492 11212 22532
rect 11252 22492 11596 22532
rect 11636 22492 11645 22532
rect 12355 22240 12364 22280
rect 12404 22240 13324 22280
rect 13364 22240 13373 22280
rect 23683 22240 23692 22280
rect 23732 22240 25132 22280
rect 25172 22240 27436 22280
rect 27476 22240 27485 22280
rect 12835 22156 12844 22196
rect 12884 22156 15244 22196
rect 15284 22156 18988 22196
rect 19028 22156 19660 22196
rect 19700 22156 19709 22196
rect 4343 21904 4352 21944
rect 4720 21904 4729 21944
rect 12117 21904 12126 21944
rect 12494 21904 12503 21944
rect 19891 21904 19900 21944
rect 20268 21904 20277 21944
rect 27665 21904 27674 21944
rect 28042 21904 28051 21944
rect 26371 21736 26380 21776
rect 26420 21736 30028 21776
rect 30068 21736 30077 21776
rect 26851 21652 26860 21692
rect 26900 21652 27052 21692
rect 27092 21652 27101 21692
rect 4675 21568 4684 21608
rect 4724 21568 5356 21608
rect 5396 21568 5405 21608
rect 27619 21568 27628 21608
rect 27668 21568 29644 21608
rect 29684 21568 29693 21608
rect 25795 21484 25804 21524
rect 25844 21484 26572 21524
rect 26612 21484 26621 21524
rect 3103 21148 3112 21188
rect 3480 21148 3489 21188
rect 10877 21148 10886 21188
rect 11254 21148 11263 21188
rect 18651 21148 18660 21188
rect 19028 21148 19037 21188
rect 26425 21148 26434 21188
rect 26802 21148 26811 21188
rect 5347 20980 5356 21020
rect 5396 20980 11500 21020
rect 11540 20980 11549 21020
rect 25507 20980 25516 21020
rect 25556 20980 26764 21020
rect 26804 20980 26813 21020
rect 2275 20812 2284 20852
rect 2324 20812 4300 20852
rect 4340 20812 4349 20852
rect 25900 20812 27244 20852
rect 27284 20812 27293 20852
rect 25900 20768 25940 20812
rect 4195 20728 4204 20768
rect 4244 20728 11884 20768
rect 11924 20728 11933 20768
rect 25411 20728 25420 20768
rect 25460 20728 25900 20768
rect 25940 20728 25949 20768
rect 27043 20728 27052 20768
rect 27092 20728 27820 20768
rect 27860 20728 27869 20768
rect 3907 20644 3916 20684
rect 3956 20644 5452 20684
rect 5492 20644 5501 20684
rect 12931 20644 12940 20684
rect 12980 20644 13324 20684
rect 13364 20644 15916 20684
rect 15956 20644 16108 20684
rect 16148 20644 16157 20684
rect 20611 20644 20620 20684
rect 20660 20644 23500 20684
rect 23540 20644 23549 20684
rect 25507 20560 25516 20600
rect 25556 20560 26476 20600
rect 26516 20560 27148 20600
rect 27188 20560 27197 20600
rect 547 20476 556 20516
rect 596 20476 14092 20516
rect 14132 20476 14141 20516
rect 4343 20392 4352 20432
rect 4720 20392 4729 20432
rect 12117 20392 12126 20432
rect 12494 20392 12503 20432
rect 19891 20392 19900 20432
rect 20268 20392 20277 20432
rect 27665 20392 27674 20432
rect 28042 20392 28051 20432
rect 26755 20308 26764 20348
rect 26804 20308 27436 20348
rect 27476 20308 27485 20348
rect 3139 20224 3148 20264
rect 3188 20224 10100 20264
rect 10060 20180 10100 20224
rect 10051 20140 10060 20180
rect 10100 20140 10109 20180
rect 3331 20056 3340 20096
rect 3380 20056 4204 20096
rect 4244 20056 4253 20096
rect 5731 20056 5740 20096
rect 5780 20056 6700 20096
rect 6740 20056 7756 20096
rect 7796 20056 7805 20096
rect 15907 20056 15916 20096
rect 15956 20056 17068 20096
rect 17108 20056 18124 20096
rect 18164 20056 18173 20096
rect 4291 19972 4300 20012
rect 4340 19972 7372 20012
rect 7412 19972 7421 20012
rect 26659 19804 26668 19844
rect 26708 19804 27244 19844
rect 27284 19804 28588 19844
rect 28628 19804 28637 19844
rect 2851 19720 2860 19760
rect 2900 19720 4588 19760
rect 4628 19720 4637 19760
rect 3103 19636 3112 19676
rect 3480 19636 3489 19676
rect 10877 19636 10886 19676
rect 11254 19636 11263 19676
rect 18651 19636 18660 19676
rect 19028 19636 19037 19676
rect 26425 19636 26434 19676
rect 26802 19636 26811 19676
rect 2179 19300 2188 19340
rect 2228 19300 2668 19340
rect 2708 19300 3148 19340
rect 3188 19300 3197 19340
rect 11491 19300 11500 19340
rect 11540 19300 12460 19340
rect 12500 19300 12509 19340
rect 1699 19216 1708 19256
rect 1748 19216 2092 19256
rect 2132 19216 2141 19256
rect 11875 19216 11884 19256
rect 11924 19216 17548 19256
rect 17588 19216 17597 19256
rect 9283 19132 9292 19172
rect 9332 19132 9964 19172
rect 10004 19132 10013 19172
rect 16867 19132 16876 19172
rect 16916 19132 17356 19172
rect 17396 19132 17405 19172
rect 22819 19048 22828 19088
rect 22868 19048 24076 19088
rect 24116 19048 24125 19088
rect 4343 18880 4352 18920
rect 4720 18880 4729 18920
rect 12117 18880 12126 18920
rect 12494 18880 12503 18920
rect 19891 18880 19900 18920
rect 20268 18880 20277 18920
rect 27665 18880 27674 18920
rect 28042 18880 28051 18920
rect 2083 18796 2092 18836
rect 2132 18796 3148 18836
rect 3188 18796 3197 18836
rect 5635 18628 5644 18668
rect 5684 18628 6604 18668
rect 6644 18628 6653 18668
rect 2467 18544 2476 18584
rect 2516 18544 2668 18584
rect 2708 18544 2717 18584
rect 11203 18544 11212 18584
rect 11252 18544 11500 18584
rect 11540 18544 11549 18584
rect 16675 18544 16684 18584
rect 16724 18544 17548 18584
rect 17588 18544 17597 18584
rect 18979 18544 18988 18584
rect 19028 18544 19180 18584
rect 19220 18544 19229 18584
rect 19459 18544 19468 18584
rect 19508 18544 19852 18584
rect 19892 18544 19901 18584
rect 6883 18460 6892 18500
rect 6932 18460 9772 18500
rect 9812 18460 9821 18500
rect 16099 18460 16108 18500
rect 16148 18460 16876 18500
rect 16916 18460 17164 18500
rect 17204 18460 17356 18500
rect 17396 18460 17932 18500
rect 17972 18460 17981 18500
rect 19651 18460 19660 18500
rect 19700 18460 19948 18500
rect 19988 18460 19997 18500
rect 18499 18376 18508 18416
rect 18548 18376 19276 18416
rect 19316 18376 20140 18416
rect 20180 18376 20189 18416
rect 3103 18124 3112 18164
rect 3480 18124 3489 18164
rect 10877 18124 10886 18164
rect 11254 18124 11263 18164
rect 18651 18124 18660 18164
rect 19028 18124 19037 18164
rect 26425 18124 26434 18164
rect 26802 18124 26811 18164
rect 2947 18040 2956 18080
rect 2996 18040 5164 18080
rect 5204 18040 5213 18080
rect 2659 17788 2668 17828
rect 2708 17788 5260 17828
rect 5300 17788 6892 17828
rect 6932 17788 6941 17828
rect 3523 17704 3532 17744
rect 3572 17704 3916 17744
rect 3956 17704 3965 17744
rect 22915 17704 22924 17744
rect 22964 17704 24940 17744
rect 24980 17704 24989 17744
rect 4675 17536 4684 17576
rect 4724 17536 4733 17576
rect 8995 17536 9004 17576
rect 9044 17536 14476 17576
rect 14516 17536 14525 17576
rect 17933 17536 18028 17576
rect 18068 17536 18077 17576
rect 4684 17492 4724 17536
rect 4684 17452 4820 17492
rect 4343 17368 4352 17408
rect 4720 17368 4729 17408
rect 4780 17240 4820 17452
rect 9475 17368 9484 17408
rect 9524 17368 10444 17408
rect 10484 17368 10636 17408
rect 10676 17368 10828 17408
rect 10868 17368 10877 17408
rect 12117 17368 12126 17408
rect 12494 17368 12503 17408
rect 19891 17368 19900 17408
rect 20268 17368 20277 17408
rect 27665 17368 27674 17408
rect 28042 17368 28051 17408
rect 2179 17200 2188 17240
rect 2228 17200 4492 17240
rect 4532 17200 4820 17240
rect 10051 17200 10060 17240
rect 10100 17200 10540 17240
rect 10580 17200 11404 17240
rect 11444 17200 11453 17240
rect 15619 17200 15628 17240
rect 15668 17200 18220 17240
rect 18260 17200 18269 17240
rect 10819 17032 10828 17072
rect 10868 17032 11884 17072
rect 11924 17032 11933 17072
rect 12835 17032 12844 17072
rect 12884 17032 19948 17072
rect 19988 17032 19997 17072
rect 11203 16948 11212 16988
rect 11252 16948 14380 16988
rect 14420 16948 14429 16988
rect 17731 16948 17740 16988
rect 17780 16948 19564 16988
rect 19604 16948 19613 16988
rect 8899 16864 8908 16904
rect 8948 16864 9004 16904
rect 9044 16864 9053 16904
rect 11011 16864 11020 16904
rect 11060 16864 11404 16904
rect 11444 16864 11453 16904
rect 17923 16864 17932 16904
rect 17972 16864 19276 16904
rect 19316 16864 19325 16904
rect 9475 16780 9484 16820
rect 9524 16780 9964 16820
rect 10004 16780 11692 16820
rect 11732 16780 11741 16820
rect 12643 16780 12652 16820
rect 12692 16780 15532 16820
rect 15572 16780 20140 16820
rect 20180 16780 20189 16820
rect 23971 16780 23980 16820
rect 24020 16780 24460 16820
rect 24500 16780 24509 16820
rect 12547 16696 12556 16736
rect 12596 16696 16012 16736
rect 16052 16696 16061 16736
rect 3103 16612 3112 16652
rect 3480 16612 3489 16652
rect 10877 16612 10886 16652
rect 11254 16612 11263 16652
rect 18651 16612 18660 16652
rect 19028 16612 19037 16652
rect 26425 16612 26434 16652
rect 26802 16612 26811 16652
rect 259 16444 268 16484
rect 308 16444 8524 16484
rect 8564 16444 8573 16484
rect 10060 16360 13612 16400
rect 13652 16360 13661 16400
rect 19171 16360 19180 16400
rect 19220 16360 20140 16400
rect 20180 16360 20189 16400
rect 10060 16316 10100 16360
rect 1603 16276 1612 16316
rect 1652 16276 1804 16316
rect 1844 16276 1853 16316
rect 6787 16276 6796 16316
rect 6836 16276 6988 16316
rect 7028 16276 10100 16316
rect 19555 16276 19564 16316
rect 19604 16276 19660 16316
rect 19700 16276 19709 16316
rect 1027 16192 1036 16232
rect 1076 16192 2188 16232
rect 2228 16192 2237 16232
rect 5443 16192 5452 16232
rect 5492 16192 7564 16232
rect 7604 16192 8428 16232
rect 8468 16192 9964 16232
rect 10004 16192 10013 16232
rect 10349 16192 10444 16232
rect 10484 16192 10493 16232
rect 15811 16192 15820 16232
rect 15860 16192 17548 16232
rect 17588 16192 18220 16232
rect 18260 16192 18269 16232
rect 4675 16024 4684 16064
rect 4724 16024 6316 16064
rect 6356 16024 6365 16064
rect 8429 16024 8524 16064
rect 8564 16024 8573 16064
rect 10051 16024 10060 16064
rect 10100 16024 14476 16064
rect 14516 16024 14525 16064
rect 7075 15940 7084 15980
rect 7124 15940 7756 15980
rect 7796 15940 7805 15980
rect 4343 15856 4352 15896
rect 4720 15856 4729 15896
rect 6883 15856 6892 15896
rect 6932 15856 7564 15896
rect 7604 15856 7613 15896
rect 12117 15856 12126 15896
rect 12494 15856 12503 15896
rect 19891 15856 19900 15896
rect 20268 15856 20277 15896
rect 27665 15856 27674 15896
rect 28042 15856 28051 15896
rect 3715 15772 3724 15812
rect 3764 15772 8044 15812
rect 8084 15772 8093 15812
rect 9772 15772 17356 15812
rect 17396 15772 17405 15812
rect 4483 15688 4492 15728
rect 4532 15688 9196 15728
rect 9236 15688 9245 15728
rect 9772 15644 9812 15772
rect 10531 15688 10540 15728
rect 10580 15688 13132 15728
rect 13172 15688 13181 15728
rect 8035 15604 8044 15644
rect 8084 15604 9812 15644
rect 9869 15604 9964 15644
rect 10004 15604 10013 15644
rect 7267 15520 7276 15560
rect 7316 15520 9772 15560
rect 9812 15520 9821 15560
rect 10445 15520 10540 15560
rect 10580 15520 12940 15560
rect 12980 15520 14764 15560
rect 14804 15520 14813 15560
rect 17731 15520 17740 15560
rect 17780 15520 18316 15560
rect 18356 15520 18365 15560
rect 5443 15436 5452 15476
rect 5492 15436 6508 15476
rect 6548 15436 6557 15476
rect 6883 15436 6892 15476
rect 6932 15436 8908 15476
rect 8948 15436 8957 15476
rect 9091 15436 9100 15476
rect 9140 15436 19564 15476
rect 19604 15436 19613 15476
rect 6019 15352 6028 15392
rect 6068 15352 8044 15392
rect 8084 15352 8093 15392
rect 8323 15352 8332 15392
rect 8372 15352 9964 15392
rect 10004 15352 10732 15392
rect 10772 15352 10781 15392
rect 11107 15268 11116 15308
rect 11156 15268 18700 15308
rect 18740 15268 18749 15308
rect 3103 15100 3112 15140
rect 3480 15100 3489 15140
rect 10877 15100 10886 15140
rect 11254 15100 11263 15140
rect 18651 15100 18660 15140
rect 19028 15100 19037 15140
rect 26425 15100 26434 15140
rect 26802 15100 26811 15140
rect 11683 15016 11692 15056
rect 11732 15016 19852 15056
rect 19892 15016 19901 15056
rect 10243 14932 10252 14972
rect 10292 14932 10732 14972
rect 10772 14932 10781 14972
rect 24355 14848 24364 14888
rect 24404 14848 25612 14888
rect 25652 14848 27820 14888
rect 27860 14848 28396 14888
rect 28436 14848 28445 14888
rect 10051 14764 10060 14804
rect 10100 14764 10252 14804
rect 10292 14764 10301 14804
rect 14083 14764 14092 14804
rect 14132 14764 16108 14804
rect 16148 14764 16157 14804
rect 18499 14764 18508 14804
rect 18548 14764 18604 14804
rect 18644 14764 18653 14804
rect 21571 14764 21580 14804
rect 21620 14764 24652 14804
rect 24692 14764 28972 14804
rect 29012 14764 29021 14804
rect 10252 14720 10292 14764
rect 5731 14680 5740 14720
rect 5780 14680 9676 14720
rect 9716 14680 9725 14720
rect 10252 14680 13996 14720
rect 14036 14680 14572 14720
rect 14612 14680 14621 14720
rect 17155 14680 17164 14720
rect 17204 14680 18700 14720
rect 18740 14680 18749 14720
rect 19555 14680 19564 14720
rect 19604 14680 19660 14720
rect 19700 14680 19709 14720
rect 23971 14680 23980 14720
rect 24020 14680 24172 14720
rect 24212 14680 24221 14720
rect 27139 14680 27148 14720
rect 27188 14680 28492 14720
rect 28532 14680 28876 14720
rect 28916 14680 28925 14720
rect 3427 14596 3436 14636
rect 3476 14596 5932 14636
rect 5972 14596 5981 14636
rect 6211 14596 6220 14636
rect 6260 14596 7084 14636
rect 7124 14596 9580 14636
rect 9620 14596 9629 14636
rect 17635 14596 17644 14636
rect 17684 14596 18604 14636
rect 18644 14596 18653 14636
rect 23779 14596 23788 14636
rect 23828 14596 24268 14636
rect 24308 14596 24317 14636
rect 13123 14512 13132 14552
rect 13172 14512 13804 14552
rect 13844 14512 13853 14552
rect 15715 14512 15724 14552
rect 15764 14512 17932 14552
rect 17972 14512 18124 14552
rect 18164 14512 18173 14552
rect 4099 14428 4108 14468
rect 4148 14428 7852 14468
rect 7892 14428 8524 14468
rect 8564 14428 8573 14468
rect 4343 14344 4352 14384
rect 4720 14344 4729 14384
rect 12117 14344 12126 14384
rect 12494 14344 12503 14384
rect 19891 14344 19900 14384
rect 20268 14344 20277 14384
rect 27665 14344 27674 14384
rect 28042 14344 28051 14384
rect 5443 14260 5452 14300
rect 5492 14260 12652 14300
rect 12692 14260 12701 14300
rect 4099 14176 4108 14216
rect 4148 14176 5644 14216
rect 5684 14176 6028 14216
rect 6068 14176 6077 14216
rect 15043 14092 15052 14132
rect 15092 14092 18796 14132
rect 18836 14092 19564 14132
rect 19604 14092 19613 14132
rect 20803 14008 20812 14048
rect 20852 14008 21388 14048
rect 21428 14008 22444 14048
rect 22484 14008 22493 14048
rect 23971 14008 23980 14048
rect 24020 14008 24652 14048
rect 24692 14008 25516 14048
rect 25556 14008 27628 14048
rect 27668 14008 27677 14048
rect 23971 13924 23980 13964
rect 24020 13924 24460 13964
rect 24500 13924 24509 13964
rect 25123 13924 25132 13964
rect 25172 13924 25804 13964
rect 25844 13924 25853 13964
rect 23405 13840 23500 13880
rect 23540 13840 23549 13880
rect 3103 13588 3112 13628
rect 3480 13588 3489 13628
rect 10877 13588 10886 13628
rect 11254 13588 11263 13628
rect 18651 13588 18660 13628
rect 19028 13588 19037 13628
rect 26425 13588 26434 13628
rect 26802 13588 26811 13628
rect 4867 13504 4876 13544
rect 4916 13504 8044 13544
rect 8084 13504 8093 13544
rect 15715 13504 15724 13544
rect 15764 13504 17836 13544
rect 17876 13504 18316 13544
rect 18356 13504 18365 13544
rect 22627 13504 22636 13544
rect 22676 13504 23500 13544
rect 23540 13504 23549 13544
rect 6211 13420 6220 13460
rect 6260 13420 7564 13460
rect 7604 13420 7613 13460
rect 11107 13420 11116 13460
rect 11156 13420 20140 13460
rect 20180 13420 20189 13460
rect 5827 13336 5836 13376
rect 5876 13336 6124 13376
rect 6164 13336 6173 13376
rect 8707 13336 8716 13376
rect 8756 13336 8908 13376
rect 8948 13336 8957 13376
rect 4867 13252 4876 13292
rect 4916 13252 5260 13292
rect 5300 13252 5644 13292
rect 5684 13252 6892 13292
rect 6932 13252 8524 13292
rect 8564 13252 8573 13292
rect 11779 13252 11788 13292
rect 11828 13252 12940 13292
rect 12980 13252 12989 13292
rect 14083 13252 14092 13292
rect 14132 13252 15244 13292
rect 15284 13252 15293 13292
rect 15523 13252 15532 13292
rect 15572 13252 17932 13292
rect 17972 13252 17981 13292
rect 24163 13252 24172 13292
rect 24212 13252 24221 13292
rect 12940 13208 12980 13252
rect 5539 13168 5548 13208
rect 5588 13168 6412 13208
rect 6452 13168 6461 13208
rect 7555 13168 7564 13208
rect 7604 13168 8140 13208
rect 8180 13168 8189 13208
rect 8323 13168 8332 13208
rect 8372 13168 8908 13208
rect 8948 13168 8957 13208
rect 12940 13168 15628 13208
rect 15668 13168 15677 13208
rect 16291 13168 16300 13208
rect 16340 13168 18508 13208
rect 18548 13168 18557 13208
rect 19565 13168 19660 13208
rect 19700 13168 19709 13208
rect 6412 13124 6452 13168
rect 24172 13124 24212 13252
rect 6412 13084 9100 13124
rect 9140 13084 9149 13124
rect 13219 13084 13228 13124
rect 13268 13084 14476 13124
rect 14516 13084 14525 13124
rect 17443 13084 17452 13124
rect 17492 13084 18220 13124
rect 18260 13084 18269 13124
rect 23683 13084 23692 13124
rect 23732 13084 25804 13124
rect 25844 13084 25853 13124
rect 7075 13000 7084 13040
rect 7124 13000 7180 13040
rect 7220 13000 7229 13040
rect 13603 13000 13612 13040
rect 13652 13000 13804 13040
rect 13844 13000 14668 13040
rect 14708 13000 14717 13040
rect 21571 13000 21580 13040
rect 21620 13000 22828 13040
rect 22868 13000 22877 13040
rect 23011 13000 23020 13040
rect 23060 13000 23924 13040
rect 23981 13000 24076 13040
rect 24116 13000 24125 13040
rect 23884 12956 23924 13000
rect 6595 12916 6604 12956
rect 6644 12916 8716 12956
rect 8756 12916 8765 12956
rect 22915 12916 22924 12956
rect 22964 12916 23692 12956
rect 23732 12916 23741 12956
rect 23884 12916 27052 12956
rect 27092 12916 27101 12956
rect 4343 12832 4352 12872
rect 4720 12832 4729 12872
rect 12117 12832 12126 12872
rect 12494 12832 12503 12872
rect 19891 12832 19900 12872
rect 20268 12832 20277 12872
rect 23981 12832 24076 12872
rect 24116 12832 24125 12872
rect 25027 12832 25036 12872
rect 25076 12832 27436 12872
rect 27476 12832 27485 12872
rect 27665 12832 27674 12872
rect 28042 12832 28051 12872
rect 18019 12748 18028 12788
rect 18068 12748 18124 12788
rect 18164 12748 18173 12788
rect 23299 12748 23308 12788
rect 23348 12748 23884 12788
rect 23924 12748 23933 12788
rect 25699 12664 25708 12704
rect 25748 12664 25900 12704
rect 25940 12664 25949 12704
rect 26851 12664 26860 12704
rect 26900 12664 28396 12704
rect 28436 12664 28445 12704
rect 8323 12580 8332 12620
rect 8372 12580 13612 12620
rect 13652 12580 13661 12620
rect 13987 12580 13996 12620
rect 14036 12580 16588 12620
rect 16628 12580 16637 12620
rect 22627 12580 22636 12620
rect 22676 12580 26956 12620
rect 26996 12580 27005 12620
rect 7651 12496 7660 12536
rect 7700 12496 7709 12536
rect 8323 12496 8332 12536
rect 8372 12496 9676 12536
rect 9716 12496 9725 12536
rect 14563 12496 14572 12536
rect 14612 12496 15244 12536
rect 15284 12496 15293 12536
rect 23587 12496 23596 12536
rect 23636 12496 23732 12536
rect 23779 12496 23788 12536
rect 23828 12496 26764 12536
rect 26804 12496 26813 12536
rect 7660 12452 7700 12496
rect 7555 12412 7564 12452
rect 7604 12412 7613 12452
rect 7660 12412 8524 12452
rect 8564 12412 8573 12452
rect 10723 12412 10732 12452
rect 10772 12412 10828 12452
rect 10868 12412 11020 12452
rect 11060 12412 11069 12452
rect 12643 12412 12652 12452
rect 12692 12412 12940 12452
rect 12980 12412 12989 12452
rect 13603 12412 13612 12452
rect 13652 12412 15148 12452
rect 15188 12412 15197 12452
rect 7564 12368 7604 12412
rect 7564 12328 8332 12368
rect 8372 12328 8381 12368
rect 8813 12328 8908 12368
rect 8948 12328 8957 12368
rect 11107 12244 11116 12284
rect 11156 12244 11165 12284
rect 18499 12244 18508 12284
rect 18548 12244 20140 12284
rect 20180 12244 20189 12284
rect 11116 12200 11156 12244
rect 10723 12160 10732 12200
rect 10772 12160 11156 12200
rect 3103 12076 3112 12116
rect 3480 12076 3489 12116
rect 10877 12076 10886 12116
rect 11254 12076 11263 12116
rect 14755 12076 14764 12116
rect 14804 12076 15436 12116
rect 15476 12076 15485 12116
rect 18651 12076 18660 12116
rect 19028 12076 19037 12116
rect 23692 12032 23732 12496
rect 23875 12412 23884 12452
rect 23924 12412 28396 12452
rect 28436 12412 28445 12452
rect 26425 12076 26434 12116
rect 26802 12076 26811 12116
rect 13219 11992 13228 12032
rect 13268 11992 13516 12032
rect 13556 11992 13565 12032
rect 23683 11992 23692 12032
rect 23732 11992 23741 12032
rect 13891 11908 13900 11948
rect 13940 11908 14668 11948
rect 14708 11908 14717 11948
rect 16483 11908 16492 11948
rect 16532 11908 16780 11948
rect 16820 11908 16829 11948
rect 12931 11824 12940 11864
rect 12980 11824 15244 11864
rect 15284 11824 15293 11864
rect 22627 11824 22636 11864
rect 22676 11824 23980 11864
rect 24020 11824 24029 11864
rect 5827 11740 5836 11780
rect 5876 11740 6028 11780
rect 6068 11740 6077 11780
rect 6691 11740 6700 11780
rect 6740 11740 9964 11780
rect 10004 11740 10013 11780
rect 15139 11740 15148 11780
rect 15188 11740 18124 11780
rect 18164 11740 18173 11780
rect 20611 11740 20620 11780
rect 20660 11740 23884 11780
rect 23924 11740 23933 11780
rect 7075 11656 7084 11696
rect 7124 11656 8236 11696
rect 8276 11656 8285 11696
rect 10531 11656 10540 11696
rect 10580 11656 11884 11696
rect 11924 11656 11933 11696
rect 14275 11656 14284 11696
rect 14324 11656 16300 11696
rect 16340 11656 16349 11696
rect 16579 11656 16588 11696
rect 16628 11656 17644 11696
rect 17684 11656 17693 11696
rect 20419 11656 20428 11696
rect 20468 11656 22060 11696
rect 22100 11656 22109 11696
rect 22723 11656 22732 11696
rect 22772 11656 25516 11696
rect 25556 11656 26188 11696
rect 26228 11656 26237 11696
rect 27331 11656 27340 11696
rect 27380 11656 27389 11696
rect 27340 11612 27380 11656
rect 15235 11572 15244 11612
rect 15284 11572 16396 11612
rect 16436 11572 16445 11612
rect 17347 11572 17356 11612
rect 17396 11572 18220 11612
rect 18260 11572 18269 11612
rect 27340 11572 28204 11612
rect 28244 11572 28253 11612
rect 7267 11488 7276 11528
rect 7316 11488 8620 11528
rect 8660 11488 8669 11528
rect 13507 11488 13516 11528
rect 13556 11488 19180 11528
rect 19220 11488 19229 11528
rect 15907 11404 15916 11444
rect 15956 11404 16780 11444
rect 16820 11404 16829 11444
rect 4343 11320 4352 11360
rect 4720 11320 4729 11360
rect 6307 11320 6316 11360
rect 6356 11320 6796 11360
rect 6836 11320 6845 11360
rect 12117 11320 12126 11360
rect 12494 11320 12503 11360
rect 16387 11320 16396 11360
rect 16436 11320 19660 11360
rect 19700 11320 19709 11360
rect 19891 11320 19900 11360
rect 20268 11320 20277 11360
rect 27665 11320 27674 11360
rect 28042 11320 28051 11360
rect 2563 11236 2572 11276
rect 2612 11236 6508 11276
rect 6548 11236 6557 11276
rect 15331 11236 15340 11276
rect 15380 11236 17260 11276
rect 17300 11236 17309 11276
rect 4195 11152 4204 11192
rect 4244 11152 8716 11192
rect 8756 11152 8765 11192
rect 14275 11152 14284 11192
rect 14324 11152 14333 11192
rect 22819 11152 22828 11192
rect 22868 11152 22908 11192
rect 4291 11068 4300 11108
rect 4340 11068 4876 11108
rect 4916 11068 4925 11108
rect 14284 11024 14324 11152
rect 22828 11108 22868 11152
rect 22243 11068 22252 11108
rect 22292 11068 23500 11108
rect 23540 11068 24748 11108
rect 24788 11068 24797 11108
rect 4387 10984 4396 11024
rect 4436 10984 5164 11024
rect 5204 10984 5213 11024
rect 8237 10984 8332 11024
rect 8372 10984 8381 11024
rect 10243 10984 10252 11024
rect 10292 10984 10732 11024
rect 10772 10984 11020 11024
rect 11060 10984 11069 11024
rect 13891 10984 13900 11024
rect 13940 10984 14324 11024
rect 15235 10984 15244 11024
rect 15284 10984 17356 11024
rect 17396 10984 17405 11024
rect 22051 10984 22060 11024
rect 22100 10984 28108 11024
rect 28148 10984 28157 11024
rect 4483 10900 4492 10940
rect 4532 10900 9772 10940
rect 9812 10900 9821 10940
rect 11299 10900 11308 10940
rect 11348 10900 11500 10940
rect 11540 10900 11549 10940
rect 14563 10900 14572 10940
rect 14612 10900 17836 10940
rect 17876 10900 17885 10940
rect 18499 10900 18508 10940
rect 18548 10900 18892 10940
rect 18932 10900 18941 10940
rect 7651 10816 7660 10856
rect 7700 10816 9100 10856
rect 9140 10816 9149 10856
rect 10147 10816 10156 10856
rect 10196 10816 11884 10856
rect 11924 10816 11933 10856
rect 13987 10732 13996 10772
rect 14036 10732 19180 10772
rect 19220 10732 19229 10772
rect 10531 10648 10540 10688
rect 10580 10648 13324 10688
rect 13364 10648 14956 10688
rect 14996 10648 17644 10688
rect 17684 10648 17693 10688
rect 3103 10564 3112 10604
rect 3480 10564 3489 10604
rect 7075 10564 7084 10604
rect 7124 10564 7564 10604
rect 7604 10564 7613 10604
rect 10877 10564 10886 10604
rect 11254 10564 11263 10604
rect 18651 10564 18660 10604
rect 19028 10564 19037 10604
rect 26425 10564 26434 10604
rect 26802 10564 26811 10604
rect 8611 10480 8620 10520
rect 8660 10480 14668 10520
rect 14708 10480 14717 10520
rect 2275 10396 2284 10436
rect 2324 10396 9292 10436
rect 9332 10396 9341 10436
rect 15811 10396 15820 10436
rect 15860 10396 17548 10436
rect 17588 10396 19564 10436
rect 19604 10396 19613 10436
rect 6787 10312 6796 10352
rect 6836 10312 8524 10352
rect 8564 10312 8573 10352
rect 8909 10312 9004 10352
rect 9044 10312 9053 10352
rect 16099 10312 16108 10352
rect 16148 10312 17836 10352
rect 17876 10312 17885 10352
rect 4675 10228 4684 10268
rect 4724 10228 6508 10268
rect 6548 10228 6557 10268
rect 6979 10228 6988 10268
rect 7028 10228 8620 10268
rect 8660 10228 8669 10268
rect 11309 10228 11404 10268
rect 11444 10228 11453 10268
rect 3523 10144 3532 10184
rect 3572 10144 4588 10184
rect 4628 10144 4637 10184
rect 4963 10144 4972 10184
rect 5012 10144 6892 10184
rect 6932 10144 6941 10184
rect 8995 10144 9004 10184
rect 9044 10144 9196 10184
rect 9236 10144 9245 10184
rect 10060 10144 10156 10184
rect 10196 10144 10205 10184
rect 15437 10144 15532 10184
rect 15572 10144 15724 10184
rect 15764 10144 15773 10184
rect 10060 10100 10100 10144
rect 10051 10060 10060 10100
rect 10100 10060 10109 10100
rect 18029 10060 18124 10100
rect 18164 10060 18173 10100
rect 23885 10060 23980 10100
rect 24020 10060 24029 10100
rect 6307 9976 6316 10016
rect 6356 9976 6988 10016
rect 7028 9976 7037 10016
rect 8419 9976 8428 10016
rect 8468 9976 9004 10016
rect 9044 9976 9053 10016
rect 12355 9976 12364 10016
rect 12404 9976 12413 10016
rect 13027 9976 13036 10016
rect 13076 9976 13228 10016
rect 13268 9976 14188 10016
rect 14228 9976 18508 10016
rect 18548 9976 18557 10016
rect 12364 9932 12404 9976
rect 6691 9892 6700 9932
rect 6740 9892 6892 9932
rect 6932 9892 8332 9932
rect 8372 9892 8381 9932
rect 9868 9892 12404 9932
rect 14947 9892 14956 9932
rect 14996 9892 16108 9932
rect 16148 9892 16157 9932
rect 4343 9808 4352 9848
rect 4720 9808 4729 9848
rect 7363 9808 7372 9848
rect 7412 9808 9388 9848
rect 9428 9808 9437 9848
rect 9868 9764 9908 9892
rect 12117 9808 12126 9848
rect 12494 9808 12503 9848
rect 19891 9808 19900 9848
rect 20268 9808 20277 9848
rect 27427 9808 27436 9848
rect 27476 9808 27485 9848
rect 27665 9808 27674 9848
rect 28042 9808 28051 9848
rect 8035 9724 8044 9764
rect 8084 9724 8716 9764
rect 8756 9724 9908 9764
rect 27436 9680 27476 9808
rect 2371 9640 2380 9680
rect 2420 9640 5548 9680
rect 5588 9640 9196 9680
rect 9236 9640 9245 9680
rect 10627 9640 10636 9680
rect 10676 9640 10828 9680
rect 10868 9640 10877 9680
rect 12931 9640 12940 9680
rect 12980 9640 20620 9680
rect 20660 9640 20669 9680
rect 27436 9640 27628 9680
rect 27668 9640 27677 9680
rect 5635 9556 5644 9596
rect 5684 9556 7948 9596
rect 7988 9556 7997 9596
rect 11203 9556 11212 9596
rect 11252 9556 13612 9596
rect 13652 9556 13661 9596
rect 19555 9556 19564 9596
rect 19604 9556 20140 9596
rect 20180 9556 20189 9596
rect 24355 9556 24364 9596
rect 24404 9556 30220 9596
rect 30260 9556 30269 9596
rect 10243 9472 10252 9512
rect 10292 9472 10924 9512
rect 10964 9472 10973 9512
rect 12739 9472 12748 9512
rect 12788 9472 15820 9512
rect 15860 9472 15869 9512
rect 23491 9472 23500 9512
rect 23540 9472 25036 9512
rect 25076 9472 25085 9512
rect 25891 9472 25900 9512
rect 25940 9472 26860 9512
rect 26900 9472 26909 9512
rect 10924 9428 10964 9472
rect 10924 9388 13036 9428
rect 13076 9388 13085 9428
rect 17635 9388 17644 9428
rect 17684 9388 19948 9428
rect 19988 9388 19997 9428
rect 11683 9304 11692 9344
rect 11732 9304 15724 9344
rect 15764 9304 20140 9344
rect 20180 9304 20189 9344
rect 13411 9220 13420 9260
rect 13460 9220 17260 9260
rect 17300 9220 17309 9260
rect 10627 9136 10636 9176
rect 10676 9136 20428 9176
rect 20468 9136 20477 9176
rect 3103 9052 3112 9092
rect 3480 9052 3489 9092
rect 10877 9052 10886 9092
rect 11254 9052 11263 9092
rect 18651 9052 18660 9092
rect 19028 9052 19037 9092
rect 26425 9052 26434 9092
rect 26802 9052 26811 9092
rect 11395 8968 11404 9008
rect 11444 8968 19852 9008
rect 19892 8968 19901 9008
rect 13219 8884 13228 8924
rect 13268 8884 14956 8924
rect 14996 8884 15005 8924
rect 16675 8884 16684 8924
rect 16724 8884 18124 8924
rect 18164 8884 18173 8924
rect 23395 8632 23404 8672
rect 23444 8632 24940 8672
rect 24980 8632 24989 8672
rect 10435 8464 10444 8504
rect 10484 8464 16012 8504
rect 16052 8464 16061 8504
rect 4343 8296 4352 8336
rect 4720 8296 4729 8336
rect 12117 8296 12126 8336
rect 12494 8296 12503 8336
rect 19891 8296 19900 8336
rect 20268 8296 20277 8336
rect 27665 8296 27674 8336
rect 28042 8296 28051 8336
rect 18115 8128 18124 8168
rect 18164 8128 19468 8168
rect 19508 8128 19517 8168
rect 6691 7960 6700 8000
rect 6740 7960 7852 8000
rect 7892 7960 7901 8000
rect 14083 7960 14092 8000
rect 14132 7960 19852 8000
rect 19892 7960 19901 8000
rect 18595 7876 18604 7916
rect 18644 7876 19084 7916
rect 19124 7876 19133 7916
rect 3103 7540 3112 7580
rect 3480 7540 3489 7580
rect 10877 7540 10886 7580
rect 11254 7540 11263 7580
rect 18651 7540 18660 7580
rect 19028 7540 19037 7580
rect 26425 7540 26434 7580
rect 26802 7540 26811 7580
rect 2851 7120 2860 7160
rect 2900 7120 4972 7160
rect 5012 7120 5021 7160
rect 18115 7120 18124 7160
rect 18164 7120 18604 7160
rect 18644 7120 18653 7160
rect 20131 7120 20140 7160
rect 20180 7120 20428 7160
rect 20468 7120 20477 7160
rect 17923 7036 17932 7076
rect 17972 7036 18412 7076
rect 18452 7036 18461 7076
rect 23107 7036 23116 7076
rect 23156 7036 28300 7076
rect 28340 7036 28780 7076
rect 28820 7036 28829 7076
rect 4099 6952 4108 6992
rect 4148 6952 4492 6992
rect 4532 6952 4780 6992
rect 4820 6952 4829 6992
rect 4343 6784 4352 6824
rect 4720 6784 4729 6824
rect 12117 6784 12126 6824
rect 12494 6784 12503 6824
rect 19891 6784 19900 6824
rect 20268 6784 20277 6824
rect 27665 6784 27674 6824
rect 28042 6784 28051 6824
rect 16483 6532 16492 6572
rect 16532 6532 16684 6572
rect 16724 6532 16733 6572
rect 11971 6448 11980 6488
rect 12020 6448 13900 6488
rect 13940 6448 13949 6488
rect 12931 6364 12940 6404
rect 12980 6364 13516 6404
rect 13556 6364 14188 6404
rect 14228 6364 14237 6404
rect 17635 6364 17644 6404
rect 17684 6364 22060 6404
rect 22100 6364 22109 6404
rect 16387 6280 16396 6320
rect 16436 6280 20140 6320
rect 20180 6280 20189 6320
rect 3103 6028 3112 6068
rect 3480 6028 3489 6068
rect 10877 6028 10886 6068
rect 11254 6028 11263 6068
rect 18651 6028 18660 6068
rect 19028 6028 19037 6068
rect 26425 6028 26434 6068
rect 26802 6028 26811 6068
rect 12451 5608 12460 5648
rect 12500 5608 13036 5648
rect 13076 5608 13085 5648
rect 14851 5608 14860 5648
rect 14900 5608 16684 5648
rect 16724 5608 16733 5648
rect 25507 5608 25516 5648
rect 25556 5608 28012 5648
rect 28052 5608 29644 5648
rect 29684 5608 30124 5648
rect 30164 5608 30173 5648
rect 4343 5272 4352 5312
rect 4720 5272 4729 5312
rect 12117 5272 12126 5312
rect 12494 5272 12503 5312
rect 19891 5272 19900 5312
rect 20268 5272 20277 5312
rect 27665 5272 27674 5312
rect 28042 5272 28051 5312
rect 8611 5020 8620 5060
rect 8660 5020 10924 5060
rect 10964 5020 13228 5060
rect 13268 5020 13277 5060
rect 6307 4936 6316 4976
rect 6356 4936 8428 4976
rect 8468 4936 9484 4976
rect 9524 4936 9533 4976
rect 16771 4936 16780 4976
rect 16820 4936 17356 4976
rect 17396 4936 17405 4976
rect 3103 4516 3112 4556
rect 3480 4516 3489 4556
rect 10877 4516 10886 4556
rect 11254 4516 11263 4556
rect 18651 4516 18660 4556
rect 19028 4516 19037 4556
rect 26425 4516 26434 4556
rect 26802 4516 26811 4556
rect 5251 4096 5260 4136
rect 5300 4096 7276 4136
rect 7316 4096 7325 4136
rect 26467 4096 26476 4136
rect 26516 4096 27436 4136
rect 27476 4096 27485 4136
rect 4343 3760 4352 3800
rect 4720 3760 4729 3800
rect 12117 3760 12126 3800
rect 12494 3760 12503 3800
rect 19891 3760 19900 3800
rect 20268 3760 20277 3800
rect 27665 3760 27674 3800
rect 28042 3760 28051 3800
rect 3103 3004 3112 3044
rect 3480 3004 3489 3044
rect 10877 3004 10886 3044
rect 11254 3004 11263 3044
rect 18651 3004 18660 3044
rect 19028 3004 19037 3044
rect 26425 3004 26434 3044
rect 26802 3004 26811 3044
rect 16195 2584 16204 2624
rect 16244 2584 17164 2624
rect 17204 2584 17213 2624
rect 4343 2248 4352 2288
rect 4720 2248 4729 2288
rect 12117 2248 12126 2288
rect 12494 2248 12503 2288
rect 19891 2248 19900 2288
rect 20268 2248 20277 2288
rect 27665 2248 27674 2288
rect 28042 2248 28051 2288
rect 12163 1912 12172 1952
rect 12212 1912 12652 1952
rect 12692 1912 13516 1952
rect 13556 1912 13565 1952
rect 3103 1492 3112 1532
rect 3480 1492 3489 1532
rect 10877 1492 10886 1532
rect 11254 1492 11263 1532
rect 18651 1492 18660 1532
rect 19028 1492 19037 1532
rect 26425 1492 26434 1532
rect 26802 1492 26811 1532
rect 8429 1072 8524 1112
rect 8564 1072 8573 1112
rect 4343 736 4352 776
rect 4720 736 4729 776
rect 12117 736 12126 776
rect 12494 736 12503 776
rect 19891 736 19900 776
rect 20268 736 20277 776
rect 27665 736 27674 776
rect 28042 736 28051 776
<< via4 >>
rect 4352 27952 4720 27992
rect 12126 27952 12494 27992
rect 19900 27952 20268 27992
rect 27674 27952 28042 27992
rect 3112 27196 3480 27236
rect 10886 27196 11254 27236
rect 18660 27196 19028 27236
rect 26434 27196 26802 27236
rect 4352 26440 4720 26480
rect 12126 26440 12494 26480
rect 19900 26440 20268 26480
rect 27674 26440 28042 26480
rect 3112 25684 3480 25724
rect 10540 25684 10580 25724
rect 10886 25684 11254 25724
rect 18660 25684 19028 25724
rect 26434 25684 26802 25724
rect 10540 25264 10580 25304
rect 4352 24928 4720 24968
rect 12126 24928 12494 24968
rect 19900 24928 20268 24968
rect 27674 24928 28042 24968
rect 25804 24676 25844 24716
rect 3112 24172 3480 24212
rect 10886 24172 11254 24212
rect 18660 24172 19028 24212
rect 26434 24172 26802 24212
rect 4352 23416 4720 23456
rect 12126 23416 12494 23456
rect 19900 23416 20268 23456
rect 27674 23416 28042 23456
rect 25804 22828 25844 22868
rect 3112 22660 3480 22700
rect 10886 22660 11254 22700
rect 18660 22660 19028 22700
rect 26434 22660 26802 22700
rect 4352 21904 4720 21944
rect 12126 21904 12494 21944
rect 19900 21904 20268 21944
rect 27674 21904 28042 21944
rect 3112 21148 3480 21188
rect 10886 21148 11254 21188
rect 18660 21148 19028 21188
rect 26434 21148 26802 21188
rect 23500 20644 23540 20684
rect 4352 20392 4720 20432
rect 12126 20392 12494 20432
rect 19900 20392 20268 20432
rect 27674 20392 28042 20432
rect 3112 19636 3480 19676
rect 10886 19636 11254 19676
rect 18660 19636 19028 19676
rect 26434 19636 26802 19676
rect 4352 18880 4720 18920
rect 12126 18880 12494 18920
rect 19900 18880 20268 18920
rect 27674 18880 28042 18920
rect 19180 18544 19220 18584
rect 3112 18124 3480 18164
rect 10886 18124 11254 18164
rect 18660 18124 19028 18164
rect 26434 18124 26802 18164
rect 9004 17536 9044 17576
rect 18028 17536 18068 17576
rect 4352 17368 4720 17408
rect 10444 17368 10484 17408
rect 12126 17368 12494 17408
rect 19900 17368 20268 17408
rect 27674 17368 28042 17408
rect 10540 17200 10580 17240
rect 9004 16864 9044 16904
rect 11404 16864 11444 16904
rect 9964 16780 10004 16820
rect 15532 16780 15572 16820
rect 3112 16612 3480 16652
rect 10886 16612 11254 16652
rect 18660 16612 19028 16652
rect 26434 16612 26802 16652
rect 19180 16360 19220 16400
rect 19564 16276 19604 16316
rect 10444 16192 10484 16232
rect 8524 16024 8564 16064
rect 4352 15856 4720 15896
rect 12126 15856 12494 15896
rect 19900 15856 20268 15896
rect 27674 15856 28042 15896
rect 9964 15604 10004 15644
rect 9772 15520 9812 15560
rect 10540 15520 10580 15560
rect 8332 15352 8372 15392
rect 3112 15100 3480 15140
rect 10886 15100 11254 15140
rect 18660 15100 19028 15140
rect 26434 15100 26802 15140
rect 18508 14764 18548 14804
rect 19660 14680 19700 14720
rect 18124 14512 18164 14552
rect 4352 14344 4720 14384
rect 12126 14344 12494 14384
rect 19900 14344 20268 14384
rect 27674 14344 28042 14384
rect 19564 14092 19604 14132
rect 23980 14008 24020 14048
rect 23500 13840 23540 13880
rect 3112 13588 3480 13628
rect 10886 13588 11254 13628
rect 18660 13588 19028 13628
rect 26434 13588 26802 13628
rect 8908 13168 8948 13208
rect 19660 13168 19700 13208
rect 7084 13000 7124 13040
rect 24076 13000 24116 13040
rect 4352 12832 4720 12872
rect 12126 12832 12494 12872
rect 19900 12832 20268 12872
rect 24076 12832 24116 12872
rect 27674 12832 28042 12872
rect 18028 12748 18068 12788
rect 8332 12580 8372 12620
rect 10732 12412 10772 12452
rect 8908 12328 8948 12368
rect 18508 12244 18548 12284
rect 3112 12076 3480 12116
rect 10886 12076 11254 12116
rect 18660 12076 19028 12116
rect 26434 12076 26802 12116
rect 4352 11320 4720 11360
rect 12126 11320 12494 11360
rect 19900 11320 20268 11360
rect 27674 11320 28042 11360
rect 8332 10984 8372 11024
rect 10252 10984 10292 11024
rect 10732 10984 10772 11024
rect 9772 10900 9812 10940
rect 18508 10900 18548 10940
rect 3112 10564 3480 10604
rect 7084 10564 7124 10604
rect 10886 10564 11254 10604
rect 18660 10564 19028 10604
rect 26434 10564 26802 10604
rect 9004 10312 9044 10352
rect 11404 10228 11444 10268
rect 10156 10144 10196 10184
rect 15532 10144 15572 10184
rect 18124 10060 18164 10100
rect 23980 10060 24020 10100
rect 4352 9808 4720 9848
rect 12126 9808 12494 9848
rect 19900 9808 20268 9848
rect 27674 9808 28042 9848
rect 3112 9052 3480 9092
rect 10886 9052 11254 9092
rect 18660 9052 19028 9092
rect 26434 9052 26802 9092
rect 4352 8296 4720 8336
rect 12126 8296 12494 8336
rect 19900 8296 20268 8336
rect 27674 8296 28042 8336
rect 3112 7540 3480 7580
rect 10886 7540 11254 7580
rect 18660 7540 19028 7580
rect 26434 7540 26802 7580
rect 4352 6784 4720 6824
rect 12126 6784 12494 6824
rect 19900 6784 20268 6824
rect 27674 6784 28042 6824
rect 3112 6028 3480 6068
rect 10886 6028 11254 6068
rect 18660 6028 19028 6068
rect 26434 6028 26802 6068
rect 4352 5272 4720 5312
rect 12126 5272 12494 5312
rect 19900 5272 20268 5312
rect 27674 5272 28042 5312
rect 3112 4516 3480 4556
rect 10886 4516 11254 4556
rect 18660 4516 19028 4556
rect 26434 4516 26802 4556
rect 4352 3760 4720 3800
rect 12126 3760 12494 3800
rect 19900 3760 20268 3800
rect 27674 3760 28042 3800
rect 3112 3004 3480 3044
rect 10886 3004 11254 3044
rect 18660 3004 19028 3044
rect 26434 3004 26802 3044
rect 4352 2248 4720 2288
rect 12126 2248 12494 2288
rect 19900 2248 20268 2288
rect 27674 2248 28042 2288
rect 3112 1492 3480 1532
rect 10886 1492 11254 1532
rect 18660 1492 19028 1532
rect 26434 1492 26802 1532
rect 8524 1072 8564 1112
rect 4352 736 4720 776
rect 12126 736 12494 776
rect 19900 736 20268 776
rect 27674 736 28042 776
<< metal5 >>
rect 3076 27236 3516 28016
rect 3076 27196 3112 27236
rect 3480 27196 3516 27236
rect 3076 25724 3516 27196
rect 3076 25684 3112 25724
rect 3480 25684 3516 25724
rect 3076 24212 3516 25684
rect 3076 24172 3112 24212
rect 3480 24172 3516 24212
rect 3076 22700 3516 24172
rect 3076 22660 3112 22700
rect 3480 22660 3516 22700
rect 3076 21188 3516 22660
rect 3076 21148 3112 21188
rect 3480 21148 3516 21188
rect 3076 19676 3516 21148
rect 3076 19636 3112 19676
rect 3480 19636 3516 19676
rect 3076 18164 3516 19636
rect 3076 18124 3112 18164
rect 3480 18124 3516 18164
rect 3076 16652 3516 18124
rect 3076 16612 3112 16652
rect 3480 16612 3516 16652
rect 3076 15140 3516 16612
rect 3076 15100 3112 15140
rect 3480 15100 3516 15140
rect 3076 13628 3516 15100
rect 3076 13588 3112 13628
rect 3480 13588 3516 13628
rect 3076 12116 3516 13588
rect 3076 12076 3112 12116
rect 3480 12076 3516 12116
rect 3076 10604 3516 12076
rect 3076 10564 3112 10604
rect 3480 10564 3516 10604
rect 3076 9092 3516 10564
rect 3076 9052 3112 9092
rect 3480 9052 3516 9092
rect 3076 7580 3516 9052
rect 3076 7540 3112 7580
rect 3480 7540 3516 7580
rect 3076 6068 3516 7540
rect 3076 6028 3112 6068
rect 3480 6028 3516 6068
rect 3076 4556 3516 6028
rect 3076 4516 3112 4556
rect 3480 4516 3516 4556
rect 3076 3044 3516 4516
rect 3076 3004 3112 3044
rect 3480 3004 3516 3044
rect 3076 1532 3516 3004
rect 3076 1492 3112 1532
rect 3480 1492 3516 1532
rect 3076 712 3516 1492
rect 4316 27992 4756 28016
rect 4316 27952 4352 27992
rect 4720 27952 4756 27992
rect 4316 26480 4756 27952
rect 4316 26440 4352 26480
rect 4720 26440 4756 26480
rect 4316 24968 4756 26440
rect 10850 27236 11290 28016
rect 10850 27196 10886 27236
rect 11254 27196 11290 27236
rect 10540 25724 10580 25733
rect 10540 25304 10580 25684
rect 10540 25255 10580 25264
rect 10850 25724 11290 27196
rect 10850 25684 10886 25724
rect 11254 25684 11290 25724
rect 4316 24928 4352 24968
rect 4720 24928 4756 24968
rect 4316 23456 4756 24928
rect 4316 23416 4352 23456
rect 4720 23416 4756 23456
rect 4316 21944 4756 23416
rect 4316 21904 4352 21944
rect 4720 21904 4756 21944
rect 4316 20432 4756 21904
rect 4316 20392 4352 20432
rect 4720 20392 4756 20432
rect 4316 18920 4756 20392
rect 4316 18880 4352 18920
rect 4720 18880 4756 18920
rect 4316 17408 4756 18880
rect 10850 24212 11290 25684
rect 10850 24172 10886 24212
rect 11254 24172 11290 24212
rect 10850 22700 11290 24172
rect 10850 22660 10886 22700
rect 11254 22660 11290 22700
rect 10850 21188 11290 22660
rect 10850 21148 10886 21188
rect 11254 21148 11290 21188
rect 10850 19676 11290 21148
rect 10850 19636 10886 19676
rect 11254 19636 11290 19676
rect 10850 18164 11290 19636
rect 10850 18124 10886 18164
rect 11254 18124 11290 18164
rect 4316 17368 4352 17408
rect 4720 17368 4756 17408
rect 4316 15896 4756 17368
rect 9004 17576 9044 17585
rect 9004 16904 9044 17536
rect 4316 15856 4352 15896
rect 4720 15856 4756 15896
rect 4316 14384 4756 15856
rect 8524 16064 8564 16073
rect 4316 14344 4352 14384
rect 4720 14344 4756 14384
rect 4316 12872 4756 14344
rect 8332 15392 8372 15401
rect 4316 12832 4352 12872
rect 4720 12832 4756 12872
rect 4316 11360 4756 12832
rect 4316 11320 4352 11360
rect 4720 11320 4756 11360
rect 4316 9848 4756 11320
rect 7084 13040 7124 13049
rect 7084 10604 7124 13000
rect 8332 12620 8372 15352
rect 8332 11024 8372 12580
rect 8332 10975 8372 10984
rect 7084 10555 7124 10564
rect 4316 9808 4352 9848
rect 4720 9808 4756 9848
rect 4316 8336 4756 9808
rect 4316 8296 4352 8336
rect 4720 8296 4756 8336
rect 4316 6824 4756 8296
rect 4316 6784 4352 6824
rect 4720 6784 4756 6824
rect 4316 5312 4756 6784
rect 4316 5272 4352 5312
rect 4720 5272 4756 5312
rect 4316 3800 4756 5272
rect 4316 3760 4352 3800
rect 4720 3760 4756 3800
rect 4316 2288 4756 3760
rect 4316 2248 4352 2288
rect 4720 2248 4756 2288
rect 4316 776 4756 2248
rect 8524 1112 8564 16024
rect 8908 13208 8948 13217
rect 8908 12368 8948 13168
rect 8908 12319 8948 12328
rect 9004 10352 9044 16864
rect 10444 17408 10484 17417
rect 9964 16820 10004 16829
rect 9964 15644 10004 16780
rect 10444 16232 10484 17368
rect 10444 16183 10484 16192
rect 10540 17240 10580 17249
rect 9964 15595 10004 15604
rect 9772 15560 9812 15569
rect 9772 10940 9812 15520
rect 10540 15560 10580 17200
rect 10540 15511 10580 15520
rect 10850 16652 11290 18124
rect 12090 27992 12530 28016
rect 12090 27952 12126 27992
rect 12494 27952 12530 27992
rect 12090 26480 12530 27952
rect 12090 26440 12126 26480
rect 12494 26440 12530 26480
rect 12090 24968 12530 26440
rect 12090 24928 12126 24968
rect 12494 24928 12530 24968
rect 12090 23456 12530 24928
rect 12090 23416 12126 23456
rect 12494 23416 12530 23456
rect 12090 21944 12530 23416
rect 12090 21904 12126 21944
rect 12494 21904 12530 21944
rect 12090 20432 12530 21904
rect 12090 20392 12126 20432
rect 12494 20392 12530 20432
rect 12090 18920 12530 20392
rect 12090 18880 12126 18920
rect 12494 18880 12530 18920
rect 12090 17408 12530 18880
rect 18624 27236 19064 28016
rect 18624 27196 18660 27236
rect 19028 27196 19064 27236
rect 18624 25724 19064 27196
rect 18624 25684 18660 25724
rect 19028 25684 19064 25724
rect 18624 24212 19064 25684
rect 18624 24172 18660 24212
rect 19028 24172 19064 24212
rect 18624 22700 19064 24172
rect 18624 22660 18660 22700
rect 19028 22660 19064 22700
rect 18624 21188 19064 22660
rect 18624 21148 18660 21188
rect 19028 21148 19064 21188
rect 18624 19676 19064 21148
rect 18624 19636 18660 19676
rect 19028 19636 19064 19676
rect 18624 18164 19064 19636
rect 19864 27992 20304 28016
rect 19864 27952 19900 27992
rect 20268 27952 20304 27992
rect 19864 26480 20304 27952
rect 19864 26440 19900 26480
rect 20268 26440 20304 26480
rect 19864 24968 20304 26440
rect 19864 24928 19900 24968
rect 20268 24928 20304 24968
rect 19864 23456 20304 24928
rect 26398 27236 26838 28016
rect 26398 27196 26434 27236
rect 26802 27196 26838 27236
rect 26398 25724 26838 27196
rect 26398 25684 26434 25724
rect 26802 25684 26838 25724
rect 19864 23416 19900 23456
rect 20268 23416 20304 23456
rect 19864 21944 20304 23416
rect 25804 24716 25844 24725
rect 25804 22868 25844 24676
rect 25804 22819 25844 22828
rect 26398 24212 26838 25684
rect 26398 24172 26434 24212
rect 26802 24172 26838 24212
rect 19864 21904 19900 21944
rect 20268 21904 20304 21944
rect 19864 20432 20304 21904
rect 26398 22700 26838 24172
rect 26398 22660 26434 22700
rect 26802 22660 26838 22700
rect 26398 21188 26838 22660
rect 26398 21148 26434 21188
rect 26802 21148 26838 21188
rect 19864 20392 19900 20432
rect 20268 20392 20304 20432
rect 19864 18920 20304 20392
rect 19864 18880 19900 18920
rect 20268 18880 20304 18920
rect 18624 18124 18660 18164
rect 19028 18124 19064 18164
rect 12090 17368 12126 17408
rect 12494 17368 12530 17408
rect 10850 16612 10886 16652
rect 11254 16612 11290 16652
rect 10850 15140 11290 16612
rect 10850 15100 10886 15140
rect 11254 15100 11290 15140
rect 10850 13628 11290 15100
rect 10850 13588 10886 13628
rect 11254 13588 11290 13628
rect 10732 12452 10772 12461
rect 9772 10891 9812 10900
rect 10252 11024 10292 11033
rect 10252 10344 10292 10984
rect 10732 11024 10772 12412
rect 10732 10975 10772 10984
rect 10850 12116 11290 13588
rect 10850 12076 10886 12116
rect 11254 12076 11290 12116
rect 9004 10303 9044 10312
rect 10156 10304 10292 10344
rect 10850 10604 11290 12076
rect 10850 10564 10886 10604
rect 11254 10564 11290 10604
rect 10156 10184 10196 10304
rect 10156 10135 10196 10144
rect 8524 1063 8564 1072
rect 10850 9092 11290 10564
rect 11404 16904 11444 16913
rect 11404 10268 11444 16864
rect 11404 10219 11444 10228
rect 12090 15896 12530 17368
rect 18028 17576 18068 17585
rect 12090 15856 12126 15896
rect 12494 15856 12530 15896
rect 12090 14384 12530 15856
rect 12090 14344 12126 14384
rect 12494 14344 12530 14384
rect 12090 12872 12530 14344
rect 12090 12832 12126 12872
rect 12494 12832 12530 12872
rect 12090 11360 12530 12832
rect 12090 11320 12126 11360
rect 12494 11320 12530 11360
rect 10850 9052 10886 9092
rect 11254 9052 11290 9092
rect 10850 7580 11290 9052
rect 10850 7540 10886 7580
rect 11254 7540 11290 7580
rect 10850 6068 11290 7540
rect 10850 6028 10886 6068
rect 11254 6028 11290 6068
rect 10850 4556 11290 6028
rect 10850 4516 10886 4556
rect 11254 4516 11290 4556
rect 10850 3044 11290 4516
rect 10850 3004 10886 3044
rect 11254 3004 11290 3044
rect 10850 1532 11290 3004
rect 10850 1492 10886 1532
rect 11254 1492 11290 1532
rect 4316 736 4352 776
rect 4720 736 4756 776
rect 4316 712 4756 736
rect 10850 712 11290 1492
rect 12090 9848 12530 11320
rect 15532 16820 15572 16829
rect 15532 10184 15572 16780
rect 18028 12788 18068 17536
rect 18624 16652 19064 18124
rect 18624 16612 18660 16652
rect 19028 16612 19064 16652
rect 18624 15140 19064 16612
rect 19180 18584 19220 18593
rect 19180 16400 19220 18544
rect 19180 16351 19220 16360
rect 19864 17408 20304 18880
rect 19864 17368 19900 17408
rect 20268 17368 20304 17408
rect 18624 15100 18660 15140
rect 19028 15100 19064 15140
rect 18508 14804 18548 14813
rect 18028 12739 18068 12748
rect 18124 14552 18164 14561
rect 15532 10135 15572 10144
rect 18124 10100 18164 14512
rect 18508 12284 18548 14764
rect 18508 10940 18548 12244
rect 18508 10891 18548 10900
rect 18624 13628 19064 15100
rect 19564 16316 19604 16325
rect 19564 14132 19604 16276
rect 19864 15896 20304 17368
rect 19864 15856 19900 15896
rect 20268 15856 20304 15896
rect 19564 14083 19604 14092
rect 19660 14720 19700 14729
rect 18624 13588 18660 13628
rect 19028 13588 19064 13628
rect 18624 12116 19064 13588
rect 19660 13208 19700 14680
rect 19660 13159 19700 13168
rect 19864 14384 20304 15856
rect 19864 14344 19900 14384
rect 20268 14344 20304 14384
rect 18624 12076 18660 12116
rect 19028 12076 19064 12116
rect 18124 10051 18164 10060
rect 18624 10604 19064 12076
rect 18624 10564 18660 10604
rect 19028 10564 19064 10604
rect 12090 9808 12126 9848
rect 12494 9808 12530 9848
rect 12090 8336 12530 9808
rect 12090 8296 12126 8336
rect 12494 8296 12530 8336
rect 12090 6824 12530 8296
rect 12090 6784 12126 6824
rect 12494 6784 12530 6824
rect 12090 5312 12530 6784
rect 12090 5272 12126 5312
rect 12494 5272 12530 5312
rect 12090 3800 12530 5272
rect 12090 3760 12126 3800
rect 12494 3760 12530 3800
rect 12090 2288 12530 3760
rect 12090 2248 12126 2288
rect 12494 2248 12530 2288
rect 12090 776 12530 2248
rect 12090 736 12126 776
rect 12494 736 12530 776
rect 12090 712 12530 736
rect 18624 9092 19064 10564
rect 18624 9052 18660 9092
rect 19028 9052 19064 9092
rect 18624 7580 19064 9052
rect 18624 7540 18660 7580
rect 19028 7540 19064 7580
rect 18624 6068 19064 7540
rect 18624 6028 18660 6068
rect 19028 6028 19064 6068
rect 18624 4556 19064 6028
rect 18624 4516 18660 4556
rect 19028 4516 19064 4556
rect 18624 3044 19064 4516
rect 18624 3004 18660 3044
rect 19028 3004 19064 3044
rect 18624 1532 19064 3004
rect 18624 1492 18660 1532
rect 19028 1492 19064 1532
rect 18624 712 19064 1492
rect 19864 12872 20304 14344
rect 23500 20684 23540 20693
rect 23500 13880 23540 20644
rect 26398 19676 26838 21148
rect 26398 19636 26434 19676
rect 26802 19636 26838 19676
rect 26398 18164 26838 19636
rect 26398 18124 26434 18164
rect 26802 18124 26838 18164
rect 26398 16652 26838 18124
rect 26398 16612 26434 16652
rect 26802 16612 26838 16652
rect 26398 15140 26838 16612
rect 26398 15100 26434 15140
rect 26802 15100 26838 15140
rect 23500 13831 23540 13840
rect 23980 14048 24020 14057
rect 19864 12832 19900 12872
rect 20268 12832 20304 12872
rect 19864 11360 20304 12832
rect 19864 11320 19900 11360
rect 20268 11320 20304 11360
rect 19864 9848 20304 11320
rect 23980 10100 24020 14008
rect 26398 13628 26838 15100
rect 26398 13588 26434 13628
rect 26802 13588 26838 13628
rect 24076 13040 24116 13049
rect 24076 12872 24116 13000
rect 24076 12823 24116 12832
rect 23980 10051 24020 10060
rect 26398 12116 26838 13588
rect 26398 12076 26434 12116
rect 26802 12076 26838 12116
rect 26398 10604 26838 12076
rect 26398 10564 26434 10604
rect 26802 10564 26838 10604
rect 19864 9808 19900 9848
rect 20268 9808 20304 9848
rect 19864 8336 20304 9808
rect 19864 8296 19900 8336
rect 20268 8296 20304 8336
rect 19864 6824 20304 8296
rect 19864 6784 19900 6824
rect 20268 6784 20304 6824
rect 19864 5312 20304 6784
rect 19864 5272 19900 5312
rect 20268 5272 20304 5312
rect 19864 3800 20304 5272
rect 19864 3760 19900 3800
rect 20268 3760 20304 3800
rect 19864 2288 20304 3760
rect 19864 2248 19900 2288
rect 20268 2248 20304 2288
rect 19864 776 20304 2248
rect 19864 736 19900 776
rect 20268 736 20304 776
rect 19864 712 20304 736
rect 26398 9092 26838 10564
rect 26398 9052 26434 9092
rect 26802 9052 26838 9092
rect 26398 7580 26838 9052
rect 26398 7540 26434 7580
rect 26802 7540 26838 7580
rect 26398 6068 26838 7540
rect 26398 6028 26434 6068
rect 26802 6028 26838 6068
rect 26398 4556 26838 6028
rect 26398 4516 26434 4556
rect 26802 4516 26838 4556
rect 26398 3044 26838 4516
rect 26398 3004 26434 3044
rect 26802 3004 26838 3044
rect 26398 1532 26838 3004
rect 26398 1492 26434 1532
rect 26802 1492 26838 1532
rect 26398 712 26838 1492
rect 27638 27992 28078 28016
rect 27638 27952 27674 27992
rect 28042 27952 28078 27992
rect 27638 26480 28078 27952
rect 27638 26440 27674 26480
rect 28042 26440 28078 26480
rect 27638 24968 28078 26440
rect 27638 24928 27674 24968
rect 28042 24928 28078 24968
rect 27638 23456 28078 24928
rect 27638 23416 27674 23456
rect 28042 23416 28078 23456
rect 27638 21944 28078 23416
rect 27638 21904 27674 21944
rect 28042 21904 28078 21944
rect 27638 20432 28078 21904
rect 27638 20392 27674 20432
rect 28042 20392 28078 20432
rect 27638 18920 28078 20392
rect 27638 18880 27674 18920
rect 28042 18880 28078 18920
rect 27638 17408 28078 18880
rect 27638 17368 27674 17408
rect 28042 17368 28078 17408
rect 27638 15896 28078 17368
rect 27638 15856 27674 15896
rect 28042 15856 28078 15896
rect 27638 14384 28078 15856
rect 27638 14344 27674 14384
rect 28042 14344 28078 14384
rect 27638 12872 28078 14344
rect 27638 12832 27674 12872
rect 28042 12832 28078 12872
rect 27638 11360 28078 12832
rect 27638 11320 27674 11360
rect 28042 11320 28078 11360
rect 27638 9848 28078 11320
rect 27638 9808 27674 9848
rect 28042 9808 28078 9848
rect 27638 8336 28078 9808
rect 27638 8296 27674 8336
rect 28042 8296 28078 8336
rect 27638 6824 28078 8296
rect 27638 6784 27674 6824
rect 28042 6784 28078 6824
rect 27638 5312 28078 6784
rect 27638 5272 27674 5312
rect 28042 5272 28078 5312
rect 27638 3800 28078 5272
rect 27638 3760 27674 3800
rect 28042 3760 28078 3800
rect 27638 2288 28078 3760
rect 27638 2248 27674 2288
rect 28042 2248 28078 2288
rect 27638 776 28078 2248
rect 27638 736 27674 776
rect 28042 736 28078 776
rect 27638 712 28078 736
use sg13g2_inv_2  _1056_
timestamp 1747537721
transform -1 0 23712 0 -1 24948
box -48 -56 432 834
use sg13g2_inv_1  _1057_
timestamp 1747537721
transform -1 0 25824 0 1 2268
box -48 -56 336 834
use sg13g2_inv_1  _1058_
timestamp 1747537721
transform -1 0 23424 0 1 2268
box -48 -56 336 834
use sg13g2_inv_1  _1059_
timestamp 1747537721
transform -1 0 9696 0 -1 8316
box -48 -56 336 834
use sg13g2_inv_1  _1060_
timestamp 1747537721
transform 1 0 7968 0 -1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1061_
timestamp 1747537721
transform -1 0 11616 0 1 21924
box -48 -56 336 834
use sg13g2_inv_2  _1062_
timestamp 1747537721
transform 1 0 24384 0 1 15876
box -48 -56 432 834
use sg13g2_inv_2  _1063_
timestamp 1747537721
transform 1 0 24192 0 1 6804
box -48 -56 432 834
use sg13g2_inv_2  _1064_
timestamp 1747537721
transform 1 0 24864 0 1 9828
box -48 -56 432 834
use sg13g2_inv_1  _1065_
timestamp 1747537721
transform 1 0 23232 0 1 14364
box -48 -56 336 834
use sg13g2_inv_2  _1066_
timestamp 1747537721
transform 1 0 26976 0 1 9828
box -48 -56 432 834
use sg13g2_inv_1  _1067_
timestamp 1747537721
transform -1 0 26880 0 -1 12852
box -48 -56 336 834
use sg13g2_inv_1  _1068_
timestamp 1747537721
transform 1 0 27456 0 1 12852
box -48 -56 336 834
use sg13g2_inv_1  _1069_
timestamp 1747537721
transform -1 0 24096 0 -1 12852
box -48 -56 336 834
use sg13g2_inv_2  _1070_
timestamp 1747537721
transform 1 0 11328 0 1 14364
box -48 -56 432 834
use sg13g2_inv_1  _1071_
timestamp 1747537721
transform -1 0 7776 0 1 21924
box -48 -56 336 834
use sg13g2_inv_1  _1072_
timestamp 1747537721
transform 1 0 20160 0 -1 20412
box -48 -56 336 834
use sg13g2_inv_1  _1073_
timestamp 1747537721
transform -1 0 20160 0 1 24948
box -48 -56 336 834
use sg13g2_inv_1  _1074_
timestamp 1747537721
transform -1 0 14304 0 -1 27972
box -48 -56 336 834
use sg13g2_inv_1  _1075_
timestamp 1747537721
transform -1 0 17184 0 -1 27972
box -48 -56 336 834
use sg13g2_inv_1  _1076_
timestamp 1747537721
transform 1 0 10176 0 1 26460
box -48 -56 336 834
use sg13g2_inv_1  _1077_
timestamp 1747537721
transform 1 0 8736 0 -1 5292
box -48 -56 336 834
use sg13g2_inv_2  _1078_
timestamp 1747537721
transform -1 0 16416 0 -1 2268
box -48 -56 432 834
use sg13g2_o21ai_1  _1079_
timestamp 1747537721
transform -1 0 24288 0 -1 14364
box -48 -56 538 834
use sg13g2_nand3_1  _1080_
timestamp 1747537721
transform -1 0 28128 0 -1 12852
box -48 -56 528 834
use sg13g2_nor2_1  _1081_
timestamp 1747537721
transform -1 0 25632 0 -1 12852
box -48 -56 432 834
use sg13g2_a21oi_1  _1082_
timestamp 1747537721
transform -1 0 23616 0 1 12852
box -48 -56 528 834
use sg13g2_a21oi_1  _1083_
timestamp 1747537721
transform 1 0 23616 0 1 12852
box -48 -56 528 834
use sg13g2_nor2_1  _1084_
timestamp 1747537721
transform 1 0 21696 0 -1 11340
box -48 -56 432 834
use sg13g2_nand2b_1  _1085_
timestamp 1747537721
transform 1 0 25248 0 -1 14364
box -48 -56 528 834
use sg13g2_nor3_1  _1086_
timestamp 1747537721
transform 1 0 25152 0 1 12852
box -48 -56 528 834
use sg13g2_nor2_1  _1087_
timestamp 1747537721
transform -1 0 23808 0 -1 12852
box -48 -56 432 834
use sg13g2_nand3_1  _1088_
timestamp 1747537721
transform 1 0 24096 0 1 12852
box -48 -56 528 834
use sg13g2_a21oi_1  _1089_
timestamp 1747537721
transform -1 0 24768 0 -1 14364
box -48 -56 528 834
use sg13g2_a22oi_1  _1090_
timestamp 1747537721
transform 1 0 23232 0 -1 14364
box -48 -56 624 834
use sg13g2_inv_1  _1091_
timestamp 1747537721
transform 1 0 12096 0 1 21924
box -48 -56 336 834
use sg13g2_and2_2  _1092_
timestamp 1747537721
transform -1 0 27264 0 -1 20412
box -48 -56 624 834
use sg13g2_nand2_1  _1093_
timestamp 1747537721
transform -1 0 26496 0 1 23436
box -48 -56 432 834
use sg13g2_nor2_1  _1094_
timestamp 1747537721
transform 1 0 26880 0 -1 24948
box -48 -56 432 834
use sg13g2_or2_1  _1095_
timestamp 1747537721
transform 1 0 24864 0 1 21924
box -48 -56 528 834
use sg13g2_nor2_1  _1096_
timestamp 1747537721
transform -1 0 26112 0 -1 23436
box -48 -56 432 834
use sg13g2_a21o_1  _1097_
timestamp 1747537721
transform 1 0 25536 0 1 21924
box -48 -56 720 834
use sg13g2_nand2_1  _1098_
timestamp 1747537721
transform 1 0 27072 0 -1 23436
box -48 -56 432 834
use sg13g2_nand3_1  _1099_
timestamp 1747537721
transform -1 0 27744 0 1 21924
box -48 -56 528 834
use sg13g2_nor3_2  _1100_
timestamp 1747537721
transform 1 0 26400 0 1 21924
box -48 -56 912 834
use sg13g2_inv_1  _1101_
timestamp 1747537721
transform 1 0 24096 0 -1 23436
box -48 -56 336 834
use sg13g2_nor2_1  _1102_
timestamp 1747537721
transform -1 0 27168 0 -1 26460
box -48 -56 432 834
use sg13g2_and2_1  _1103_
timestamp 1747537721
transform 1 0 26496 0 1 23436
box -48 -56 528 834
use sg13g2_nor2b_1  _1104_
timestamp 1747537721
transform 1 0 27456 0 -1 21924
box -54 -56 528 834
use sg13g2_a221oi_1  _1105_
timestamp 1747537721
transform 1 0 26208 0 -1 23436
box -48 -56 816 834
use sg13g2_a21oi_2  _1106_
timestamp 1747537721
transform 1 0 24960 0 -1 23436
box -48 -56 816 834
use sg13g2_and2_2  _1107_
timestamp 1747537721
transform 1 0 20160 0 -1 21924
box -48 -56 624 834
use sg13g2_nand2_1  _1108_
timestamp 1747537721
transform -1 0 19968 0 1 20412
box -48 -56 432 834
use sg13g2_nor2_1  _1109_
timestamp 1747537721
transform -1 0 9600 0 1 23436
box -48 -56 432 834
use sg13g2_a21oi_1  _1110_
timestamp 1747537721
transform 1 0 7872 0 1 23436
box -48 -56 528 834
use sg13g2_nand2_1  _1111_
timestamp 1747537721
transform 1 0 4608 0 -1 23436
box -48 -56 432 834
use sg13g2_nor2_1  _1112_
timestamp 1747537721
transform -1 0 4896 0 -1 24948
box -48 -56 432 834
use sg13g2_a21oi_1  _1113_
timestamp 1747537721
transform 1 0 5184 0 1 23436
box -48 -56 528 834
use sg13g2_o21ai_1  _1114_
timestamp 1747537721
transform -1 0 5184 0 1 23436
box -48 -56 538 834
use sg13g2_nor2_1  _1115_
timestamp 1747537721
transform -1 0 9984 0 1 23436
box -48 -56 432 834
use sg13g2_a21oi_2  _1116_
timestamp 1747537721
transform -1 0 11232 0 -1 24948
box -48 -56 816 834
use sg13g2_nor2_1  _1117_
timestamp 1747537721
transform 1 0 5376 0 -1 24948
box -48 -56 432 834
use sg13g2_or2_1  _1118_
timestamp 1747537721
transform -1 0 5376 0 -1 24948
box -48 -56 528 834
use sg13g2_inv_1  _1119_
timestamp 1747537721
transform 1 0 8064 0 -1 26460
box -48 -56 336 834
use sg13g2_nor2_1  _1120_
timestamp 1747537721
transform -1 0 4032 0 1 26460
box -48 -56 432 834
use sg13g2_nor2_1  _1121_
timestamp 1747537721
transform 1 0 4896 0 1 24948
box -48 -56 432 834
use sg13g2_a21oi_1  _1122_
timestamp 1747537721
transform 1 0 4416 0 1 24948
box -48 -56 528 834
use sg13g2_nor2_1  _1123_
timestamp 1747537721
transform -1 0 5376 0 -1 26460
box -48 -56 432 834
use sg13g2_xnor2_1  _1124_
timestamp 1747537721
transform -1 0 24000 0 1 23436
box -48 -56 816 834
use sg13g2_nor2_2  _1125_
timestamp 1747537721
transform 1 0 12960 0 1 18900
box -48 -56 624 834
use sg13g2_and2_1  _1126_
timestamp 1747537721
transform 1 0 15648 0 -1 20412
box -48 -56 528 834
use sg13g2_nand2_1  _1127_
timestamp 1747537721
transform -1 0 14976 0 -1 18900
box -48 -56 432 834
use sg13g2_nand2_2  _1128_
timestamp 1747537721
transform -1 0 12096 0 -1 21924
box -48 -56 624 834
use sg13g2_o21ai_1  _1129_
timestamp 1747537721
transform -1 0 20832 0 1 20412
box -48 -56 538 834
use sg13g2_and2_2  _1130_
timestamp 1747537721
transform -1 0 20160 0 -1 21924
box -48 -56 624 834
use sg13g2_o21ai_1  _1131_
timestamp 1747537721
transform 1 0 7968 0 1 20412
box -48 -56 538 834
use sg13g2_nand3b_1  _1132_
timestamp 1747537721
transform -1 0 27840 0 -1 14364
box -48 -56 720 834
use sg13g2_nor2_2  _1133_
timestamp 1747537721
transform -1 0 27648 0 1 14364
box -48 -56 624 834
use sg13g2_nor2_2  _1134_
timestamp 1747537721
transform -1 0 7488 0 -1 20412
box -48 -56 624 834
use sg13g2_xnor2_1  _1135_
timestamp 1747537721
transform 1 0 22464 0 1 18900
box -48 -56 816 834
use sg13g2_nand2_1  _1136_
timestamp 1747537721
transform 1 0 23424 0 1 21924
box -48 -56 432 834
use sg13g2_xnor2_1  _1137_
timestamp 1747537721
transform -1 0 23424 0 1 21924
box -48 -56 816 834
use sg13g2_inv_1  _1138_
timestamp 1747537721
transform -1 0 23040 0 -1 21924
box -48 -56 336 834
use sg13g2_nand2_1  _1139_
timestamp 1747537721
transform 1 0 15360 0 -1 26460
box -48 -56 432 834
use sg13g2_nand2_1  _1140_
timestamp 1747537721
transform 1 0 14208 0 1 24948
box -48 -56 432 834
use sg13g2_xnor2_1  _1141_
timestamp 1747537721
transform 1 0 15744 0 -1 26460
box -48 -56 816 834
use sg13g2_o21ai_1  _1142_
timestamp 1747537721
transform 1 0 16512 0 -1 26460
box -48 -56 538 834
use sg13g2_and2_1  _1143_
timestamp 1747537721
transform 1 0 18048 0 -1 26460
box -48 -56 528 834
use sg13g2_xor2_1  _1144_
timestamp 1747537721
transform -1 0 18048 0 -1 26460
box -48 -56 816 834
use sg13g2_nand2_1  _1145_
timestamp 1747537721
transform 1 0 18624 0 1 24948
box -48 -56 432 834
use sg13g2_a21oi_1  _1146_
timestamp 1747537721
transform 1 0 19008 0 -1 26460
box -48 -56 528 834
use sg13g2_a22oi_1  _1147_
timestamp 1747537721
transform -1 0 20544 0 -1 24948
box -48 -56 624 834
use sg13g2_and2_1  _1148_
timestamp 1747537721
transform 1 0 18528 0 1 21924
box -48 -56 528 834
use sg13g2_or2_1  _1149_
timestamp 1747537721
transform 1 0 18720 0 1 23436
box -48 -56 528 834
use sg13g2_xnor2_1  _1150_
timestamp 1747537721
transform 1 0 18048 0 -1 23436
box -48 -56 816 834
use sg13g2_nand2_1  _1151_
timestamp 1747537721
transform 1 0 21600 0 -1 23436
box -48 -56 432 834
use sg13g2_xnor2_1  _1152_
timestamp 1747537721
transform -1 0 21120 0 -1 23436
box -48 -56 816 834
use sg13g2_nor2_1  _1153_
timestamp 1747537721
transform 1 0 19200 0 1 23436
box -48 -56 432 834
use sg13g2_inv_1  _1154_
timestamp 1747537721
transform 1 0 18912 0 -1 24948
box -48 -56 336 834
use sg13g2_a221oi_1  _1155_
timestamp 1747537721
transform 1 0 19200 0 -1 24948
box -48 -56 816 834
use sg13g2_o21ai_1  _1156_
timestamp 1747537721
transform -1 0 21600 0 -1 23436
box -48 -56 538 834
use sg13g2_nand2_1  _1157_
timestamp 1747537721
transform 1 0 21024 0 1 21924
box -48 -56 432 834
use sg13g2_nor2_1  _1158_
timestamp 1747537721
transform 1 0 21792 0 -1 21924
box -48 -56 432 834
use sg13g2_o21ai_1  _1159_
timestamp 1747537721
transform 1 0 21408 0 1 21924
box -48 -56 538 834
use sg13g2_a21oi_2  _1160_
timestamp 1747537721
transform -1 0 24000 0 1 18900
box -48 -56 816 834
use sg13g2_a21o_1  _1161_
timestamp 1747537721
transform -1 0 24672 0 1 18900
box -48 -56 720 834
use sg13g2_a21oi_1  _1162_
timestamp 1747537721
transform -1 0 24576 0 -1 17388
box -48 -56 528 834
use sg13g2_and3_1  _1163_
timestamp 1747537721
transform -1 0 25248 0 1 17388
box -48 -56 720 834
use sg13g2_nor3_1  _1164_
timestamp 1747537721
transform 1 0 23616 0 -1 17388
box -48 -56 528 834
use sg13g2_xor2_1  _1165_
timestamp 1747537721
transform -1 0 24576 0 1 17388
box -48 -56 816 834
use sg13g2_nor2_1  _1166_
timestamp 1747537721
transform -1 0 23904 0 -1 15876
box -48 -56 432 834
use sg13g2_o21ai_1  _1167_
timestamp 1747537721
transform 1 0 23424 0 1 15876
box -48 -56 538 834
use sg13g2_o21ai_1  _1168_
timestamp 1747537721
transform 1 0 23904 0 1 15876
box -48 -56 538 834
use sg13g2_xor2_1  _1169_
timestamp 1747537721
transform -1 0 19776 0 1 24948
box -48 -56 816 834
use sg13g2_a21oi_1  _1170_
timestamp 1747537721
transform -1 0 18144 0 -1 24948
box -48 -56 528 834
use sg13g2_xnor2_1  _1171_
timestamp 1747537721
transform -1 0 18624 0 1 24948
box -48 -56 816 834
use sg13g2_nor2_1  _1172_
timestamp 1747537721
transform 1 0 21792 0 1 11340
box -48 -56 432 834
use sg13g2_xnor2_1  _1173_
timestamp 1747537721
transform 1 0 17088 0 1 24948
box -48 -56 816 834
use sg13g2_inv_2  _1174_
timestamp 1747537721
transform 1 0 7104 0 1 5292
box -48 -56 432 834
use sg13g2_nor2b_1  _1175_
timestamp 1747537721
transform -1 0 24576 0 -1 12852
box -54 -56 528 834
use sg13g2_xor2_1  _1176_
timestamp 1747537721
transform -1 0 16896 0 1 24948
box -48 -56 816 834
use sg13g2_xor2_1  _1177_
timestamp 1747537721
transform -1 0 10560 0 1 21924
box -48 -56 816 834
use sg13g2_xnor2_1  _1178_
timestamp 1747537721
transform -1 0 11328 0 1 21924
box -48 -56 816 834
use sg13g2_and2_1  _1179_
timestamp 1747537721
transform 1 0 24384 0 1 9828
box -48 -56 528 834
use sg13g2_nand2_1  _1180_
timestamp 1747537721
transform 1 0 22080 0 -1 11340
box -48 -56 432 834
use sg13g2_mux4_1  _1181_
timestamp 1747537721
transform 1 0 8544 0 1 8316
box -48 -56 2064 834
use sg13g2_nand3_1  _1182_
timestamp 1747537721
transform 1 0 26016 0 -1 9828
box -48 -56 528 834
use sg13g2_inv_1  _1183_
timestamp 1747537721
transform 1 0 26880 0 1 8316
box -48 -56 336 834
use sg13g2_nand3b_1  _1184_
timestamp 1747537721
transform 1 0 21504 0 -1 8316
box -48 -56 720 834
use sg13g2_and3_2  _1185_
timestamp 1747537721
transform 1 0 22656 0 -1 18900
box -48 -56 720 834
use sg13g2_nor2_2  _1186_
timestamp 1747537721
transform -1 0 23712 0 1 6804
box -48 -56 624 834
use sg13g2_nor2b_1  _1187_
timestamp 1747537721
transform -1 0 23712 0 1 11340
box -54 -56 528 834
use sg13g2_xnor2_1  _1188_
timestamp 1747537721
transform 1 0 21888 0 1 21924
box -48 -56 816 834
use sg13g2_inv_1  _1189_
timestamp 1747537721
transform 1 0 22272 0 -1 6804
box -48 -56 336 834
use sg13g2_a21oi_1  _1190_
timestamp 1747537721
transform -1 0 19488 0 1 21924
box -48 -56 528 834
use sg13g2_xnor2_1  _1191_
timestamp 1747537721
transform 1 0 19584 0 -1 23436
box -48 -56 816 834
use sg13g2_xnor2_1  _1192_
timestamp 1747537721
transform -1 0 19584 0 -1 23436
box -48 -56 816 834
use sg13g2_a22oi_1  _1193_
timestamp 1747537721
transform 1 0 22176 0 1 11340
box -48 -56 624 834
use sg13g2_o21ai_1  _1194_
timestamp 1747537721
transform 1 0 22752 0 1 11340
box -48 -56 538 834
use sg13g2_o21ai_1  _1195_
timestamp 1747537721
transform -1 0 23424 0 -1 12852
box -48 -56 538 834
use sg13g2_nand3_1  _1196_
timestamp 1747537721
transform -1 0 23232 0 1 15876
box -48 -56 528 834
use sg13g2_o21ai_1  _1197_
timestamp 1747537721
transform 1 0 9696 0 1 18900
box -48 -56 538 834
use sg13g2_mux4_1  _1198_
timestamp 1747537721
transform -1 0 22272 0 1 15876
box -48 -56 2064 834
use sg13g2_nor2b_1  _1199_
timestamp 1747537721
transform -1 0 11712 0 1 12852
box -54 -56 528 834
use sg13g2_nand2_2  _1200_
timestamp 1747537721
transform 1 0 9984 0 1 11340
box -48 -56 624 834
use sg13g2_nor2_2  _1201_
timestamp 1747537721
transform -1 0 9696 0 1 12852
box -48 -56 624 834
use sg13g2_or2_2  _1202_
timestamp 1747537721
transform 1 0 11040 0 -1 14364
box -48 -56 624 834
use sg13g2_nor2_1  _1203_
timestamp 1747537721
transform 1 0 9600 0 1 14364
box -48 -56 432 834
use sg13g2_a221oi_1  _1204_
timestamp 1747537721
transform -1 0 9888 0 -1 15876
box -48 -56 816 834
use sg13g2_nor2b_2  _1205_
timestamp 1747537721
transform 1 0 13344 0 -1 20412
box -54 -56 720 834
use sg13g2_and2_1  _1206_
timestamp 1747537721
transform -1 0 14016 0 -1 18900
box -48 -56 528 834
use sg13g2_nand2_2  _1207_
timestamp 1747537721
transform 1 0 12288 0 -1 17388
box -48 -56 624 834
use sg13g2_nor2_1  _1208_
timestamp 1747537721
transform -1 0 26208 0 1 17388
box -48 -56 432 834
use sg13g2_mux2_2  _1209_
timestamp 1747537721
transform -1 0 21984 0 -1 17388
box -48 -56 1104 834
use sg13g2_and2_2  _1210_
timestamp 1747537721
transform -1 0 16992 0 -1 17388
box -48 -56 624 834
use sg13g2_nand2_2  _1211_
timestamp 1747537721
transform 1 0 17184 0 -1 17388
box -48 -56 624 834
use sg13g2_nand2_1  _1212_
timestamp 1747537721
transform -1 0 9984 0 1 17388
box -48 -56 432 834
use sg13g2_nor2_1  _1213_
timestamp 1747537721
transform 1 0 20544 0 -1 17388
box -48 -56 432 834
use sg13g2_nand2b_2  _1214_
timestamp 1747537721
transform -1 0 16416 0 -1 17388
box -48 -56 816 834
use sg13g2_o21ai_1  _1215_
timestamp 1747537721
transform -1 0 9600 0 1 17388
box -48 -56 538 834
use sg13g2_inv_1  _1216_
timestamp 1747537721
transform -1 0 9120 0 1 17388
box -48 -56 336 834
use sg13g2_nor2b_2  _1217_
timestamp 1747537721
transform 1 0 12672 0 -1 20412
box -54 -56 720 834
use sg13g2_and2_1  _1218_
timestamp 1747537721
transform -1 0 14016 0 1 18900
box -48 -56 528 834
use sg13g2_nand2_2  _1219_
timestamp 1747537721
transform -1 0 14112 0 -1 17388
box -48 -56 624 834
use sg13g2_xnor2_1  _1220_
timestamp 1747537721
transform -1 0 10176 0 -1 21924
box -48 -56 816 834
use sg13g2_nand2b_2  _1221_
timestamp 1747537721
transform -1 0 9600 0 1 15876
box -48 -56 816 834
use sg13g2_and2_2  _1222_
timestamp 1747537721
transform 1 0 15264 0 1 18900
box -48 -56 624 834
use sg13g2_nand2_2  _1223_
timestamp 1747537721
transform -1 0 15264 0 1 18900
box -48 -56 624 834
use sg13g2_a21oi_1  _1224_
timestamp 1747537721
transform -1 0 10080 0 1 15876
box -48 -56 528 834
use sg13g2_a221oi_1  _1225_
timestamp 1747537721
transform 1 0 8832 0 -1 17388
box -48 -56 816 834
use sg13g2_a21oi_1  _1226_
timestamp 1747537721
transform 1 0 8736 0 -1 18900
box -48 -56 528 834
use sg13g2_o21ai_1  _1227_
timestamp 1747537721
transform -1 0 9120 0 1 18900
box -48 -56 538 834
use sg13g2_a21oi_2  _1228_
timestamp 1747537721
transform -1 0 9312 0 -1 20412
box -48 -56 816 834
use sg13g2_o21ai_1  _1229_
timestamp 1747537721
transform 1 0 5280 0 1 20412
box -48 -56 538 834
use sg13g2_nor2_2  _1230_
timestamp 1747537721
transform -1 0 6528 0 1 18900
box -48 -56 624 834
use sg13g2_o21ai_1  _1231_
timestamp 1747537721
transform -1 0 6816 0 -1 18900
box -48 -56 538 834
use sg13g2_nand2_1  _1232_
timestamp 1747537721
transform 1 0 2016 0 1 8316
box -48 -56 432 834
use sg13g2_nor2_1  _1233_
timestamp 1747537721
transform 1 0 2304 0 -1 8316
box -48 -56 432 834
use sg13g2_xor2_1  _1234_
timestamp 1747537721
transform 1 0 2784 0 -1 12852
box -48 -56 816 834
use sg13g2_xnor2_1  _1235_
timestamp 1747537721
transform 1 0 3360 0 1 12852
box -48 -56 816 834
use sg13g2_nand2_1  _1236_
timestamp 1747537721
transform 1 0 4704 0 1 14364
box -48 -56 432 834
use sg13g2_nand2_1  _1237_
timestamp 1747537721
transform 1 0 3456 0 -1 14364
box -48 -56 432 834
use sg13g2_xnor2_1  _1238_
timestamp 1747537721
transform 1 0 3456 0 1 14364
box -48 -56 816 834
use sg13g2_xnor2_1  _1239_
timestamp 1747537721
transform 1 0 3936 0 -1 15876
box -48 -56 816 834
use sg13g2_xnor2_1  _1240_
timestamp 1747537721
transform -1 0 4992 0 1 11340
box -48 -56 816 834
use sg13g2_xnor2_1  _1241_
timestamp 1747537721
transform -1 0 9984 0 1 11340
box -48 -56 816 834
use sg13g2_and2_1  _1242_
timestamp 1747537721
transform -1 0 15360 0 1 17388
box -48 -56 528 834
use sg13g2_nand2_1  _1243_
timestamp 1747537721
transform -1 0 15744 0 1 17388
box -48 -56 432 834
use sg13g2_a21oi_1  _1244_
timestamp 1747537721
transform 1 0 4608 0 -1 12852
box -48 -56 528 834
use sg13g2_o21ai_1  _1245_
timestamp 1747537721
transform -1 0 4608 0 -1 12852
box -48 -56 538 834
use sg13g2_nor2b_2  _1246_
timestamp 1747537721
transform -1 0 13536 0 -1 17388
box -54 -56 720 834
use sg13g2_nand2b_2  _1247_
timestamp 1747537721
transform -1 0 13536 0 1 17388
box -48 -56 816 834
use sg13g2_a21o_1  _1248_
timestamp 1747537721
transform 1 0 9984 0 -1 11340
box -48 -56 720 834
use sg13g2_nor2_1  _1249_
timestamp 1747537721
transform 1 0 7296 0 -1 12852
box -48 -56 432 834
use sg13g2_mux2_1  _1250_
timestamp 1747537721
transform -1 0 21696 0 -1 12852
box -48 -56 1008 834
use sg13g2_mux2_1  _1251_
timestamp 1747537721
transform 1 0 19200 0 1 14364
box -48 -56 1008 834
use sg13g2_mux2_2  _1252_
timestamp 1747537721
transform -1 0 20544 0 1 12852
box -48 -56 1104 834
use sg13g2_a221oi_1  _1253_
timestamp 1747537721
transform -1 0 8064 0 1 12852
box -48 -56 816 834
use sg13g2_inv_1  _1254_
timestamp 1747537721
transform 1 0 5376 0 -1 15876
box -48 -56 336 834
use sg13g2_a22oi_1  _1255_
timestamp 1747537721
transform 1 0 5664 0 -1 15876
box -48 -56 624 834
use sg13g2_o21ai_1  _1256_
timestamp 1747537721
transform -1 0 6720 0 -1 15876
box -48 -56 538 834
use sg13g2_nor2_2  _1257_
timestamp 1747537721
transform -1 0 10464 0 -1 15876
box -48 -56 624 834
use sg13g2_nand2_2  _1258_
timestamp 1747537721
transform 1 0 15072 0 1 15876
box -48 -56 624 834
use sg13g2_a221oi_1  _1259_
timestamp 1747537721
transform -1 0 6432 0 1 15876
box -48 -56 816 834
use sg13g2_nor2_1  _1260_
timestamp 1747537721
transform -1 0 6048 0 1 17388
box -48 -56 432 834
use sg13g2_o21ai_1  _1261_
timestamp 1747537721
transform 1 0 4896 0 -1 18900
box -48 -56 538 834
use sg13g2_a21oi_2  _1262_
timestamp 1747537721
transform 1 0 4896 0 -1 20412
box -48 -56 816 834
use sg13g2_o21ai_1  _1263_
timestamp 1747537721
transform -1 0 4128 0 -1 20412
box -48 -56 538 834
use sg13g2_nor2_2  _1264_
timestamp 1747537721
transform 1 0 4128 0 -1 20412
box -48 -56 624 834
use sg13g2_o21ai_1  _1265_
timestamp 1747537721
transform -1 0 5184 0 1 17388
box -48 -56 538 834
use sg13g2_mux4_1  _1266_
timestamp 1747537721
transform -1 0 21408 0 -1 11340
box -48 -56 2064 834
use sg13g2_inv_1  _1267_
timestamp 1747537721
transform -1 0 7200 0 -1 11340
box -48 -56 336 834
use sg13g2_nor2_1  _1268_
timestamp 1747537721
transform 1 0 6336 0 1 11340
box -48 -56 432 834
use sg13g2_a221oi_1  _1269_
timestamp 1747537721
transform -1 0 6336 0 1 11340
box -48 -56 816 834
use sg13g2_and2_1  _1270_
timestamp 1747537721
transform -1 0 4320 0 -1 11340
box -48 -56 528 834
use sg13g2_o21ai_1  _1271_
timestamp 1747537721
transform -1 0 4704 0 1 14364
box -48 -56 538 834
use sg13g2_and2_1  _1272_
timestamp 1747537721
transform 1 0 4128 0 -1 8316
box -48 -56 528 834
use sg13g2_xor2_1  _1273_
timestamp 1747537721
transform 1 0 4608 0 -1 8316
box -48 -56 816 834
use sg13g2_xnor2_1  _1274_
timestamp 1747537721
transform -1 0 5472 0 1 8316
box -48 -56 816 834
use sg13g2_o21ai_1  _1275_
timestamp 1747537721
transform 1 0 2400 0 1 8316
box -48 -56 538 834
use sg13g2_nor2b_1  _1276_
timestamp 1747537721
transform 1 0 2880 0 1 8316
box -54 -56 528 834
use sg13g2_xnor2_1  _1277_
timestamp 1747537721
transform 1 0 3360 0 1 8316
box -48 -56 816 834
use sg13g2_xor2_1  _1278_
timestamp 1747537721
transform 1 0 3456 0 1 9828
box -48 -56 816 834
use sg13g2_xnor2_1  _1279_
timestamp 1747537721
transform 1 0 5184 0 1 9828
box -48 -56 816 834
use sg13g2_o21ai_1  _1280_
timestamp 1747537721
transform -1 0 7104 0 1 9828
box -48 -56 538 834
use sg13g2_nand2_1  _1281_
timestamp 1747537721
transform 1 0 864 0 -1 8316
box -48 -56 432 834
use sg13g2_nand2_1  _1282_
timestamp 1747537721
transform -1 0 2592 0 1 6804
box -48 -56 432 834
use sg13g2_xnor2_1  _1283_
timestamp 1747537721
transform 1 0 960 0 1 6804
box -48 -56 816 834
use sg13g2_xnor2_1  _1284_
timestamp 1747537721
transform 1 0 1248 0 -1 8316
box -48 -56 816 834
use sg13g2_nand2_1  _1285_
timestamp 1747537721
transform -1 0 3168 0 1 5292
box -48 -56 432 834
use sg13g2_xnor2_1  _1286_
timestamp 1747537721
transform 1 0 1248 0 -1 6804
box -48 -56 816 834
use sg13g2_nand2_1  _1287_
timestamp 1747537721
transform -1 0 3264 0 -1 6804
box -48 -56 432 834
use sg13g2_xor2_1  _1288_
timestamp 1747537721
transform 1 0 2112 0 -1 6804
box -48 -56 816 834
use sg13g2_a21oi_1  _1289_
timestamp 1747537721
transform -1 0 3264 0 1 6804
box -48 -56 528 834
use sg13g2_o21ai_1  _1290_
timestamp 1747537721
transform 1 0 2880 0 -1 8316
box -48 -56 538 834
use sg13g2_a221oi_1  _1291_
timestamp 1747537721
transform -1 0 4992 0 1 9828
box -48 -56 816 834
use sg13g2_o21ai_1  _1292_
timestamp 1747537721
transform 1 0 5088 0 1 11340
box -48 -56 538 834
use sg13g2_o21ai_1  _1293_
timestamp 1747537721
transform -1 0 5568 0 -1 11340
box -48 -56 538 834
use sg13g2_a21oi_1  _1294_
timestamp 1747537721
transform -1 0 4416 0 1 15876
box -48 -56 528 834
use sg13g2_o21ai_1  _1295_
timestamp 1747537721
transform 1 0 4512 0 -1 17388
box -48 -56 538 834
use sg13g2_a21oi_2  _1296_
timestamp 1747537721
transform -1 0 4512 0 -1 17388
box -48 -56 816 834
use sg13g2_o21ai_1  _1297_
timestamp 1747537721
transform -1 0 10752 0 1 20412
box -48 -56 538 834
use sg13g2_nor2_1  _1298_
timestamp 1747537721
transform -1 0 10752 0 -1 20412
box -48 -56 432 834
use sg13g2_nand2_1  _1299_
timestamp 1747537721
transform 1 0 10656 0 1 17388
box -48 -56 432 834
use sg13g2_o21ai_1  _1300_
timestamp 1747537721
transform -1 0 11808 0 1 18900
box -48 -56 538 834
use sg13g2_nand2_1  _1301_
timestamp 1747537721
transform 1 0 21792 0 -1 12852
box -48 -56 432 834
use sg13g2_o21ai_1  _1302_
timestamp 1747537721
transform -1 0 22848 0 1 12852
box -48 -56 538 834
use sg13g2_mux2_2  _1303_
timestamp 1747537721
transform -1 0 21600 0 1 12852
box -48 -56 1104 834
use sg13g2_a22oi_1  _1304_
timestamp 1747537721
transform -1 0 11136 0 1 12852
box -48 -56 624 834
use sg13g2_o21ai_1  _1305_
timestamp 1747537721
transform -1 0 10560 0 1 12852
box -48 -56 538 834
use sg13g2_a21oi_1  _1306_
timestamp 1747537721
transform -1 0 4608 0 1 8316
box -48 -56 528 834
use sg13g2_xor2_1  _1307_
timestamp 1747537721
transform 1 0 9600 0 -1 6804
box -48 -56 816 834
use sg13g2_nand2b_1  _1308_
timestamp 1747537721
transform 1 0 10464 0 -1 6804
box -48 -56 528 834
use sg13g2_xnor2_1  _1309_
timestamp 1747537721
transform -1 0 10560 0 1 6804
box -48 -56 816 834
use sg13g2_a21o_1  _1310_
timestamp 1747537721
transform -1 0 6048 0 -1 8316
box -48 -56 720 834
use sg13g2_nand2_1  _1311_
timestamp 1747537721
transform 1 0 7584 0 -1 8316
box -48 -56 432 834
use sg13g2_nor2_1  _1312_
timestamp 1747537721
transform 1 0 6624 0 1 6804
box -48 -56 432 834
use sg13g2_xnor2_1  _1313_
timestamp 1747537721
transform 1 0 6336 0 -1 8316
box -48 -56 816 834
use sg13g2_xnor2_1  _1314_
timestamp 1747537721
transform 1 0 6624 0 1 8316
box -48 -56 816 834
use sg13g2_xnor2_1  _1315_
timestamp 1747537721
transform 1 0 7776 0 1 8316
box -48 -56 816 834
use sg13g2_o21ai_1  _1316_
timestamp 1747537721
transform -1 0 8256 0 -1 9828
box -48 -56 538 834
use sg13g2_o21ai_1  _1317_
timestamp 1747537721
transform 1 0 2304 0 1 5292
box -48 -56 538 834
use sg13g2_xnor2_1  _1318_
timestamp 1747537721
transform -1 0 9312 0 1 5292
box -48 -56 816 834
use sg13g2_xor2_1  _1319_
timestamp 1747537721
transform 1 0 7776 0 1 5292
box -48 -56 816 834
use sg13g2_nor2_1  _1320_
timestamp 1747537721
transform -1 0 9504 0 -1 6804
box -48 -56 432 834
use sg13g2_xor2_1  _1321_
timestamp 1747537721
transform 1 0 6912 0 -1 6804
box -48 -56 816 834
use sg13g2_o21ai_1  _1322_
timestamp 1747537721
transform 1 0 1728 0 1 6804
box -48 -56 538 834
use sg13g2_xnor2_1  _1323_
timestamp 1747537721
transform 1 0 7584 0 1 6804
box -48 -56 816 834
use sg13g2_a21oi_1  _1324_
timestamp 1747537721
transform 1 0 7872 0 -1 6804
box -48 -56 528 834
use sg13g2_o21ai_1  _1325_
timestamp 1747537721
transform 1 0 8352 0 1 6804
box -48 -56 538 834
use sg13g2_a21oi_1  _1326_
timestamp 1747537721
transform 1 0 8256 0 -1 9828
box -48 -56 528 834
use sg13g2_o21ai_1  _1327_
timestamp 1747537721
transform 1 0 7488 0 1 9828
box -48 -56 538 834
use sg13g2_o21ai_1  _1328_
timestamp 1747537721
transform -1 0 10368 0 -1 14364
box -48 -56 538 834
use sg13g2_a22oi_1  _1329_
timestamp 1747537721
transform -1 0 10656 0 1 14364
box -48 -56 624 834
use sg13g2_nor2_1  _1330_
timestamp 1747537721
transform -1 0 10656 0 1 17388
box -48 -56 432 834
use sg13g2_nor2_1  _1331_
timestamp 1747537721
transform -1 0 12576 0 1 18900
box -48 -56 432 834
use sg13g2_o21ai_1  _1332_
timestamp 1747537721
transform 1 0 10368 0 1 18900
box -48 -56 538 834
use sg13g2_a21oi_2  _1333_
timestamp 1747537721
transform -1 0 12288 0 1 20412
box -48 -56 816 834
use sg13g2_o21ai_1  _1334_
timestamp 1747537721
transform -1 0 2112 0 -1 20412
box -48 -56 538 834
use sg13g2_nor2_1  _1335_
timestamp 1747537721
transform 1 0 3360 0 1 18900
box -48 -56 432 834
use sg13g2_o21ai_1  _1336_
timestamp 1747537721
transform -1 0 2496 0 -1 18900
box -48 -56 538 834
use sg13g2_mux4_1  _1337_
timestamp 1747537721
transform -1 0 21120 0 1 11340
box -48 -56 2064 834
use sg13g2_a22oi_1  _1338_
timestamp 1747537721
transform 1 0 13440 0 1 12852
box -48 -56 624 834
use sg13g2_o21ai_1  _1339_
timestamp 1747537721
transform 1 0 12672 0 -1 12852
box -48 -56 538 834
use sg13g2_o21ai_1  _1340_
timestamp 1747537721
transform 1 0 7104 0 -1 8316
box -48 -56 538 834
use sg13g2_nand2_1  _1341_
timestamp 1747537721
transform 1 0 13152 0 1 6804
box -48 -56 432 834
use sg13g2_nor2_1  _1342_
timestamp 1747537721
transform 1 0 13920 0 -1 6804
box -48 -56 432 834
use sg13g2_xor2_1  _1343_
timestamp 1747537721
transform -1 0 13152 0 -1 6804
box -48 -56 816 834
use sg13g2_xnor2_1  _1344_
timestamp 1747537721
transform 1 0 11616 0 -1 6804
box -48 -56 816 834
use sg13g2_o21ai_1  _1345_
timestamp 1747537721
transform 1 0 10944 0 1 6804
box -48 -56 538 834
use sg13g2_and2_1  _1346_
timestamp 1747537721
transform -1 0 12384 0 1 6804
box -48 -56 528 834
use sg13g2_or2_1  _1347_
timestamp 1747537721
transform 1 0 12384 0 1 6804
box -48 -56 528 834
use sg13g2_nand2b_1  _1348_
timestamp 1747537721
transform 1 0 12960 0 -1 8316
box -48 -56 528 834
use sg13g2_xnor2_1  _1349_
timestamp 1747537721
transform -1 0 12960 0 -1 8316
box -48 -56 816 834
use sg13g2_xnor2_1  _1350_
timestamp 1747537721
transform 1 0 10656 0 1 8316
box -48 -56 816 834
use sg13g2_inv_1  _1351_
timestamp 1747537721
transform -1 0 12192 0 -1 9828
box -48 -56 336 834
use sg13g2_a21oi_1  _1352_
timestamp 1747537721
transform 1 0 10944 0 -1 9828
box -48 -56 528 834
use sg13g2_a22oi_1  _1353_
timestamp 1747537721
transform -1 0 9888 0 1 5292
box -48 -56 624 834
use sg13g2_nand2b_1  _1354_
timestamp 1747537721
transform -1 0 11712 0 1 3780
box -48 -56 528 834
use sg13g2_nor2b_1  _1355_
timestamp 1747537721
transform 1 0 10272 0 1 3780
box -54 -56 528 834
use sg13g2_xnor2_1  _1356_
timestamp 1747537721
transform 1 0 9120 0 -1 5292
box -48 -56 816 834
use sg13g2_xnor2_1  _1357_
timestamp 1747537721
transform 1 0 9888 0 -1 5292
box -48 -56 816 834
use sg13g2_nand2_1  _1358_
timestamp 1747537721
transform -1 0 9312 0 -1 2268
box -48 -56 432 834
use sg13g2_xnor2_1  _1359_
timestamp 1747537721
transform 1 0 8160 0 1 2268
box -48 -56 816 834
use sg13g2_a21oi_2  _1360_
timestamp 1747537721
transform 1 0 8832 0 1 6804
box -48 -56 816 834
use sg13g2_xnor2_1  _1361_
timestamp 1747537721
transform 1 0 8928 0 1 2268
box -48 -56 816 834
use sg13g2_o21ai_1  _1362_
timestamp 1747537721
transform 1 0 10656 0 -1 5292
box -48 -56 538 834
use sg13g2_a21oi_1  _1363_
timestamp 1747537721
transform -1 0 11616 0 1 5292
box -48 -56 528 834
use sg13g2_o21ai_1  _1364_
timestamp 1747537721
transform 1 0 11424 0 1 8316
box -48 -56 538 834
use sg13g2_a21o_1  _1365_
timestamp 1747537721
transform -1 0 12768 0 1 8316
box -48 -56 720 834
use sg13g2_o21ai_1  _1366_
timestamp 1747537721
transform -1 0 13152 0 -1 15876
box -48 -56 538 834
use sg13g2_a22oi_1  _1367_
timestamp 1747537721
transform 1 0 12096 0 -1 15876
box -48 -56 624 834
use sg13g2_nor2_1  _1368_
timestamp 1747537721
transform 1 0 6912 0 1 17388
box -48 -56 432 834
use sg13g2_nor2_1  _1369_
timestamp 1747537721
transform 1 0 2688 0 -1 17388
box -48 -56 432 834
use sg13g2_o21ai_1  _1370_
timestamp 1747537721
transform 1 0 1056 0 -1 18900
box -48 -56 538 834
use sg13g2_a21oi_2  _1371_
timestamp 1747537721
transform 1 0 1056 0 1 18900
box -48 -56 816 834
use sg13g2_o21ai_1  _1372_
timestamp 1747537721
transform -1 0 3360 0 1 18900
box -48 -56 538 834
use sg13g2_nor2_1  _1373_
timestamp 1747537721
transform -1 0 2688 0 -1 17388
box -48 -56 432 834
use sg13g2_o21ai_1  _1374_
timestamp 1747537721
transform -1 0 2496 0 1 15876
box -48 -56 538 834
use sg13g2_nand2_1  _1375_
timestamp 1747537721
transform 1 0 14304 0 -1 12852
box -48 -56 432 834
use sg13g2_mux2_1  _1376_
timestamp 1747537721
transform -1 0 22080 0 -1 14364
box -48 -56 1008 834
use sg13g2_mux2_2  _1377_
timestamp 1747537721
transform -1 0 20736 0 -1 14364
box -48 -56 1104 834
use sg13g2_a22oi_1  _1378_
timestamp 1747537721
transform -1 0 15264 0 1 12852
box -48 -56 624 834
use sg13g2_a21oi_1  _1379_
timestamp 1747537721
transform -1 0 15552 0 -1 14364
box -48 -56 528 834
use sg13g2_nand3_1  _1380_
timestamp 1747537721
transform -1 0 14592 0 -1 14364
box -48 -56 528 834
use sg13g2_a21oi_1  _1381_
timestamp 1747537721
transform -1 0 12192 0 -1 8316
box -48 -56 528 834
use sg13g2_and2_1  _1382_
timestamp 1747537721
transform 1 0 20352 0 -1 5292
box -48 -56 528 834
use sg13g2_xor2_1  _1383_
timestamp 1747537721
transform 1 0 19584 0 -1 5292
box -48 -56 816 834
use sg13g2_xor2_1  _1384_
timestamp 1747537721
transform -1 0 20544 0 1 5292
box -48 -56 816 834
use sg13g2_o21ai_1  _1385_
timestamp 1747537721
transform -1 0 13920 0 -1 6804
box -48 -56 538 834
use sg13g2_nand2_1  _1386_
timestamp 1747537721
transform 1 0 14592 0 -1 8316
box -48 -56 432 834
use sg13g2_xnor2_1  _1387_
timestamp 1747537721
transform -1 0 15744 0 1 6804
box -48 -56 816 834
use sg13g2_xnor2_1  _1388_
timestamp 1747537721
transform 1 0 14208 0 1 6804
box -48 -56 816 834
use sg13g2_xor2_1  _1389_
timestamp 1747537721
transform 1 0 12768 0 -1 9828
box -48 -56 816 834
use sg13g2_a21o_1  _1390_
timestamp 1747537721
transform -1 0 14208 0 -1 9828
box -48 -56 720 834
use sg13g2_o21ai_1  _1391_
timestamp 1747537721
transform 1 0 10752 0 1 3780
box -48 -56 538 834
use sg13g2_xor2_1  _1392_
timestamp 1747537721
transform 1 0 14016 0 1 3780
box -48 -56 816 834
use sg13g2_xnor2_1  _1393_
timestamp 1747537721
transform -1 0 14976 0 -1 3780
box -48 -56 816 834
use sg13g2_and2_1  _1394_
timestamp 1747537721
transform 1 0 13632 0 -1 2268
box -48 -56 528 834
use sg13g2_xor2_1  _1395_
timestamp 1747537721
transform 1 0 11712 0 -1 2268
box -48 -56 816 834
use sg13g2_o21ai_1  _1396_
timestamp 1747537721
transform 1 0 9696 0 1 2268
box -48 -56 538 834
use sg13g2_xor2_1  _1397_
timestamp 1747537721
transform -1 0 14880 0 -1 2268
box -48 -56 816 834
use sg13g2_a21oi_1  _1398_
timestamp 1747537721
transform 1 0 13728 0 -1 3780
box -48 -56 528 834
use sg13g2_o21ai_1  _1399_
timestamp 1747537721
transform 1 0 14592 0 1 2268
box -48 -56 538 834
use sg13g2_a21oi_1  _1400_
timestamp 1747537721
transform 1 0 14400 0 1 8316
box -48 -56 528 834
use sg13g2_o21ai_1  _1401_
timestamp 1747537721
transform -1 0 15936 0 1 8316
box -48 -56 538 834
use sg13g2_a21oi_1  _1402_
timestamp 1747537721
transform 1 0 14592 0 -1 14364
box -48 -56 528 834
use sg13g2_o21ai_1  _1403_
timestamp 1747537721
transform -1 0 14976 0 1 14364
box -48 -56 538 834
use sg13g2_nor2b_1  _1404_
timestamp 1747537721
transform -1 0 2208 0 -1 15876
box -54 -56 528 834
use sg13g2_o21ai_1  _1405_
timestamp 1747537721
transform 1 0 1056 0 1 15876
box -48 -56 538 834
use sg13g2_a21oi_2  _1406_
timestamp 1747537721
transform 1 0 1056 0 -1 17388
box -48 -56 816 834
use sg13g2_o21ai_1  _1407_
timestamp 1747537721
transform 1 0 15936 0 1 20412
box -48 -56 538 834
use sg13g2_nor2_1  _1408_
timestamp 1747537721
transform 1 0 15936 0 1 18900
box -48 -56 432 834
use sg13g2_o21ai_1  _1409_
timestamp 1747537721
transform -1 0 17568 0 1 18900
box -48 -56 538 834
use sg13g2_o21ai_1  _1410_
timestamp 1747537721
transform 1 0 14688 0 -1 6804
box -48 -56 538 834
use sg13g2_and2_1  _1411_
timestamp 1747537721
transform 1 0 21504 0 -1 5292
box -48 -56 528 834
use sg13g2_xor2_1  _1412_
timestamp 1747537721
transform -1 0 22848 0 -1 3780
box -48 -56 816 834
use sg13g2_xor2_1  _1413_
timestamp 1747537721
transform -1 0 22176 0 -1 6804
box -48 -56 816 834
use sg13g2_a21oi_1  _1414_
timestamp 1747537721
transform -1 0 21024 0 1 5292
box -48 -56 528 834
use sg13g2_nor2_1  _1415_
timestamp 1747537721
transform 1 0 19200 0 1 6804
box -48 -56 432 834
use sg13g2_xor2_1  _1416_
timestamp 1747537721
transform -1 0 20352 0 1 6804
box -48 -56 816 834
use sg13g2_nor2_1  _1417_
timestamp 1747537721
transform -1 0 17568 0 -1 8316
box -48 -56 432 834
use sg13g2_nand2_1  _1418_
timestamp 1747537721
transform -1 0 17184 0 -1 8316
box -48 -56 432 834
use sg13g2_nor2_1  _1419_
timestamp 1747537721
transform 1 0 16416 0 -1 8316
box -48 -56 432 834
use sg13g2_xnor2_1  _1420_
timestamp 1747537721
transform -1 0 21696 0 1 9828
box -48 -56 816 834
use sg13g2_o21ai_1  _1421_
timestamp 1747537721
transform -1 0 17376 0 1 9828
box -48 -56 538 834
use sg13g2_a22oi_1  _1422_
timestamp 1747537721
transform -1 0 15552 0 -1 3780
box -48 -56 624 834
use sg13g2_xor2_1  _1423_
timestamp 1747537721
transform 1 0 16032 0 -1 3780
box -48 -56 816 834
use sg13g2_nand2b_1  _1424_
timestamp 1747537721
transform 1 0 16320 0 1 2268
box -48 -56 528 834
use sg13g2_xor2_1  _1425_
timestamp 1747537721
transform 1 0 16800 0 -1 3780
box -48 -56 816 834
use sg13g2_xnor2_1  _1426_
timestamp 1747537721
transform -1 0 19104 0 1 2268
box -48 -56 816 834
use sg13g2_a21o_1  _1427_
timestamp 1747537721
transform -1 0 15552 0 -1 2268
box -48 -56 720 834
use sg13g2_nor2b_1  _1428_
timestamp 1747537721
transform 1 0 18240 0 -1 3780
box -54 -56 528 834
use sg13g2_xnor2_1  _1429_
timestamp 1747537721
transform -1 0 18240 0 1 2268
box -48 -56 816 834
use sg13g2_a21oi_1  _1430_
timestamp 1747537721
transform 1 0 16800 0 1 2268
box -48 -56 528 834
use sg13g2_o21ai_1  _1431_
timestamp 1747537721
transform -1 0 16320 0 1 2268
box -48 -56 538 834
use sg13g2_a221oi_1  _1432_
timestamp 1747537721
transform 1 0 16128 0 1 8316
box -48 -56 816 834
use sg13g2_nor2_1  _1433_
timestamp 1747537721
transform 1 0 16224 0 1 12852
box -48 -56 432 834
use sg13g2_mux4_1  _1434_
timestamp 1747537721
transform 1 0 20832 0 1 14364
box -48 -56 2064 834
use sg13g2_a221oi_1  _1435_
timestamp 1747537721
transform 1 0 16416 0 -1 14364
box -48 -56 816 834
use sg13g2_nor2_1  _1436_
timestamp 1747537721
transform -1 0 16800 0 1 17388
box -48 -56 432 834
use sg13g2_a21oi_1  _1437_
timestamp 1747537721
transform -1 0 16416 0 1 17388
box -48 -56 528 834
use sg13g2_or3_1  _1438_
timestamp 1747537721
transform 1 0 16128 0 -1 18900
box -48 -56 720 834
use sg13g2_a21oi_1  _1439_
timestamp 1747537721
transform -1 0 17280 0 -1 18900
box -48 -56 528 834
use sg13g2_a21oi_1  _1440_
timestamp 1747537721
transform 1 0 16608 0 1 18900
box -48 -56 528 834
use sg13g2_o21ai_1  _1441_
timestamp 1747537721
transform 1 0 17184 0 -1 20412
box -48 -56 538 834
use sg13g2_a21oi_2  _1442_
timestamp 1747537721
transform 1 0 17184 0 1 20412
box -48 -56 816 834
use sg13g2_o21ai_1  _1443_
timestamp 1747537721
transform 1 0 19680 0 -1 20412
box -48 -56 538 834
use sg13g2_nor2_1  _1444_
timestamp 1747537721
transform -1 0 19584 0 -1 20412
box -48 -56 432 834
use sg13g2_o21ai_1  _1445_
timestamp 1747537721
transform 1 0 19008 0 -1 18900
box -48 -56 538 834
use sg13g2_xnor2_1  _1446_
timestamp 1747537721
transform -1 0 27648 0 -1 12852
box -48 -56 816 834
use sg13g2_a21oi_2  _1447_
timestamp 1747537721
transform -1 0 19008 0 -1 11340
box -48 -56 816 834
use sg13g2_o21ai_1  _1448_
timestamp 1747537721
transform 1 0 17472 0 1 3780
box -48 -56 538 834
use sg13g2_xor2_1  _1449_
timestamp 1747537721
transform -1 0 23520 0 -1 5292
box -48 -56 816 834
use sg13g2_a21oi_1  _1450_
timestamp 1747537721
transform 1 0 21120 0 1 2268
box -48 -56 528 834
use sg13g2_xor2_1  _1451_
timestamp 1747537721
transform -1 0 22080 0 -1 3780
box -48 -56 816 834
use sg13g2_xnor2_1  _1452_
timestamp 1747537721
transform 1 0 20736 0 1 3780
box -48 -56 816 834
use sg13g2_xnor2_1  _1453_
timestamp 1747537721
transform -1 0 22272 0 1 3780
box -48 -56 816 834
use sg13g2_xnor2_1  _1454_
timestamp 1747537721
transform -1 0 20160 0 1 3780
box -48 -56 816 834
use sg13g2_a21oi_1  _1455_
timestamp 1747537721
transform 1 0 19200 0 -1 8316
box -48 -56 528 834
use sg13g2_a21oi_1  _1456_
timestamp 1747537721
transform 1 0 20352 0 1 6804
box -48 -56 528 834
use sg13g2_a21o_1  _1457_
timestamp 1747537721
transform 1 0 21984 0 1 5292
box -48 -56 720 834
use sg13g2_xnor2_1  _1458_
timestamp 1747537721
transform -1 0 21984 0 1 5292
box -48 -56 816 834
use sg13g2_xnor2_1  _1459_
timestamp 1747537721
transform -1 0 22656 0 1 6804
box -48 -56 816 834
use sg13g2_xnor2_1  _1460_
timestamp 1747537721
transform -1 0 21888 0 1 6804
box -48 -56 816 834
use sg13g2_xnor2_1  _1461_
timestamp 1747537721
transform -1 0 20448 0 -1 8316
box -48 -56 816 834
use sg13g2_mux2_1  _1462_
timestamp 1747537721
transform 1 0 19008 0 1 8316
box -48 -56 1008 834
use sg13g2_nor2_1  _1463_
timestamp 1747537721
transform -1 0 16992 0 1 12852
box -48 -56 432 834
use sg13g2_nor2b_1  _1464_
timestamp 1747537721
transform -1 0 22368 0 1 12852
box -54 -56 528 834
use sg13g2_nor2_1  _1465_
timestamp 1747537721
transform 1 0 20736 0 -1 14364
box -48 -56 432 834
use sg13g2_a21oi_2  _1466_
timestamp 1747537721
transform -1 0 22848 0 -1 14364
box -48 -56 816 834
use sg13g2_a221oi_1  _1467_
timestamp 1747537721
transform 1 0 16992 0 1 12852
box -48 -56 816 834
use sg13g2_nor2_1  _1468_
timestamp 1747537721
transform 1 0 17472 0 1 17388
box -48 -56 432 834
use sg13g2_a221oi_1  _1469_
timestamp 1747537721
transform -1 0 19296 0 -1 17388
box -48 -56 816 834
use sg13g2_o21ai_1  _1470_
timestamp 1747537721
transform 1 0 20064 0 -1 17388
box -48 -56 538 834
use sg13g2_a21oi_1  _1471_
timestamp 1747537721
transform -1 0 18240 0 -1 18900
box -48 -56 528 834
use sg13g2_a21oi_1  _1472_
timestamp 1747537721
transform -1 0 19872 0 1 17388
box -48 -56 528 834
use sg13g2_o21ai_1  _1473_
timestamp 1747537721
transform 1 0 19776 0 1 18900
box -48 -56 538 834
use sg13g2_a21oi_2  _1474_
timestamp 1747537721
transform 1 0 20832 0 -1 18900
box -48 -56 816 834
use sg13g2_nor2_1  _1475_
timestamp 1747537721
transform -1 0 11904 0 -1 11340
box -48 -56 432 834
use sg13g2_nand2b_2  _1476_
timestamp 1747537721
transform -1 0 9600 0 1 14364
box -48 -56 816 834
use sg13g2_nor2_1  _1477_
timestamp 1747537721
transform -1 0 8448 0 1 14364
box -48 -56 432 834
use sg13g2_a221oi_1  _1478_
timestamp 1747537721
transform -1 0 8064 0 1 14364
box -48 -56 816 834
use sg13g2_nand2b_1  _1479_
timestamp 1747537721
transform 1 0 8064 0 -1 15876
box -48 -56 528 834
use sg13g2_nor2_1  _1480_
timestamp 1747537721
transform -1 0 9120 0 -1 15876
box -48 -56 432 834
use sg13g2_nand2_2  _1481_
timestamp 1747537721
transform -1 0 15360 0 1 9828
box -48 -56 624 834
use sg13g2_nor2_1  _1482_
timestamp 1747537721
transform 1 0 6432 0 1 14364
box -48 -56 432 834
use sg13g2_or2_1  _1483_
timestamp 1747537721
transform 1 0 6816 0 1 14364
box -48 -56 528 834
use sg13g2_a22oi_1  _1484_
timestamp 1747537721
transform 1 0 7296 0 -1 15876
box -48 -56 624 834
use sg13g2_o21ai_1  _1485_
timestamp 1747537721
transform 1 0 6816 0 1 15876
box -48 -56 538 834
use sg13g2_a221oi_1  _1486_
timestamp 1747537721
transform 1 0 7296 0 1 15876
box -48 -56 816 834
use sg13g2_nor2_1  _1487_
timestamp 1747537721
transform 1 0 7104 0 -1 18900
box -48 -56 432 834
use sg13g2_o21ai_1  _1488_
timestamp 1747537721
transform 1 0 6624 0 1 18900
box -48 -56 538 834
use sg13g2_a21oi_2  _1489_
timestamp 1747537721
transform 1 0 7488 0 -1 20412
box -48 -56 816 834
use sg13g2_a22oi_1  _1490_
timestamp 1747537721
transform -1 0 8640 0 -1 12852
box -48 -56 624 834
use sg13g2_o21ai_1  _1491_
timestamp 1747537721
transform 1 0 8064 0 1 12852
box -48 -56 538 834
use sg13g2_nor2_1  _1492_
timestamp 1747537721
transform 1 0 6336 0 -1 11340
box -48 -56 432 834
use sg13g2_and2_1  _1493_
timestamp 1747537721
transform 1 0 1536 0 -1 9828
box -48 -56 528 834
use sg13g2_xnor2_1  _1494_
timestamp 1747537721
transform 1 0 1056 0 1 9828
box -48 -56 816 834
use sg13g2_xnor2_1  _1495_
timestamp 1747537721
transform 1 0 1824 0 1 9828
box -48 -56 816 834
use sg13g2_nand2_1  _1496_
timestamp 1747537721
transform -1 0 1920 0 -1 5292
box -48 -56 432 834
use sg13g2_nand2_1  _1497_
timestamp 1747537721
transform -1 0 2496 0 1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _1498_
timestamp 1747537721
transform 1 0 672 0 1 3780
box -48 -56 432 834
use sg13g2_xor2_1  _1499_
timestamp 1747537721
transform 1 0 576 0 1 5292
box -48 -56 816 834
use sg13g2_xnor2_1  _1500_
timestamp 1747537721
transform 1 0 1344 0 1 5292
box -48 -56 816 834
use sg13g2_a21oi_1  _1501_
timestamp 1747537721
transform -1 0 3168 0 -1 9828
box -48 -56 528 834
use sg13g2_o21ai_1  _1502_
timestamp 1747537721
transform 1 0 2688 0 1 9828
box -48 -56 538 834
use sg13g2_o21ai_1  _1503_
timestamp 1747537721
transform -1 0 6624 0 1 9828
box -48 -56 538 834
use sg13g2_nand3b_1  _1504_
timestamp 1747537721
transform -1 0 9696 0 -1 11340
box -48 -56 720 834
use sg13g2_nand3_1  _1505_
timestamp 1747537721
transform 1 0 8544 0 -1 11340
box -48 -56 528 834
use sg13g2_o21ai_1  _1506_
timestamp 1747537721
transform -1 0 9408 0 -1 12852
box -48 -56 538 834
use sg13g2_a22oi_1  _1507_
timestamp 1747537721
transform -1 0 9120 0 1 12852
box -48 -56 624 834
use sg13g2_nor2_1  _1508_
timestamp 1747537721
transform 1 0 7296 0 1 17388
box -48 -56 432 834
use sg13g2_nor2_1  _1509_
timestamp 1747537721
transform 1 0 6528 0 1 17388
box -48 -56 432 834
use sg13g2_o21ai_1  _1510_
timestamp 1747537721
transform 1 0 5472 0 1 18900
box -48 -56 538 834
use sg13g2_a21oi_2  _1511_
timestamp 1747537721
transform 1 0 5664 0 -1 20412
box -48 -56 816 834
use sg13g2_a22oi_1  _1512_
timestamp 1747537721
transform -1 0 7872 0 1 11340
box -48 -56 624 834
use sg13g2_o21ai_1  _1513_
timestamp 1747537721
transform -1 0 7680 0 -1 11340
box -48 -56 538 834
use sg13g2_nor2_1  _1514_
timestamp 1747537721
transform -1 0 7488 0 1 9828
box -48 -56 432 834
use sg13g2_nor2_1  _1515_
timestamp 1747537721
transform 1 0 6720 0 -1 9828
box -48 -56 432 834
use sg13g2_a22oi_1  _1516_
timestamp 1747537721
transform -1 0 2592 0 -1 9828
box -48 -56 624 834
use sg13g2_xor2_1  _1517_
timestamp 1747537721
transform 1 0 6144 0 1 3780
box -48 -56 816 834
use sg13g2_xnor2_1  _1518_
timestamp 1747537721
transform 1 0 6912 0 1 3780
box -48 -56 816 834
use sg13g2_and2_1  _1519_
timestamp 1747537721
transform 1 0 5856 0 -1 3780
box -48 -56 528 834
use sg13g2_or2_1  _1520_
timestamp 1747537721
transform -1 0 7200 0 -1 2268
box -48 -56 528 834
use sg13g2_nand2b_1  _1521_
timestamp 1747537721
transform 1 0 7584 0 1 2268
box -48 -56 528 834
use sg13g2_o21ai_1  _1522_
timestamp 1747537721
transform 1 0 1632 0 1 3780
box -48 -56 538 834
use sg13g2_xnor2_1  _1523_
timestamp 1747537721
transform 1 0 6816 0 1 2268
box -48 -56 816 834
use sg13g2_o21ai_1  _1524_
timestamp 1747537721
transform 1 0 7296 0 -1 5292
box -48 -56 538 834
use sg13g2_a21oi_1  _1525_
timestamp 1747537721
transform 1 0 7776 0 -1 5292
box -48 -56 528 834
use sg13g2_nor3_1  _1526_
timestamp 1747537721
transform -1 0 16992 0 -1 9828
box -48 -56 528 834
use sg13g2_nor2_1  _1527_
timestamp 1747537721
transform 1 0 15360 0 -1 9828
box -48 -56 432 834
use sg13g2_o21ai_1  _1528_
timestamp 1747537721
transform 1 0 7104 0 -1 9828
box -48 -56 538 834
use sg13g2_o21ai_1  _1529_
timestamp 1747537721
transform -1 0 7296 0 -1 12852
box -48 -56 538 834
use sg13g2_a22oi_1  _1530_
timestamp 1747537721
transform 1 0 6528 0 1 12852
box -48 -56 624 834
use sg13g2_nor2_1  _1531_
timestamp 1747537721
transform 1 0 6432 0 1 15876
box -48 -56 432 834
use sg13g2_nor2_1  _1532_
timestamp 1747537721
transform 1 0 4992 0 -1 17388
box -48 -56 432 834
use sg13g2_o21ai_1  _1533_
timestamp 1747537721
transform -1 0 4704 0 1 17388
box -48 -56 538 834
use sg13g2_a21oi_1  _1534_
timestamp 1747537721
transform 1 0 3264 0 1 17388
box -48 -56 528 834
use sg13g2_a22oi_1  _1535_
timestamp 1747537721
transform 1 0 10464 0 -1 12852
box -48 -56 624 834
use sg13g2_o21ai_1  _1536_
timestamp 1747537721
transform -1 0 11040 0 -1 14364
box -48 -56 538 834
use sg13g2_o21ai_1  _1537_
timestamp 1747537721
transform -1 0 10944 0 1 9828
box -48 -56 538 834
use sg13g2_and2_1  _1538_
timestamp 1747537721
transform 1 0 10560 0 1 2268
box -48 -56 528 834
use sg13g2_xor2_1  _1539_
timestamp 1747537721
transform 1 0 9792 0 -1 2268
box -48 -56 816 834
use sg13g2_a21o_1  _1540_
timestamp 1747537721
transform -1 0 6816 0 1 2268
box -48 -56 720 834
use sg13g2_xor2_1  _1541_
timestamp 1747537721
transform -1 0 11328 0 -1 2268
box -48 -56 816 834
use sg13g2_or2_1  _1542_
timestamp 1747537721
transform 1 0 7392 0 -1 3780
box -48 -56 528 834
use sg13g2_o21ai_1  _1543_
timestamp 1747537721
transform 1 0 7680 0 1 3780
box -48 -56 538 834
use sg13g2_and2_1  _1544_
timestamp 1747537721
transform -1 0 10176 0 1 3780
box -48 -56 528 834
use sg13g2_xnor2_1  _1545_
timestamp 1747537721
transform -1 0 9696 0 1 3780
box -48 -56 816 834
use sg13g2_xnor2_1  _1546_
timestamp 1747537721
transform 1 0 9216 0 -1 3780
box -48 -56 816 834
use sg13g2_xnor2_1  _1547_
timestamp 1747537721
transform 1 0 10368 0 -1 3780
box -48 -56 816 834
use sg13g2_o21ai_1  _1548_
timestamp 1747537721
transform 1 0 10944 0 1 9828
box -48 -56 538 834
use sg13g2_nor2_1  _1549_
timestamp 1747537721
transform -1 0 19968 0 1 15876
box -48 -56 432 834
use sg13g2_a21oi_1  _1550_
timestamp 1747537721
transform 1 0 16032 0 1 15876
box -48 -56 528 834
use sg13g2_a21oi_1  _1551_
timestamp 1747537721
transform -1 0 11904 0 -1 17388
box -48 -56 528 834
use sg13g2_o21ai_1  _1552_
timestamp 1747537721
transform 1 0 10464 0 -1 17388
box -48 -56 538 834
use sg13g2_a21oi_1  _1553_
timestamp 1747537721
transform 1 0 10944 0 -1 17388
box -48 -56 528 834
use sg13g2_o21ai_1  _1554_
timestamp 1747537721
transform 1 0 10368 0 1 15876
box -48 -56 538 834
use sg13g2_o21ai_1  _1555_
timestamp 1747537721
transform 1 0 11040 0 1 17388
box -48 -56 538 834
use sg13g2_nand2b_1  _1556_
timestamp 1747537721
transform 1 0 10656 0 -1 18900
box -48 -56 528 834
use sg13g2_nand2_1  _1557_
timestamp 1747537721
transform -1 0 12192 0 1 18900
box -48 -56 432 834
use sg13g2_a21oi_2  _1558_
timestamp 1747537721
transform -1 0 11520 0 1 20412
box -48 -56 816 834
use sg13g2_nor2_1  _1559_
timestamp 1747537721
transform 1 0 12576 0 1 11340
box -48 -56 432 834
use sg13g2_a221oi_1  _1560_
timestamp 1747537721
transform 1 0 12960 0 1 11340
box -48 -56 816 834
use sg13g2_or2_1  _1561_
timestamp 1747537721
transform -1 0 13920 0 -1 12852
box -48 -56 528 834
use sg13g2_nor2_1  _1562_
timestamp 1747537721
transform 1 0 13056 0 -1 11340
box -48 -56 432 834
use sg13g2_a21oi_1  _1563_
timestamp 1747537721
transform -1 0 8928 0 1 3780
box -48 -56 528 834
use sg13g2_xnor2_1  _1564_
timestamp 1747537721
transform 1 0 11328 0 -1 3780
box -48 -56 816 834
use sg13g2_xor2_1  _1565_
timestamp 1747537721
transform 1 0 12096 0 -1 3780
box -48 -56 816 834
use sg13g2_nand2_1  _1566_
timestamp 1747537721
transform -1 0 13632 0 -1 2268
box -48 -56 432 834
use sg13g2_xnor2_1  _1567_
timestamp 1747537721
transform 1 0 12384 0 1 756
box -48 -56 816 834
use sg13g2_a21oi_1  _1568_
timestamp 1747537721
transform -1 0 11328 0 1 756
box -48 -56 528 834
use sg13g2_xnor2_1  _1569_
timestamp 1747537721
transform 1 0 12480 0 -1 2268
box -48 -56 816 834
use sg13g2_a21oi_1  _1570_
timestamp 1747537721
transform -1 0 13536 0 1 2268
box -48 -56 528 834
use sg13g2_o21ai_1  _1571_
timestamp 1747537721
transform 1 0 12960 0 -1 3780
box -48 -56 538 834
use sg13g2_o21ai_1  _1572_
timestamp 1747537721
transform 1 0 13152 0 1 9828
box -48 -56 538 834
use sg13g2_nor2_1  _1573_
timestamp 1747537721
transform -1 0 19392 0 1 9828
box -48 -56 432 834
use sg13g2_a21oi_1  _1574_
timestamp 1747537721
transform 1 0 14208 0 -1 11340
box -48 -56 528 834
use sg13g2_a22oi_1  _1575_
timestamp 1747537721
transform -1 0 14304 0 1 11340
box -48 -56 624 834
use sg13g2_o21ai_1  _1576_
timestamp 1747537721
transform -1 0 13920 0 -1 11340
box -48 -56 538 834
use sg13g2_a21oi_1  _1577_
timestamp 1747537721
transform 1 0 2112 0 1 17388
box -48 -56 528 834
use sg13g2_o21ai_1  _1578_
timestamp 1747537721
transform 1 0 1536 0 -1 18900
box -48 -56 538 834
use sg13g2_a21oi_1  _1579_
timestamp 1747537721
transform -1 0 2304 0 1 18900
box -48 -56 528 834
use sg13g2_and2_1  _1580_
timestamp 1747537721
transform 1 0 14400 0 1 11340
box -48 -56 528 834
use sg13g2_a221oi_1  _1581_
timestamp 1747537721
transform 1 0 14880 0 1 11340
box -48 -56 816 834
use sg13g2_or2_1  _1582_
timestamp 1747537721
transform 1 0 15264 0 -1 11340
box -48 -56 528 834
use sg13g2_nor2_1  _1583_
timestamp 1747537721
transform -1 0 18048 0 -1 11340
box -48 -56 432 834
use sg13g2_nand2b_1  _1584_
timestamp 1747537721
transform 1 0 12288 0 1 3780
box -48 -56 528 834
use sg13g2_o21ai_1  _1585_
timestamp 1747537721
transform 1 0 12288 0 1 2268
box -48 -56 538 834
use sg13g2_nor2_1  _1586_
timestamp 1747537721
transform -1 0 16800 0 1 3780
box -48 -56 432 834
use sg13g2_xnor2_1  _1587_
timestamp 1747537721
transform 1 0 15072 0 -1 5292
box -48 -56 816 834
use sg13g2_xnor2_1  _1588_
timestamp 1747537721
transform 1 0 15840 0 -1 5292
box -48 -56 816 834
use sg13g2_and2_1  _1589_
timestamp 1747537721
transform 1 0 19104 0 -1 3780
box -48 -56 528 834
use sg13g2_xor2_1  _1590_
timestamp 1747537721
transform -1 0 21120 0 -1 3780
box -48 -56 816 834
use sg13g2_o21ai_1  _1591_
timestamp 1747537721
transform 1 0 13152 0 1 756
box -48 -56 538 834
use sg13g2_xor2_1  _1592_
timestamp 1747537721
transform -1 0 20352 0 -1 3780
box -48 -56 816 834
use sg13g2_a21oi_1  _1593_
timestamp 1747537721
transform 1 0 17088 0 -1 5292
box -48 -56 528 834
use sg13g2_o21ai_1  _1594_
timestamp 1747537721
transform -1 0 17088 0 -1 5292
box -48 -56 538 834
use sg13g2_o21ai_1  _1595_
timestamp 1747537721
transform -1 0 16896 0 1 9828
box -48 -56 538 834
use sg13g2_nor3_1  _1596_
timestamp 1747537721
transform -1 0 19008 0 1 9828
box -48 -56 528 834
use sg13g2_nor2_1  _1597_
timestamp 1747537721
transform -1 0 19392 0 -1 11340
box -48 -56 432 834
use sg13g2_a22oi_1  _1598_
timestamp 1747537721
transform -1 0 16320 0 -1 11340
box -48 -56 624 834
use sg13g2_o21ai_1  _1599_
timestamp 1747537721
transform -1 0 16128 0 1 11340
box -48 -56 538 834
use sg13g2_a21oi_1  _1600_
timestamp 1747537721
transform 1 0 2592 0 1 15876
box -48 -56 528 834
use sg13g2_o21ai_1  _1601_
timestamp 1747537721
transform -1 0 2304 0 -1 17388
box -48 -56 538 834
use sg13g2_a21oi_1  _1602_
timestamp 1747537721
transform 1 0 576 0 -1 17388
box -48 -56 528 834
use sg13g2_o21ai_1  _1603_
timestamp 1747537721
transform -1 0 17664 0 -1 11340
box -48 -56 538 834
use sg13g2_nand2_1  _1604_
timestamp 1747537721
transform -1 0 24768 0 -1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _1605_
timestamp 1747537721
transform -1 0 23808 0 1 3780
box -48 -56 432 834
use sg13g2_xnor2_1  _1606_
timestamp 1747537721
transform -1 0 24384 0 -1 3780
box -48 -56 816 834
use sg13g2_a21oi_1  _1607_
timestamp 1747537721
transform -1 0 20352 0 1 2268
box -48 -56 528 834
use sg13g2_xnor2_1  _1608_
timestamp 1747537721
transform -1 0 23616 0 -1 3780
box -48 -56 816 834
use sg13g2_a21oi_1  _1609_
timestamp 1747537721
transform -1 0 16416 0 1 3780
box -48 -56 528 834
use sg13g2_nand2b_1  _1610_
timestamp 1747537721
transform 1 0 17472 0 1 5292
box -48 -56 528 834
use sg13g2_nor2b_1  _1611_
timestamp 1747537721
transform 1 0 17376 0 -1 6804
box -54 -56 528 834
use sg13g2_xnor2_1  _1612_
timestamp 1747537721
transform 1 0 15552 0 -1 6804
box -48 -56 816 834
use sg13g2_xnor2_1  _1613_
timestamp 1747537721
transform 1 0 15936 0 1 5292
box -48 -56 816 834
use sg13g2_xnor2_1  _1614_
timestamp 1747537721
transform 1 0 16320 0 -1 6804
box -48 -56 816 834
use sg13g2_o21ai_1  _1615_
timestamp 1747537721
transform -1 0 17088 0 -1 11340
box -48 -56 538 834
use sg13g2_nor2_1  _1616_
timestamp 1747537721
transform -1 0 19584 0 -1 14364
box -48 -56 432 834
use sg13g2_a21oi_1  _1617_
timestamp 1747537721
transform 1 0 18432 0 1 14364
box -48 -56 528 834
use sg13g2_a22oi_1  _1618_
timestamp 1747537721
transform 1 0 16128 0 1 11340
box -48 -56 624 834
use sg13g2_o21ai_1  _1619_
timestamp 1747537721
transform -1 0 16800 0 1 14364
box -48 -56 538 834
use sg13g2_o21ai_1  _1620_
timestamp 1747537721
transform 1 0 15264 0 -1 15876
box -48 -56 538 834
use sg13g2_a221oi_1  _1621_
timestamp 1747537721
transform 1 0 16224 0 -1 15876
box -48 -56 816 834
use sg13g2_o21ai_1  _1622_
timestamp 1747537721
transform 1 0 15744 0 -1 15876
box -48 -56 538 834
use sg13g2_nor2_1  _1623_
timestamp 1747537721
transform -1 0 16896 0 1 15876
box -48 -56 432 834
use sg13g2_nor2_1  _1624_
timestamp 1747537721
transform 1 0 16320 0 -1 20412
box -48 -56 432 834
use sg13g2_o21ai_1  _1625_
timestamp 1747537721
transform -1 0 18144 0 -1 20412
box -48 -56 538 834
use sg13g2_a21oi_2  _1626_
timestamp 1747537721
transform -1 0 17952 0 -1 21924
box -48 -56 816 834
use sg13g2_nor2_1  _1627_
timestamp 1747537721
transform -1 0 16896 0 -1 12852
box -48 -56 432 834
use sg13g2_a221oi_1  _1628_
timestamp 1747537721
transform 1 0 16704 0 1 11340
box -48 -56 816 834
use sg13g2_or2_1  _1629_
timestamp 1747537721
transform 1 0 17952 0 1 11340
box -48 -56 528 834
use sg13g2_o21ai_1  _1630_
timestamp 1747537721
transform 1 0 17568 0 -1 9828
box -48 -56 538 834
use sg13g2_nor2_1  _1631_
timestamp 1747537721
transform 1 0 17376 0 1 9828
box -48 -56 432 834
use sg13g2_or2_1  _1632_
timestamp 1747537721
transform 1 0 17664 0 1 8316
box -48 -56 528 834
use sg13g2_o21ai_1  _1633_
timestamp 1747537721
transform 1 0 17856 0 -1 6804
box -48 -56 538 834
use sg13g2_xnor2_1  _1634_
timestamp 1747537721
transform 1 0 22848 0 -1 6804
box -48 -56 816 834
use sg13g2_o21ai_1  _1635_
timestamp 1747537721
transform 1 0 23424 0 1 2268
box -48 -56 538 834
use sg13g2_xnor2_1  _1636_
timestamp 1747537721
transform -1 0 25056 0 -1 5292
box -48 -56 816 834
use sg13g2_xnor2_1  _1637_
timestamp 1747537721
transform 1 0 23520 0 -1 5292
box -48 -56 816 834
use sg13g2_xnor2_1  _1638_
timestamp 1747537721
transform -1 0 24384 0 -1 6804
box -48 -56 816 834
use sg13g2_and2_1  _1639_
timestamp 1747537721
transform 1 0 17856 0 1 6804
box -48 -56 528 834
use sg13g2_o21ai_1  _1640_
timestamp 1747537721
transform 1 0 18336 0 1 6804
box -48 -56 538 834
use sg13g2_o21ai_1  _1641_
timestamp 1747537721
transform -1 0 18816 0 -1 8316
box -48 -56 538 834
use sg13g2_nor2_1  _1642_
timestamp 1747537721
transform -1 0 19200 0 -1 14364
box -48 -56 432 834
use sg13g2_a21oi_1  _1643_
timestamp 1747537721
transform 1 0 18624 0 1 12852
box -48 -56 528 834
use sg13g2_a22oi_1  _1644_
timestamp 1747537721
transform -1 0 18720 0 -1 12852
box -48 -56 624 834
use sg13g2_o21ai_1  _1645_
timestamp 1747537721
transform 1 0 18720 0 -1 12852
box -48 -56 538 834
use sg13g2_a21oi_1  _1646_
timestamp 1747537721
transform -1 0 19584 0 1 18900
box -48 -56 528 834
use sg13g2_o21ai_1  _1647_
timestamp 1747537721
transform 1 0 20256 0 1 18900
box -48 -56 538 834
use sg13g2_a21oi_2  _1648_
timestamp 1747537721
transform 1 0 20448 0 -1 20412
box -48 -56 816 834
use sg13g2_nor2_2  _1649_
timestamp 1747537721
transform 1 0 12480 0 -1 14364
box -48 -56 624 834
use sg13g2_nor2_1  _1650_
timestamp 1747537721
transform -1 0 6624 0 -1 14364
box -48 -56 432 834
use sg13g2_a221oi_1  _1651_
timestamp 1747537721
transform -1 0 6432 0 1 14364
box -48 -56 816 834
use sg13g2_and2_1  _1652_
timestamp 1747537721
transform -1 0 5760 0 -1 14364
box -48 -56 528 834
use sg13g2_nand2_1  _1653_
timestamp 1747537721
transform -1 0 5184 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  _1654_
timestamp 1747537721
transform 1 0 4128 0 1 5292
box -48 -56 336 834
use sg13g2_xnor2_1  _1655_
timestamp 1747537721
transform 1 0 3264 0 -1 6804
box -48 -56 816 834
use sg13g2_xnor2_1  _1656_
timestamp 1747537721
transform 1 0 4032 0 -1 6804
box -48 -56 816 834
use sg13g2_nand2_1  _1657_
timestamp 1747537721
transform 1 0 3264 0 1 3780
box -48 -56 432 834
use sg13g2_nand2_1  _1658_
timestamp 1747537721
transform 1 0 3360 0 1 5292
box -48 -56 432 834
use sg13g2_xnor2_1  _1659_
timestamp 1747537721
transform 1 0 2592 0 -1 5292
box -48 -56 816 834
use sg13g2_xor2_1  _1660_
timestamp 1747537721
transform 1 0 3360 0 -1 5292
box -48 -56 816 834
use sg13g2_a21oi_1  _1661_
timestamp 1747537721
transform -1 0 5088 0 1 6804
box -48 -56 528 834
use sg13g2_o21ai_1  _1662_
timestamp 1747537721
transform -1 0 4608 0 1 6804
box -48 -56 538 834
use sg13g2_a221oi_1  _1663_
timestamp 1747537721
transform -1 0 5088 0 -1 11340
box -48 -56 816 834
use sg13g2_o21ai_1  _1664_
timestamp 1747537721
transform 1 0 4608 0 1 12852
box -48 -56 538 834
use sg13g2_o21ai_1  _1665_
timestamp 1747537721
transform -1 0 5280 0 -1 14364
box -48 -56 538 834
use sg13g2_a21oi_1  _1666_
timestamp 1747537721
transform -1 0 7968 0 -1 18900
box -48 -56 528 834
use sg13g2_o21ai_1  _1667_
timestamp 1747537721
transform 1 0 7104 0 1 18900
box -48 -56 538 834
use sg13g2_a21oi_2  _1668_
timestamp 1747537721
transform 1 0 7584 0 1 18900
box -48 -56 816 834
use sg13g2_a22oi_1  _1669_
timestamp 1747537721
transform -1 0 6432 0 1 12852
box -48 -56 624 834
use sg13g2_o21ai_1  _1670_
timestamp 1747537721
transform -1 0 6144 0 -1 12852
box -48 -56 538 834
use sg13g2_a22oi_1  _1671_
timestamp 1747537721
transform -1 0 4992 0 1 5292
box -48 -56 624 834
use sg13g2_xor2_1  _1672_
timestamp 1747537721
transform 1 0 5088 0 -1 3780
box -48 -56 816 834
use sg13g2_xor2_1  _1673_
timestamp 1747537721
transform 1 0 5376 0 1 5292
box -48 -56 816 834
use sg13g2_and2_1  _1674_
timestamp 1747537721
transform 1 0 4704 0 1 3780
box -48 -56 528 834
use sg13g2_xor2_1  _1675_
timestamp 1747537721
transform 1 0 4320 0 -1 3780
box -48 -56 816 834
use sg13g2_o21ai_1  _1676_
timestamp 1747537721
transform 1 0 4128 0 -1 5292
box -48 -56 538 834
use sg13g2_xnor2_1  _1677_
timestamp 1747537721
transform 1 0 5088 0 -1 5292
box -48 -56 816 834
use sg13g2_a21oi_1  _1678_
timestamp 1747537721
transform -1 0 6816 0 -1 6804
box -48 -56 528 834
use sg13g2_o21ai_1  _1679_
timestamp 1747537721
transform 1 0 5856 0 -1 6804
box -48 -56 538 834
use sg13g2_a21oi_1  _1680_
timestamp 1747537721
transform -1 0 6720 0 -1 9828
box -48 -56 528 834
use sg13g2_o21ai_1  _1681_
timestamp 1747537721
transform -1 0 6240 0 -1 9828
box -48 -56 538 834
use sg13g2_o21ai_1  _1682_
timestamp 1747537721
transform -1 0 6240 0 -1 14364
box -48 -56 538 834
use sg13g2_a22oi_1  _1683_
timestamp 1747537721
transform 1 0 5280 0 1 12852
box -48 -56 624 834
use sg13g2_inv_1  _1684_
timestamp 1747537721
transform 1 0 5952 0 -1 17388
box -48 -56 336 834
use sg13g2_a21oi_1  _1685_
timestamp 1747537721
transform 1 0 5856 0 -1 18900
box -48 -56 528 834
use sg13g2_o21ai_1  _1686_
timestamp 1747537721
transform -1 0 5856 0 -1 18900
box -48 -56 538 834
use sg13g2_a21oi_1  _1687_
timestamp 1747537721
transform 1 0 6432 0 -1 20412
box -48 -56 528 834
use sg13g2_a22oi_1  _1688_
timestamp 1747537721
transform -1 0 8448 0 1 11340
box -48 -56 624 834
use sg13g2_o21ai_1  _1689_
timestamp 1747537721
transform 1 0 6816 0 1 11340
box -48 -56 538 834
use sg13g2_nand2_1  _1690_
timestamp 1747537721
transform 1 0 7968 0 1 9828
box -48 -56 432 834
use sg13g2_nand2_1  _1691_
timestamp 1747537721
transform 1 0 12960 0 1 3780
box -48 -56 432 834
use sg13g2_xnor2_1  _1692_
timestamp 1747537721
transform -1 0 13152 0 -1 5292
box -48 -56 816 834
use sg13g2_a21oi_2  _1693_
timestamp 1747537721
transform -1 0 5952 0 1 3780
box -48 -56 816 834
use sg13g2_xnor2_1  _1694_
timestamp 1747537721
transform 1 0 11616 0 -1 5292
box -48 -56 816 834
use sg13g2_or2_1  _1695_
timestamp 1747537721
transform 1 0 6144 0 1 5292
box -48 -56 528 834
use sg13g2_o21ai_1  _1696_
timestamp 1747537721
transform 1 0 6624 0 1 5292
box -48 -56 538 834
use sg13g2_and2_1  _1697_
timestamp 1747537721
transform 1 0 14400 0 -1 5292
box -48 -56 528 834
use sg13g2_xnor2_1  _1698_
timestamp 1747537721
transform -1 0 15168 0 1 5292
box -48 -56 816 834
use sg13g2_xor2_1  _1699_
timestamp 1747537721
transform -1 0 14400 0 1 5292
box -48 -56 816 834
use sg13g2_o21ai_1  _1700_
timestamp 1747537721
transform 1 0 12864 0 1 5292
box -48 -56 538 834
use sg13g2_a21oi_1  _1701_
timestamp 1747537721
transform 1 0 12384 0 1 5292
box -48 -56 528 834
use sg13g2_nor2_1  _1702_
timestamp 1747537721
transform -1 0 9120 0 -1 9828
box -48 -56 432 834
use sg13g2_o21ai_1  _1703_
timestamp 1747537721
transform 1 0 11424 0 -1 9828
box -48 -56 538 834
use sg13g2_o21ai_1  _1704_
timestamp 1747537721
transform -1 0 8832 0 1 9828
box -48 -56 538 834
use sg13g2_nand2_1  _1705_
timestamp 1747537721
transform -1 0 8064 0 -1 12852
box -48 -56 432 834
use sg13g2_o21ai_1  _1706_
timestamp 1747537721
transform -1 0 8448 0 -1 11340
box -48 -56 538 834
use sg13g2_a21oi_1  _1707_
timestamp 1747537721
transform 1 0 4416 0 1 15876
box -48 -56 528 834
use sg13g2_o21ai_1  _1708_
timestamp 1747537721
transform 1 0 3744 0 1 17388
box -48 -56 538 834
use sg13g2_a21oi_1  _1709_
timestamp 1747537721
transform 1 0 3936 0 -1 18900
box -48 -56 528 834
use sg13g2_a21oi_1  _1710_
timestamp 1747537721
transform -1 0 15648 0 1 5292
box -48 -56 528 834
use sg13g2_xnor2_1  _1711_
timestamp 1747537721
transform 1 0 17952 0 1 3780
box -48 -56 816 834
use sg13g2_xnor2_1  _1712_
timestamp 1747537721
transform 1 0 17760 0 -1 5292
box -48 -56 816 834
use sg13g2_and2_1  _1713_
timestamp 1747537721
transform 1 0 25632 0 -1 3780
box -48 -56 528 834
use sg13g2_xor2_1  _1714_
timestamp 1747537721
transform 1 0 24864 0 -1 3780
box -48 -56 816 834
use sg13g2_o21ai_1  _1715_
timestamp 1747537721
transform 1 0 13152 0 -1 5292
box -48 -56 538 834
use sg13g2_xor2_1  _1716_
timestamp 1747537721
transform -1 0 25440 0 1 3780
box -48 -56 816 834
use sg13g2_a21oi_1  _1717_
timestamp 1747537721
transform 1 0 19008 0 -1 5292
box -48 -56 528 834
use sg13g2_o21ai_1  _1718_
timestamp 1747537721
transform -1 0 19008 0 -1 5292
box -48 -56 538 834
use sg13g2_nand2b_1  _1719_
timestamp 1747537721
transform 1 0 11040 0 -1 12852
box -48 -56 528 834
use sg13g2_o21ai_1  _1720_
timestamp 1747537721
transform 1 0 11040 0 -1 11340
box -48 -56 538 834
use sg13g2_a21oi_2  _1721_
timestamp 1747537721
transform 1 0 10848 0 1 11340
box -48 -56 816 834
use sg13g2_a22oi_1  _1722_
timestamp 1747537721
transform 1 0 12000 0 1 9828
box -48 -56 624 834
use sg13g2_o21ai_1  _1723_
timestamp 1747537721
transform 1 0 11520 0 1 9828
box -48 -56 538 834
use sg13g2_o21ai_1  _1724_
timestamp 1747537721
transform 1 0 11328 0 -1 15876
box -48 -56 538 834
use sg13g2_a21oi_1  _1725_
timestamp 1747537721
transform 1 0 12000 0 1 15876
box -48 -56 528 834
use sg13g2_nor2_1  _1726_
timestamp 1747537721
transform 1 0 11136 0 -1 18900
box -48 -56 432 834
use sg13g2_o21ai_1  _1727_
timestamp 1747537721
transform -1 0 11328 0 1 18900
box -48 -56 538 834
use sg13g2_a21oi_2  _1728_
timestamp 1747537721
transform 1 0 10752 0 -1 20412
box -48 -56 816 834
use sg13g2_nand2b_1  _1729_
timestamp 1747537721
transform 1 0 18048 0 1 5292
box -48 -56 528 834
use sg13g2_o21ai_1  _1730_
timestamp 1747537721
transform 1 0 18528 0 1 5292
box -48 -56 538 834
use sg13g2_nor2_1  _1731_
timestamp 1747537721
transform 1 0 25152 0 1 5292
box -48 -56 432 834
use sg13g2_xor2_1  _1732_
timestamp 1747537721
transform 1 0 24384 0 1 5292
box -48 -56 816 834
use sg13g2_xnor2_1  _1733_
timestamp 1747537721
transform -1 0 26496 0 -1 6804
box -48 -56 816 834
use sg13g2_a21oi_1  _1734_
timestamp 1747537721
transform 1 0 26592 0 1 3780
box -48 -56 528 834
use sg13g2_nor2_1  _1735_
timestamp 1747537721
transform 1 0 27072 0 1 3780
box -48 -56 432 834
use sg13g2_xor2_1  _1736_
timestamp 1747537721
transform -1 0 27264 0 -1 5292
box -48 -56 816 834
use sg13g2_xnor2_1  _1737_
timestamp 1747537721
transform -1 0 26496 0 -1 5292
box -48 -56 816 834
use sg13g2_xnor2_1  _1738_
timestamp 1747537721
transform -1 0 26304 0 1 5292
box -48 -56 816 834
use sg13g2_o21ai_1  _1739_
timestamp 1747537721
transform -1 0 17376 0 1 8316
box -48 -56 538 834
use sg13g2_a21oi_1  _1740_
timestamp 1747537721
transform -1 0 14016 0 1 8316
box -48 -56 528 834
use sg13g2_a22oi_1  _1741_
timestamp 1747537721
transform -1 0 13440 0 1 12852
box -48 -56 624 834
use sg13g2_o21ai_1  _1742_
timestamp 1747537721
transform -1 0 12864 0 1 12852
box -48 -56 538 834
use sg13g2_inv_1  _1743_
timestamp 1747537721
transform 1 0 12768 0 1 14364
box -48 -56 336 834
use sg13g2_o21ai_1  _1744_
timestamp 1747537721
transform -1 0 14304 0 1 14364
box -48 -56 538 834
use sg13g2_a221oi_1  _1745_
timestamp 1747537721
transform 1 0 13056 0 1 14364
box -48 -56 816 834
use sg13g2_a21oi_1  _1746_
timestamp 1747537721
transform -1 0 13632 0 -1 15876
box -48 -56 528 834
use sg13g2_a21oi_1  _1747_
timestamp 1747537721
transform 1 0 2496 0 -1 18900
box -48 -56 528 834
use sg13g2_o21ai_1  _1748_
timestamp 1747537721
transform -1 0 3456 0 -1 18900
box -48 -56 538 834
use sg13g2_a21oi_1  _1749_
timestamp 1747537721
transform 1 0 2400 0 1 18900
box -48 -56 528 834
use sg13g2_a21oi_2  _1750_
timestamp 1747537721
transform 1 0 24960 0 -1 6804
box -48 -56 816 834
use sg13g2_nor2b_1  _1751_
timestamp 1747537721
transform 1 0 27744 0 -1 5292
box -54 -56 528 834
use sg13g2_xnor2_1  _1752_
timestamp 1747537721
transform 1 0 27360 0 1 5292
box -48 -56 816 834
use sg13g2_nand2b_1  _1753_
timestamp 1747537721
transform 1 0 30048 0 1 5292
box -48 -56 528 834
use sg13g2_xor2_1  _1754_
timestamp 1747537721
transform -1 0 28224 0 -1 6804
box -48 -56 816 834
use sg13g2_xnor2_1  _1755_
timestamp 1747537721
transform 1 0 27168 0 -1 3780
box -48 -56 816 834
use sg13g2_a221oi_1  _1756_
timestamp 1747537721
transform 1 0 25824 0 1 3780
box -48 -56 816 834
use sg13g2_nor3_1  _1757_
timestamp 1747537721
transform -1 0 28416 0 1 3780
box -48 -56 528 834
use sg13g2_o21ai_1  _1758_
timestamp 1747537721
transform 1 0 29472 0 1 3780
box -48 -56 538 834
use sg13g2_nand2b_1  _1759_
timestamp 1747537721
transform -1 0 27936 0 1 3780
box -48 -56 528 834
use sg13g2_xnor2_1  _1760_
timestamp 1747537721
transform -1 0 27456 0 -1 6804
box -48 -56 816 834
use sg13g2_a21oi_1  _1761_
timestamp 1747537721
transform 1 0 17856 0 -1 8316
box -48 -56 528 834
use sg13g2_o21ai_1  _1762_
timestamp 1747537721
transform -1 0 15840 0 1 9828
box -48 -56 538 834
use sg13g2_nand2_1  _1763_
timestamp 1747537721
transform 1 0 14688 0 -1 12852
box -48 -56 432 834
use sg13g2_a22oi_1  _1764_
timestamp 1747537721
transform 1 0 15264 0 1 12852
box -48 -56 624 834
use sg13g2_nand2_1  _1765_
timestamp 1747537721
transform -1 0 14688 0 1 12852
box -48 -56 432 834
use sg13g2_o21ai_1  _1766_
timestamp 1747537721
transform 1 0 14304 0 -1 15876
box -48 -56 538 834
use sg13g2_a21oi_1  _1767_
timestamp 1747537721
transform 1 0 14784 0 -1 15876
box -48 -56 528 834
use sg13g2_o21ai_1  _1768_
timestamp 1747537721
transform -1 0 15264 0 -1 11340
box -48 -56 538 834
use sg13g2_o21ai_1  _1769_
timestamp 1747537721
transform -1 0 13344 0 1 15876
box -48 -56 538 834
use sg13g2_inv_1  _1770_
timestamp 1747537721
transform -1 0 3936 0 -1 15876
box -48 -56 336 834
use sg13g2_a21oi_1  _1771_
timestamp 1747537721
transform 1 0 2688 0 -1 15876
box -48 -56 528 834
use sg13g2_o21ai_1  _1772_
timestamp 1747537721
transform -1 0 2016 0 1 15876
box -48 -56 538 834
use sg13g2_a21oi_1  _1773_
timestamp 1747537721
transform 1 0 1344 0 1 17388
box -48 -56 528 834
use sg13g2_nor3_1  _1774_
timestamp 1747537721
transform -1 0 29280 0 1 6804
box -48 -56 528 834
use sg13g2_or3_1  _1775_
timestamp 1747537721
transform 1 0 28224 0 -1 6804
box -48 -56 720 834
use sg13g2_o21ai_1  _1776_
timestamp 1747537721
transform 1 0 28896 0 -1 6804
box -48 -56 538 834
use sg13g2_a21oi_1  _1777_
timestamp 1747537721
transform -1 0 29856 0 -1 6804
box -48 -56 528 834
use sg13g2_nand3_1  _1778_
timestamp 1747537721
transform 1 0 29280 0 1 6804
box -48 -56 528 834
use sg13g2_nand3_1  _1779_
timestamp 1747537721
transform 1 0 28896 0 1 5292
box -48 -56 528 834
use sg13g2_o21ai_1  _1780_
timestamp 1747537721
transform 1 0 29760 0 1 6804
box -48 -56 538 834
use sg13g2_a21oi_1  _1781_
timestamp 1747537721
transform 1 0 30528 0 1 5292
box -48 -56 528 834
use sg13g2_nand2_1  _1782_
timestamp 1747537721
transform 1 0 30816 0 1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _1783_
timestamp 1747537721
transform 1 0 29280 0 -1 5292
box -48 -56 432 834
use sg13g2_xnor2_1  _1784_
timestamp 1747537721
transform 1 0 29664 0 -1 5292
box -48 -56 816 834
use sg13g2_a21oi_1  _1785_
timestamp 1747537721
transform 1 0 28224 0 -1 5292
box -48 -56 528 834
use sg13g2_xnor2_1  _1786_
timestamp 1747537721
transform -1 0 31200 0 -1 5292
box -48 -56 816 834
use sg13g2_xnor2_1  _1787_
timestamp 1747537721
transform -1 0 31008 0 -1 6804
box -48 -56 816 834
use sg13g2_o21ai_1  _1788_
timestamp 1747537721
transform -1 0 18624 0 1 8316
box -48 -56 538 834
use sg13g2_a21oi_1  _1789_
timestamp 1747537721
transform 1 0 17952 0 1 14364
box -48 -56 528 834
use sg13g2_nor2_1  _1790_
timestamp 1747537721
transform -1 0 17184 0 1 14364
box -48 -56 432 834
use sg13g2_a221oi_1  _1791_
timestamp 1747537721
transform 1 0 17184 0 1 14364
box -48 -56 816 834
use sg13g2_a21oi_1  _1792_
timestamp 1747537721
transform 1 0 17088 0 -1 15876
box -48 -56 528 834
use sg13g2_o21ai_1  _1793_
timestamp 1747537721
transform 1 0 18240 0 -1 15876
box -48 -56 538 834
use sg13g2_a21o_1  _1794_
timestamp 1747537721
transform 1 0 17568 0 -1 15876
box -48 -56 720 834
use sg13g2_a21oi_1  _1795_
timestamp 1747537721
transform 1 0 18240 0 -1 18900
box -48 -56 528 834
use sg13g2_a21oi_1  _1796_
timestamp 1747537721
transform 1 0 17568 0 1 18900
box -48 -56 528 834
use sg13g2_o21ai_1  _1797_
timestamp 1747537721
transform -1 0 17184 0 -1 20412
box -48 -56 538 834
use sg13g2_a21oi_2  _1798_
timestamp 1747537721
transform -1 0 17184 0 -1 21924
box -48 -56 816 834
use sg13g2_xor2_1  _1799_
timestamp 1747537721
transform -1 0 24192 0 1 8316
box -48 -56 816 834
use sg13g2_a21oi_1  _1800_
timestamp 1747537721
transform 1 0 19680 0 1 9828
box -48 -56 528 834
use sg13g2_o21ai_1  _1801_
timestamp 1747537721
transform 1 0 30336 0 1 3780
box -48 -56 538 834
use sg13g2_xnor2_1  _1802_
timestamp 1747537721
transform 1 0 30240 0 -1 8316
box -48 -56 816 834
use sg13g2_xnor2_1  _1803_
timestamp 1747537721
transform -1 0 31104 0 1 6804
box -48 -56 816 834
use sg13g2_xnor2_1  _1804_
timestamp 1747537721
transform 1 0 28512 0 -1 8316
box -48 -56 816 834
use sg13g2_a21oi_1  _1805_
timestamp 1747537721
transform -1 0 28896 0 1 5292
box -48 -56 528 834
use sg13g2_o21ai_1  _1806_
timestamp 1747537721
transform 1 0 29568 0 1 5292
box -48 -56 538 834
use sg13g2_xnor2_1  _1807_
timestamp 1747537721
transform 1 0 29472 0 -1 8316
box -48 -56 816 834
use sg13g2_xnor2_1  _1808_
timestamp 1747537721
transform -1 0 30528 0 1 8316
box -48 -56 816 834
use sg13g2_a21oi_1  _1809_
timestamp 1747537721
transform 1 0 19968 0 1 8316
box -48 -56 528 834
use sg13g2_o21ai_1  _1810_
timestamp 1747537721
transform 1 0 19776 0 -1 9828
box -48 -56 538 834
use sg13g2_nor2_1  _1811_
timestamp 1747537721
transform -1 0 17280 0 -1 12852
box -48 -56 432 834
use sg13g2_a221oi_1  _1812_
timestamp 1747537721
transform 1 0 17760 0 1 12852
box -48 -56 816 834
use sg13g2_nor2_1  _1813_
timestamp 1747537721
transform 1 0 17568 0 1 15876
box -48 -56 432 834
use sg13g2_a221oi_1  _1814_
timestamp 1747537721
transform 1 0 17760 0 -1 17388
box -48 -56 816 834
use sg13g2_o21ai_1  _1815_
timestamp 1747537721
transform -1 0 19776 0 -1 9828
box -48 -56 538 834
use sg13g2_a21oi_1  _1816_
timestamp 1747537721
transform -1 0 18336 0 1 17388
box -48 -56 528 834
use sg13g2_a21oi_1  _1817_
timestamp 1747537721
transform -1 0 19968 0 -1 18900
box -48 -56 528 834
use sg13g2_o21ai_1  _1818_
timestamp 1747537721
transform 1 0 19968 0 -1 18900
box -48 -56 538 834
use sg13g2_a21oi_2  _1819_
timestamp 1747537721
transform 1 0 20736 0 1 18900
box -48 -56 816 834
use sg13g2_a21o_1  _1820_
timestamp 1747537721
transform 1 0 4128 0 -1 26460
box -48 -56 720 834
use sg13g2_nand3_1  _1821_
timestamp 1747537721
transform -1 0 27072 0 1 14364
box -48 -56 528 834
use sg13g2_o21ai_1  _1822_
timestamp 1747537721
transform -1 0 25728 0 1 14364
box -48 -56 538 834
use sg13g2_nand2_1  _1823_
timestamp 1747537721
transform -1 0 25248 0 -1 14364
box -48 -56 432 834
use sg13g2_nor4_1  _1824_
timestamp 1747537721
transform 1 0 24480 0 1 14364
box -48 -56 624 834
use sg13g2_nand3_1  _1825_
timestamp 1747537721
transform 1 0 23904 0 1 14364
box -48 -56 528 834
use sg13g2_o21ai_1  _1826_
timestamp 1747537721
transform 1 0 24000 0 -1 15876
box -48 -56 538 834
use sg13g2_and3_2  _1827_
timestamp 1747537721
transform -1 0 25248 0 -1 15876
box -48 -56 720 834
use sg13g2_nand3_1  _1828_
timestamp 1747537721
transform -1 0 25728 0 -1 15876
box -48 -56 528 834
use sg13g2_nor2_2  _1829_
timestamp 1747537721
transform 1 0 27264 0 -1 24948
box -48 -56 624 834
use sg13g2_nand2_2  _1830_
timestamp 1747537721
transform -1 0 23616 0 1 17388
box -48 -56 624 834
use sg13g2_and2_1  _1831_
timestamp 1747537721
transform 1 0 29088 0 1 17388
box -48 -56 528 834
use sg13g2_nor3_1  _1832_
timestamp 1747537721
transform 1 0 23808 0 -1 11340
box -48 -56 528 834
use sg13g2_xnor2_1  _1833_
timestamp 1747537721
transform -1 0 25248 0 -1 9828
box -48 -56 816 834
use sg13g2_nor2_1  _1834_
timestamp 1747537721
transform 1 0 24384 0 1 8316
box -48 -56 432 834
use sg13g2_nor2_1  _1835_
timestamp 1747537721
transform 1 0 23232 0 -1 11340
box -48 -56 432 834
use sg13g2_xnor2_1  _1836_
timestamp 1747537721
transform 1 0 22464 0 -1 11340
box -48 -56 816 834
use sg13g2_nor2_1  _1837_
timestamp 1747537721
transform 1 0 23520 0 -1 9828
box -48 -56 432 834
use sg13g2_xnor2_1  _1838_
timestamp 1747537721
transform 1 0 28128 0 -1 9828
box -48 -56 816 834
use sg13g2_nor2_1  _1839_
timestamp 1747537721
transform -1 0 30432 0 1 11340
box -48 -56 432 834
use sg13g2_nand2_1  _1840_
timestamp 1747537721
transform 1 0 26592 0 1 9828
box -48 -56 432 834
use sg13g2_nor2_2  _1841_
timestamp 1747537721
transform -1 0 28800 0 1 9828
box -48 -56 624 834
use sg13g2_a21oi_1  _1842_
timestamp 1747537721
transform -1 0 27936 0 -1 9828
box -48 -56 528 834
use sg13g2_nor3_1  _1843_
timestamp 1747537721
transform 1 0 26496 0 -1 9828
box -48 -56 528 834
use sg13g2_o21ai_1  _1844_
timestamp 1747537721
transform -1 0 28608 0 1 11340
box -48 -56 538 834
use sg13g2_a21oi_1  _1845_
timestamp 1747537721
transform -1 0 28128 0 1 11340
box -48 -56 528 834
use sg13g2_nor3_1  _1846_
timestamp 1747537721
transform -1 0 30336 0 1 9828
box -48 -56 528 834
use sg13g2_xnor2_1  _1847_
timestamp 1747537721
transform 1 0 27264 0 -1 11340
box -48 -56 816 834
use sg13g2_nor2_1  _1848_
timestamp 1747537721
transform -1 0 30048 0 1 11340
box -48 -56 432 834
use sg13g2_nand3_1  _1849_
timestamp 1747537721
transform 1 0 28128 0 -1 12852
box -48 -56 528 834
use sg13g2_xor2_1  _1850_
timestamp 1747537721
transform 1 0 28128 0 -1 14364
box -48 -56 816 834
use sg13g2_nor2_1  _1851_
timestamp 1747537721
transform -1 0 29088 0 1 12852
box -48 -56 432 834
use sg13g2_nor2_1  _1852_
timestamp 1747537721
transform -1 0 31008 0 1 14364
box -48 -56 432 834
use sg13g2_xnor2_1  _1853_
timestamp 1747537721
transform -1 0 28896 0 1 14364
box -48 -56 816 834
use sg13g2_nor2_1  _1854_
timestamp 1747537721
transform 1 0 27744 0 1 14364
box -48 -56 432 834
use sg13g2_nand3_1  _1855_
timestamp 1747537721
transform 1 0 26784 0 1 24948
box -48 -56 528 834
use sg13g2_nor4_1  _1856_
timestamp 1747537721
transform 1 0 25440 0 1 20412
box -48 -56 624 834
use sg13g2_nor2_1  _1857_
timestamp 1747537721
transform -1 0 26304 0 -1 21924
box -48 -56 432 834
use sg13g2_and3_1  _1858_
timestamp 1747537721
transform 1 0 26112 0 1 24948
box -48 -56 720 834
use sg13g2_nand3_1  _1859_
timestamp 1747537721
transform -1 0 27264 0 1 20412
box -48 -56 528 834
use sg13g2_and2_1  _1860_
timestamp 1747537721
transform 1 0 25440 0 -1 21924
box -48 -56 528 834
use sg13g2_nor4_2  _1861_
timestamp 1747537721
transform 1 0 24864 0 -1 20412
box -48 -56 1200 834
use sg13g2_or4_1  _1862_
timestamp 1747537721
transform 1 0 26016 0 1 20412
box -48 -56 816 834
use sg13g2_nand4_1  _1863_
timestamp 1747537721
transform 1 0 26304 0 -1 21924
box -48 -56 624 834
use sg13g2_o21ai_1  _1864_
timestamp 1747537721
transform 1 0 27264 0 1 20412
box -48 -56 538 834
use sg13g2_inv_1  _1865_
timestamp 1747537721
transform -1 0 26688 0 -1 20412
box -48 -56 336 834
use sg13g2_nor3_1  _1866_
timestamp 1747537721
transform 1 0 24384 0 -1 20412
box -48 -56 528 834
use sg13g2_nor2b_2  _1867_
timestamp 1747537721
transform 1 0 24672 0 1 18900
box -54 -56 720 834
use sg13g2_nor2_1  _1868_
timestamp 1747537721
transform -1 0 5376 0 -1 21924
box -48 -56 432 834
use sg13g2_nor2b_1  _1869_
timestamp 1747537721
transform 1 0 4512 0 -1 21924
box -54 -56 528 834
use sg13g2_nor3_1  _1870_
timestamp 1747537721
transform 1 0 4032 0 -1 21924
box -48 -56 528 834
use sg13g2_a21oi_1  _1871_
timestamp 1747537721
transform -1 0 2112 0 -1 14364
box -48 -56 528 834
use sg13g2_and4_1  _1872_
timestamp 1747537721
transform -1 0 3264 0 1 14364
box -48 -56 816 834
use sg13g2_and3_1  _1873_
timestamp 1747537721
transform -1 0 1632 0 1 14364
box -48 -56 720 834
use sg13g2_nor3_1  _1874_
timestamp 1747537721
transform 1 0 960 0 -1 14364
box -48 -56 528 834
use sg13g2_nor2_1  _1875_
timestamp 1747537721
transform -1 0 1632 0 -1 12852
box -48 -56 432 834
use sg13g2_and2_1  _1876_
timestamp 1747537721
transform -1 0 1056 0 1 9828
box -48 -56 528 834
use sg13g2_nor3_1  _1877_
timestamp 1747537721
transform -1 0 1536 0 -1 11340
box -48 -56 528 834
use sg13g2_nor2b_1  _1878_
timestamp 1747537721
transform 1 0 1056 0 -1 9828
box -54 -56 528 834
use sg13g2_a21oi_1  _1879_
timestamp 1747537721
transform -1 0 2016 0 1 2268
box -48 -56 528 834
use sg13g2_o21ai_1  _1880_
timestamp 1747537721
transform -1 0 1536 0 1 2268
box -48 -56 538 834
use sg13g2_inv_1  _1881_
timestamp 1747537721
transform 1 0 1056 0 -1 3780
box -48 -56 336 834
use sg13g2_nand2_1  _1882_
timestamp 1747537721
transform 1 0 2976 0 1 2268
box -48 -56 432 834
use sg13g2_xor2_1  _1883_
timestamp 1747537721
transform -1 0 4800 0 -1 2268
box -48 -56 816 834
use sg13g2_nor2_1  _1884_
timestamp 1747537721
transform 1 0 1152 0 -1 2268
box -48 -56 432 834
use sg13g2_nor2_1  _1885_
timestamp 1747537721
transform 1 0 4128 0 1 756
box -48 -56 432 834
use sg13g2_a21oi_1  _1886_
timestamp 1747537721
transform -1 0 5856 0 1 756
box -48 -56 528 834
use sg13g2_o21ai_1  _1887_
timestamp 1747537721
transform 1 0 4896 0 1 756
box -48 -56 538 834
use sg13g2_inv_1  _1888_
timestamp 1747537721
transform 1 0 4608 0 1 756
box -48 -56 336 834
use sg13g2_and4_2  _1889_
timestamp 1747537721
transform 1 0 4416 0 1 2268
box -48 -56 912 834
use sg13g2_xnor2_1  _1890_
timestamp 1747537721
transform -1 0 15360 0 1 756
box -48 -56 816 834
use sg13g2_nor2_1  _1891_
timestamp 1747537721
transform 1 0 14208 0 1 756
box -48 -56 432 834
use sg13g2_a21oi_1  _1892_
timestamp 1747537721
transform -1 0 18336 0 -1 2268
box -48 -56 528 834
use sg13g2_and3_1  _1893_
timestamp 1747537721
transform 1 0 18336 0 -1 2268
box -48 -56 720 834
use sg13g2_nor3_1  _1894_
timestamp 1747537721
transform -1 0 19200 0 1 756
box -48 -56 528 834
use sg13g2_nand3_1  _1895_
timestamp 1747537721
transform 1 0 22464 0 1 2268
box -48 -56 528 834
use sg13g2_xnor2_1  _1896_
timestamp 1747537721
transform 1 0 22464 0 -1 2268
box -48 -56 816 834
use sg13g2_nor2_1  _1897_
timestamp 1747537721
transform -1 0 23616 0 -1 2268
box -48 -56 432 834
use sg13g2_nor2_1  _1898_
timestamp 1747537721
transform 1 0 23904 0 1 2268
box -48 -56 432 834
use sg13g2_nor2_1  _1899_
timestamp 1747537721
transform -1 0 26400 0 1 756
box -48 -56 432 834
use sg13g2_a21oi_1  _1900_
timestamp 1747537721
transform 1 0 25056 0 1 2268
box -48 -56 528 834
use sg13g2_nor2b_1  _1901_
timestamp 1747537721
transform 1 0 24096 0 -1 2268
box -54 -56 528 834
use sg13g2_or3_1  _1902_
timestamp 1747537721
transform 1 0 24288 0 1 2268
box -48 -56 720 834
use sg13g2_xor2_1  _1903_
timestamp 1747537721
transform -1 0 28896 0 -1 3780
box -48 -56 816 834
use sg13g2_nor2_1  _1904_
timestamp 1747537721
transform 1 0 28512 0 1 2268
box -48 -56 432 834
use sg13g2_nor2_1  _1905_
timestamp 1747537721
transform -1 0 28512 0 1 2268
box -48 -56 432 834
use sg13g2_nor2_1  _1906_
timestamp 1747537721
transform -1 0 31296 0 -1 2268
box -48 -56 432 834
use sg13g2_a21oi_1  _1907_
timestamp 1747537721
transform 1 0 28416 0 -1 2268
box -48 -56 528 834
use sg13g2_nor2b_1  _1908_
timestamp 1747537721
transform 1 0 28896 0 1 2268
box -54 -56 528 834
use sg13g2_xor2_1  _1909_
timestamp 1747537721
transform -1 0 13728 0 -1 21924
box -48 -56 816 834
use sg13g2_xor2_1  _1910_
timestamp 1747537721
transform 1 0 3072 0 -1 23436
box -48 -56 816 834
use sg13g2_xor2_1  _1911_
timestamp 1747537721
transform 1 0 3072 0 1 20412
box -48 -56 816 834
use sg13g2_nor3_1  _1912_
timestamp 1747537721
transform -1 0 12192 0 -1 23436
box -48 -56 528 834
use sg13g2_nor3_1  _1913_
timestamp 1747537721
transform -1 0 13344 0 1 21924
box -48 -56 528 834
use sg13g2_nor2_1  _1914_
timestamp 1747537721
transform 1 0 11712 0 1 23436
box -48 -56 432 834
use sg13g2_nand2_2  _1915_
timestamp 1747537721
transform 1 0 7968 0 -1 17388
box -48 -56 624 834
use sg13g2_and2_1  _1916_
timestamp 1747537721
transform 1 0 4032 0 -1 24948
box -48 -56 528 834
use sg13g2_a221oi_1  _1917_
timestamp 1747537721
transform 1 0 9696 0 -1 24948
box -48 -56 816 834
use sg13g2_a21oi_1  _1918_
timestamp 1747537721
transform 1 0 10464 0 1 26460
box -48 -56 528 834
use sg13g2_and2_1  _1919_
timestamp 1747537721
transform 1 0 9600 0 -1 26460
box -48 -56 528 834
use sg13g2_a221oi_1  _1920_
timestamp 1747537721
transform 1 0 10080 0 -1 26460
box -48 -56 816 834
use sg13g2_a21oi_1  _1921_
timestamp 1747537721
transform 1 0 14016 0 1 26460
box -48 -56 528 834
use sg13g2_nand3_1  _1922_
timestamp 1747537721
transform 1 0 8832 0 -1 26460
box -48 -56 528 834
use sg13g2_a21oi_1  _1923_
timestamp 1747537721
transform -1 0 12768 0 1 24948
box -48 -56 528 834
use sg13g2_a22oi_1  _1924_
timestamp 1747537721
transform 1 0 12192 0 -1 26460
box -48 -56 624 834
use sg13g2_and2_1  _1925_
timestamp 1747537721
transform 1 0 8832 0 -1 24948
box -48 -56 528 834
use sg13g2_a221oi_1  _1926_
timestamp 1747537721
transform 1 0 9216 0 1 24948
box -48 -56 816 834
use sg13g2_a21oi_1  _1927_
timestamp 1747537721
transform 1 0 18528 0 -1 26460
box -48 -56 528 834
use sg13g2_nand2_1  _1928_
timestamp 1747537721
transform 1 0 14976 0 1 23436
box -48 -56 432 834
use sg13g2_nand3_1  _1929_
timestamp 1747537721
transform 1 0 12192 0 -1 23436
box -48 -56 528 834
use sg13g2_nand3_1  _1930_
timestamp 1747537721
transform 1 0 12672 0 -1 23436
box -48 -56 528 834
use sg13g2_and2_1  _1931_
timestamp 1747537721
transform 1 0 8064 0 1 24948
box -48 -56 528 834
use sg13g2_a22oi_1  _1932_
timestamp 1747537721
transform 1 0 8256 0 -1 24948
box -48 -56 624 834
use sg13g2_nand2_1  _1933_
timestamp 1747537721
transform 1 0 18144 0 -1 24948
box -48 -56 432 834
use sg13g2_o21ai_1  _1934_
timestamp 1747537721
transform 1 0 14400 0 -1 24948
box -48 -56 538 834
use sg13g2_nand3_1  _1935_
timestamp 1747537721
transform 1 0 10464 0 1 24948
box -48 -56 528 834
use sg13g2_o21ai_1  _1936_
timestamp 1747537721
transform 1 0 11040 0 -1 26460
box -48 -56 538 834
use sg13g2_mux2_1  _1937_
timestamp 1747537721
transform 1 0 16896 0 1 26460
box -48 -56 1008 834
use sg13g2_nand3_1  _1938_
timestamp 1747537721
transform 1 0 8352 0 -1 26460
box -48 -56 528 834
use sg13g2_o21ai_1  _1939_
timestamp 1747537721
transform -1 0 21024 0 -1 26460
box -48 -56 538 834
use sg13g2_mux2_1  _1940_
timestamp 1747537721
transform 1 0 20160 0 1 24948
box -48 -56 1008 834
use sg13g2_nor2_1  _1941_
timestamp 1747537721
transform -1 0 26688 0 1 11340
box -48 -56 432 834
use sg13g2_nand4_1  _1942_
timestamp 1747537721
transform 1 0 26016 0 -1 12852
box -48 -56 624 834
use sg13g2_nor4_1  _1943_
timestamp 1747537721
transform 1 0 25728 0 -1 14364
box -48 -56 624 834
use sg13g2_nand2_2  _1944_
timestamp 1747537721
transform 1 0 22464 0 1 17388
box -48 -56 624 834
use sg13g2_nand3_1  _1945_
timestamp 1747537721
transform 1 0 25248 0 1 11340
box -48 -56 528 834
use sg13g2_nor2_1  _1946_
timestamp 1747537721
transform -1 0 26016 0 -1 12852
box -48 -56 432 834
use sg13g2_nand2_1  _1947_
timestamp 1747537721
transform -1 0 26016 0 1 12852
box -48 -56 432 834
use sg13g2_nor2_1  _1948_
timestamp 1747537721
transform -1 0 27072 0 1 15876
box -48 -56 432 834
use sg13g2_and2_1  _1949_
timestamp 1747537721
transform 1 0 25824 0 1 11340
box -48 -56 528 834
use sg13g2_nor4_1  _1950_
timestamp 1747537721
transform 1 0 26592 0 -1 14364
box -48 -56 624 834
use sg13g2_a21oi_1  _1951_
timestamp 1747537721
transform -1 0 27552 0 -1 15876
box -48 -56 528 834
use sg13g2_nor4_1  _1952_
timestamp 1747537721
transform -1 0 27456 0 1 12852
box -48 -56 624 834
use sg13g2_a21oi_1  _1953_
timestamp 1747537721
transform 1 0 26592 0 -1 15876
box -48 -56 528 834
use sg13g2_a22oi_1  _1954_
timestamp 1747537721
transform 1 0 26016 0 -1 15876
box -48 -56 624 834
use sg13g2_nor2_1  _1955_
timestamp 1747537721
transform -1 0 28320 0 1 15876
box -48 -56 432 834
use sg13g2_nand2b_1  _1956_
timestamp 1747537721
transform -1 0 26688 0 1 15876
box -48 -56 528 834
use sg13g2_a21oi_1  _1957_
timestamp 1747537721
transform -1 0 26208 0 1 15876
box -48 -56 528 834
use sg13g2_nor2_2  _1958_
timestamp 1747537721
transform 1 0 24192 0 -1 18900
box -48 -56 624 834
use sg13g2_o21ai_1  _1959_
timestamp 1747537721
transform -1 0 24288 0 1 24948
box -48 -56 538 834
use sg13g2_a21oi_1  _1960_
timestamp 1747537721
transform 1 0 23808 0 -1 26460
box -48 -56 528 834
use sg13g2_a21oi_1  _1961_
timestamp 1747537721
transform 1 0 26784 0 1 26460
box -48 -56 528 834
use sg13g2_and3_1  _1962_
timestamp 1747537721
transform -1 0 26304 0 1 26460
box -48 -56 720 834
use sg13g2_nor3_1  _1963_
timestamp 1747537721
transform 1 0 24960 0 -1 27972
box -48 -56 528 834
use sg13g2_nand2b_1  _1964_
timestamp 1747537721
transform 1 0 24576 0 -1 21924
box -48 -56 528 834
use sg13g2_nand2_1  _1965_
timestamp 1747537721
transform -1 0 26688 0 -1 24948
box -48 -56 432 834
use sg13g2_nand3_1  _1966_
timestamp 1747537721
transform 1 0 27168 0 -1 26460
box -48 -56 528 834
use sg13g2_xnor2_1  _1967_
timestamp 1747537721
transform 1 0 28128 0 1 26460
box -48 -56 816 834
use sg13g2_nor2_1  _1968_
timestamp 1747537721
transform -1 0 30720 0 -1 26460
box -48 -56 432 834
use sg13g2_nand2_1  _1969_
timestamp 1747537721
transform 1 0 27840 0 -1 24948
box -48 -56 432 834
use sg13g2_nand2_2  _1970_
timestamp 1747537721
transform 1 0 24288 0 1 21924
box -48 -56 624 834
use sg13g2_inv_1  _1971_
timestamp 1747537721
transform -1 0 28896 0 -1 18900
box -48 -56 336 834
use sg13g2_nor2_1  _1972_
timestamp 1747537721
transform 1 0 28128 0 -1 26460
box -48 -56 432 834
use sg13g2_xnor2_1  _1973_
timestamp 1747537721
transform 1 0 27552 0 1 24948
box -48 -56 816 834
use sg13g2_o21ai_1  _1974_
timestamp 1747537721
transform 1 0 28416 0 1 24948
box -48 -56 538 834
use sg13g2_a21oi_1  _1975_
timestamp 1747537721
transform -1 0 28800 0 1 23436
box -48 -56 528 834
use sg13g2_and3_1  _1976_
timestamp 1747537721
transform 1 0 27648 0 1 23436
box -48 -56 720 834
use sg13g2_nand2_1  _1977_
timestamp 1747537721
transform 1 0 28224 0 -1 24948
box -48 -56 432 834
use sg13g2_nor3_1  _1978_
timestamp 1747537721
transform 1 0 27168 0 1 23436
box -48 -56 528 834
use sg13g2_nand2_1  _1979_
timestamp 1747537721
transform -1 0 31392 0 1 21924
box -48 -56 432 834
use sg13g2_xnor2_1  _1980_
timestamp 1747537721
transform 1 0 27936 0 1 21924
box -48 -56 816 834
use sg13g2_o21ai_1  _1981_
timestamp 1747537721
transform 1 0 30528 0 1 21924
box -48 -56 538 834
use sg13g2_a21oi_1  _1982_
timestamp 1747537721
transform 1 0 29760 0 -1 21924
box -48 -56 528 834
use sg13g2_nor2b_1  _1983_
timestamp 1747537721
transform -1 0 28608 0 1 20412
box -54 -56 528 834
use sg13g2_nor2_1  _1984_
timestamp 1747537721
transform 1 0 27072 0 -1 21924
box -48 -56 432 834
use sg13g2_nor3_1  _1985_
timestamp 1747537721
transform 1 0 28224 0 -1 21924
box -48 -56 528 834
use sg13g2_xnor2_1  _1986_
timestamp 1747537721
transform 1 0 27936 0 -1 20412
box -48 -56 816 834
use sg13g2_nor2_1  _1987_
timestamp 1747537721
transform -1 0 31296 0 -1 20412
box -48 -56 432 834
use sg13g2_nand2_1  _1988_
timestamp 1747537721
transform -1 0 28128 0 1 20412
box -48 -56 432 834
use sg13g2_a22oi_1  _1989_
timestamp 1747537721
transform -1 0 28608 0 -1 18900
box -48 -56 624 834
use sg13g2_a21oi_1  _1990_
timestamp 1747537721
transform -1 0 28704 0 1 18900
box -48 -56 528 834
use sg13g2_nor2_1  _1991_
timestamp 1747537721
transform 1 0 28320 0 1 17388
box -48 -56 432 834
use sg13g2_nand2_1  _1992_
timestamp 1747537721
transform -1 0 27936 0 1 17388
box -48 -56 432 834
use sg13g2_xnor2_1  _1993_
timestamp 1747537721
transform 1 0 25632 0 1 18900
box -48 -56 816 834
use sg13g2_o21ai_1  _1994_
timestamp 1747537721
transform 1 0 27264 0 -1 20412
box -48 -56 538 834
use sg13g2_o21ai_1  _1995_
timestamp 1747537721
transform 1 0 24960 0 1 23436
box -48 -56 538 834
use sg13g2_nor3_1  _1996_
timestamp 1747537721
transform -1 0 25248 0 1 24948
box -48 -56 528 834
use sg13g2_nand3_1  _1997_
timestamp 1747537721
transform -1 0 24768 0 1 24948
box -48 -56 528 834
use sg13g2_nor2_1  _1998_
timestamp 1747537721
transform 1 0 24384 0 -1 23436
box -48 -56 432 834
use sg13g2_nor4_1  _1999_
timestamp 1747537721
transform 1 0 25248 0 1 24948
box -48 -56 624 834
use sg13g2_nor2_1  _2000_
timestamp 1747537721
transform 1 0 25920 0 -1 26460
box -48 -56 432 834
use sg13g2_nand4_1  _2001_
timestamp 1747537721
transform -1 0 26304 0 -1 24948
box -48 -56 624 834
use sg13g2_a21oi_1  _2002_
timestamp 1747537721
transform 1 0 25056 0 -1 24948
box -48 -56 528 834
use sg13g2_a22oi_1  _2003_
timestamp 1747537721
transform 1 0 24288 0 -1 24948
box -48 -56 624 834
use sg13g2_nor2_1  _2004_
timestamp 1747537721
transform 1 0 23424 0 -1 23436
box -48 -56 432 834
use sg13g2_nand2b_1  _2005_
timestamp 1747537721
transform 1 0 25440 0 1 23436
box -48 -56 528 834
use sg13g2_a21oi_1  _2006_
timestamp 1747537721
transform 1 0 24000 0 1 23436
box -48 -56 528 834
use sg13g2_nor2_1  _2007_
timestamp 1747537721
transform 1 0 5280 0 1 24948
box -48 -56 432 834
use sg13g2_nor2_1  _2008_
timestamp 1747537721
transform -1 0 6144 0 1 21924
box -48 -56 432 834
use sg13g2_a21oi_1  _2009_
timestamp 1747537721
transform -1 0 4704 0 1 21924
box -48 -56 528 834
use sg13g2_o21ai_1  _2010_
timestamp 1747537721
transform -1 0 5472 0 -1 23436
box -48 -56 538 834
use sg13g2_nand2_1  _2011_
timestamp 1747537721
transform 1 0 8448 0 1 23436
box -48 -56 432 834
use sg13g2_o21ai_1  _2012_
timestamp 1747537721
transform 1 0 8352 0 1 21924
box -48 -56 538 834
use sg13g2_nand2_1  _2013_
timestamp 1747537721
transform 1 0 12096 0 1 23436
box -48 -56 432 834
use sg13g2_o21ai_1  _2014_
timestamp 1747537721
transform 1 0 11424 0 -1 24948
box -48 -56 538 834
use sg13g2_mux2_1  _2015_
timestamp 1747537721
transform 1 0 2112 0 -1 20412
box -48 -56 1008 834
use sg13g2_mux2_1  _2016_
timestamp 1747537721
transform -1 0 4032 0 1 23436
box -48 -56 1008 834
use sg13g2_mux2_1  _2017_
timestamp 1747537721
transform 1 0 12384 0 1 20412
box -48 -56 1008 834
use sg13g2_o21ai_1  _2018_
timestamp 1747537721
transform 1 0 20832 0 1 20412
box -48 -56 538 834
use sg13g2_dfrbp_1  _2019_
timestamp 1747537721
transform -1 0 3648 0 1 24948
box -60 -56 2556 834
use sg13g2_tiehi  _2019__26
timestamp 1747537721
transform -1 0 3360 0 -1 24948
box -48 -56 432 834
use sg13g2_dfrbp_1  _2020_
timestamp 1747537721
transform 1 0 5664 0 -1 27972
box -60 -56 2556 834
use sg13g2_tiehi  _2020__18
timestamp 1747537721
transform -1 0 7008 0 1 26460
box -48 -56 432 834
use sg13g2_tiehi  _2021__58
timestamp 1747537721
transform -1 0 7200 0 1 24948
box -48 -56 432 834
use sg13g2_dfrbp_1  _2021_
timestamp 1747537721
transform 1 0 5760 0 -1 24948
box -60 -56 2556 834
use sg13g2_tiehi  _2022__57
timestamp 1747537721
transform 1 0 2496 0 1 26460
box -48 -56 432 834
use sg13g2_dfrbp_1  _2022_
timestamp 1747537721
transform -1 0 4128 0 -1 26460
box -60 -56 2556 834
use sg13g2_dfrbp_1  _2023_
timestamp 1747537721
transform 1 0 8160 0 -1 27972
box -60 -56 2556 834
use sg13g2_tiehi  _2023__56
timestamp 1747537721
transform -1 0 9600 0 1 26460
box -48 -56 432 834
use sg13g2_tiehi  _2024__55
timestamp 1747537721
transform -1 0 30912 0 -1 17388
box -48 -56 432 834
use sg13g2_dfrbp_1  _2024_
timestamp 1747537721
transform -1 0 31392 0 1 15876
box -60 -56 2556 834
use sg13g2_dfrbp_1  _2025_
timestamp 1747537721
transform 1 0 24288 0 -1 11340
box -60 -56 2556 834
use sg13g2_tiehi  _2025__54
timestamp 1747537721
transform -1 0 25728 0 1 9828
box -48 -56 432 834
use sg13g2_dfrbp_1  _2026_
timestamp 1747537721
transform -1 0 22944 0 -1 9828
box -60 -56 2556 834
use sg13g2_tiehi  _2026__53
timestamp 1747537721
transform 1 0 21504 0 1 8316
box -48 -56 432 834
use sg13g2_dfrbp_1  _2027_
timestamp 1747537721
transform 1 0 23040 0 -1 8316
box -60 -56 2556 834
use sg13g2_tiehi  _2027__52
timestamp 1747537721
transform -1 0 24960 0 1 6804
box -48 -56 432 834
use sg13g2_dfrbp_1  _2028_
timestamp 1747537721
transform -1 0 31392 0 -1 9828
box -60 -56 2556 834
use sg13g2_tiehi  _2028__51
timestamp 1747537721
transform -1 0 31392 0 -1 8316
box -48 -56 432 834
use sg13g2_tiehi  _2029__50
timestamp 1747537721
transform -1 0 26880 0 1 8316
box -48 -56 432 834
use sg13g2_dfrbp_1  _2029_
timestamp 1747537721
transform 1 0 25536 0 -1 8316
box -60 -56 2556 834
use sg13g2_dfrbp_1  _2030_
timestamp 1747537721
transform -1 0 31392 0 -1 11340
box -60 -56 2556 834
use sg13g2_tiehi  _2030__49
timestamp 1747537721
transform -1 0 31392 0 1 8316
box -48 -56 432 834
use sg13g2_tiehi  _2031__48
timestamp 1747537721
transform 1 0 29664 0 1 12852
box -48 -56 432 834
use sg13g2_dfrbp_1  _2031_
timestamp 1747537721
transform -1 0 31104 0 -1 12852
box -60 -56 2556 834
use sg13g2_tiehi  _2032__47
timestamp 1747537721
transform -1 0 31392 0 1 14364
box -48 -56 432 834
use sg13g2_dfrbp_1  _2032_
timestamp 1747537721
transform -1 0 31392 0 -1 14364
box -60 -56 2556 834
use sg13g2_tiehi  _2033__46
timestamp 1747537721
transform 1 0 30144 0 -1 17388
box -48 -56 432 834
use sg13g2_dfrbp_1  _2033_
timestamp 1747537721
transform -1 0 31392 0 -1 15876
box -60 -56 2556 834
use sg13g2_tiehi  _2034__45
timestamp 1747537721
transform -1 0 6816 0 1 21924
box -48 -56 432 834
use sg13g2_dfrbp_1  _2034_
timestamp 1747537721
transform 1 0 5376 0 -1 21924
box -60 -56 2556 834
use sg13g2_tiehi  _2035__43
timestamp 1747537721
transform 1 0 576 0 -1 14364
box -48 -56 432 834
use sg13g2_dfrbp_1  _2035_
timestamp 1747537721
transform 1 0 576 0 1 12852
box -60 -56 2556 834
use sg13g2_tiehi  _2036__41
timestamp 1747537721
transform -1 0 2208 0 -1 12852
box -48 -56 432 834
use sg13g2_dfrbp_1  _2036_
timestamp 1747537721
transform 1 0 864 0 1 11340
box -60 -56 2556 834
use sg13g2_dfrbp_1  _2037_
timestamp 1747537721
transform 1 0 1344 0 -1 3780
box -60 -56 2556 834
use sg13g2_tiehi  _2037__39
timestamp 1747537721
transform -1 0 2784 0 1 2268
box -48 -56 432 834
use sg13g2_dfrbp_1  _2038_
timestamp 1747537721
transform 1 0 1536 0 -1 2268
box -60 -56 2556 834
use sg13g2_tiehi  _2038__37
timestamp 1747537721
transform -1 0 2976 0 1 756
box -48 -56 432 834
use sg13g2_dfrbp_1  _2039_
timestamp 1747537721
transform 1 0 6432 0 1 756
box -60 -56 2556 834
use sg13g2_tiehi  _2039__35
timestamp 1747537721
transform -1 0 7872 0 -1 2268
box -48 -56 432 834
use sg13g2_tiehi  _2040__33
timestamp 1747537721
transform -1 0 17088 0 -1 2268
box -48 -56 432 834
use sg13g2_dfrbp_1  _2040_
timestamp 1747537721
transform 1 0 15648 0 1 756
box -60 -56 2556 834
use sg13g2_dfrbp_1  _2041_
timestamp 1747537721
transform 1 0 19104 0 -1 2268
box -60 -56 2556 834
use sg13g2_tiehi  _2041__31
timestamp 1747537721
transform -1 0 21216 0 1 756
box -48 -56 432 834
use sg13g2_dfrbp_1  _2042_
timestamp 1747537721
transform 1 0 22656 0 1 756
box -60 -56 2556 834
use sg13g2_tiehi  _2042__29
timestamp 1747537721
transform -1 0 24096 0 -1 2268
box -48 -56 432 834
use sg13g2_tiehi  _2043__27
timestamp 1747537721
transform -1 0 27168 0 1 2268
box -48 -56 432 834
use sg13g2_dfrbp_1  _2043_
timestamp 1747537721
transform 1 0 25728 0 -1 2268
box -60 -56 2556 834
use sg13g2_tiehi  _2044__25
timestamp 1747537721
transform 1 0 29952 0 1 3780
box -48 -56 432 834
use sg13g2_dfrbp_1  _2044_
timestamp 1747537721
transform -1 0 31392 0 -1 3780
box -60 -56 2556 834
use sg13g2_tiehi  _2045__23
timestamp 1747537721
transform -1 0 30624 0 1 2268
box -48 -56 432 834
use sg13g2_dfrbp_1  _2045_
timestamp 1747537721
transform -1 0 30912 0 1 756
box -60 -56 2556 834
use sg13g2_dfrbp_1  _2046_
timestamp 1747537721
transform 1 0 11136 0 -1 27972
box -60 -56 2556 834
use sg13g2_tiehi  _2046__21
timestamp 1747537721
transform -1 0 14016 0 -1 27972
box -48 -56 432 834
use sg13g2_dfrbp_1  _2047_
timestamp 1747537721
transform -1 0 16896 0 -1 27972
box -60 -56 2556 834
use sg13g2_tiehi  _2047__20
timestamp 1747537721
transform 1 0 15456 0 1 26460
box -48 -56 432 834
use sg13g2_tiehi  _2048__19
timestamp 1747537721
transform -1 0 14016 0 1 26460
box -48 -56 432 834
use sg13g2_dfrbp_1  _2048_
timestamp 1747537721
transform 1 0 12768 0 -1 26460
box -60 -56 2556 834
use sg13g2_tiehi  _2049__17
timestamp 1747537721
transform -1 0 21120 0 -1 27972
box -48 -56 432 834
use sg13g2_dfrbp_1  _2049_
timestamp 1747537721
transform 1 0 19680 0 1 26460
box -60 -56 2556 834
use sg13g2_tiehi  _2050__73
timestamp 1747537721
transform -1 0 14976 0 1 24948
box -48 -56 432 834
use sg13g2_dfrbp_1  _2050_
timestamp 1747537721
transform 1 0 13152 0 -1 23436
box -60 -56 2556 834
use sg13g2_tiehi  _2051__72
timestamp 1747537721
transform -1 0 17472 0 -1 24948
box -48 -56 432 834
use sg13g2_dfrbp_1  _2051_
timestamp 1747537721
transform 1 0 15360 0 1 23436
box -60 -56 2556 834
use sg13g2_tiehi  _2052__71
timestamp 1747537721
transform -1 0 20544 0 -1 27972
box -48 -56 432 834
use sg13g2_dfrbp_1  _2052_
timestamp 1747537721
transform 1 0 17664 0 -1 27972
box -60 -56 2556 834
use sg13g2_tiehi  _2053__70
timestamp 1747537721
transform -1 0 22560 0 -1 26460
box -48 -56 432 834
use sg13g2_dfrbp_1  _2053_
timestamp 1747537721
transform 1 0 21120 0 1 24948
box -60 -56 2556 834
use sg13g2_dfrbp_1  _2054_
timestamp 1747537721
transform -1 0 29088 0 -1 17388
box -60 -56 2556 834
use sg13g2_tiehi  _2054__69
timestamp 1747537721
transform -1 0 28704 0 1 15876
box -48 -56 432 834
use sg13g2_dfrbp_1  _2055_
timestamp 1747537721
transform 1 0 22272 0 -1 27972
box -60 -56 2556 834
use sg13g2_tiehi  _2055__68
timestamp 1747537721
transform -1 0 24768 0 1 26460
box -48 -56 432 834
use sg13g2_dfrbp_1  _2056_
timestamp 1747537721
transform 1 0 25440 0 -1 27972
box -60 -56 2556 834
use sg13g2_tiehi  _2056__66
timestamp 1747537721
transform -1 0 28128 0 1 26460
box -48 -56 432 834
use sg13g2_tiehi  _2057__64
timestamp 1747537721
transform -1 0 31392 0 -1 27972
box -48 -56 432 834
use sg13g2_dfrbp_1  _2057_
timestamp 1747537721
transform -1 0 31392 0 1 26460
box -60 -56 2556 834
use sg13g2_tiehi  _2058__62
timestamp 1747537721
transform -1 0 30624 0 -1 27972
box -48 -56 432 834
use sg13g2_dfrbp_1  _2058_
timestamp 1747537721
transform 1 0 28896 0 1 24948
box -60 -56 2556 834
use sg13g2_tiehi  _2059__60
timestamp 1747537721
transform -1 0 30336 0 -1 26460
box -48 -56 432 834
use sg13g2_dfrbp_1  _2059_
timestamp 1747537721
transform 1 0 28896 0 1 23436
box -60 -56 2556 834
use sg13g2_tiehi  _2060__44
timestamp 1747537721
transform 1 0 29664 0 -1 24948
box -48 -56 432 834
use sg13g2_dfrbp_1  _2060_
timestamp 1747537721
transform 1 0 28896 0 -1 23436
box -60 -56 2556 834
use sg13g2_tiehi  _2061__40
timestamp 1747537721
transform -1 0 31296 0 -1 24948
box -48 -56 432 834
use sg13g2_dfrbp_1  _2061_
timestamp 1747537721
transform 1 0 28896 0 1 20412
box -60 -56 2556 834
use sg13g2_dfrbp_1  _2062_
timestamp 1747537721
transform -1 0 31392 0 1 18900
box -60 -56 2556 834
use sg13g2_tiehi  _2062__36
timestamp 1747537721
transform 1 0 29568 0 1 17388
box -48 -56 432 834
use sg13g2_dfrbp_1  _2063_
timestamp 1747537721
transform -1 0 31392 0 -1 18900
box -60 -56 2556 834
use sg13g2_tiehi  _2063__32
timestamp 1747537721
transform -1 0 31200 0 1 17388
box -48 -56 432 834
use sg13g2_tiehi  _2064__28
timestamp 1747537721
transform 1 0 26016 0 -1 20412
box -48 -56 432 834
use sg13g2_dfrbp_1  _2064_
timestamp 1747537721
transform -1 0 27456 0 -1 18900
box -60 -56 2556 834
use sg13g2_tiehi  _2065__24
timestamp 1747537721
transform -1 0 23328 0 -1 24948
box -48 -56 432 834
use sg13g2_dfrbp_1  _2065_
timestamp 1747537721
transform -1 0 23232 0 1 23436
box -60 -56 2556 834
use sg13g2_tiehi  _2066__22
timestamp 1747537721
transform 1 0 5184 0 1 26460
box -48 -56 432 834
use sg13g2_dfrbp_1  _2066_
timestamp 1747537721
transform 1 0 5568 0 -1 26460
box -60 -56 2556 834
use sg13g2_dfrbp_1  _2067_
timestamp 1747537721
transform 1 0 3168 0 -1 27972
box -60 -56 2556 834
use sg13g2_tiehi  _2067__67
timestamp 1747537721
transform 1 0 3264 0 1 26460
box -48 -56 432 834
use sg13g2_tiehi  _2068__65
timestamp 1747537721
transform 1 0 1824 0 -1 23436
box -48 -56 432 834
use sg13g2_dfrbp_1  _2068_
timestamp 1747537721
transform -1 0 3264 0 1 21924
box -60 -56 2556 834
use sg13g2_tiehi  _2069__63
timestamp 1747537721
transform -1 0 7392 0 1 23436
box -48 -56 432 834
use sg13g2_dfrbp_1  _2069_
timestamp 1747537721
transform 1 0 5472 0 -1 23436
box -60 -56 2556 834
use sg13g2_tiehi  _2070__61
timestamp 1747537721
transform 1 0 8832 0 1 23436
box -48 -56 432 834
use sg13g2_dfrbp_1  _2070_
timestamp 1747537721
transform 1 0 8352 0 -1 23436
box -60 -56 2556 834
use sg13g2_tiehi  _2071__59
timestamp 1747537721
transform -1 0 13344 0 1 24948
box -48 -56 432 834
use sg13g2_dfrbp_1  _2071_
timestamp 1747537721
transform 1 0 11904 0 -1 24948
box -60 -56 2556 834
use sg13g2_dfrbp_1  _2072_
timestamp 1747537721
transform -1 0 3072 0 1 20412
box -60 -56 2556 834
use sg13g2_tiehi  _2072__42
timestamp 1747537721
transform -1 0 2880 0 -1 21924
box -48 -56 432 834
use sg13g2_tiehi  _2073__38
timestamp 1747537721
transform 1 0 1632 0 -1 24948
box -48 -56 432 834
use sg13g2_dfrbp_1  _2073_
timestamp 1747537721
transform -1 0 3072 0 1 23436
box -60 -56 2556 834
use sg13g2_tiehi  _2074__34
timestamp 1747537721
transform -1 0 14784 0 -1 21924
box -48 -56 432 834
use sg13g2_dfrbp_1  _2074_
timestamp 1747537721
transform 1 0 13344 0 1 20412
box -60 -56 2556 834
use sg13g2_tiehi  _2075__30
timestamp 1747537721
transform -1 0 22752 0 -1 21924
box -48 -56 432 834
use sg13g2_dfrbp_1  _2075_
timestamp 1747537721
transform 1 0 21312 0 1 20412
box -60 -56 2556 834
use sg13g2_buf_2  _2141_
timestamp 1747537721
transform -1 0 18432 0 1 20412
box -48 -56 528 834
use sg13g2_buf_2  _2142_
timestamp 1747537721
transform -1 0 21984 0 1 18900
box -48 -56 528 834
use sg13g2_buf_2  _2143_
timestamp 1747537721
transform -1 0 18432 0 -1 21924
box -48 -56 528 834
use sg13g2_buf_2  _2144_
timestamp 1747537721
transform -1 0 21696 0 -1 20412
box -48 -56 528 834
use sg13g2_buf_1  _2145_
timestamp 1747537721
transform -1 0 16416 0 -1 21924
box -48 -56 432 834
use sg13g2_buf_1  _2146_
timestamp 1747537721
transform -1 0 21984 0 -1 18900
box -48 -56 432 834
use sg13g2_buf_2  clkbuf_0_clk
timestamp 1747537721
transform 1 0 15840 0 1 14364
box -48 -56 528 834
use sg13g2_buf_2  clkbuf_4_0_0_clk
timestamp 1747537721
transform 1 0 3168 0 -1 15876
box -48 -56 528 834
use sg13g2_buf_2  clkbuf_4_1_0_clk
timestamp 1747537721
transform 1 0 2784 0 1 17388
box -48 -56 528 834
use sg13g2_buf_2  clkbuf_4_2_0_clk
timestamp 1747537721
transform 1 0 8352 0 1 15876
box -48 -56 528 834
use sg13g2_buf_2  clkbuf_4_3_0_clk
timestamp 1747537721
transform 1 0 7968 0 -1 18900
box -48 -56 528 834
use sg13g2_buf_2  clkbuf_4_4_0_clk
timestamp 1747537721
transform -1 0 8736 0 1 26460
box -48 -56 528 834
use sg13g2_buf_2  clkbuf_4_5_0_clk
timestamp 1747537721
transform 1 0 11712 0 -1 26460
box -48 -56 528 834
use sg13g2_buf_2  clkbuf_4_6_0_clk
timestamp 1747537721
transform 1 0 16320 0 -1 23436
box -48 -56 528 834
use sg13g2_buf_2  clkbuf_4_7_0_clk
timestamp 1747537721
transform 1 0 16608 0 -1 24948
box -48 -56 528 834
use sg13g2_buf_2  clkbuf_4_8_0_clk
timestamp 1747537721
transform -1 0 24192 0 1 6804
box -48 -56 528 834
use sg13g2_buf_2  clkbuf_4_9_0_clk
timestamp 1747537721
transform 1 0 24000 0 -1 9828
box -48 -56 528 834
use sg13g2_buf_2  clkbuf_4_10_0_clk
timestamp 1747537721
transform -1 0 31008 0 1 8316
box -48 -56 528 834
use sg13g2_buf_2  clkbuf_4_11_0_clk
timestamp 1747537721
transform -1 0 31296 0 1 9828
box -48 -56 528 834
use sg13g2_buf_2  clkbuf_4_12_0_clk
timestamp 1747537721
transform 1 0 27552 0 -1 23436
box -48 -56 528 834
use sg13g2_buf_2  clkbuf_4_13_0_clk
timestamp 1747537721
transform -1 0 24960 0 1 23436
box -48 -56 528 834
use sg13g2_buf_2  clkbuf_4_14_0_clk
timestamp 1747537721
transform -1 0 30912 0 -1 20412
box -48 -56 528 834
use sg13g2_buf_2  clkbuf_4_15_0_clk
timestamp 1747537721
transform -1 0 30720 0 -1 21924
box -48 -56 528 834
use sg13g2_inv_1  clkload0
timestamp 1747537721
transform 1 0 8448 0 -1 18900
box -48 -56 336 834
use sg13g2_inv_1  clkload1
timestamp 1747537721
transform 1 0 11904 0 1 24948
box -48 -56 336 834
use sg13g2_inv_1  clkload2
timestamp 1747537721
transform -1 0 18816 0 -1 24948
box -48 -56 336 834
use sg13g2_inv_1  clkload3
timestamp 1747537721
transform 1 0 24768 0 1 8316
box -48 -56 336 834
use sg13g2_inv_1  clkload4
timestamp 1747537721
transform 1 0 30048 0 1 12852
box -48 -56 336 834
use sg13g2_inv_1  clkload5
timestamp 1747537721
transform 1 0 25824 0 1 24948
box -48 -56 336 834
use sg13g2_inv_1  clkload6
timestamp 1747537721
transform -1 0 28224 0 -1 21924
box -48 -56 336 834
use sg13g2_tielo  controller_11
timestamp 1747537721
transform -1 0 9120 0 1 26460
box -48 -56 432 834
use sg13g2_tielo  controller_12
timestamp 1747537721
transform 1 0 7008 0 1 26460
box -48 -56 432 834
use sg13g2_tielo  controller_13
timestamp 1747537721
transform -1 0 7584 0 1 24948
box -48 -56 432 834
use sg13g2_tielo  controller_14
timestamp 1747537721
transform 1 0 4800 0 1 26460
box -48 -56 432 834
use sg13g2_tielo  controller_15
timestamp 1747537721
transform 1 0 4416 0 1 26460
box -48 -56 432 834
use sg13g2_tielo  controller_16
timestamp 1747537721
transform 1 0 4032 0 1 26460
box -48 -56 432 834
use sg13g2_tiehi  controller_74
timestamp 1747537721
transform 1 0 2880 0 1 26460
box -48 -56 432 834
use sg13g2_tiehi  controller_75
timestamp 1747537721
transform 1 0 2784 0 -1 27972
box -48 -56 432 834
use sg13g2_buf_2  fanout319
timestamp 1747537721
transform 1 0 14304 0 1 23436
box -48 -56 528 834
use sg13g2_buf_2  fanout320
timestamp 1747537721
transform -1 0 15360 0 -1 24948
box -48 -56 528 834
use sg13g2_buf_4  fanout321
timestamp 1747537721
transform -1 0 20928 0 -1 6804
box -48 -56 816 834
use sg13g2_buf_2  fanout322
timestamp 1747537721
transform -1 0 20736 0 1 9828
box -48 -56 528 834
use sg13g2_buf_4  fanout323
timestamp 1747537721
transform 1 0 21984 0 -1 17388
box -48 -56 816 834
use sg13g2_buf_2  fanout324
timestamp 1747537721
transform -1 0 23232 0 -1 17388
box -48 -56 528 834
use sg13g2_buf_4  fanout325
timestamp 1747537721
transform 1 0 18528 0 -1 6804
box -48 -56 816 834
use sg13g2_buf_2  fanout326
timestamp 1747537721
transform 1 0 18624 0 -1 9828
box -48 -56 528 834
use sg13g2_buf_2  fanout327
timestamp 1747537721
transform 1 0 10656 0 1 5292
box -48 -56 528 834
use sg13g2_buf_4  fanout328
timestamp 1747537721
transform 1 0 16800 0 -1 23436
box -48 -56 816 834
use sg13g2_buf_2  fanout329
timestamp 1747537721
transform 1 0 13344 0 1 15876
box -48 -56 528 834
use sg13g2_buf_4  fanout330
timestamp 1747537721
transform 1 0 19296 0 -1 17388
box -48 -56 816 834
use sg13g2_buf_2  fanout331
timestamp 1747537721
transform 1 0 19104 0 1 15876
box -48 -56 528 834
use sg13g2_buf_4  fanout332
timestamp 1747537721
transform 1 0 5472 0 1 8316
box -48 -56 816 834
use sg13g2_buf_2  fanout333
timestamp 1747537721
transform -1 0 18048 0 -1 23436
box -48 -56 528 834
use sg13g2_buf_2  fanout334
timestamp 1747537721
transform 1 0 4416 0 -1 18900
box -48 -56 528 834
use sg13g2_buf_1  fanout335
timestamp 1747537721
transform -1 0 3936 0 -1 18900
box -48 -56 432 834
use sg13g2_buf_2  fanout336
timestamp 1747537721
transform -1 0 9696 0 1 18900
box -48 -56 528 834
use sg13g2_buf_1  fanout337
timestamp 1747537721
transform -1 0 9600 0 -1 18900
box -48 -56 432 834
use sg13g2_buf_2  fanout338
timestamp 1747537721
transform -1 0 18912 0 -1 20412
box -48 -56 528 834
use sg13g2_buf_2  fanout339
timestamp 1747537721
transform 1 0 3168 0 -1 20412
box -48 -56 528 834
use sg13g2_buf_1  fanout340
timestamp 1747537721
transform -1 0 4512 0 1 18900
box -48 -56 432 834
use sg13g2_buf_4  fanout341
timestamp 1747537721
transform 1 0 4128 0 1 20412
box -48 -56 816 834
use sg13g2_buf_1  fanout342
timestamp 1747537721
transform 1 0 8928 0 1 20412
box -48 -56 432 834
use sg13g2_buf_1  fanout343
timestamp 1747537721
transform -1 0 12480 0 -1 21924
box -48 -56 432 834
use sg13g2_buf_4  fanout344
timestamp 1747537721
transform -1 0 16704 0 1 21924
box -48 -56 816 834
use sg13g2_buf_4  fanout345
timestamp 1747537721
transform -1 0 12384 0 1 11340
box -48 -56 816 834
use sg13g2_buf_1  fanout346
timestamp 1747537721
transform 1 0 12288 0 -1 11340
box -48 -56 432 834
use sg13g2_buf_4  fanout347
timestamp 1747537721
transform 1 0 6432 0 -1 17388
box -48 -56 816 834
use sg13g2_buf_2  fanout348
timestamp 1747537721
transform -1 0 16224 0 -1 9828
box -48 -56 528 834
use sg13g2_buf_2  fanout349
timestamp 1747537721
transform 1 0 14400 0 1 17388
box -48 -56 528 834
use sg13g2_buf_2  fanout350
timestamp 1747537721
transform -1 0 15168 0 -1 9828
box -48 -56 528 834
use sg13g2_buf_2  fanout351
timestamp 1747537721
transform 1 0 14208 0 1 9828
box -48 -56 528 834
use sg13g2_buf_2  fanout352
timestamp 1747537721
transform -1 0 14688 0 -1 9828
box -48 -56 528 834
use sg13g2_buf_4  fanout353
timestamp 1747537721
transform 1 0 14304 0 1 15876
box -48 -56 816 834
use sg13g2_buf_2  fanout354
timestamp 1747537721
transform 1 0 5184 0 1 15876
box -48 -56 528 834
use sg13g2_buf_2  fanout355
timestamp 1747537721
transform 1 0 11520 0 1 15876
box -48 -56 528 834
use sg13g2_buf_2  fanout356
timestamp 1747537721
transform -1 0 17760 0 -1 18900
box -48 -56 528 834
use sg13g2_buf_2  fanout357
timestamp 1747537721
transform 1 0 12288 0 -1 18900
box -48 -56 528 834
use sg13g2_buf_2  fanout358
timestamp 1747537721
transform -1 0 15456 0 1 8316
box -48 -56 528 834
use sg13g2_buf_2  fanout359
timestamp 1747537721
transform -1 0 15648 0 -1 17388
box -48 -56 528 834
use sg13g2_buf_4  fanout360
timestamp 1747537721
transform 1 0 12768 0 -1 18900
box -48 -56 816 834
use sg13g2_buf_4  fanout361
timestamp 1747537721
transform 1 0 9312 0 1 9828
box -48 -56 816 834
use sg13g2_buf_2  fanout362
timestamp 1747537721
transform 1 0 8832 0 1 9828
box -48 -56 528 834
use sg13g2_buf_2  fanout363
timestamp 1747537721
transform 1 0 7872 0 1 17388
box -48 -56 528 834
use sg13g2_buf_2  fanout364
timestamp 1747537721
transform -1 0 9792 0 -1 20412
box -48 -56 528 834
use sg13g2_buf_2  fanout365
timestamp 1747537721
transform 1 0 14496 0 -1 17388
box -48 -56 528 834
use sg13g2_buf_2  fanout366
timestamp 1747537721
transform 1 0 11520 0 1 17388
box -48 -56 528 834
use sg13g2_buf_2  fanout367
timestamp 1747537721
transform 1 0 15168 0 -1 20412
box -48 -56 528 834
use sg13g2_buf_2  fanout368
timestamp 1747537721
transform 1 0 11904 0 1 12852
box -48 -56 528 834
use sg13g2_buf_4  fanout369
timestamp 1747537721
transform 1 0 8640 0 -1 21924
box -48 -56 816 834
use sg13g2_buf_4  fanout370
timestamp 1747537721
transform -1 0 25440 0 1 20412
box -48 -56 816 834
use sg13g2_buf_1  fanout371
timestamp 1747537721
transform 1 0 25056 0 -1 21924
box -48 -56 432 834
use sg13g2_buf_2  fanout372
timestamp 1747537721
transform 1 0 14208 0 1 18900
box -48 -56 528 834
use sg13g2_buf_4  fanout373
timestamp 1747537721
transform -1 0 20256 0 -1 15876
box -48 -56 816 834
use sg13g2_buf_4  fanout374
timestamp 1747537721
transform -1 0 21504 0 -1 15876
box -48 -56 816 834
use sg13g2_buf_2  fanout375
timestamp 1747537721
transform 1 0 10848 0 -1 23436
box -48 -56 528 834
use sg13g2_buf_2  fanout376
timestamp 1747537721
transform 1 0 10848 0 1 14364
box -48 -56 528 834
use sg13g2_buf_1  fanout377
timestamp 1747537721
transform 1 0 11616 0 -1 14364
box -48 -56 432 834
use sg13g2_buf_2  fanout378
timestamp 1747537721
transform 1 0 8736 0 1 11340
box -48 -56 528 834
use sg13g2_buf_4  fanout379
timestamp 1747537721
transform -1 0 4224 0 1 21924
box -48 -56 816 834
use sg13g2_buf_2  fanout380
timestamp 1747537721
transform 1 0 27552 0 -1 18900
box -48 -56 528 834
use sg13g2_buf_2  fanout381
timestamp 1747537721
transform 1 0 30720 0 -1 21924
box -48 -56 528 834
use sg13g2_buf_1  fanout382
timestamp 1747537721
transform -1 0 31104 0 -1 26460
box -48 -56 432 834
use sg13g2_buf_2  fanout383
timestamp 1747537721
transform 1 0 28608 0 -1 26460
box -48 -56 528 834
use sg13g2_buf_2  fanout384
timestamp 1747537721
transform 1 0 27648 0 -1 26460
box -48 -56 528 834
use sg13g2_buf_2  fanout385
timestamp 1747537721
transform -1 0 24384 0 1 26460
box -48 -56 528 834
use sg13g2_buf_2  fanout386
timestamp 1747537721
transform 1 0 23424 0 1 26460
box -48 -56 528 834
use sg13g2_buf_2  fanout387
timestamp 1747537721
transform 1 0 17760 0 -1 3780
box -48 -56 528 834
use sg13g2_buf_2  fanout388
timestamp 1747537721
transform 1 0 21600 0 -1 2268
box -48 -56 528 834
use sg13g2_buf_4  fanout389
timestamp 1747537721
transform -1 0 22080 0 1 756
box -48 -56 816 834
use sg13g2_buf_4  fanout390
timestamp 1747537721
transform -1 0 10752 0 1 756
box -48 -56 816 834
use sg13g2_buf_2  fanout391
timestamp 1747537721
transform -1 0 11808 0 1 756
box -48 -56 528 834
use sg13g2_buf_4  fanout392
timestamp 1747537721
transform 1 0 4896 0 -1 2268
box -48 -56 816 834
use sg13g2_buf_2  fanout393
timestamp 1747537721
transform -1 0 6336 0 1 756
box -48 -56 528 834
use sg13g2_buf_2  fanout394
timestamp 1747537721
transform 1 0 1056 0 1 3780
box -48 -56 528 834
use sg13g2_buf_4  fanout395
timestamp 1747537721
transform -1 0 4128 0 1 2268
box -48 -56 816 834
use sg13g2_buf_2  fanout396
timestamp 1747537721
transform 1 0 3072 0 -1 11340
box -48 -56 528 834
use sg13g2_buf_2  fanout397
timestamp 1747537721
transform 1 0 2112 0 -1 14364
box -48 -56 528 834
use sg13g2_buf_4  fanout398
timestamp 1747537721
transform -1 0 31296 0 1 11340
box -48 -56 816 834
use sg13g2_buf_1  fanout399
timestamp 1747537721
transform -1 0 30912 0 1 12852
box -48 -56 432 834
use sg13g2_buf_2  fanout400
timestamp 1747537721
transform 1 0 28704 0 -1 5292
box -48 -56 528 834
use sg13g2_buf_2  fanout401
timestamp 1747537721
transform -1 0 30816 0 1 9828
box -48 -56 528 834
use sg13g2_buf_4  fanout402
timestamp 1747537721
transform 1 0 28032 0 1 6804
box -48 -56 816 834
use sg13g2_buf_2  fanout403
timestamp 1747537721
transform 1 0 27360 0 1 6804
box -48 -56 528 834
use sg13g2_buf_2  fanout404
timestamp 1747537721
transform 1 0 26976 0 -1 9828
box -48 -56 528 834
use sg13g2_buf_4  fanout405
timestamp 1747537721
transform 1 0 25248 0 -1 9828
box -48 -56 816 834
use sg13g2_buf_4  fanout406
timestamp 1747537721
transform 1 0 13536 0 -1 8316
box -48 -56 816 834
use sg13g2_buf_2  fanout407
timestamp 1747537721
transform -1 0 25440 0 1 6804
box -48 -56 528 834
use sg13g2_buf_4  fanout408
timestamp 1747537721
transform 1 0 22176 0 -1 8316
box -48 -56 816 834
use sg13g2_buf_2  fanout409
timestamp 1747537721
transform 1 0 23040 0 -1 9828
box -48 -56 528 834
use sg13g2_buf_4  fanout410
timestamp 1747537721
transform 1 0 1056 0 1 8316
box -48 -56 816 834
use sg13g2_buf_2  fanout411
timestamp 1747537721
transform 1 0 10272 0 -1 9828
box -48 -56 528 834
use sg13g2_buf_2  fanout412
timestamp 1747537721
transform 1 0 26784 0 -1 11340
box -48 -56 528 834
use sg13g2_buf_4  fanout413
timestamp 1747537721
transform 1 0 24768 0 -1 17388
box -48 -56 816 834
use sg13g2_buf_2  fanout414
timestamp 1747537721
transform 1 0 25536 0 -1 17388
box -48 -56 528 834
use sg13g2_buf_2  fanout415
timestamp 1747537721
transform 1 0 4032 0 1 23436
box -48 -56 528 834
use sg13g2_buf_2  fanout416
timestamp 1747537721
transform 1 0 12384 0 1 21924
box -48 -56 528 834
use sg13g2_buf_2  fanout417
timestamp 1747537721
transform 1 0 10944 0 1 24948
box -48 -56 528 834
use sg13g2_buf_1  fanout418
timestamp 1747537721
transform -1 0 11712 0 -1 23436
box -48 -56 432 834
use sg13g2_buf_4  fanout419
timestamp 1747537721
transform 1 0 14688 0 1 21924
box -48 -56 816 834
use sg13g2_buf_4  fanout420
timestamp 1747537721
transform 1 0 18816 0 -1 21924
box -48 -56 816 834
use sg13g2_buf_2  fanout421
timestamp 1747537721
transform -1 0 20064 0 1 23436
box -48 -56 528 834
use sg13g2_buf_2  fanout422
timestamp 1747537721
transform 1 0 19104 0 1 20412
box -48 -56 528 834
use sg13g2_buf_2  fanout423
timestamp 1747537721
transform -1 0 11904 0 1 24948
box -48 -56 528 834
use sg13g2_buf_4  fanout424
timestamp 1747537721
transform -1 0 21600 0 -1 21924
box -48 -56 816 834
use sg13g2_decap_8  FILLER_0_0
timestamp 1747537721
transform 1 0 576 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_7
timestamp 1747537721
transform 1 0 1248 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_14
timestamp 1747537721
transform 1 0 1920 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_25
timestamp 1747537721
transform 1 0 2976 0 1 756
box -48 -56 720 834
use sg13g2_decap_4  FILLER_0_32
timestamp 1747537721
transform 1 0 3648 0 1 756
box -48 -56 432 834
use sg13g2_fill_1  FILLER_0_36
timestamp 1747537721
transform 1 0 4032 0 1 756
box -48 -56 144 834
use sg13g2_fill_1  FILLER_0_41
timestamp 1747537721
transform 1 0 4512 0 1 756
box -48 -56 144 834
use sg13g2_fill_1  FILLER_0_60
timestamp 1747537721
transform 1 0 6336 0 1 756
box -48 -56 144 834
use sg13g2_fill_2  FILLER_0_87
timestamp 1747537721
transform 1 0 8928 0 1 756
box -48 -56 240 834
use sg13g2_fill_1  FILLER_0_106
timestamp 1747537721
transform 1 0 10752 0 1 756
box -48 -56 144 834
use sg13g2_decap_4  FILLER_0_117
timestamp 1747537721
transform 1 0 11808 0 1 756
box -48 -56 432 834
use sg13g2_fill_2  FILLER_0_121
timestamp 1747537721
transform 1 0 12192 0 1 756
box -48 -56 240 834
use sg13g2_decap_4  FILLER_0_136
timestamp 1747537721
transform 1 0 13632 0 1 756
box -48 -56 432 834
use sg13g2_fill_2  FILLER_0_140
timestamp 1747537721
transform 1 0 14016 0 1 756
box -48 -56 240 834
use sg13g2_fill_2  FILLER_0_154
timestamp 1747537721
transform 1 0 15360 0 1 756
box -48 -56 240 834
use sg13g2_fill_1  FILLER_0_156
timestamp 1747537721
transform 1 0 15552 0 1 756
box -48 -56 144 834
use sg13g2_decap_4  FILLER_0_183
timestamp 1747537721
transform 1 0 18144 0 1 756
box -48 -56 432 834
use sg13g2_fill_2  FILLER_0_187
timestamp 1747537721
transform 1 0 18528 0 1 756
box -48 -56 240 834
use sg13g2_decap_8  FILLER_0_194
timestamp 1747537721
transform 1 0 19200 0 1 756
box -48 -56 720 834
use sg13g2_fill_1  FILLER_0_201
timestamp 1747537721
transform 1 0 19872 0 1 756
box -48 -56 144 834
use sg13g2_fill_1  FILLER_0_215
timestamp 1747537721
transform 1 0 21216 0 1 756
box -48 -56 144 834
use sg13g2_decap_4  FILLER_0_224
timestamp 1747537721
transform 1 0 22080 0 1 756
box -48 -56 432 834
use sg13g2_fill_2  FILLER_0_228
timestamp 1747537721
transform 1 0 22464 0 1 756
box -48 -56 240 834
use sg13g2_decap_4  FILLER_0_269
timestamp 1747537721
transform 1 0 26400 0 1 756
box -48 -56 432 834
use sg13g2_decap_8  FILLER_0_282
timestamp 1747537721
transform 1 0 27648 0 1 756
box -48 -56 720 834
use sg13g2_fill_1  FILLER_0_289
timestamp 1747537721
transform 1 0 28320 0 1 756
box -48 -56 144 834
use sg13g2_decap_4  FILLER_0_316
timestamp 1747537721
transform 1 0 30912 0 1 756
box -48 -56 432 834
use sg13g2_fill_1  FILLER_0_320
timestamp 1747537721
transform 1 0 31296 0 1 756
box -48 -56 144 834
use sg13g2_decap_4  FILLER_1_0
timestamp 1747537721
transform 1 0 576 0 -1 2268
box -48 -56 432 834
use sg13g2_fill_2  FILLER_1_4
timestamp 1747537721
transform 1 0 960 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_44
timestamp 1747537721
transform 1 0 4800 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_1_62
timestamp 1747537721
transform 1 0 6528 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_2  FILLER_1_69
timestamp 1747537721
transform 1 0 7200 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_71
timestamp 1747537721
transform 1 0 7392 0 -1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_76
timestamp 1747537721
transform 1 0 7872 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_1_83
timestamp 1747537721
transform 1 0 8544 0 -1 2268
box -48 -56 432 834
use sg13g2_decap_4  FILLER_1_91
timestamp 1747537721
transform 1 0 9312 0 -1 2268
box -48 -56 432 834
use sg13g2_fill_1  FILLER_1_95
timestamp 1747537721
transform 1 0 9696 0 -1 2268
box -48 -56 144 834
use sg13g2_decap_4  FILLER_1_112
timestamp 1747537721
transform 1 0 11328 0 -1 2268
box -48 -56 432 834
use sg13g2_decap_4  FILLER_1_156
timestamp 1747537721
transform 1 0 15552 0 -1 2268
box -48 -56 432 834
use sg13g2_fill_1  FILLER_1_160
timestamp 1747537721
transform 1 0 15936 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_1_165
timestamp 1747537721
transform 1 0 16416 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_167
timestamp 1747537721
transform 1 0 16608 0 -1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_172
timestamp 1747537721
transform 1 0 17088 0 -1 2268
box -48 -56 720 834
use sg13g2_fill_1  FILLER_1_179
timestamp 1747537721
transform 1 0 17760 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_1  FILLER_1_192
timestamp 1747537721
transform 1 0 19008 0 -1 2268
box -48 -56 144 834
use sg13g2_decap_4  FILLER_1_224
timestamp 1747537721
transform 1 0 22080 0 -1 2268
box -48 -56 432 834
use sg13g2_fill_1  FILLER_1_240
timestamp 1747537721
transform 1 0 23616 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_1_259
timestamp 1747537721
transform 1 0 25440 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_261
timestamp 1747537721
transform 1 0 25632 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_1_288
timestamp 1747537721
transform 1 0 28224 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_2  FILLER_1_295
timestamp 1747537721
transform 1 0 28896 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_306
timestamp 1747537721
transform 1 0 29952 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_1  FILLER_1_320
timestamp 1747537721
transform 1 0 31296 0 -1 2268
box -48 -56 144 834
use sg13g2_decap_4  FILLER_2_0
timestamp 1747537721
transform 1 0 576 0 1 2268
box -48 -56 432 834
use sg13g2_fill_1  FILLER_2_4
timestamp 1747537721
transform 1 0 960 0 1 2268
box -48 -56 144 834
use sg13g2_decap_4  FILLER_2_15
timestamp 1747537721
transform 1 0 2016 0 1 2268
box -48 -56 432 834
use sg13g2_fill_2  FILLER_2_23
timestamp 1747537721
transform 1 0 2784 0 1 2268
box -48 -56 240 834
use sg13g2_fill_2  FILLER_2_37
timestamp 1747537721
transform 1 0 4128 0 1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_39
timestamp 1747537721
transform 1 0 4320 0 1 2268
box -48 -56 144 834
use sg13g2_fill_1  FILLER_2_78
timestamp 1747537721
transform 1 0 8064 0 1 2268
box -48 -56 144 834
use sg13g2_decap_4  FILLER_2_100
timestamp 1747537721
transform 1 0 10176 0 1 2268
box -48 -56 432 834
use sg13g2_decap_8  FILLER_2_109
timestamp 1747537721
transform 1 0 11040 0 1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_116
timestamp 1747537721
transform 1 0 11712 0 1 2268
box -48 -56 432 834
use sg13g2_fill_2  FILLER_2_120
timestamp 1747537721
transform 1 0 12096 0 1 2268
box -48 -56 240 834
use sg13g2_fill_2  FILLER_2_127
timestamp 1747537721
transform 1 0 12768 0 1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_129
timestamp 1747537721
transform 1 0 12960 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_135
timestamp 1747537721
transform 1 0 13536 0 1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_142
timestamp 1747537721
transform 1 0 14208 0 1 2268
box -48 -56 432 834
use sg13g2_decap_8  FILLER_2_151
timestamp 1747537721
transform 1 0 15072 0 1 2268
box -48 -56 720 834
use sg13g2_fill_1  FILLER_2_158
timestamp 1747537721
transform 1 0 15744 0 1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_2_174
timestamp 1747537721
transform 1 0 17280 0 1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_184
timestamp 1747537721
transform 1 0 18240 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_193
timestamp 1747537721
transform 1 0 19104 0 1 2268
box -48 -56 720 834
use sg13g2_fill_1  FILLER_2_200
timestamp 1747537721
transform 1 0 19776 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_206
timestamp 1747537721
transform 1 0 20352 0 1 2268
box -48 -56 720 834
use sg13g2_fill_1  FILLER_2_213
timestamp 1747537721
transform 1 0 21024 0 1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_2_233
timestamp 1747537721
transform 1 0 22944 0 1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_254
timestamp 1747537721
transform 1 0 24960 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_263
timestamp 1747537721
transform 1 0 25824 0 1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_2_270
timestamp 1747537721
transform 1 0 26496 0 1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_272
timestamp 1747537721
transform 1 0 26688 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_277
timestamp 1747537721
transform 1 0 27168 0 1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_2_284
timestamp 1747537721
transform 1 0 27840 0 1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_286
timestamp 1747537721
transform 1 0 28032 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_313
timestamp 1747537721
transform 1 0 30624 0 1 2268
box -48 -56 720 834
use sg13g2_fill_1  FILLER_2_320
timestamp 1747537721
transform 1 0 31296 0 1 2268
box -48 -56 144 834
use sg13g2_decap_4  FILLER_3_0
timestamp 1747537721
transform 1 0 576 0 -1 3780
box -48 -56 432 834
use sg13g2_fill_1  FILLER_3_4
timestamp 1747537721
transform 1 0 960 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_4  FILLER_3_34
timestamp 1747537721
transform 1 0 3840 0 -1 3780
box -48 -56 432 834
use sg13g2_fill_1  FILLER_3_38
timestamp 1747537721
transform 1 0 4224 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_60
timestamp 1747537721
transform 1 0 6336 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_67
timestamp 1747537721
transform 1 0 7008 0 -1 3780
box -48 -56 432 834
use sg13g2_decap_8  FILLER_3_76
timestamp 1747537721
transform 1 0 7872 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_83
timestamp 1747537721
transform 1 0 8544 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_98
timestamp 1747537721
transform 1 0 9984 0 -1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_3_110
timestamp 1747537721
transform 1 0 11136 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_128
timestamp 1747537721
transform 1 0 12864 0 -1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_3_134
timestamp 1747537721
transform 1 0 13440 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_136
timestamp 1747537721
transform 1 0 13632 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_4  FILLER_3_156
timestamp 1747537721
transform 1 0 15552 0 -1 3780
box -48 -56 432 834
use sg13g2_fill_1  FILLER_3_160
timestamp 1747537721
transform 1 0 15936 0 -1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_3_177
timestamp 1747537721
transform 1 0 17568 0 -1 3780
box -48 -56 240 834
use sg13g2_decap_4  FILLER_3_189
timestamp 1747537721
transform 1 0 18720 0 -1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_3_214
timestamp 1747537721
transform 1 0 21120 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_252
timestamp 1747537721
transform 1 0 24768 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_266
timestamp 1747537721
transform 1 0 26112 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_273
timestamp 1747537721
transform 1 0 26784 0 -1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_3_285
timestamp 1747537721
transform 1 0 27936 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_0
timestamp 1747537721
transform 1 0 576 0 1 3780
box -48 -56 144 834
use sg13g2_fill_1  FILLER_4_10
timestamp 1747537721
transform 1 0 1536 0 1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_20
timestamp 1747537721
transform 1 0 2496 0 1 3780
box -48 -56 720 834
use sg13g2_fill_1  FILLER_4_27
timestamp 1747537721
transform 1 0 3168 0 1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_32
timestamp 1747537721
transform 1 0 3648 0 1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_39
timestamp 1747537721
transform 1 0 4320 0 1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_4_56
timestamp 1747537721
transform 1 0 5952 0 1 3780
box -48 -56 240 834
use sg13g2_fill_2  FILLER_4_79
timestamp 1747537721
transform 1 0 8160 0 1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_81
timestamp 1747537721
transform 1 0 8352 0 1 3780
box -48 -56 144 834
use sg13g2_fill_1  FILLER_4_100
timestamp 1747537721
transform 1 0 10176 0 1 3780
box -48 -56 144 834
use sg13g2_decap_4  FILLER_4_116
timestamp 1747537721
transform 1 0 11712 0 1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_4_120
timestamp 1747537721
transform 1 0 12096 0 1 3780
box -48 -56 240 834
use sg13g2_fill_2  FILLER_4_127
timestamp 1747537721
transform 1 0 12768 0 1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_4_133
timestamp 1747537721
transform 1 0 13344 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_148
timestamp 1747537721
transform 1 0 14784 0 1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_155
timestamp 1747537721
transform 1 0 15456 0 1 3780
box -48 -56 432 834
use sg13g2_fill_1  FILLER_4_159
timestamp 1747537721
transform 1 0 15840 0 1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_169
timestamp 1747537721
transform 1 0 16800 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_189
timestamp 1747537721
transform 1 0 18720 0 1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_204
timestamp 1747537721
transform 1 0 20160 0 1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_4_208
timestamp 1747537721
transform 1 0 20544 0 1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_4_226
timestamp 1747537721
transform 1 0 22272 0 1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_233
timestamp 1747537721
transform 1 0 22944 0 1 3780
box -48 -56 432 834
use sg13g2_fill_1  FILLER_4_237
timestamp 1747537721
transform 1 0 23328 0 1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_242
timestamp 1747537721
transform 1 0 23808 0 1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_4_249
timestamp 1747537721
transform 1 0 24480 0 1 3780
box -48 -56 240 834
use sg13g2_decap_4  FILLER_4_259
timestamp 1747537721
transform 1 0 25440 0 1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_4_290
timestamp 1747537721
transform 1 0 28416 0 1 3780
box -48 -56 240 834
use sg13g2_fill_2  FILLER_4_319
timestamp 1747537721
transform 1 0 31200 0 1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_5_0
timestamp 1747537721
transform 1 0 576 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_7
timestamp 1747537721
transform 1 0 1248 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_9
timestamp 1747537721
transform 1 0 1440 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_14
timestamp 1747537721
transform 1 0 1920 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_42
timestamp 1747537721
transform 1 0 4608 0 -1 5292
box -48 -56 432 834
use sg13g2_fill_1  FILLER_5_46
timestamp 1747537721
transform 1 0 4992 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_55
timestamp 1747537721
transform 1 0 5856 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_62
timestamp 1747537721
transform 1 0 6528 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_1  FILLER_5_69
timestamp 1747537721
transform 1 0 7200 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_4  FILLER_5_80
timestamp 1747537721
transform 1 0 8256 0 -1 5292
box -48 -56 432 834
use sg13g2_fill_1  FILLER_5_84
timestamp 1747537721
transform 1 0 8640 0 -1 5292
box -48 -56 144 834
use sg13g2_fill_1  FILLER_5_88
timestamp 1747537721
transform 1 0 9024 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_4  FILLER_5_110
timestamp 1747537721
transform 1 0 11136 0 -1 5292
box -48 -56 432 834
use sg13g2_fill_1  FILLER_5_114
timestamp 1747537721
transform 1 0 11520 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_136
timestamp 1747537721
transform 1 0 13632 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_1  FILLER_5_143
timestamp 1747537721
transform 1 0 14304 0 -1 5292
box -48 -56 144 834
use sg13g2_fill_2  FILLER_5_149
timestamp 1747537721
transform 1 0 14880 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_2  FILLER_5_177
timestamp 1747537721
transform 1 0 17568 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_197
timestamp 1747537721
transform 1 0 19488 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_211
timestamp 1747537721
transform 1 0 20832 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_223
timestamp 1747537721
transform 1 0 21984 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_1  FILLER_5_230
timestamp 1747537721
transform 1 0 22656 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_255
timestamp 1747537721
transform 1 0 25056 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_278
timestamp 1747537721
transform 1 0 27264 0 -1 5292
box -48 -56 432 834
use sg13g2_fill_1  FILLER_5_282
timestamp 1747537721
transform 1 0 27648 0 -1 5292
box -48 -56 144 834
use sg13g2_fill_1  FILLER_5_298
timestamp 1747537721
transform 1 0 29184 0 -1 5292
box -48 -56 144 834
use sg13g2_fill_2  FILLER_5_319
timestamp 1747537721
transform 1 0 31200 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_2  FILLER_6_16
timestamp 1747537721
transform 1 0 2112 0 1 5292
box -48 -56 240 834
use sg13g2_fill_2  FILLER_6_27
timestamp 1747537721
transform 1 0 3168 0 1 5292
box -48 -56 240 834
use sg13g2_decap_4  FILLER_6_33
timestamp 1747537721
transform 1 0 3744 0 1 5292
box -48 -56 432 834
use sg13g2_decap_4  FILLER_6_46
timestamp 1747537721
transform 1 0 4992 0 1 5292
box -48 -56 432 834
use sg13g2_fill_2  FILLER_6_72
timestamp 1747537721
transform 1 0 7488 0 1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_74
timestamp 1747537721
transform 1 0 7680 0 1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_97
timestamp 1747537721
transform 1 0 9888 0 1 5292
box -48 -56 720 834
use sg13g2_fill_1  FILLER_6_104
timestamp 1747537721
transform 1 0 10560 0 1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_115
timestamp 1747537721
transform 1 0 11616 0 1 5292
box -48 -56 720 834
use sg13g2_fill_1  FILLER_6_122
timestamp 1747537721
transform 1 0 12288 0 1 5292
box -48 -56 144 834
use sg13g2_fill_2  FILLER_6_133
timestamp 1747537721
transform 1 0 13344 0 1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_135
timestamp 1747537721
transform 1 0 13536 0 1 5292
box -48 -56 144 834
use sg13g2_fill_2  FILLER_6_157
timestamp 1747537721
transform 1 0 15648 0 1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_159
timestamp 1747537721
transform 1 0 15840 0 1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_168
timestamp 1747537721
transform 1 0 16704 0 1 5292
box -48 -56 720 834
use sg13g2_fill_1  FILLER_6_175
timestamp 1747537721
transform 1 0 17376 0 1 5292
box -48 -56 144 834
use sg13g2_fill_1  FILLER_6_181
timestamp 1747537721
transform 1 0 17952 0 1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_192
timestamp 1747537721
transform 1 0 19008 0 1 5292
box -48 -56 720 834
use sg13g2_fill_1  FILLER_6_199
timestamp 1747537721
transform 1 0 19680 0 1 5292
box -48 -56 144 834
use sg13g2_fill_2  FILLER_6_213
timestamp 1747537721
transform 1 0 21024 0 1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_6_230
timestamp 1747537721
transform 1 0 22656 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_237
timestamp 1747537721
transform 1 0 23328 0 1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_244
timestamp 1747537721
transform 1 0 24000 0 1 5292
box -48 -56 432 834
use sg13g2_decap_8  FILLER_6_268
timestamp 1747537721
transform 1 0 26304 0 1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_275
timestamp 1747537721
transform 1 0 26976 0 1 5292
box -48 -56 432 834
use sg13g2_fill_2  FILLER_6_287
timestamp 1747537721
transform 1 0 28128 0 1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_289
timestamp 1747537721
transform 1 0 28320 0 1 5292
box -48 -56 144 834
use sg13g2_fill_2  FILLER_6_300
timestamp 1747537721
transform 1 0 29376 0 1 5292
box -48 -56 240 834
use sg13g2_decap_4  FILLER_6_317
timestamp 1747537721
transform 1 0 31008 0 1 5292
box -48 -56 432 834
use sg13g2_decap_8  FILLER_7_0
timestamp 1747537721
transform 1 0 576 0 -1 6804
box -48 -56 720 834
use sg13g2_fill_1  FILLER_7_15
timestamp 1747537721
transform 1 0 2016 0 -1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_48
timestamp 1747537721
transform 1 0 5184 0 -1 6804
box -48 -56 720 834
use sg13g2_fill_1  FILLER_7_65
timestamp 1747537721
transform 1 0 6816 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_7_74
timestamp 1747537721
transform 1 0 7680 0 -1 6804
box -48 -56 240 834
use sg13g2_decap_8  FILLER_7_81
timestamp 1747537721
transform 1 0 8352 0 -1 6804
box -48 -56 720 834
use sg13g2_fill_1  FILLER_7_88
timestamp 1747537721
transform 1 0 9024 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_7_93
timestamp 1747537721
transform 1 0 9504 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_7_102
timestamp 1747537721
transform 1 0 10368 0 -1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_108
timestamp 1747537721
transform 1 0 10944 0 -1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_7_131
timestamp 1747537721
transform 1 0 13152 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_133
timestamp 1747537721
transform 1 0 13344 0 -1 6804
box -48 -56 144 834
use sg13g2_decap_4  FILLER_7_143
timestamp 1747537721
transform 1 0 14304 0 -1 6804
box -48 -56 432 834
use sg13g2_decap_4  FILLER_7_152
timestamp 1747537721
transform 1 0 15168 0 -1 6804
box -48 -56 432 834
use sg13g2_fill_2  FILLER_7_172
timestamp 1747537721
transform 1 0 17088 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_174
timestamp 1747537721
transform 1 0 17280 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_7_185
timestamp 1747537721
transform 1 0 18336 0 -1 6804
box -48 -56 240 834
use sg13g2_decap_8  FILLER_7_195
timestamp 1747537721
transform 1 0 19296 0 -1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_7_202
timestamp 1747537721
transform 1 0 19968 0 -1 6804
box -48 -56 240 834
use sg13g2_decap_4  FILLER_7_212
timestamp 1747537721
transform 1 0 20928 0 -1 6804
box -48 -56 432 834
use sg13g2_fill_1  FILLER_7_216
timestamp 1747537721
transform 1 0 21312 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_7_225
timestamp 1747537721
transform 1 0 22176 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_7_229
timestamp 1747537721
transform 1 0 22560 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_231
timestamp 1747537721
transform 1 0 22752 0 -1 6804
box -48 -56 144 834
use sg13g2_decap_4  FILLER_7_248
timestamp 1747537721
transform 1 0 24384 0 -1 6804
box -48 -56 432 834
use sg13g2_fill_2  FILLER_7_252
timestamp 1747537721
transform 1 0 24768 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_2  FILLER_7_270
timestamp 1747537721
transform 1 0 26496 0 -1 6804
box -48 -56 240 834
use sg13g2_decap_4  FILLER_7_305
timestamp 1747537721
transform 1 0 29856 0 -1 6804
box -48 -56 432 834
use sg13g2_decap_4  FILLER_7_317
timestamp 1747537721
transform 1 0 31008 0 -1 6804
box -48 -56 432 834
use sg13g2_decap_4  FILLER_8_0
timestamp 1747537721
transform 1 0 576 0 1 6804
box -48 -56 432 834
use sg13g2_fill_2  FILLER_8_21
timestamp 1747537721
transform 1 0 2592 0 1 6804
box -48 -56 240 834
use sg13g2_decap_8  FILLER_8_28
timestamp 1747537721
transform 1 0 3264 0 1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_8_35
timestamp 1747537721
transform 1 0 3936 0 1 6804
box -48 -56 240 834
use sg13g2_decap_8  FILLER_8_47
timestamp 1747537721
transform 1 0 5088 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_54
timestamp 1747537721
transform 1 0 5760 0 1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_8_61
timestamp 1747537721
transform 1 0 6432 0 1 6804
box -48 -56 240 834
use sg13g2_decap_4  FILLER_8_67
timestamp 1747537721
transform 1 0 7008 0 1 6804
box -48 -56 432 834
use sg13g2_fill_2  FILLER_8_71
timestamp 1747537721
transform 1 0 7392 0 1 6804
box -48 -56 240 834
use sg13g2_fill_2  FILLER_8_94
timestamp 1747537721
transform 1 0 9600 0 1 6804
box -48 -56 240 834
use sg13g2_decap_4  FILLER_8_104
timestamp 1747537721
transform 1 0 10560 0 1 6804
box -48 -56 432 834
use sg13g2_decap_4  FILLER_8_113
timestamp 1747537721
transform 1 0 11424 0 1 6804
box -48 -56 432 834
use sg13g2_fill_1  FILLER_8_117
timestamp 1747537721
transform 1 0 11808 0 1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_8_128
timestamp 1747537721
transform 1 0 12864 0 1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_130
timestamp 1747537721
transform 1 0 13056 0 1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_135
timestamp 1747537721
transform 1 0 13536 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_158
timestamp 1747537721
transform 1 0 15744 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_165
timestamp 1747537721
transform 1 0 16416 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_172
timestamp 1747537721
transform 1 0 17088 0 1 6804
box -48 -56 720 834
use sg13g2_fill_1  FILLER_8_179
timestamp 1747537721
transform 1 0 17760 0 1 6804
box -48 -56 144 834
use sg13g2_decap_4  FILLER_8_190
timestamp 1747537721
transform 1 0 18816 0 1 6804
box -48 -56 432 834
use sg13g2_fill_2  FILLER_8_211
timestamp 1747537721
transform 1 0 20832 0 1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_213
timestamp 1747537721
transform 1 0 21024 0 1 6804
box -48 -56 144 834
use sg13g2_decap_4  FILLER_8_230
timestamp 1747537721
transform 1 0 22656 0 1 6804
box -48 -56 432 834
use sg13g2_fill_1  FILLER_8_234
timestamp 1747537721
transform 1 0 23040 0 1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_259
timestamp 1747537721
transform 1 0 25440 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_266
timestamp 1747537721
transform 1 0 26112 0 1 6804
box -48 -56 720 834
use sg13g2_decap_4  FILLER_8_273
timestamp 1747537721
transform 1 0 26784 0 1 6804
box -48 -56 432 834
use sg13g2_fill_2  FILLER_8_277
timestamp 1747537721
transform 1 0 27168 0 1 6804
box -48 -56 240 834
use sg13g2_fill_2  FILLER_8_284
timestamp 1747537721
transform 1 0 27840 0 1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_309
timestamp 1747537721
transform 1 0 30240 0 1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_8_318
timestamp 1747537721
transform 1 0 31104 0 1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_320
timestamp 1747537721
transform 1 0 31296 0 1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_9_0
timestamp 1747537721
transform 1 0 576 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_2
timestamp 1747537721
transform 1 0 768 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_9_15
timestamp 1747537721
transform 1 0 2016 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_17
timestamp 1747537721
transform 1 0 2208 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_9_22
timestamp 1747537721
transform 1 0 2688 0 -1 8316
box -48 -56 240 834
use sg13g2_decap_8  FILLER_9_29
timestamp 1747537721
transform 1 0 3360 0 -1 8316
box -48 -56 720 834
use sg13g2_fill_1  FILLER_9_36
timestamp 1747537721
transform 1 0 4032 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_9_57
timestamp 1747537721
transform 1 0 6048 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_59
timestamp 1747537721
transform 1 0 6240 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_77
timestamp 1747537721
transform 1 0 7968 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_84
timestamp 1747537721
transform 1 0 8640 0 -1 8316
box -48 -56 720 834
use sg13g2_fill_1  FILLER_9_91
timestamp 1747537721
transform 1 0 9312 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_95
timestamp 1747537721
transform 1 0 9696 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_102
timestamp 1747537721
transform 1 0 10368 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_109
timestamp 1747537721
transform 1 0 11040 0 -1 8316
box -48 -56 720 834
use sg13g2_fill_1  FILLER_9_134
timestamp 1747537721
transform 1 0 13440 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_9_143
timestamp 1747537721
transform 1 0 14304 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_145
timestamp 1747537721
transform 1 0 14496 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_150
timestamp 1747537721
transform 1 0 14976 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_157
timestamp 1747537721
transform 1 0 15648 0 -1 8316
box -48 -56 720 834
use sg13g2_fill_1  FILLER_9_164
timestamp 1747537721
transform 1 0 16320 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_9_177
timestamp 1747537721
transform 1 0 17568 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_179
timestamp 1747537721
transform 1 0 17760 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_4  FILLER_9_190
timestamp 1747537721
transform 1 0 18816 0 -1 8316
box -48 -56 432 834
use sg13g2_decap_8  FILLER_9_207
timestamp 1747537721
transform 1 0 20448 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_4  FILLER_9_214
timestamp 1747537721
transform 1 0 21120 0 -1 8316
box -48 -56 432 834
use sg13g2_fill_1  FILLER_9_233
timestamp 1747537721
transform 1 0 22944 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_4  FILLER_9_286
timestamp 1747537721
transform 1 0 28032 0 -1 8316
box -48 -56 432 834
use sg13g2_fill_1  FILLER_9_290
timestamp 1747537721
transform 1 0 28416 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_9_299
timestamp 1747537721
transform 1 0 29280 0 -1 8316
box -48 -56 240 834
use sg13g2_decap_4  FILLER_10_0
timestamp 1747537721
transform 1 0 576 0 1 8316
box -48 -56 432 834
use sg13g2_fill_1  FILLER_10_4
timestamp 1747537721
transform 1 0 960 0 1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_10_13
timestamp 1747537721
transform 1 0 1824 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_42
timestamp 1747537721
transform 1 0 4608 0 1 8316
box -48 -56 144 834
use sg13g2_decap_4  FILLER_10_59
timestamp 1747537721
transform 1 0 6240 0 1 8316
box -48 -56 432 834
use sg13g2_decap_4  FILLER_10_71
timestamp 1747537721
transform 1 0 7392 0 1 8316
box -48 -56 432 834
use sg13g2_fill_1  FILLER_10_104
timestamp 1747537721
transform 1 0 10560 0 1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_10_118
timestamp 1747537721
transform 1 0 11904 0 1 8316
box -48 -56 240 834
use sg13g2_decap_8  FILLER_10_127
timestamp 1747537721
transform 1 0 12768 0 1 8316
box -48 -56 720 834
use sg13g2_fill_1  FILLER_10_134
timestamp 1747537721
transform 1 0 13440 0 1 8316
box -48 -56 144 834
use sg13g2_decap_4  FILLER_10_140
timestamp 1747537721
transform 1 0 14016 0 1 8316
box -48 -56 432 834
use sg13g2_fill_1  FILLER_10_149
timestamp 1747537721
transform 1 0 14880 0 1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_10_160
timestamp 1747537721
transform 1 0 15936 0 1 8316
box -48 -56 240 834
use sg13g2_fill_2  FILLER_10_175
timestamp 1747537721
transform 1 0 17376 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_177
timestamp 1747537721
transform 1 0 17568 0 1 8316
box -48 -56 144 834
use sg13g2_decap_4  FILLER_10_188
timestamp 1747537721
transform 1 0 18624 0 1 8316
box -48 -56 432 834
use sg13g2_decap_8  FILLER_10_207
timestamp 1747537721
transform 1 0 20448 0 1 8316
box -48 -56 720 834
use sg13g2_decap_4  FILLER_10_214
timestamp 1747537721
transform 1 0 21120 0 1 8316
box -48 -56 432 834
use sg13g2_decap_8  FILLER_10_222
timestamp 1747537721
transform 1 0 21888 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_229
timestamp 1747537721
transform 1 0 22560 0 1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_10_236
timestamp 1747537721
transform 1 0 23232 0 1 8316
box -48 -56 240 834
use sg13g2_fill_2  FILLER_10_246
timestamp 1747537721
transform 1 0 24192 0 1 8316
box -48 -56 240 834
use sg13g2_decap_8  FILLER_10_255
timestamp 1747537721
transform 1 0 25056 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_262
timestamp 1747537721
transform 1 0 25728 0 1 8316
box -48 -56 720 834
use sg13g2_fill_1  FILLER_10_269
timestamp 1747537721
transform 1 0 26400 0 1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_277
timestamp 1747537721
transform 1 0 27168 0 1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_10_284
timestamp 1747537721
transform 1 0 27840 0 1 8316
box -48 -56 240 834
use sg13g2_decap_4  FILLER_11_0
timestamp 1747537721
transform 1 0 576 0 -1 9828
box -48 -56 432 834
use sg13g2_fill_1  FILLER_11_4
timestamp 1747537721
transform 1 0 960 0 -1 9828
box -48 -56 144 834
use sg13g2_fill_1  FILLER_11_21
timestamp 1747537721
transform 1 0 2592 0 -1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_27
timestamp 1747537721
transform 1 0 3168 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_34
timestamp 1747537721
transform 1 0 3840 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_41
timestamp 1747537721
transform 1 0 4512 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_11_48
timestamp 1747537721
transform 1 0 5184 0 -1 9828
box -48 -56 432 834
use sg13g2_fill_2  FILLER_11_52
timestamp 1747537721
transform 1 0 5568 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_2  FILLER_11_73
timestamp 1747537721
transform 1 0 7584 0 -1 9828
box -48 -56 240 834
use sg13g2_decap_8  FILLER_11_89
timestamp 1747537721
transform 1 0 9120 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_11_96
timestamp 1747537721
transform 1 0 9792 0 -1 9828
box -48 -56 432 834
use sg13g2_fill_1  FILLER_11_100
timestamp 1747537721
transform 1 0 10176 0 -1 9828
box -48 -56 144 834
use sg13g2_fill_2  FILLER_11_106
timestamp 1747537721
transform 1 0 10752 0 -1 9828
box -48 -56 240 834
use sg13g2_decap_4  FILLER_11_121
timestamp 1747537721
transform 1 0 12192 0 -1 9828
box -48 -56 432 834
use sg13g2_fill_2  FILLER_11_125
timestamp 1747537721
transform 1 0 12576 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_2  FILLER_11_152
timestamp 1747537721
transform 1 0 15168 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_2  FILLER_11_163
timestamp 1747537721
transform 1 0 16224 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_165
timestamp 1747537721
transform 1 0 16416 0 -1 9828
box -48 -56 144 834
use sg13g2_decap_4  FILLER_11_171
timestamp 1747537721
transform 1 0 16992 0 -1 9828
box -48 -56 432 834
use sg13g2_fill_2  FILLER_11_175
timestamp 1747537721
transform 1 0 17376 0 -1 9828
box -48 -56 240 834
use sg13g2_decap_4  FILLER_11_182
timestamp 1747537721
transform 1 0 18048 0 -1 9828
box -48 -56 432 834
use sg13g2_fill_2  FILLER_11_186
timestamp 1747537721
transform 1 0 18432 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_2  FILLER_11_193
timestamp 1747537721
transform 1 0 19104 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_2  FILLER_11_205
timestamp 1747537721
transform 1 0 20256 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_233
timestamp 1747537721
transform 1 0 22944 0 -1 9828
box -48 -56 144 834
use sg13g2_fill_1  FILLER_11_243
timestamp 1747537721
transform 1 0 23904 0 -1 9828
box -48 -56 144 834
use sg13g2_fill_2  FILLER_11_285
timestamp 1747537721
transform 1 0 27936 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_12_21
timestamp 1747537721
transform 1 0 2592 0 1 9828
box -48 -56 144 834
use sg13g2_fill_2  FILLER_12_27
timestamp 1747537721
transform 1 0 3168 0 1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_12_29
timestamp 1747537721
transform 1 0 3360 0 1 9828
box -48 -56 144 834
use sg13g2_fill_2  FILLER_12_46
timestamp 1747537721
transform 1 0 4992 0 1 9828
box -48 -56 240 834
use sg13g2_fill_2  FILLER_12_56
timestamp 1747537721
transform 1 0 5952 0 1 9828
box -48 -56 240 834
use sg13g2_decap_4  FILLER_12_99
timestamp 1747537721
transform 1 0 10080 0 1 9828
box -48 -56 432 834
use sg13g2_fill_1  FILLER_12_113
timestamp 1747537721
transform 1 0 11424 0 1 9828
box -48 -56 144 834
use sg13g2_decap_4  FILLER_12_125
timestamp 1747537721
transform 1 0 12576 0 1 9828
box -48 -56 432 834
use sg13g2_fill_2  FILLER_12_129
timestamp 1747537721
transform 1 0 12960 0 1 9828
box -48 -56 240 834
use sg13g2_decap_4  FILLER_12_136
timestamp 1747537721
transform 1 0 13632 0 1 9828
box -48 -56 432 834
use sg13g2_fill_2  FILLER_12_140
timestamp 1747537721
transform 1 0 14016 0 1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_12_147
timestamp 1747537721
transform 1 0 14688 0 1 9828
box -48 -56 144 834
use sg13g2_decap_4  FILLER_12_159
timestamp 1747537721
transform 1 0 15840 0 1 9828
box -48 -56 432 834
use sg13g2_fill_2  FILLER_12_163
timestamp 1747537721
transform 1 0 16224 0 1 9828
box -48 -56 240 834
use sg13g2_decap_8  FILLER_12_179
timestamp 1747537721
transform 1 0 17760 0 1 9828
box -48 -56 720 834
use sg13g2_fill_1  FILLER_12_186
timestamp 1747537721
transform 1 0 18432 0 1 9828
box -48 -56 144 834
use sg13g2_fill_2  FILLER_12_196
timestamp 1747537721
transform 1 0 19392 0 1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_12_198
timestamp 1747537721
transform 1 0 19584 0 1 9828
box -48 -56 144 834
use sg13g2_fill_1  FILLER_12_204
timestamp 1747537721
transform 1 0 20160 0 1 9828
box -48 -56 144 834
use sg13g2_fill_2  FILLER_12_210
timestamp 1747537721
transform 1 0 20736 0 1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_12_247
timestamp 1747537721
transform 1 0 24288 0 1 9828
box -48 -56 144 834
use sg13g2_fill_1  FILLER_12_257
timestamp 1747537721
transform 1 0 25248 0 1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_12_262
timestamp 1747537721
transform 1 0 25728 0 1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_12_269
timestamp 1747537721
transform 1 0 26400 0 1 9828
box -48 -56 240 834
use sg13g2_fill_2  FILLER_12_294
timestamp 1747537721
transform 1 0 28800 0 1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_12_320
timestamp 1747537721
transform 1 0 31296 0 1 9828
box -48 -56 144 834
use sg13g2_decap_4  FILLER_13_0
timestamp 1747537721
transform 1 0 576 0 -1 11340
box -48 -56 432 834
use sg13g2_fill_1  FILLER_13_4
timestamp 1747537721
transform 1 0 960 0 -1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_13_10
timestamp 1747537721
transform 1 0 1536 0 -1 11340
box -48 -56 720 834
use sg13g2_fill_2  FILLER_13_31
timestamp 1747537721
transform 1 0 3552 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_13_33
timestamp 1747537721
transform 1 0 3744 0 -1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_13_52
timestamp 1747537721
transform 1 0 5568 0 -1 11340
box -48 -56 720 834
use sg13g2_fill_1  FILLER_13_59
timestamp 1747537721
transform 1 0 6240 0 -1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_13_64
timestamp 1747537721
transform 1 0 6720 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_2  FILLER_13_74
timestamp 1747537721
transform 1 0 7680 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_13_76
timestamp 1747537721
transform 1 0 7872 0 -1 11340
box -48 -56 144 834
use sg13g2_fill_1  FILLER_13_82
timestamp 1747537721
transform 1 0 8448 0 -1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_13_95
timestamp 1747537721
transform 1 0 9696 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_13_97
timestamp 1747537721
transform 1 0 9888 0 -1 11340
box -48 -56 144 834
use sg13g2_decap_4  FILLER_13_105
timestamp 1747537721
transform 1 0 10656 0 -1 11340
box -48 -56 432 834
use sg13g2_decap_4  FILLER_13_118
timestamp 1747537721
transform 1 0 11904 0 -1 11340
box -48 -56 432 834
use sg13g2_decap_4  FILLER_13_126
timestamp 1747537721
transform 1 0 12672 0 -1 11340
box -48 -56 432 834
use sg13g2_fill_2  FILLER_13_139
timestamp 1747537721
transform 1 0 13920 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_13_141
timestamp 1747537721
transform 1 0 14112 0 -1 11340
box -48 -56 144 834
use sg13g2_fill_1  FILLER_13_147
timestamp 1747537721
transform 1 0 14688 0 -1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_13_164
timestamp 1747537721
transform 1 0 16320 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_13_166
timestamp 1747537721
transform 1 0 16512 0 -1 11340
box -48 -56 144 834
use sg13g2_fill_1  FILLER_13_172
timestamp 1747537721
transform 1 0 17088 0 -1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_13_182
timestamp 1747537721
transform 1 0 18048 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_2  FILLER_13_217
timestamp 1747537721
transform 1 0 21408 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_13_219
timestamp 1747537721
transform 1 0 21600 0 -1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_13_240
timestamp 1747537721
transform 1 0 23616 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_2  FILLER_14_0
timestamp 1747537721
transform 1 0 576 0 1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_14_2
timestamp 1747537721
transform 1 0 768 0 1 11340
box -48 -56 144 834
use sg13g2_fill_1  FILLER_14_46
timestamp 1747537721
transform 1 0 4992 0 1 11340
box -48 -56 144 834
use sg13g2_fill_1  FILLER_14_64
timestamp 1747537721
transform 1 0 6720 0 1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_14_82
timestamp 1747537721
transform 1 0 8448 0 1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_14_84
timestamp 1747537721
transform 1 0 8640 0 1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_14_104
timestamp 1747537721
transform 1 0 10560 0 1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_14_106
timestamp 1747537721
transform 1 0 10752 0 1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_14_123
timestamp 1747537721
transform 1 0 12384 0 1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_14_143
timestamp 1747537721
transform 1 0 14304 0 1 11340
box -48 -56 144 834
use sg13g2_decap_4  FILLER_14_176
timestamp 1747537721
transform 1 0 17472 0 1 11340
box -48 -56 432 834
use sg13g2_fill_1  FILLER_14_180
timestamp 1747537721
transform 1 0 17856 0 1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_14_186
timestamp 1747537721
transform 1 0 18432 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_214
timestamp 1747537721
transform 1 0 21120 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_250
timestamp 1747537721
transform 1 0 24576 0 1 11340
box -48 -56 720 834
use sg13g2_fill_1  FILLER_14_262
timestamp 1747537721
transform 1 0 25728 0 1 11340
box -48 -56 144 834
use sg13g2_fill_1  FILLER_14_272
timestamp 1747537721
transform 1 0 26688 0 1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_14_292
timestamp 1747537721
transform 1 0 28608 0 1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_14_311
timestamp 1747537721
transform 1 0 30432 0 1 11340
box -48 -56 144 834
use sg13g2_fill_1  FILLER_14_320
timestamp 1747537721
transform 1 0 31296 0 1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_15_0
timestamp 1747537721
transform 1 0 576 0 -1 12852
box -48 -56 720 834
use sg13g2_fill_2  FILLER_15_11
timestamp 1747537721
transform 1 0 1632 0 -1 12852
box -48 -56 240 834
use sg13g2_decap_4  FILLER_15_17
timestamp 1747537721
transform 1 0 2208 0 -1 12852
box -48 -56 432 834
use sg13g2_fill_2  FILLER_15_21
timestamp 1747537721
transform 1 0 2592 0 -1 12852
box -48 -56 240 834
use sg13g2_decap_4  FILLER_15_31
timestamp 1747537721
transform 1 0 3552 0 -1 12852
box -48 -56 432 834
use sg13g2_fill_2  FILLER_15_35
timestamp 1747537721
transform 1 0 3936 0 -1 12852
box -48 -56 240 834
use sg13g2_decap_4  FILLER_15_47
timestamp 1747537721
transform 1 0 5088 0 -1 12852
box -48 -56 432 834
use sg13g2_fill_2  FILLER_15_51
timestamp 1747537721
transform 1 0 5472 0 -1 12852
box -48 -56 240 834
use sg13g2_decap_8  FILLER_15_58
timestamp 1747537721
transform 1 0 6144 0 -1 12852
box -48 -56 720 834
use sg13g2_fill_2  FILLER_15_84
timestamp 1747537721
transform 1 0 8640 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_15_86
timestamp 1747537721
transform 1 0 8832 0 -1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_15_92
timestamp 1747537721
transform 1 0 9408 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_15_99
timestamp 1747537721
transform 1 0 10080 0 -1 12852
box -48 -56 432 834
use sg13g2_decap_8  FILLER_15_114
timestamp 1747537721
transform 1 0 11520 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_15_121
timestamp 1747537721
transform 1 0 12192 0 -1 12852
box -48 -56 432 834
use sg13g2_fill_1  FILLER_15_125
timestamp 1747537721
transform 1 0 12576 0 -1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_15_131
timestamp 1747537721
transform 1 0 13152 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_15_133
timestamp 1747537721
transform 1 0 13344 0 -1 12852
box -48 -56 144 834
use sg13g2_decap_4  FILLER_15_139
timestamp 1747537721
transform 1 0 13920 0 -1 12852
box -48 -56 432 834
use sg13g2_decap_8  FILLER_15_151
timestamp 1747537721
transform 1 0 15072 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_158
timestamp 1747537721
transform 1 0 15744 0 -1 12852
box -48 -56 720 834
use sg13g2_fill_1  FILLER_15_165
timestamp 1747537721
transform 1 0 16416 0 -1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_15_174
timestamp 1747537721
transform 1 0 17280 0 -1 12852
box -48 -56 720 834
use sg13g2_fill_2  FILLER_15_181
timestamp 1747537721
transform 1 0 17952 0 -1 12852
box -48 -56 240 834
use sg13g2_decap_8  FILLER_15_194
timestamp 1747537721
transform 1 0 19200 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_201
timestamp 1747537721
transform 1 0 19872 0 -1 12852
box -48 -56 720 834
use sg13g2_fill_2  FILLER_15_208
timestamp 1747537721
transform 1 0 20544 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_15_220
timestamp 1747537721
transform 1 0 21696 0 -1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_15_225
timestamp 1747537721
transform 1 0 22176 0 -1 12852
box -48 -56 720 834
use sg13g2_fill_1  FILLER_15_232
timestamp 1747537721
transform 1 0 22848 0 -1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_15_250
timestamp 1747537721
transform 1 0 24576 0 -1 12852
box -48 -56 720 834
use sg13g2_fill_2  FILLER_15_318
timestamp 1747537721
transform 1 0 31104 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_15_320
timestamp 1747537721
transform 1 0 31296 0 -1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_16_26
timestamp 1747537721
transform 1 0 3072 0 1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_16_28
timestamp 1747537721
transform 1 0 3264 0 1 12852
box -48 -56 144 834
use sg13g2_decap_4  FILLER_16_37
timestamp 1747537721
transform 1 0 4128 0 1 12852
box -48 -56 432 834
use sg13g2_fill_1  FILLER_16_41
timestamp 1747537721
transform 1 0 4512 0 1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_16_47
timestamp 1747537721
transform 1 0 5088 0 1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_16_61
timestamp 1747537721
transform 1 0 6432 0 1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_16_68
timestamp 1747537721
transform 1 0 7104 0 1 12852
box -48 -56 240 834
use sg13g2_decap_4  FILLER_16_95
timestamp 1747537721
transform 1 0 9696 0 1 12852
box -48 -56 432 834
use sg13g2_fill_1  FILLER_16_110
timestamp 1747537721
transform 1 0 11136 0 1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_16_116
timestamp 1747537721
transform 1 0 11712 0 1 12852
box -48 -56 240 834
use sg13g2_fill_2  FILLER_16_140
timestamp 1747537721
transform 1 0 14016 0 1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_16_142
timestamp 1747537721
transform 1 0 14208 0 1 12852
box -48 -56 144 834
use sg13g2_decap_4  FILLER_16_159
timestamp 1747537721
transform 1 0 15840 0 1 12852
box -48 -56 432 834
use sg13g2_fill_1  FILLER_16_187
timestamp 1747537721
transform 1 0 18528 0 1 12852
box -48 -56 144 834
use sg13g2_decap_4  FILLER_16_193
timestamp 1747537721
transform 1 0 19104 0 1 12852
box -48 -56 432 834
use sg13g2_fill_2  FILLER_16_219
timestamp 1747537721
transform 1 0 21600 0 1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_16_221
timestamp 1747537721
transform 1 0 21792 0 1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_16_232
timestamp 1747537721
transform 1 0 22848 0 1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_16_234
timestamp 1747537721
transform 1 0 23040 0 1 12852
box -48 -56 144 834
use sg13g2_decap_4  FILLER_16_250
timestamp 1747537721
transform 1 0 24576 0 1 12852
box -48 -56 432 834
use sg13g2_fill_2  FILLER_16_254
timestamp 1747537721
transform 1 0 24960 0 1 12852
box -48 -56 240 834
use sg13g2_decap_8  FILLER_16_265
timestamp 1747537721
transform 1 0 26016 0 1 12852
box -48 -56 720 834
use sg13g2_fill_2  FILLER_16_272
timestamp 1747537721
transform 1 0 26688 0 1 12852
box -48 -56 240 834
use sg13g2_decap_8  FILLER_16_283
timestamp 1747537721
transform 1 0 27744 0 1 12852
box -48 -56 720 834
use sg13g2_fill_2  FILLER_16_290
timestamp 1747537721
transform 1 0 28416 0 1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_16_292
timestamp 1747537721
transform 1 0 28608 0 1 12852
box -48 -56 144 834
use sg13g2_decap_4  FILLER_16_297
timestamp 1747537721
transform 1 0 29088 0 1 12852
box -48 -56 432 834
use sg13g2_fill_2  FILLER_16_301
timestamp 1747537721
transform 1 0 29472 0 1 12852
box -48 -56 240 834
use sg13g2_fill_2  FILLER_16_310
timestamp 1747537721
transform 1 0 30336 0 1 12852
box -48 -56 240 834
use sg13g2_decap_4  FILLER_16_316
timestamp 1747537721
transform 1 0 30912 0 1 12852
box -48 -56 432 834
use sg13g2_fill_1  FILLER_16_320
timestamp 1747537721
transform 1 0 31296 0 1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_17_9
timestamp 1747537721
transform 1 0 1440 0 -1 14364
box -48 -56 240 834
use sg13g2_decap_8  FILLER_17_34
timestamp 1747537721
transform 1 0 3840 0 -1 14364
box -48 -56 720 834
use sg13g2_fill_2  FILLER_17_41
timestamp 1747537721
transform 1 0 4512 0 -1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_17_43
timestamp 1747537721
transform 1 0 4704 0 -1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_17_63
timestamp 1747537721
transform 1 0 6624 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_70
timestamp 1747537721
transform 1 0 7296 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_77
timestamp 1747537721
transform 1 0 7968 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_84
timestamp 1747537721
transform 1 0 8640 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_4  FILLER_17_91
timestamp 1747537721
transform 1 0 9312 0 -1 14364
box -48 -56 432 834
use sg13g2_fill_2  FILLER_17_95
timestamp 1747537721
transform 1 0 9696 0 -1 14364
box -48 -56 240 834
use sg13g2_fill_2  FILLER_17_102
timestamp 1747537721
transform 1 0 10368 0 -1 14364
box -48 -56 240 834
use sg13g2_decap_4  FILLER_17_119
timestamp 1747537721
transform 1 0 12000 0 -1 14364
box -48 -56 432 834
use sg13g2_fill_1  FILLER_17_123
timestamp 1747537721
transform 1 0 12384 0 -1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_17_130
timestamp 1747537721
transform 1 0 13056 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_4  FILLER_17_137
timestamp 1747537721
transform 1 0 13728 0 -1 14364
box -48 -56 432 834
use sg13g2_decap_8  FILLER_17_156
timestamp 1747537721
transform 1 0 15552 0 -1 14364
box -48 -56 720 834
use sg13g2_fill_2  FILLER_17_163
timestamp 1747537721
transform 1 0 16224 0 -1 14364
box -48 -56 240 834
use sg13g2_decap_8  FILLER_17_173
timestamp 1747537721
transform 1 0 17184 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_180
timestamp 1747537721
transform 1 0 17856 0 -1 14364
box -48 -56 720 834
use sg13g2_fill_2  FILLER_17_187
timestamp 1747537721
transform 1 0 18528 0 -1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_17_189
timestamp 1747537721
transform 1 0 18720 0 -1 14364
box -48 -56 144 834
use sg13g2_fill_1  FILLER_17_198
timestamp 1747537721
transform 1 0 19584 0 -1 14364
box -48 -56 144 834
use sg13g2_decap_4  FILLER_17_232
timestamp 1747537721
transform 1 0 22848 0 -1 14364
box -48 -56 432 834
use sg13g2_fill_1  FILLER_17_252
timestamp 1747537721
transform 1 0 24768 0 -1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_17_268
timestamp 1747537721
transform 1 0 26304 0 -1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_17_270
timestamp 1747537721
transform 1 0 26496 0 -1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_17_284
timestamp 1747537721
transform 1 0 27840 0 -1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_17_286
timestamp 1747537721
transform 1 0 28032 0 -1 14364
box -48 -56 144 834
use sg13g2_decap_4  FILLER_18_0
timestamp 1747537721
transform 1 0 576 0 1 14364
box -48 -56 432 834
use sg13g2_fill_2  FILLER_18_28
timestamp 1747537721
transform 1 0 3264 0 1 14364
box -48 -56 240 834
use sg13g2_decap_4  FILLER_18_47
timestamp 1747537721
transform 1 0 5088 0 1 14364
box -48 -56 432 834
use sg13g2_fill_2  FILLER_18_51
timestamp 1747537721
transform 1 0 5472 0 1 14364
box -48 -56 240 834
use sg13g2_decap_4  FILLER_18_82
timestamp 1747537721
transform 1 0 8448 0 1 14364
box -48 -56 432 834
use sg13g2_fill_1  FILLER_18_98
timestamp 1747537721
transform 1 0 9984 0 1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_18_105
timestamp 1747537721
transform 1 0 10656 0 1 14364
box -48 -56 240 834
use sg13g2_decap_8  FILLER_18_116
timestamp 1747537721
transform 1 0 11712 0 1 14364
box -48 -56 720 834
use sg13g2_decap_4  FILLER_18_123
timestamp 1747537721
transform 1 0 12384 0 1 14364
box -48 -56 432 834
use sg13g2_fill_2  FILLER_18_143
timestamp 1747537721
transform 1 0 14304 0 1 14364
box -48 -56 240 834
use sg13g2_decap_8  FILLER_18_150
timestamp 1747537721
transform 1 0 14976 0 1 14364
box -48 -56 720 834
use sg13g2_fill_2  FILLER_18_157
timestamp 1747537721
transform 1 0 15648 0 1 14364
box -48 -56 240 834
use sg13g2_fill_2  FILLER_18_191
timestamp 1747537721
transform 1 0 18912 0 1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_18_193
timestamp 1747537721
transform 1 0 19104 0 1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_18_204
timestamp 1747537721
transform 1 0 20160 0 1 14364
box -48 -56 720 834
use sg13g2_decap_4  FILLER_18_232
timestamp 1747537721
transform 1 0 22848 0 1 14364
box -48 -56 432 834
use sg13g2_decap_4  FILLER_18_239
timestamp 1747537721
transform 1 0 23520 0 1 14364
box -48 -56 432 834
use sg13g2_fill_1  FILLER_18_248
timestamp 1747537721
transform 1 0 24384 0 1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_18_255
timestamp 1747537721
transform 1 0 25056 0 1 14364
box -48 -56 240 834
use sg13g2_decap_8  FILLER_18_262
timestamp 1747537721
transform 1 0 25728 0 1 14364
box -48 -56 720 834
use sg13g2_fill_2  FILLER_18_269
timestamp 1747537721
transform 1 0 26400 0 1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_18_282
timestamp 1747537721
transform 1 0 27648 0 1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_19_0
timestamp 1747537721
transform 1 0 576 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_4  FILLER_19_7
timestamp 1747537721
transform 1 0 1248 0 -1 15876
box -48 -56 432 834
use sg13g2_fill_1  FILLER_19_11
timestamp 1747537721
transform 1 0 1632 0 -1 15876
box -48 -56 144 834
use sg13g2_decap_4  FILLER_19_17
timestamp 1747537721
transform 1 0 2208 0 -1 15876
box -48 -56 432 834
use sg13g2_fill_1  FILLER_19_21
timestamp 1747537721
transform 1 0 2592 0 -1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_19_43
timestamp 1747537721
transform 1 0 4704 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_4  FILLER_19_64
timestamp 1747537721
transform 1 0 6720 0 -1 15876
box -48 -56 432 834
use sg13g2_fill_2  FILLER_19_68
timestamp 1747537721
transform 1 0 7104 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_2  FILLER_19_76
timestamp 1747537721
transform 1 0 7872 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_2  FILLER_19_83
timestamp 1747537721
transform 1 0 8544 0 -1 15876
box -48 -56 240 834
use sg13g2_decap_8  FILLER_19_103
timestamp 1747537721
transform 1 0 10464 0 -1 15876
box -48 -56 720 834
use sg13g2_fill_2  FILLER_19_110
timestamp 1747537721
transform 1 0 11136 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_2  FILLER_19_117
timestamp 1747537721
transform 1 0 11808 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_19_119
timestamp 1747537721
transform 1 0 12000 0 -1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_19_136
timestamp 1747537721
transform 1 0 13632 0 -1 15876
box -48 -56 720 834
use sg13g2_fill_1  FILLER_19_171
timestamp 1747537721
transform 1 0 16992 0 -1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_19_189
timestamp 1747537721
transform 1 0 18720 0 -1 15876
box -48 -56 720 834
use sg13g2_fill_1  FILLER_19_196
timestamp 1747537721
transform 1 0 19392 0 -1 15876
box -48 -56 144 834
use sg13g2_decap_4  FILLER_19_205
timestamp 1747537721
transform 1 0 20256 0 -1 15876
box -48 -56 432 834
use sg13g2_fill_1  FILLER_19_209
timestamp 1747537721
transform 1 0 20640 0 -1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_19_218
timestamp 1747537721
transform 1 0 21504 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_225
timestamp 1747537721
transform 1 0 22176 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_232
timestamp 1747537721
transform 1 0 22848 0 -1 15876
box -48 -56 720 834
use sg13g2_fill_1  FILLER_19_243
timestamp 1747537721
transform 1 0 23904 0 -1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_19_249
timestamp 1747537721
transform 1 0 24480 0 -1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_19_262
timestamp 1747537721
transform 1 0 25728 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_19_264
timestamp 1747537721
transform 1 0 25920 0 -1 15876
box -48 -56 144 834
use sg13g2_decap_4  FILLER_19_281
timestamp 1747537721
transform 1 0 27552 0 -1 15876
box -48 -56 432 834
use sg13g2_fill_1  FILLER_19_285
timestamp 1747537721
transform 1 0 27936 0 -1 15876
box -48 -56 144 834
use sg13g2_decap_4  FILLER_20_0
timestamp 1747537721
transform 1 0 576 0 1 15876
box -48 -56 432 834
use sg13g2_fill_1  FILLER_20_4
timestamp 1747537721
transform 1 0 960 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_20
timestamp 1747537721
transform 1 0 2496 0 1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_20_26
timestamp 1747537721
transform 1 0 3072 0 1 15876
box -48 -56 720 834
use sg13g2_fill_2  FILLER_20_33
timestamp 1747537721
transform 1 0 3744 0 1 15876
box -48 -56 240 834
use sg13g2_fill_2  FILLER_20_45
timestamp 1747537721
transform 1 0 4896 0 1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_20_47
timestamp 1747537721
transform 1 0 5088 0 1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_20_78
timestamp 1747537721
transform 1 0 8064 0 1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_20_80
timestamp 1747537721
transform 1 0 8256 0 1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_20_99
timestamp 1747537721
transform 1 0 10080 0 1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_20_101
timestamp 1747537721
transform 1 0 10272 0 1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_20_107
timestamp 1747537721
transform 1 0 10848 0 1 15876
box -48 -56 720 834
use sg13g2_decap_4  FILLER_20_124
timestamp 1747537721
transform 1 0 12480 0 1 15876
box -48 -56 432 834
use sg13g2_decap_4  FILLER_20_138
timestamp 1747537721
transform 1 0 13824 0 1 15876
box -48 -56 432 834
use sg13g2_fill_1  FILLER_20_142
timestamp 1747537721
transform 1 0 14208 0 1 15876
box -48 -56 144 834
use sg13g2_decap_4  FILLER_20_157
timestamp 1747537721
transform 1 0 15648 0 1 15876
box -48 -56 432 834
use sg13g2_decap_8  FILLER_20_170
timestamp 1747537721
transform 1 0 16896 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_181
timestamp 1747537721
transform 1 0 17952 0 1 15876
box -48 -56 720 834
use sg13g2_decap_4  FILLER_20_188
timestamp 1747537721
transform 1 0 18624 0 1 15876
box -48 -56 432 834
use sg13g2_fill_1  FILLER_20_192
timestamp 1747537721
transform 1 0 19008 0 1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_20_202
timestamp 1747537721
transform 1 0 19968 0 1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_20_204
timestamp 1747537721
transform 1 0 20160 0 1 15876
box -48 -56 144 834
use sg13g2_decap_4  FILLER_20_226
timestamp 1747537721
transform 1 0 22272 0 1 15876
box -48 -56 432 834
use sg13g2_fill_1  FILLER_20_230
timestamp 1747537721
transform 1 0 22656 0 1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_20_236
timestamp 1747537721
transform 1 0 23232 0 1 15876
box -48 -56 240 834
use sg13g2_decap_8  FILLER_20_252
timestamp 1747537721
transform 1 0 24768 0 1 15876
box -48 -56 720 834
use sg13g2_fill_2  FILLER_20_259
timestamp 1747537721
transform 1 0 25440 0 1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_20_261
timestamp 1747537721
transform 1 0 25632 0 1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_20_293
timestamp 1747537721
transform 1 0 28704 0 1 15876
box -48 -56 240 834
use sg13g2_decap_8  FILLER_21_26
timestamp 1747537721
transform 1 0 3072 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_21_50
timestamp 1747537721
transform 1 0 5376 0 -1 17388
box -48 -56 432 834
use sg13g2_fill_2  FILLER_21_54
timestamp 1747537721
transform 1 0 5760 0 -1 17388
box -48 -56 240 834
use sg13g2_fill_2  FILLER_21_59
timestamp 1747537721
transform 1 0 6240 0 -1 17388
box -48 -56 240 834
use sg13g2_decap_8  FILLER_21_69
timestamp 1747537721
transform 1 0 7200 0 -1 17388
box -48 -56 720 834
use sg13g2_fill_1  FILLER_21_76
timestamp 1747537721
transform 1 0 7872 0 -1 17388
box -48 -56 144 834
use sg13g2_fill_2  FILLER_21_83
timestamp 1747537721
transform 1 0 8544 0 -1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_21_85
timestamp 1747537721
transform 1 0 8736 0 -1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_21_94
timestamp 1747537721
transform 1 0 9600 0 -1 17388
box -48 -56 720 834
use sg13g2_fill_2  FILLER_21_101
timestamp 1747537721
transform 1 0 10272 0 -1 17388
box -48 -56 240 834
use sg13g2_decap_4  FILLER_21_118
timestamp 1747537721
transform 1 0 11904 0 -1 17388
box -48 -56 432 834
use sg13g2_decap_4  FILLER_21_141
timestamp 1747537721
transform 1 0 14112 0 -1 17388
box -48 -56 432 834
use sg13g2_fill_2  FILLER_21_150
timestamp 1747537721
transform 1 0 14976 0 -1 17388
box -48 -56 240 834
use sg13g2_fill_2  FILLER_21_171
timestamp 1747537721
transform 1 0 16992 0 -1 17388
box -48 -56 240 834
use sg13g2_decap_4  FILLER_21_236
timestamp 1747537721
transform 1 0 23232 0 -1 17388
box -48 -56 432 834
use sg13g2_fill_2  FILLER_21_250
timestamp 1747537721
transform 1 0 24576 0 -1 17388
box -48 -56 240 834
use sg13g2_decap_4  FILLER_21_265
timestamp 1747537721
transform 1 0 26016 0 -1 17388
box -48 -56 432 834
use sg13g2_fill_2  FILLER_21_269
timestamp 1747537721
transform 1 0 26400 0 -1 17388
box -48 -56 240 834
use sg13g2_fill_2  FILLER_21_297
timestamp 1747537721
transform 1 0 29088 0 -1 17388
box -48 -56 240 834
use sg13g2_decap_4  FILLER_21_316
timestamp 1747537721
transform 1 0 30912 0 -1 17388
box -48 -56 432 834
use sg13g2_fill_1  FILLER_21_320
timestamp 1747537721
transform 1 0 31296 0 -1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_22_0
timestamp 1747537721
transform 1 0 576 0 1 17388
box -48 -56 720 834
use sg13g2_fill_1  FILLER_22_7
timestamp 1747537721
transform 1 0 1248 0 1 17388
box -48 -56 144 834
use sg13g2_fill_2  FILLER_22_13
timestamp 1747537721
transform 1 0 1824 0 1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_22_15
timestamp 1747537721
transform 1 0 2016 0 1 17388
box -48 -56 144 834
use sg13g2_fill_2  FILLER_22_21
timestamp 1747537721
transform 1 0 2592 0 1 17388
box -48 -56 240 834
use sg13g2_decap_4  FILLER_22_48
timestamp 1747537721
transform 1 0 5184 0 1 17388
box -48 -56 432 834
use sg13g2_fill_1  FILLER_22_52
timestamp 1747537721
transform 1 0 5568 0 1 17388
box -48 -56 144 834
use sg13g2_decap_4  FILLER_22_57
timestamp 1747537721
transform 1 0 6048 0 1 17388
box -48 -56 432 834
use sg13g2_fill_1  FILLER_22_61
timestamp 1747537721
transform 1 0 6432 0 1 17388
box -48 -56 144 834
use sg13g2_fill_2  FILLER_22_74
timestamp 1747537721
transform 1 0 7680 0 1 17388
box -48 -56 240 834
use sg13g2_decap_4  FILLER_22_81
timestamp 1747537721
transform 1 0 8352 0 1 17388
box -48 -56 432 834
use sg13g2_fill_1  FILLER_22_85
timestamp 1747537721
transform 1 0 8736 0 1 17388
box -48 -56 144 834
use sg13g2_fill_2  FILLER_22_98
timestamp 1747537721
transform 1 0 9984 0 1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_22_100
timestamp 1747537721
transform 1 0 10176 0 1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_22_119
timestamp 1747537721
transform 1 0 12000 0 1 17388
box -48 -56 720 834
use sg13g2_fill_1  FILLER_22_126
timestamp 1747537721
transform 1 0 12672 0 1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_22_135
timestamp 1747537721
transform 1 0 13536 0 1 17388
box -48 -56 720 834
use sg13g2_fill_2  FILLER_22_142
timestamp 1747537721
transform 1 0 14208 0 1 17388
box -48 -56 240 834
use sg13g2_fill_2  FILLER_22_158
timestamp 1747537721
transform 1 0 15744 0 1 17388
box -48 -56 240 834
use sg13g2_decap_8  FILLER_22_169
timestamp 1747537721
transform 1 0 16800 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_185
timestamp 1747537721
transform 1 0 18336 0 1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_22_192
timestamp 1747537721
transform 1 0 19008 0 1 17388
box -48 -56 432 834
use sg13g2_decap_8  FILLER_22_201
timestamp 1747537721
transform 1 0 19872 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_208
timestamp 1747537721
transform 1 0 20544 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_215
timestamp 1747537721
transform 1 0 21216 0 1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_22_222
timestamp 1747537721
transform 1 0 21888 0 1 17388
box -48 -56 432 834
use sg13g2_fill_2  FILLER_22_226
timestamp 1747537721
transform 1 0 22272 0 1 17388
box -48 -56 240 834
use sg13g2_fill_2  FILLER_22_240
timestamp 1747537721
transform 1 0 23616 0 1 17388
box -48 -56 240 834
use sg13g2_decap_4  FILLER_22_257
timestamp 1747537721
transform 1 0 25248 0 1 17388
box -48 -56 432 834
use sg13g2_fill_2  FILLER_22_261
timestamp 1747537721
transform 1 0 25632 0 1 17388
box -48 -56 240 834
use sg13g2_decap_8  FILLER_22_267
timestamp 1747537721
transform 1 0 26208 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_274
timestamp 1747537721
transform 1 0 26880 0 1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_22_285
timestamp 1747537721
transform 1 0 27936 0 1 17388
box -48 -56 432 834
use sg13g2_decap_4  FILLER_22_293
timestamp 1747537721
transform 1 0 28704 0 1 17388
box -48 -56 432 834
use sg13g2_fill_2  FILLER_22_319
timestamp 1747537721
transform 1 0 31200 0 1 17388
box -48 -56 240 834
use sg13g2_decap_4  FILLER_23_0
timestamp 1747537721
transform 1 0 576 0 -1 18900
box -48 -56 432 834
use sg13g2_fill_1  FILLER_23_4
timestamp 1747537721
transform 1 0 960 0 -1 18900
box -48 -56 144 834
use sg13g2_fill_1  FILLER_23_30
timestamp 1747537721
transform 1 0 3456 0 -1 18900
box -48 -56 144 834
use sg13g2_fill_2  FILLER_23_65
timestamp 1747537721
transform 1 0 6816 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_23_67
timestamp 1747537721
transform 1 0 7008 0 -1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_23_94
timestamp 1747537721
transform 1 0 9600 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_4  FILLER_23_101
timestamp 1747537721
transform 1 0 10272 0 -1 18900
box -48 -56 432 834
use sg13g2_decap_8  FILLER_23_114
timestamp 1747537721
transform 1 0 11520 0 -1 18900
box -48 -56 720 834
use sg13g2_fill_1  FILLER_23_121
timestamp 1747537721
transform 1 0 12192 0 -1 18900
box -48 -56 144 834
use sg13g2_decap_4  FILLER_23_140
timestamp 1747537721
transform 1 0 14016 0 -1 18900
box -48 -56 432 834
use sg13g2_fill_2  FILLER_23_144
timestamp 1747537721
transform 1 0 14400 0 -1 18900
box -48 -56 240 834
use sg13g2_decap_8  FILLER_23_150
timestamp 1747537721
transform 1 0 14976 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_4  FILLER_23_157
timestamp 1747537721
transform 1 0 15648 0 -1 18900
box -48 -56 432 834
use sg13g2_fill_1  FILLER_23_161
timestamp 1747537721
transform 1 0 16032 0 -1 18900
box -48 -56 144 834
use sg13g2_fill_2  FILLER_23_189
timestamp 1747537721
transform 1 0 18720 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_23_191
timestamp 1747537721
transform 1 0 18912 0 -1 18900
box -48 -56 144 834
use sg13g2_decap_4  FILLER_23_207
timestamp 1747537721
transform 1 0 20448 0 -1 18900
box -48 -56 432 834
use sg13g2_decap_8  FILLER_23_223
timestamp 1747537721
transform 1 0 21984 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_237
timestamp 1747537721
transform 1 0 23328 0 -1 18900
box -48 -56 720 834
use sg13g2_fill_2  FILLER_23_244
timestamp 1747537721
transform 1 0 24000 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_2  FILLER_23_252
timestamp 1747537721
transform 1 0 24768 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_23_280
timestamp 1747537721
transform 1 0 27456 0 -1 18900
box -48 -56 144 834
use sg13g2_decap_4  FILLER_24_0
timestamp 1747537721
transform 1 0 576 0 1 18900
box -48 -56 432 834
use sg13g2_fill_1  FILLER_24_4
timestamp 1747537721
transform 1 0 960 0 1 18900
box -48 -56 144 834
use sg13g2_fill_1  FILLER_24_18
timestamp 1747537721
transform 1 0 2304 0 1 18900
box -48 -56 144 834
use sg13g2_decap_4  FILLER_24_33
timestamp 1747537721
transform 1 0 3744 0 1 18900
box -48 -56 432 834
use sg13g2_decap_8  FILLER_24_41
timestamp 1747537721
transform 1 0 4512 0 1 18900
box -48 -56 720 834
use sg13g2_fill_2  FILLER_24_48
timestamp 1747537721
transform 1 0 5184 0 1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_24_50
timestamp 1747537721
transform 1 0 5376 0 1 18900
box -48 -56 144 834
use sg13g2_fill_1  FILLER_24_62
timestamp 1747537721
transform 1 0 6528 0 1 18900
box -48 -56 144 834
use sg13g2_fill_2  FILLER_24_81
timestamp 1747537721
transform 1 0 8352 0 1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_24_83
timestamp 1747537721
transform 1 0 8544 0 1 18900
box -48 -56 144 834
use sg13g2_fill_1  FILLER_24_89
timestamp 1747537721
transform 1 0 9120 0 1 18900
box -48 -56 144 834
use sg13g2_fill_2  FILLER_24_100
timestamp 1747537721
transform 1 0 10176 0 1 18900
box -48 -56 240 834
use sg13g2_decap_4  FILLER_24_125
timestamp 1747537721
transform 1 0 12576 0 1 18900
box -48 -56 432 834
use sg13g2_fill_2  FILLER_24_140
timestamp 1747537721
transform 1 0 14016 0 1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_24_159
timestamp 1747537721
transform 1 0 15840 0 1 18900
box -48 -56 144 834
use sg13g2_fill_2  FILLER_24_164
timestamp 1747537721
transform 1 0 16320 0 1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_24_166
timestamp 1747537721
transform 1 0 16512 0 1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_24_182
timestamp 1747537721
transform 1 0 18048 0 1 18900
box -48 -56 720 834
use sg13g2_decap_4  FILLER_24_189
timestamp 1747537721
transform 1 0 18720 0 1 18900
box -48 -56 432 834
use sg13g2_fill_2  FILLER_24_198
timestamp 1747537721
transform 1 0 19584 0 1 18900
box -48 -56 240 834
use sg13g2_decap_4  FILLER_24_223
timestamp 1747537721
transform 1 0 21984 0 1 18900
box -48 -56 432 834
use sg13g2_fill_1  FILLER_24_227
timestamp 1747537721
transform 1 0 22368 0 1 18900
box -48 -56 144 834
use sg13g2_fill_2  FILLER_24_258
timestamp 1747537721
transform 1 0 25344 0 1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_24_260
timestamp 1747537721
transform 1 0 25536 0 1 18900
box -48 -56 144 834
use sg13g2_fill_1  FILLER_24_278
timestamp 1747537721
transform 1 0 27264 0 1 18900
box -48 -56 144 834
use sg13g2_fill_2  FILLER_24_293
timestamp 1747537721
transform 1 0 28704 0 1 18900
box -48 -56 240 834
use sg13g2_decap_8  FILLER_25_0
timestamp 1747537721
transform 1 0 576 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_4  FILLER_25_7
timestamp 1747537721
transform 1 0 1248 0 -1 20412
box -48 -56 432 834
use sg13g2_fill_1  FILLER_25_26
timestamp 1747537721
transform 1 0 3072 0 -1 20412
box -48 -56 144 834
use sg13g2_fill_2  FILLER_25_43
timestamp 1747537721
transform 1 0 4704 0 -1 20412
box -48 -56 240 834
use sg13g2_fill_2  FILLER_25_80
timestamp 1747537721
transform 1 0 8256 0 -1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_25_82
timestamp 1747537721
transform 1 0 8448 0 -1 20412
box -48 -56 144 834
use sg13g2_decap_4  FILLER_25_96
timestamp 1747537721
transform 1 0 9792 0 -1 20412
box -48 -56 432 834
use sg13g2_fill_2  FILLER_25_100
timestamp 1747537721
transform 1 0 10176 0 -1 20412
box -48 -56 240 834
use sg13g2_decap_8  FILLER_25_114
timestamp 1747537721
transform 1 0 11520 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_4  FILLER_25_121
timestamp 1747537721
transform 1 0 12192 0 -1 20412
box -48 -56 432 834
use sg13g2_fill_1  FILLER_25_125
timestamp 1747537721
transform 1 0 12576 0 -1 20412
box -48 -56 144 834
use sg13g2_fill_2  FILLER_25_140
timestamp 1747537721
transform 1 0 14016 0 -1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_25_142
timestamp 1747537721
transform 1 0 14208 0 -1 20412
box -48 -56 144 834
use sg13g2_fill_2  FILLER_25_162
timestamp 1747537721
transform 1 0 16128 0 -1 20412
box -48 -56 240 834
use sg13g2_fill_2  FILLER_25_183
timestamp 1747537721
transform 1 0 18144 0 -1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_25_185
timestamp 1747537721
transform 1 0 18336 0 -1 20412
box -48 -56 144 834
use sg13g2_fill_2  FILLER_25_191
timestamp 1747537721
transform 1 0 18912 0 -1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_25_193
timestamp 1747537721
transform 1 0 19104 0 -1 20412
box -48 -56 144 834
use sg13g2_fill_1  FILLER_25_198
timestamp 1747537721
transform 1 0 19584 0 -1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_25_220
timestamp 1747537721
transform 1 0 21696 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_227
timestamp 1747537721
transform 1 0 22368 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_234
timestamp 1747537721
transform 1 0 23040 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_241
timestamp 1747537721
transform 1 0 23712 0 -1 20412
box -48 -56 720 834
use sg13g2_fill_2  FILLER_25_283
timestamp 1747537721
transform 1 0 27744 0 -1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_25_320
timestamp 1747537721
transform 1 0 31296 0 -1 20412
box -48 -56 144 834
use sg13g2_fill_2  FILLER_26_34
timestamp 1747537721
transform 1 0 3840 0 1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_26_36
timestamp 1747537721
transform 1 0 4032 0 1 20412
box -48 -56 144 834
use sg13g2_decap_4  FILLER_26_45
timestamp 1747537721
transform 1 0 4896 0 1 20412
box -48 -56 432 834
use sg13g2_decap_4  FILLER_26_54
timestamp 1747537721
transform 1 0 5760 0 1 20412
box -48 -56 432 834
use sg13g2_decap_8  FILLER_26_67
timestamp 1747537721
transform 1 0 7008 0 1 20412
box -48 -56 720 834
use sg13g2_fill_2  FILLER_26_74
timestamp 1747537721
transform 1 0 7680 0 1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_26_76
timestamp 1747537721
transform 1 0 7872 0 1 20412
box -48 -56 144 834
use sg13g2_decap_4  FILLER_26_82
timestamp 1747537721
transform 1 0 8448 0 1 20412
box -48 -56 432 834
use sg13g2_fill_1  FILLER_26_86
timestamp 1747537721
transform 1 0 8832 0 1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_26_91
timestamp 1747537721
transform 1 0 9312 0 1 20412
box -48 -56 720 834
use sg13g2_fill_2  FILLER_26_98
timestamp 1747537721
transform 1 0 9984 0 1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_26_100
timestamp 1747537721
transform 1 0 10176 0 1 20412
box -48 -56 144 834
use sg13g2_fill_1  FILLER_26_122
timestamp 1747537721
transform 1 0 12288 0 1 20412
box -48 -56 144 834
use sg13g2_fill_1  FILLER_26_159
timestamp 1747537721
transform 1 0 15840 0 1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_26_165
timestamp 1747537721
transform 1 0 16416 0 1 20412
box -48 -56 720 834
use sg13g2_fill_1  FILLER_26_172
timestamp 1747537721
transform 1 0 17088 0 1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_26_186
timestamp 1747537721
transform 1 0 18432 0 1 20412
box -48 -56 720 834
use sg13g2_decap_4  FILLER_26_202
timestamp 1747537721
transform 1 0 19968 0 1 20412
box -48 -56 432 834
use sg13g2_fill_2  FILLER_26_292
timestamp 1747537721
transform 1 0 28608 0 1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_26_294
timestamp 1747537721
transform 1 0 28800 0 1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_27_0
timestamp 1747537721
transform 1 0 576 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_27_7
timestamp 1747537721
transform 1 0 1248 0 -1 21924
box -48 -56 432 834
use sg13g2_decap_8  FILLER_27_24
timestamp 1747537721
transform 1 0 2880 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_27_31
timestamp 1747537721
transform 1 0 3552 0 -1 21924
box -48 -56 432 834
use sg13g2_fill_1  FILLER_27_35
timestamp 1747537721
transform 1 0 3936 0 -1 21924
box -48 -56 144 834
use sg13g2_decap_8  FILLER_27_76
timestamp 1747537721
transform 1 0 7872 0 -1 21924
box -48 -56 720 834
use sg13g2_fill_1  FILLER_27_83
timestamp 1747537721
transform 1 0 8544 0 -1 21924
box -48 -56 144 834
use sg13g2_decap_8  FILLER_27_100
timestamp 1747537721
transform 1 0 10176 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_107
timestamp 1747537721
transform 1 0 10848 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_27_124
timestamp 1747537721
transform 1 0 12480 0 -1 21924
box -48 -56 432 834
use sg13g2_fill_1  FILLER_27_128
timestamp 1747537721
transform 1 0 12864 0 -1 21924
box -48 -56 144 834
use sg13g2_decap_8  FILLER_27_137
timestamp 1747537721
transform 1 0 13728 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_148
timestamp 1747537721
transform 1 0 14784 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_27_155
timestamp 1747537721
transform 1 0 15456 0 -1 21924
box -48 -56 432 834
use sg13g2_fill_2  FILLER_27_159
timestamp 1747537721
transform 1 0 15840 0 -1 21924
box -48 -56 240 834
use sg13g2_decap_4  FILLER_27_186
timestamp 1747537721
transform 1 0 18432 0 -1 21924
box -48 -56 432 834
use sg13g2_fill_1  FILLER_27_210
timestamp 1747537721
transform 1 0 20736 0 -1 21924
box -48 -56 144 834
use sg13g2_fill_2  FILLER_27_219
timestamp 1747537721
transform 1 0 21600 0 -1 21924
box -48 -56 240 834
use sg13g2_fill_2  FILLER_27_225
timestamp 1747537721
transform 1 0 22176 0 -1 21924
box -48 -56 240 834
use sg13g2_decap_8  FILLER_27_234
timestamp 1747537721
transform 1 0 23040 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_241
timestamp 1747537721
transform 1 0 23712 0 -1 21924
box -48 -56 720 834
use sg13g2_fill_2  FILLER_27_248
timestamp 1747537721
transform 1 0 24384 0 -1 21924
box -48 -56 240 834
use sg13g2_fill_2  FILLER_27_274
timestamp 1747537721
transform 1 0 26880 0 -1 21924
box -48 -56 240 834
use sg13g2_fill_2  FILLER_27_293
timestamp 1747537721
transform 1 0 28704 0 -1 21924
box -48 -56 240 834
use sg13g2_fill_2  FILLER_27_319
timestamp 1747537721
transform 1 0 31200 0 -1 21924
box -48 -56 240 834
use sg13g2_fill_2  FILLER_28_0
timestamp 1747537721
transform 1 0 576 0 1 21924
box -48 -56 240 834
use sg13g2_fill_2  FILLER_28_28
timestamp 1747537721
transform 1 0 3264 0 1 21924
box -48 -56 240 834
use sg13g2_fill_2  FILLER_28_43
timestamp 1747537721
transform 1 0 4704 0 1 21924
box -48 -56 240 834
use sg13g2_fill_2  FILLER_28_58
timestamp 1747537721
transform 1 0 6144 0 1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_28_60
timestamp 1747537721
transform 1 0 6336 0 1 21924
box -48 -56 144 834
use sg13g2_decap_8  FILLER_28_65
timestamp 1747537721
transform 1 0 6816 0 1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_28_75
timestamp 1747537721
transform 1 0 7776 0 1 21924
box -48 -56 432 834
use sg13g2_fill_2  FILLER_28_79
timestamp 1747537721
transform 1 0 8160 0 1 21924
box -48 -56 240 834
use sg13g2_decap_8  FILLER_28_86
timestamp 1747537721
transform 1 0 8832 0 1 21924
box -48 -56 720 834
use sg13g2_fill_2  FILLER_28_93
timestamp 1747537721
transform 1 0 9504 0 1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_28_95
timestamp 1747537721
transform 1 0 9696 0 1 21924
box -48 -56 144 834
use sg13g2_decap_4  FILLER_28_115
timestamp 1747537721
transform 1 0 11616 0 1 21924
box -48 -56 432 834
use sg13g2_fill_1  FILLER_28_119
timestamp 1747537721
transform 1 0 12000 0 1 21924
box -48 -56 144 834
use sg13g2_decap_8  FILLER_28_133
timestamp 1747537721
transform 1 0 13344 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_140
timestamp 1747537721
transform 1 0 14016 0 1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_28_155
timestamp 1747537721
transform 1 0 15456 0 1 21924
box -48 -56 432 834
use sg13g2_fill_1  FILLER_28_159
timestamp 1747537721
transform 1 0 15840 0 1 21924
box -48 -56 144 834
use sg13g2_decap_8  FILLER_28_168
timestamp 1747537721
transform 1 0 16704 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_175
timestamp 1747537721
transform 1 0 17376 0 1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_28_182
timestamp 1747537721
transform 1 0 18048 0 1 21924
box -48 -56 432 834
use sg13g2_fill_1  FILLER_28_186
timestamp 1747537721
transform 1 0 18432 0 1 21924
box -48 -56 144 834
use sg13g2_decap_8  FILLER_28_197
timestamp 1747537721
transform 1 0 19488 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_204
timestamp 1747537721
transform 1 0 20160 0 1 21924
box -48 -56 720 834
use sg13g2_fill_2  FILLER_28_211
timestamp 1747537721
transform 1 0 20832 0 1 21924
box -48 -56 240 834
use sg13g2_decap_4  FILLER_28_242
timestamp 1747537721
transform 1 0 23808 0 1 21924
box -48 -56 432 834
use sg13g2_fill_1  FILLER_28_246
timestamp 1747537721
transform 1 0 24192 0 1 21924
box -48 -56 144 834
use sg13g2_fill_2  FILLER_28_258
timestamp 1747537721
transform 1 0 25344 0 1 21924
box -48 -56 240 834
use sg13g2_fill_2  FILLER_28_267
timestamp 1747537721
transform 1 0 26208 0 1 21924
box -48 -56 240 834
use sg13g2_fill_2  FILLER_28_283
timestamp 1747537721
transform 1 0 27744 0 1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_28_302
timestamp 1747537721
transform 1 0 29568 0 1 21924
box -48 -56 144 834
use sg13g2_decap_8  FILLER_29_0
timestamp 1747537721
transform 1 0 576 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_4  FILLER_29_7
timestamp 1747537721
transform 1 0 1248 0 -1 23436
box -48 -56 432 834
use sg13g2_fill_2  FILLER_29_11
timestamp 1747537721
transform 1 0 1632 0 -1 23436
box -48 -56 240 834
use sg13g2_decap_8  FILLER_29_34
timestamp 1747537721
transform 1 0 3840 0 -1 23436
box -48 -56 720 834
use sg13g2_fill_1  FILLER_29_41
timestamp 1747537721
transform 1 0 4512 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_29_80
timestamp 1747537721
transform 1 0 8256 0 -1 23436
box -48 -56 144 834
use sg13g2_decap_8  FILLER_29_157
timestamp 1747537721
transform 1 0 15648 0 -1 23436
box -48 -56 720 834
use sg13g2_fill_2  FILLER_29_223
timestamp 1747537721
transform 1 0 21984 0 -1 23436
box -48 -56 240 834
use sg13g2_decap_4  FILLER_29_234
timestamp 1747537721
transform 1 0 23040 0 -1 23436
box -48 -56 432 834
use sg13g2_fill_2  FILLER_29_242
timestamp 1747537721
transform 1 0 23808 0 -1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_29_244
timestamp 1747537721
transform 1 0 24000 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_29_252
timestamp 1747537721
transform 1 0 24768 0 -1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_29_266
timestamp 1747537721
transform 1 0 26112 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_29_275
timestamp 1747537721
transform 1 0 26976 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_29_280
timestamp 1747537721
transform 1 0 27456 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_30_41
timestamp 1747537721
transform 1 0 4512 0 1 23436
box -48 -56 240 834
use sg13g2_decap_4  FILLER_30_53
timestamp 1747537721
transform 1 0 5664 0 1 23436
box -48 -56 432 834
use sg13g2_fill_1  FILLER_30_57
timestamp 1747537721
transform 1 0 6048 0 1 23436
box -48 -56 144 834
use sg13g2_decap_4  FILLER_30_71
timestamp 1747537721
transform 1 0 7392 0 1 23436
box -48 -56 432 834
use sg13g2_fill_1  FILLER_30_75
timestamp 1747537721
transform 1 0 7776 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_81
timestamp 1747537721
transform 1 0 8352 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_133
timestamp 1747537721
transform 1 0 13344 0 1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_30_148
timestamp 1747537721
transform 1 0 14784 0 1 23436
box -48 -56 240 834
use sg13g2_decap_8  FILLER_30_203
timestamp 1747537721
transform 1 0 20064 0 1 23436
box -48 -56 720 834
use sg13g2_fill_2  FILLER_30_264
timestamp 1747537721
transform 1 0 25920 0 1 23436
box -48 -56 240 834
use sg13g2_fill_2  FILLER_30_275
timestamp 1747537721
transform 1 0 26976 0 1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_30_294
timestamp 1747537721
transform 1 0 28800 0 1 23436
box -48 -56 144 834
use sg13g2_decap_8  FILLER_31_0
timestamp 1747537721
transform 1 0 576 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_4  FILLER_31_7
timestamp 1747537721
transform 1 0 1248 0 -1 24948
box -48 -56 432 834
use sg13g2_fill_1  FILLER_31_15
timestamp 1747537721
transform 1 0 2016 0 -1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_31_29
timestamp 1747537721
transform 1 0 3360 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_4  FILLER_31_91
timestamp 1747537721
transform 1 0 9312 0 -1 24948
box -48 -56 432 834
use sg13g2_fill_2  FILLER_31_111
timestamp 1747537721
transform 1 0 11232 0 -1 24948
box -48 -56 240 834
use sg13g2_decap_4  FILLER_31_163
timestamp 1747537721
transform 1 0 16224 0 -1 24948
box -48 -56 432 834
use sg13g2_fill_2  FILLER_31_176
timestamp 1747537721
transform 1 0 17472 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_31_190
timestamp 1747537721
transform 1 0 18816 0 -1 24948
box -48 -56 144 834
use sg13g2_decap_4  FILLER_31_208
timestamp 1747537721
transform 1 0 20544 0 -1 24948
box -48 -56 432 834
use sg13g2_fill_2  FILLER_31_212
timestamp 1747537721
transform 1 0 20928 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_31_223
timestamp 1747537721
transform 1 0 21984 0 -1 24948
box -48 -56 144 834
use sg13g2_decap_4  FILLER_31_241
timestamp 1747537721
transform 1 0 23712 0 -1 24948
box -48 -56 432 834
use sg13g2_fill_2  FILLER_31_245
timestamp 1747537721
transform 1 0 24096 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_2  FILLER_31_253
timestamp 1747537721
transform 1 0 24864 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_2  FILLER_31_260
timestamp 1747537721
transform 1 0 25536 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_2  FILLER_31_272
timestamp 1747537721
transform 1 0 26688 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_2  FILLER_31_292
timestamp 1747537721
transform 1 0 28608 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_31_320
timestamp 1747537721
transform 1 0 31296 0 -1 24948
box -48 -56 144 834
use sg13g2_decap_4  FILLER_32_0
timestamp 1747537721
transform 1 0 576 0 1 24948
box -48 -56 432 834
use sg13g2_fill_2  FILLER_32_4
timestamp 1747537721
transform 1 0 960 0 1 24948
box -48 -56 240 834
use sg13g2_decap_8  FILLER_32_32
timestamp 1747537721
transform 1 0 3648 0 1 24948
box -48 -56 720 834
use sg13g2_fill_1  FILLER_32_39
timestamp 1747537721
transform 1 0 4320 0 1 24948
box -48 -56 144 834
use sg13g2_fill_1  FILLER_32_53
timestamp 1747537721
transform 1 0 5664 0 1 24948
box -48 -56 144 834
use sg13g2_fill_2  FILLER_32_63
timestamp 1747537721
transform 1 0 6624 0 1 24948
box -48 -56 240 834
use sg13g2_decap_4  FILLER_32_73
timestamp 1747537721
transform 1 0 7584 0 1 24948
box -48 -56 432 834
use sg13g2_fill_1  FILLER_32_77
timestamp 1747537721
transform 1 0 7968 0 1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_32_83
timestamp 1747537721
transform 1 0 8544 0 1 24948
box -48 -56 720 834
use sg13g2_decap_4  FILLER_32_98
timestamp 1747537721
transform 1 0 9984 0 1 24948
box -48 -56 432 834
use sg13g2_fill_1  FILLER_32_102
timestamp 1747537721
transform 1 0 10368 0 1 24948
box -48 -56 144 834
use sg13g2_fill_1  FILLER_32_121
timestamp 1747537721
transform 1 0 12192 0 1 24948
box -48 -56 144 834
use sg13g2_fill_2  FILLER_32_127
timestamp 1747537721
transform 1 0 12768 0 1 24948
box -48 -56 240 834
use sg13g2_decap_8  FILLER_32_133
timestamp 1747537721
transform 1 0 13344 0 1 24948
box -48 -56 720 834
use sg13g2_fill_2  FILLER_32_140
timestamp 1747537721
transform 1 0 14016 0 1 24948
box -48 -56 240 834
use sg13g2_fill_2  FILLER_32_150
timestamp 1747537721
transform 1 0 14976 0 1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_32_152
timestamp 1747537721
transform 1 0 15168 0 1 24948
box -48 -56 144 834
use sg13g2_fill_2  FILLER_32_170
timestamp 1747537721
transform 1 0 16896 0 1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_32_200
timestamp 1747537721
transform 1 0 19776 0 1 24948
box -48 -56 144 834
use sg13g2_fill_2  FILLER_32_240
timestamp 1747537721
transform 1 0 23616 0 1 24948
box -48 -56 240 834
use sg13g2_fill_2  FILLER_32_278
timestamp 1747537721
transform 1 0 27264 0 1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_32_280
timestamp 1747537721
transform 1 0 27456 0 1 24948
box -48 -56 144 834
use sg13g2_fill_1  FILLER_32_289
timestamp 1747537721
transform 1 0 28320 0 1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_33_0
timestamp 1747537721
transform 1 0 576 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_4  FILLER_33_7
timestamp 1747537721
transform 1 0 1248 0 -1 26460
box -48 -56 432 834
use sg13g2_fill_2  FILLER_33_44
timestamp 1747537721
transform 1 0 4800 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_2  FILLER_33_50
timestamp 1747537721
transform 1 0 5376 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_2  FILLER_33_91
timestamp 1747537721
transform 1 0 9312 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_33_93
timestamp 1747537721
transform 1 0 9504 0 -1 26460
box -48 -56 144 834
use sg13g2_fill_2  FILLER_33_107
timestamp 1747537721
transform 1 0 10848 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_2  FILLER_33_114
timestamp 1747537721
transform 1 0 11520 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_33_153
timestamp 1747537721
transform 1 0 15264 0 -1 26460
box -48 -56 144 834
use sg13g2_fill_2  FILLER_33_171
timestamp 1747537721
transform 1 0 16992 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_33_173
timestamp 1747537721
transform 1 0 17184 0 -1 26460
box -48 -56 144 834
use sg13g2_fill_2  FILLER_33_197
timestamp 1747537721
transform 1 0 19488 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_2  FILLER_33_222
timestamp 1747537721
transform 1 0 21888 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_33_224
timestamp 1747537721
transform 1 0 22080 0 -1 26460
box -48 -56 144 834
use sg13g2_decap_8  FILLER_33_229
timestamp 1747537721
transform 1 0 22560 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_4  FILLER_33_236
timestamp 1747537721
transform 1 0 23232 0 -1 26460
box -48 -56 432 834
use sg13g2_fill_2  FILLER_33_240
timestamp 1747537721
transform 1 0 23616 0 -1 26460
box -48 -56 240 834
use sg13g2_decap_4  FILLER_33_247
timestamp 1747537721
transform 1 0 24288 0 -1 26460
box -48 -56 432 834
use sg13g2_fill_2  FILLER_33_256
timestamp 1747537721
transform 1 0 25152 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_33_258
timestamp 1747537721
transform 1 0 25344 0 -1 26460
box -48 -56 144 834
use sg13g2_fill_1  FILLER_33_268
timestamp 1747537721
transform 1 0 26304 0 -1 26460
box -48 -56 144 834
use sg13g2_fill_1  FILLER_33_291
timestamp 1747537721
transform 1 0 28512 0 -1 26460
box -48 -56 144 834
use sg13g2_fill_2  FILLER_33_318
timestamp 1747537721
transform 1 0 31104 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_33_320
timestamp 1747537721
transform 1 0 31296 0 -1 26460
box -48 -56 144 834
use sg13g2_decap_8  FILLER_34_0
timestamp 1747537721
transform 1 0 576 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_7
timestamp 1747537721
transform 1 0 1248 0 1 26460
box -48 -56 720 834
use sg13g2_decap_4  FILLER_34_14
timestamp 1747537721
transform 1 0 1920 0 1 26460
box -48 -56 432 834
use sg13g2_fill_2  FILLER_34_18
timestamp 1747537721
transform 1 0 2304 0 1 26460
box -48 -56 240 834
use sg13g2_fill_2  FILLER_34_61
timestamp 1747537721
transform 1 0 6432 0 1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_34_89
timestamp 1747537721
transform 1 0 9120 0 1 26460
box -48 -56 144 834
use sg13g2_decap_4  FILLER_34_94
timestamp 1747537721
transform 1 0 9600 0 1 26460
box -48 -56 432 834
use sg13g2_fill_2  FILLER_34_98
timestamp 1747537721
transform 1 0 9984 0 1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_34_135
timestamp 1747537721
transform 1 0 13536 0 1 26460
box -48 -56 144 834
use sg13g2_fill_1  FILLER_34_154
timestamp 1747537721
transform 1 0 15360 0 1 26460
box -48 -56 144 834
use sg13g2_fill_2  FILLER_34_159
timestamp 1747537721
transform 1 0 15840 0 1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_34_198
timestamp 1747537721
transform 1 0 19584 0 1 26460
box -48 -56 144 834
use sg13g2_decap_8  FILLER_34_225
timestamp 1747537721
transform 1 0 22176 0 1 26460
box -48 -56 720 834
use sg13g2_fill_2  FILLER_34_232
timestamp 1747537721
transform 1 0 22848 0 1 26460
box -48 -56 240 834
use sg13g2_decap_8  FILLER_35_0
timestamp 1747537721
transform 1 0 576 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_7
timestamp 1747537721
transform 1 0 1248 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_14
timestamp 1747537721
transform 1 0 1920 0 -1 27972
box -48 -56 720 834
use sg13g2_fill_2  FILLER_35_21
timestamp 1747537721
transform 1 0 2592 0 -1 27972
box -48 -56 240 834
use sg13g2_decap_4  FILLER_35_105
timestamp 1747537721
transform 1 0 10656 0 -1 27972
box -48 -56 432 834
use sg13g2_fill_1  FILLER_35_109
timestamp 1747537721
transform 1 0 11040 0 -1 27972
box -48 -56 144 834
use sg13g2_fill_1  FILLER_35_143
timestamp 1747537721
transform 1 0 14304 0 -1 27972
box -48 -56 144 834
use sg13g2_decap_4  FILLER_35_173
timestamp 1747537721
transform 1 0 17184 0 -1 27972
box -48 -56 432 834
use sg13g2_fill_1  FILLER_35_177
timestamp 1747537721
transform 1 0 17568 0 -1 27972
box -48 -56 144 834
use sg13g2_fill_2  FILLER_35_208
timestamp 1747537721
transform 1 0 20544 0 -1 27972
box -48 -56 240 834
use sg13g2_decap_8  FILLER_35_214
timestamp 1747537721
transform 1 0 21120 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_4  FILLER_35_221
timestamp 1747537721
transform 1 0 21792 0 -1 27972
box -48 -56 432 834
use sg13g2_fill_1  FILLER_35_225
timestamp 1747537721
transform 1 0 22176 0 -1 27972
box -48 -56 144 834
use sg13g2_fill_2  FILLER_35_252
timestamp 1747537721
transform 1 0 24768 0 -1 27972
box -48 -56 240 834
use sg13g2_dlygate4sd3_1  hold1
timestamp 1747537721
transform -1 0 13344 0 1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold2
timestamp 1747537721
transform -1 0 6624 0 1 24948
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold3
timestamp 1747537721
transform 1 0 27072 0 1 15876
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold4
timestamp 1747537721
transform -1 0 3456 0 -1 14364
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold5
timestamp 1747537721
transform -1 0 2496 0 1 14364
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold6
timestamp 1747537721
transform -1 0 29568 0 -1 20412
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold7
timestamp 1747537721
transform 1 0 29952 0 1 17388
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold8
timestamp 1747537721
transform 1 0 22176 0 -1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold9
timestamp 1747537721
transform 1 0 16032 0 1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold10
timestamp 1747537721
transform 1 0 14496 0 1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold11
timestamp 1747537721
transform -1 0 30144 0 -1 17388
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold12
timestamp 1747537721
transform 1 0 7392 0 1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold13
timestamp 1747537721
transform 1 0 12672 0 1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold14
timestamp 1747537721
transform 1 0 17856 0 1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold15
timestamp 1747537721
transform 1 0 15264 0 1 24948
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold16
timestamp 1747537721
transform -1 0 30528 0 1 21924
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold17
timestamp 1747537721
transform 1 0 28032 0 -1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold18
timestamp 1747537721
transform -1 0 16224 0 -1 24948
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold19
timestamp 1747537721
transform -1 0 7008 0 1 20412
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold20
timestamp 1747537721
transform 1 0 4896 0 1 21924
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold21
timestamp 1747537721
transform 1 0 26400 0 1 18900
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold22
timestamp 1747537721
transform -1 0 28224 0 1 18900
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold23
timestamp 1747537721
transform -1 0 14304 0 1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold24
timestamp 1747537721
transform -1 0 12672 0 1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold25
timestamp 1747537721
transform 1 0 10944 0 1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold26
timestamp 1747537721
transform -1 0 7008 0 1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold27
timestamp 1747537721
transform -1 0 6432 0 1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold28
timestamp 1747537721
transform -1 0 21888 0 -1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold29
timestamp 1747537721
transform -1 0 20544 0 -1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold30
timestamp 1747537721
transform -1 0 22944 0 -1 24948
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold31
timestamp 1747537721
transform -1 0 21984 0 -1 24948
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold32
timestamp 1747537721
transform -1 0 29760 0 -1 21924
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold33
timestamp 1747537721
transform -1 0 29568 0 1 21924
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold34
timestamp 1747537721
transform -1 0 19584 0 1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold35
timestamp 1747537721
transform -1 0 18720 0 1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold36
timestamp 1747537721
transform -1 0 29952 0 -1 2268
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold37
timestamp 1747537721
transform -1 0 30240 0 1 2268
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold38
timestamp 1747537721
transform 1 0 30048 0 -1 2268
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold39
timestamp 1747537721
transform 1 0 28896 0 1 14364
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold40
timestamp 1747537721
transform -1 0 28896 0 -1 15876
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold41
timestamp 1747537721
transform -1 0 29472 0 1 3780
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold42
timestamp 1747537721
transform -1 0 15168 0 -1 20412
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold43
timestamp 1747537721
transform -1 0 29760 0 1 8316
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold44
timestamp 1747537721
transform -1 0 10848 0 1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold45
timestamp 1747537721
transform -1 0 27648 0 1 756
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold46
timestamp 1747537721
transform -1 0 26016 0 1 756
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold47
timestamp 1747537721
transform -1 0 29664 0 -1 24948
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold48
timestamp 1747537721
transform 1 0 1632 0 -1 21924
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold49
timestamp 1747537721
transform -1 0 30432 0 -1 20412
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold50
timestamp 1747537721
transform 1 0 2208 0 -1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold51
timestamp 1747537721
transform 1 0 21696 0 1 9828
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold52
timestamp 1747537721
transform 1 0 23424 0 1 9828
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold53
timestamp 1747537721
transform -1 0 30912 0 -1 24948
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold54
timestamp 1747537721
transform 1 0 2112 0 -1 24948
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold55
timestamp 1747537721
transform 1 0 28032 0 1 8316
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold56
timestamp 1747537721
transform -1 0 28224 0 1 9828
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold57
timestamp 1747537721
transform 1 0 10848 0 1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold58
timestamp 1747537721
transform 1 0 23808 0 1 20412
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold59
timestamp 1747537721
transform 1 0 28992 0 1 9828
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold60
timestamp 1747537721
transform 1 0 27936 0 -1 27972
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold61
timestamp 1747537721
transform 1 0 28032 0 -1 11340
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold62
timestamp 1747537721
transform 1 0 28800 0 1 11340
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold63
timestamp 1747537721
transform -1 0 6144 0 1 2268
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold64
timestamp 1747537721
transform -1 0 30624 0 1 14364
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold65
timestamp 1747537721
transform 1 0 9120 0 1 756
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold66
timestamp 1747537721
transform -1 0 6528 0 -1 2268
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold67
timestamp 1747537721
transform -1 0 25632 0 1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold68
timestamp 1747537721
transform -1 0 3072 0 -1 11340
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold69
timestamp 1747537721
transform 1 0 22560 0 1 9828
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold70
timestamp 1747537721
transform -1 0 29952 0 -1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold71
timestamp 1747537721
transform 1 0 26784 0 1 11340
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold72
timestamp 1747537721
transform -1 0 24576 0 1 11340
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold73
timestamp 1747537721
transform 1 0 21600 0 1 2268
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold74
timestamp 1747537721
transform -1 0 25440 0 -1 2268
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold75
timestamp 1747537721
transform -1 0 4224 0 1 11340
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold76
timestamp 1747537721
transform 1 0 19968 0 1 756
box -48 -56 912 834
use sg13g2_buf_1  input1
timestamp 1747537721
transform -1 0 26784 0 -1 26460
box -48 -56 432 834
use sg13g2_buf_1  input2
timestamp 1747537721
transform -1 0 31008 0 -1 27972
box -48 -56 432 834
use sg13g2_buf_2  input3
timestamp 1747537721
transform -1 0 30240 0 -1 27972
box -48 -56 528 834
use sg13g2_buf_2  input4
timestamp 1747537721
transform -1 0 29760 0 -1 27972
box -48 -56 528 834
use sg13g2_buf_2  input5
timestamp 1747537721
transform -1 0 29280 0 -1 27972
box -48 -56 528 834
use sg13g2_buf_2  input6
timestamp 1747537721
transform -1 0 27744 0 1 26460
box -48 -56 528 834
use sg13g2_buf_2  input7
timestamp 1747537721
transform -1 0 25920 0 -1 26460
box -48 -56 528 834
use sg13g2_buf_2  input8
timestamp 1747537721
transform -1 0 25152 0 -1 26460
box -48 -56 528 834
use sg13g2_buf_2  input9
timestamp 1747537721
transform -1 0 26784 0 1 26460
box -48 -56 528 834
use sg13g2_buf_1  input10
timestamp 1747537721
transform -1 0 23424 0 1 26460
box -48 -56 432 834
<< labels >>
flabel metal5 s 27638 712 28078 28016 0 FreeSans 3200 90 0 0 VGND
port 1 nsew
flabel metal5 s 19864 712 20304 28016 0 FreeSans 3200 90 0 0 VGND
port 1 nsew
flabel metal5 s 12090 712 12530 28016 0 FreeSans 3200 90 0 0 VGND
port 1 nsew
flabel metal5 s 4316 712 4756 28016 0 FreeSans 3200 90 0 0 VGND
port 1 nsew
flabel metal5 s 26398 712 26838 28016 0 FreeSans 3200 90 0 0 VPWR
port 2 nsew
flabel metal5 s 18624 712 19064 28016 0 FreeSans 3200 90 0 0 VPWR
port 2 nsew
flabel metal5 s 10850 712 11290 28016 0 FreeSans 3200 90 0 0 VPWR
port 2 nsew
flabel metal5 s 3076 712 3516 28016 0 FreeSans 3200 90 0 0 VPWR
port 2 nsew
flabel metal3 s 11576 28600 11656 29000 0 FreeSans 400 90 0 0 b6
port 3 nsew
flabel metal3 s 14648 28600 14728 29000 0 FreeSans 400 90 0 0 b7
port 4 nsew
flabel metal3 s 30008 28600 30088 29000 0 FreeSans 400 90 0 0 clk
port 5 nsew
flabel metal2 s 0 8864 400 8944 0 FreeSans 400 0 0 0 db[0]
port 6 nsew
flabel metal2 s 0 8444 400 8524 0 FreeSans 400 0 0 0 db[1]
port 7 nsew
flabel metal2 s 0 8024 400 8104 0 FreeSans 400 0 0 0 db[2]
port 8 nsew
flabel metal2 s 0 7604 400 7684 0 FreeSans 400 0 0 0 db[3]
port 9 nsew
flabel metal2 s 0 7184 400 7264 0 FreeSans 400 0 0 0 db[4]
port 10 nsew
flabel metal2 s 0 6764 400 6844 0 FreeSans 400 0 0 0 db[5]
port 11 nsew
flabel metal2 s 0 6344 400 6424 0 FreeSans 400 0 0 0 db[6]
port 12 nsew
flabel metal2 s 0 5924 400 6004 0 FreeSans 400 0 0 0 db[7]
port 13 nsew
flabel metal2 s 0 15584 400 15664 0 FreeSans 400 0 0 0 dg[0]
port 14 nsew
flabel metal2 s 0 15164 400 15244 0 FreeSans 400 0 0 0 dg[1]
port 15 nsew
flabel metal2 s 0 14744 400 14824 0 FreeSans 400 0 0 0 dg[2]
port 16 nsew
flabel metal2 s 0 14324 400 14404 0 FreeSans 400 0 0 0 dg[3]
port 17 nsew
flabel metal2 s 0 13904 400 13984 0 FreeSans 400 0 0 0 dg[4]
port 18 nsew
flabel metal2 s 0 13484 400 13564 0 FreeSans 400 0 0 0 dg[5]
port 19 nsew
flabel metal2 s 0 13064 400 13144 0 FreeSans 400 0 0 0 dg[6]
port 20 nsew
flabel metal2 s 0 12644 400 12724 0 FreeSans 400 0 0 0 dg[7]
port 21 nsew
flabel metal2 s 0 22304 400 22384 0 FreeSans 400 0 0 0 dr[0]
port 22 nsew
flabel metal2 s 0 21884 400 21964 0 FreeSans 400 0 0 0 dr[1]
port 23 nsew
flabel metal2 s 0 21464 400 21544 0 FreeSans 400 0 0 0 dr[2]
port 24 nsew
flabel metal2 s 0 21044 400 21124 0 FreeSans 400 0 0 0 dr[3]
port 25 nsew
flabel metal2 s 0 20624 400 20704 0 FreeSans 400 0 0 0 dr[4]
port 26 nsew
flabel metal2 s 0 20204 400 20284 0 FreeSans 400 0 0 0 dr[5]
port 27 nsew
flabel metal2 s 0 19784 400 19864 0 FreeSans 400 0 0 0 dr[6]
port 28 nsew
flabel metal2 s 0 19364 400 19444 0 FreeSans 400 0 0 0 dr[7]
port 29 nsew
flabel metal3 s 30776 28600 30856 29000 0 FreeSans 400 90 0 0 ena
port 30 nsew
flabel metal3 s 12344 28600 12424 29000 0 FreeSans 400 90 0 0 g6
port 31 nsew
flabel metal3 s 15416 28600 15496 29000 0 FreeSans 400 90 0 0 g7
port 32 nsew
flabel metal3 s 9272 28600 9352 29000 0 FreeSans 400 90 0 0 hblank
port 33 nsew
flabel metal3 s 10808 28600 10888 29000 0 FreeSans 400 90 0 0 hsync
port 34 nsew
flabel metal3 s 13112 28600 13192 29000 0 FreeSans 400 90 0 0 r6
port 35 nsew
flabel metal3 s 16184 28600 16264 29000 0 FreeSans 400 90 0 0 r7
port 36 nsew
flabel metal3 s 29240 28600 29320 29000 0 FreeSans 400 90 0 0 rst_n
port 37 nsew
flabel metal3 s 28472 28600 28552 29000 0 FreeSans 400 90 0 0 ui_in[0]
port 38 nsew
flabel metal3 s 27704 28600 27784 29000 0 FreeSans 400 90 0 0 ui_in[1]
port 39 nsew
flabel metal3 s 26936 28600 27016 29000 0 FreeSans 400 90 0 0 ui_in[2]
port 40 nsew
flabel metal3 s 26168 28600 26248 29000 0 FreeSans 400 90 0 0 ui_in[3]
port 41 nsew
flabel metal3 s 25400 28600 25480 29000 0 FreeSans 400 90 0 0 ui_in[4]
port 42 nsew
flabel metal3 s 24632 28600 24712 29000 0 FreeSans 400 90 0 0 ui_in[5]
port 43 nsew
flabel metal3 s 23864 28600 23944 29000 0 FreeSans 400 90 0 0 ui_in[6]
port 44 nsew
flabel metal3 s 23096 28600 23176 29000 0 FreeSans 400 90 0 0 ui_in[7]
port 45 nsew
flabel metal3 s 3896 28600 3976 29000 0 FreeSans 400 90 0 0 uio_oe[0]
port 46 nsew
flabel metal3 s 3128 28600 3208 29000 0 FreeSans 400 90 0 0 uio_oe[1]
port 47 nsew
flabel metal3 s 8504 28600 8584 29000 0 FreeSans 400 90 0 0 uio_out2
port 48 nsew
flabel metal3 s 7736 28600 7816 29000 0 FreeSans 400 90 0 0 uio_out3
port 49 nsew
flabel metal3 s 6968 28600 7048 29000 0 FreeSans 400 90 0 0 uio_out4
port 50 nsew
flabel metal3 s 6200 28600 6280 29000 0 FreeSans 400 90 0 0 uio_out5
port 51 nsew
flabel metal3 s 5432 28600 5512 29000 0 FreeSans 400 90 0 0 uio_out6
port 52 nsew
flabel metal3 s 4664 28600 4744 29000 0 FreeSans 400 90 0 0 uio_out7
port 53 nsew
flabel metal3 s 10040 28600 10120 29000 0 FreeSans 400 90 0 0 vblank
port 54 nsew
flabel metal3 s 13880 28600 13960 29000 0 FreeSans 400 90 0 0 vsync
port 55 nsew
<< properties >>
string FIXED_BBOX 0 0 32000 29000
string GDS_END 2194422
string GDS_FILE ../gds/controller.gds
string GDS_START 261558
<< end >>
