module controller (b6,
    b7,
    clk,
    ena,
    g6,
    g7,
    hblank,
    hsync,
    r6,
    r7,
    rst_n,
    uio_out2,
    uio_out3,
    uio_out4,
    uio_out5,
    uio_out6,
    uio_out7,
    vblank,
    vsync,
    VPWR,
    VGND,
    db,
    dg,
    dr,
    ui_in,
    uio_oe);
 output b6;
 output b7;
 input clk;
 input ena;
 output g6;
 output g7;
 output hblank;
 output hsync;
 output r6;
 output r7;
 input rst_n;
 output uio_out2;
 output uio_out3;
 output uio_out4;
 output uio_out5;
 output uio_out6;
 output uio_out7;
 output vblank;
 output vsync;
 inout VPWR;
 inout VGND;
 output [7:0] db;
 output [7:0] dg;
 output [7:0] dr;
 input [7:0] ui_in;
 output [1:0] uio_oe;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire \divider[0] ;
 wire \divider[1] ;
 wire gate;
 wire \h[0] ;
 wire \h[1] ;
 wire \h[2] ;
 wire \h[3] ;
 wire \h[4] ;
 wire \h[5] ;
 wire \h[6] ;
 wire \h[7] ;
 wire \h[8] ;
 wire \h[9] ;
 wire \mode[0] ;
 wire \mode[1] ;
 wire \mode[2] ;
 wire \rampc[0] ;
 wire \rampc[1] ;
 wire \rampc[2] ;
 wire \rampc[3] ;
 wire \rampc[4] ;
 wire \rampc[5] ;
 wire \rampc[6] ;
 wire \rampc[7] ;
 wire registered;
 wire \t[10] ;
 wire \t[11] ;
 wire \t[8] ;
 wire \t[9] ;
 wire net75;
 wire clknet_0_clk;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire \v[0] ;
 wire \v[1] ;
 wire \v[2] ;
 wire \v[3] ;
 wire \v[4] ;
 wire \v[5] ;
 wire \v[6] ;
 wire \v[7] ;
 wire \v[8] ;
 wire \v[9] ;
 wire \vga_sync.hsync ;
 wire \vga_sync.mode ;
 wire \vga_sync.vsync ;
 wire \voffset[0] ;
 wire \voffset[1] ;
 wire \voffset[2] ;
 wire \voffset[3] ;
 wire \voffset[4] ;
 wire \voffset[5] ;
 wire \voffset[6] ;
 wire \voffset[7] ;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;

 sg13g2_inv_2 _1056_ (.Y(_0194_),
    .A(\v[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _1057_ (.VDD(VPWR),
    .Y(_0195_),
    .A(\t[9] ),
    .VSS(VGND));
 sg13g2_inv_1 _1058_ (.VDD(VPWR),
    .Y(_0196_),
    .A(net149),
    .VSS(VGND));
 sg13g2_inv_1 _1059_ (.VDD(VPWR),
    .Y(_0197_),
    .A(net390),
    .VSS(VGND));
 sg13g2_inv_1 _1060_ (.VDD(VPWR),
    .Y(_0198_),
    .A(net5),
    .VSS(VGND));
 sg13g2_inv_1 _1061_ (.VDD(VPWR),
    .Y(_0199_),
    .A(net6),
    .VSS(VGND));
 sg13g2_inv_2 _1062_ (.Y(_0200_),
    .A(net408),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _1063_ (.Y(_0201_),
    .A(net402),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _1064_ (.Y(_0202_),
    .A(net404),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _1065_ (.VDD(VPWR),
    .Y(_0203_),
    .A(net365),
    .VSS(VGND));
 sg13g2_inv_1 _1066_ (.VDD(VPWR),
    .Y(_0204_),
    .A(net398),
    .VSS(VGND));
 sg13g2_inv_1 _1067_ (.VDD(VPWR),
    .Y(_0205_),
    .A(net396),
    .VSS(VGND));
 sg13g2_inv_1 _1068_ (.VDD(VPWR),
    .Y(_0206_),
    .A(net393),
    .VSS(VGND));
 sg13g2_inv_1 _1069_ (.VDD(VPWR),
    .Y(_0207_),
    .A(_0015_),
    .VSS(VGND));
 sg13g2_inv_2 _1070_ (.Y(_0208_),
    .A(net370),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _1071_ (.VDD(VPWR),
    .Y(_0209_),
    .A(net3),
    .VSS(VGND));
 sg13g2_inv_1 _1072_ (.VDD(VPWR),
    .Y(_0210_),
    .A(net10),
    .VSS(VGND));
 sg13g2_inv_1 _1073_ (.VDD(VPWR),
    .Y(_0211_),
    .A(net103),
    .VSS(VGND));
 sg13g2_inv_1 _1074_ (.VDD(VPWR),
    .Y(_0212_),
    .A(net84),
    .VSS(VGND));
 sg13g2_inv_1 _1075_ (.VDD(VPWR),
    .Y(_0213_),
    .A(net96),
    .VSS(VGND));
 sg13g2_inv_1 _1076_ (.VDD(VPWR),
    .Y(_0214_),
    .A(net101),
    .VSS(VGND));
 sg13g2_inv_1 _1077_ (.VDD(VPWR),
    .Y(_0215_),
    .A(_0027_),
    .VSS(VGND));
 sg13g2_inv_2 _1078_ (.Y(_0216_),
    .A(_0030_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1079_ (.B1(\h[9] ),
    .VDD(VPWR),
    .Y(_0217_),
    .VSS(VGND),
    .A1(net393),
    .A2(\h[8] ));
 sg13g2_nand3_1 _1080_ (.B(net396),
    .C(_0206_),
    .A(net398),
    .Y(_0218_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1081_ (.A(\h[4] ),
    .B(_0218_),
    .Y(_0219_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1082_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net396),
    .A2(_0207_),
    .Y(_0220_),
    .B1(net393));
 sg13g2_a21oi_1 _1083_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0201_),
    .A2(_0219_),
    .Y(_0221_),
    .B1(_0220_));
 sg13g2_nor2_1 _1084_ (.A(net409),
    .B(net407),
    .Y(_0222_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1085_ (.Y(_0223_),
    .B(\h[8] ),
    .A_N(\h[9] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _1086_ (.A(net408),
    .B(net407),
    .C(_0223_),
    .Y(_0224_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1087_ (.A(_0201_),
    .B(net404),
    .Y(_0225_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _1088_ (.B(_0224_),
    .C(_0225_),
    .A(_0219_),
    .Y(_0226_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1089_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\h[8] ),
    .A2(_0221_),
    .Y(_0227_),
    .B1(\h[9] ));
 sg13g2_a22oi_1 _1090_ (.Y(hblank),
    .B1(_0226_),
    .B2(_0227_),
    .A2(_0217_),
    .A1(_0203_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _1091_ (.VDD(VPWR),
    .Y(_0228_),
    .A(hblank),
    .VSS(VGND));
 sg13g2_and2_2 _1092_ (.A(\v[8] ),
    .B(\v[7] ),
    .X(_0229_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1093_ (.Y(_0230_),
    .A(\v[9] ),
    .B(_0229_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1094_ (.A(\v[3] ),
    .B(net378),
    .Y(_0231_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _1095_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0232_),
    .B(\v[4] ),
    .A(\v[6] ));
 sg13g2_nor2_1 _1096_ (.A(net376),
    .B(_0232_),
    .Y(_0233_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _1097_ (.A2(_0233_),
    .A1(_0231_),
    .B1(_0230_),
    .X(_0234_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1098_ (.Y(_0235_),
    .A(\v[6] ),
    .B(net377),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _1099_ (.B(net376),
    .C(_0229_),
    .A(\v[6] ),
    .Y(_0236_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _1100_ (.A(\v[9] ),
    .B(\v[4] ),
    .C(_0236_),
    .Y(_0237_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _1101_ (.VDD(VPWR),
    .Y(_0238_),
    .A(_0237_),
    .VSS(VGND));
 sg13g2_nor2_1 _1102_ (.A(\v[1] ),
    .B(net381),
    .Y(_0239_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _1103_ (.A(_0231_),
    .B(_0239_),
    .X(_0240_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _1104_ (.A(_0019_),
    .B_N(\v[6] ),
    .Y(_0241_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _1105_ (.VSS(VGND),
    .VDD(VPWR),
    .B2(_0229_),
    .C1(\v[9] ),
    .B1(_0241_),
    .A1(_0237_),
    .Y(_0242_),
    .A2(_0240_));
 sg13g2_a21oi_2 _1106_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_0242_),
    .Y(vblank),
    .A2(_0234_),
    .A1(net365));
 sg13g2_and2_1 _1107_ (.A(net2),
    .B(net1),
    .X(_0243_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1108_ (.Y(_0244_),
    .A(net2),
    .B(net1),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1109_ (.A(net92),
    .B(net413),
    .Y(_0245_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1110_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net5),
    .A2(net413),
    .Y(_0246_),
    .B1(_0245_));
 sg13g2_nand2_1 _1111_ (.Y(_0247_),
    .A(net4),
    .B(net410),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1112_ (.A(net111),
    .B(net412),
    .Y(_0248_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _1113_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_0248_),
    .Y(_0249_),
    .A2(net412),
    .A1(net4));
 sg13g2_o21ai_1 _1114_ (.B1(_0247_),
    .VDD(VPWR),
    .Y(_0250_),
    .VSS(VGND),
    .A1(net111),
    .A2(net412));
 sg13g2_nor2_1 _1115_ (.A(net109),
    .B(net413),
    .Y(_0251_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1116_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net6),
    .A2(net413),
    .Y(_0252_),
    .B1(_0251_));
 sg13g2_nor2_1 _1117_ (.A(_0250_),
    .B(_0252_),
    .Y(_0036_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _1118_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0253_),
    .B(_0252_),
    .A(_0246_));
 sg13g2_inv_1 _1119_ (.VDD(VPWR),
    .Y(_0038_),
    .A(_0253_),
    .VSS(VGND));
 sg13g2_nor2_1 _1120_ (.A(_0250_),
    .B(_0253_),
    .Y(_0082_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1121_ (.A(_0249_),
    .B(_0252_),
    .Y(_0254_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1122_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0249_),
    .A2(_0253_),
    .Y(_0000_),
    .B1(_0254_));
 sg13g2_nor2_1 _1123_ (.A(_0246_),
    .B(_0254_),
    .Y(_0001_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1124_ (.Y(vsync),
    .A(net365),
    .B(\vga_sync.vsync ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _1125_ (.A(\mode[1] ),
    .B(\mode[0] ),
    .Y(_0255_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _1126_ (.A(net367),
    .B(_0255_),
    .X(_0256_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1127_ (.Y(_0257_),
    .A(net367),
    .B(_0255_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1128_ (.Y(_0258_),
    .A(_0208_),
    .B(net361),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1129_ (.B1(net335),
    .VDD(VPWR),
    .Y(_0259_),
    .VSS(VGND),
    .A1(hblank),
    .A2(vblank));
 sg13g2_and2_2 _1130_ (.A(net1),
    .B(_0259_),
    .X(_0260_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1131_ (.B1(_0260_),
    .VDD(VPWR),
    .Y(_0261_),
    .VSS(VGND),
    .A1(net3),
    .A2(net334));
 sg13g2_nand3b_1 _1132_ (.B(\h[9] ),
    .C(net399),
    .Y(_0262_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(\h[8] ));
 sg13g2_nor2_2 _1133_ (.A(_0218_),
    .B(_0262_),
    .Y(_0263_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1134_ (.A(net3),
    .B(net359),
    .Y(_0264_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1135_ (.Y(_0265_),
    .A(\v[7] ),
    .B(\voffset[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1136_ (.Y(_0266_),
    .A(\v[6] ),
    .B(\voffset[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1137_ (.Y(_0267_),
    .A(\v[6] ),
    .B(\voffset[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _1138_ (.VDD(VPWR),
    .Y(_0268_),
    .A(_0267_),
    .VSS(VGND));
 sg13g2_nand2_1 _1139_ (.Y(_0269_),
    .A(net379),
    .B(\voffset[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1140_ (.Y(_0270_),
    .A(net381),
    .B(\voffset[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1141_ (.Y(_0271_),
    .A(net379),
    .B(\voffset[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1142_ (.B1(_0269_),
    .VDD(VPWR),
    .Y(_0272_),
    .VSS(VGND),
    .A1(_0270_),
    .A2(_0271_));
 sg13g2_and2_1 _1143_ (.A(net378),
    .B(\voffset[2] ),
    .X(_0273_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1144_ (.B(\voffset[2] ),
    .A(net378),
    .X(_0274_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1145_ (.Y(_0275_),
    .A(_0272_),
    .B(_0274_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1146_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\v[3] ),
    .A2(\voffset[3] ),
    .Y(_0276_),
    .B1(_0273_));
 sg13g2_a22oi_1 _1147_ (.Y(_0277_),
    .B1(_0275_),
    .B2(_0276_),
    .A2(_0211_),
    .A1(_0194_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _1148_ (.A(\v[4] ),
    .B(\voffset[4] ),
    .X(_0278_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _1149_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0279_),
    .B(\voffset[4] ),
    .A(\v[4] ));
 sg13g2_xnor2_1 _1150_ (.Y(_0280_),
    .A(\v[4] ),
    .B(\voffset[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1151_ (.Y(_0281_),
    .A(net377),
    .B(\voffset[5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1152_ (.Y(_0282_),
    .A(net377),
    .B(\voffset[5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1153_ (.A(_0280_),
    .B(_0282_),
    .Y(_0283_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _1154_ (.VDD(VPWR),
    .Y(_0284_),
    .A(_0283_),
    .VSS(VGND));
 sg13g2_a221oi_1 _1155_ (.VSS(VGND),
    .VDD(VPWR),
    .B2(_0276_),
    .C1(_0284_),
    .B1(_0275_),
    .A1(_0194_),
    .Y(_0285_),
    .A2(_0211_));
 sg13g2_o21ai_1 _1156_ (.B1(_0278_),
    .VDD(VPWR),
    .Y(_0286_),
    .VSS(VGND),
    .A1(net376),
    .A2(\voffset[5] ));
 sg13g2_nand2_1 _1157_ (.Y(_0287_),
    .A(_0281_),
    .B(_0286_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1158_ (.A(_0285_),
    .B(_0287_),
    .Y(_0288_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1159_ (.B1(_0268_),
    .VDD(VPWR),
    .Y(_0289_),
    .VSS(VGND),
    .A1(_0285_),
    .A2(_0287_));
 sg13g2_a21oi_2 _1160_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_0265_),
    .Y(_0290_),
    .A2(_0289_),
    .A1(_0266_));
 sg13g2_a21o_1 _1161_ (.A2(\voffset[7] ),
    .A1(\v[7] ),
    .B1(_0290_),
    .X(_0291_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1162_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net375),
    .A2(_0291_),
    .Y(_0292_),
    .B1(_0017_));
 sg13g2_and3_1 _1163_ (.X(_0293_),
    .A(net375),
    .B(_0017_),
    .C(_0291_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _1164_ (.A(net408),
    .B(_0292_),
    .C(_0293_),
    .Y(_0294_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1165_ (.B(_0291_),
    .A(net375),
    .X(_0295_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1166_ (.A(_0202_),
    .B(_0020_),
    .Y(_0296_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1167_ (.B1(_0296_),
    .VDD(VPWR),
    .Y(_0297_),
    .VSS(VGND),
    .A1(_0200_),
    .A2(_0295_));
 sg13g2_o21ai_1 _1168_ (.B1(_0201_),
    .VDD(VPWR),
    .Y(_0298_),
    .VSS(VGND),
    .A1(_0294_),
    .A2(_0297_));
 sg13g2_xor2_1 _1169_ (.B(\voffset[3] ),
    .A(\v[3] ),
    .X(_0299_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1170_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0272_),
    .A2(_0274_),
    .Y(_0300_),
    .B1(_0273_));
 sg13g2_xnor2_1 _1171_ (.Y(_0301_),
    .A(_0299_),
    .B(_0300_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1172_ (.A(_0200_),
    .B(net407),
    .Y(_0302_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1173_ (.Y(_0303_),
    .A(_0272_),
    .B(_0274_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _1174_ (.VDD(VPWR),
    .Y(_0304_),
    .A(net327),
    .VSS(VGND));
 sg13g2_nor2b_1 _1175_ (.A(net409),
    .B_N(net407),
    .Y(_0305_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1176_ (.B(_0271_),
    .A(_0270_),
    .X(_0306_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1177_ (.B(\voffset[0] ),
    .A(net380),
    .X(_0307_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1178_ (.Y(_0308_),
    .A(net380),
    .B(\voffset[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _1179_ (.A(net409),
    .B(net407),
    .X(_0309_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1180_ (.Y(_0310_),
    .A(net409),
    .B(net407),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1181_ (.S0(net408),
    .A0(net323),
    .A1(_0304_),
    .A2(net356),
    .A3(net364),
    .S1(net406),
    .X(_0311_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _1182_ (.B(net404),
    .C(_0309_),
    .A(net402),
    .Y(_0312_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _1183_ (.VDD(VPWR),
    .Y(_0313_),
    .A(_0312_),
    .VSS(VGND));
 sg13g2_nand3b_1 _1184_ (.B(net404),
    .C(net401),
    .Y(_0314_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_0311_));
 sg13g2_and3_2 _1185_ (.X(_0315_),
    .A(_0265_),
    .B(_0266_),
    .C(_0289_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _1186_ (.A(_0290_),
    .B(_0315_),
    .Y(_0316_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _1187_ (.A(_0316_),
    .B_N(_0222_),
    .Y(_0317_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1188_ (.Y(_0318_),
    .A(_0268_),
    .B(_0288_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _1189_ (.VDD(VPWR),
    .Y(_0319_),
    .A(net319),
    .VSS(VGND));
 sg13g2_a21oi_1 _1190_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0277_),
    .A2(_0279_),
    .Y(_0320_),
    .B1(_0278_));
 sg13g2_xnor2_1 _1191_ (.Y(_0321_),
    .A(_0282_),
    .B(_0320_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1192_ (.Y(_0322_),
    .A(_0277_),
    .B(_0280_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _1193_ (.Y(_0323_),
    .B1(net317),
    .B2(_0305_),
    .A2(_0319_),
    .A1(_0302_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1194_ (.B1(_0323_),
    .VDD(VPWR),
    .Y(_0324_),
    .VSS(VGND),
    .A1(_0310_),
    .A2(net321));
 sg13g2_o21ai_1 _1195_ (.B1(_0225_),
    .VDD(VPWR),
    .Y(_0325_),
    .VSS(VGND),
    .A1(_0317_),
    .A2(_0324_));
 sg13g2_nand3_1 _1196_ (.B(_0314_),
    .C(_0325_),
    .A(_0298_),
    .Y(_0326_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1197_ (.B1(net330),
    .VDD(VPWR),
    .Y(_0327_),
    .VSS(VGND),
    .A1(_0264_),
    .A2(_0326_));
 sg13g2_mux4_1 _1198_ (.S0(net368),
    .A0(_0035_),
    .A1(_0021_),
    .A2(_0020_),
    .A3(_0013_),
    .S1(net369),
    .X(_0328_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _1199_ (.A(net371),
    .B_N(net372),
    .Y(_0329_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _1200_ (.Y(_0330_),
    .A(_0208_),
    .B(net372),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _1201_ (.A(net370),
    .B(net373),
    .Y(_0331_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_2 _1202_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0332_),
    .B(net374),
    .A(net371));
 sg13g2_nor2_1 _1203_ (.A(\rampc[0] ),
    .B(_0332_),
    .Y(_0333_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _1204_ (.VSS(VGND),
    .VDD(VPWR),
    .B2(_0308_),
    .C1(_0333_),
    .B1(net363),
    .A1(net371),
    .Y(_0334_),
    .A2(_0328_));
 sg13g2_nor2b_2 _1205_ (.A(\mode[0] ),
    .B_N(\mode[1] ),
    .Y(_0335_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _1206_ (.A(net367),
    .B(_0335_),
    .X(_0336_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _1207_ (.Y(_0337_),
    .A(net367),
    .B(_0335_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1208_ (.A(\v[9] ),
    .B(net375),
    .Y(_0338_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_2 _1209_ (.A0(_0035_),
    .A1(_0328_),
    .S(_0338_),
    .X(_0339_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_2 _1210_ (.A(net353),
    .B(_0339_),
    .X(_0340_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _1211_ (.Y(_0341_),
    .A(net353),
    .B(_0339_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1212_ (.Y(_0342_),
    .A(_0334_),
    .B(_0340_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1213_ (.A(_0337_),
    .B(_0339_),
    .Y(_0343_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _1214_ (.Y(_0344_),
    .B(net353),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_0339_));
 sg13g2_o21ai_1 _1215_ (.B1(_0342_),
    .VDD(VPWR),
    .Y(_0345_),
    .VSS(VGND),
    .A1(_0334_),
    .A2(net324));
 sg13g2_inv_1 _1216_ (.VDD(VPWR),
    .Y(_0346_),
    .A(_0345_),
    .VSS(VGND));
 sg13g2_nor2b_2 _1217_ (.A(\mode[1] ),
    .B_N(\mode[0] ),
    .Y(_0347_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _1218_ (.A(_0016_),
    .B(_0347_),
    .X(_0348_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1219_ (.Y(_0349_),
    .A(_0016_),
    .B(_0347_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1220_ (.Y(_0350_),
    .A(\rampc[0] ),
    .B(_0307_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1221_ (.Y(_0351_),
    .B(net408),
    .A_N(_0350_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_2 _1222_ (.A(\mode[2] ),
    .B(_0255_),
    .X(_0352_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1223_ (.Y(_0353_),
    .A(\mode[2] ),
    .B(_0255_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1224_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0200_),
    .A2(_0350_),
    .Y(_0354_),
    .B1(net346));
 sg13g2_a221oi_1 _1225_ (.VSS(VGND),
    .VDD(VPWR),
    .B2(_0354_),
    .C1(net361),
    .B1(_0351_),
    .A1(_0334_),
    .Y(_0355_),
    .A2(net351));
 sg13g2_a21oi_1 _1226_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0346_),
    .A2(_0355_),
    .Y(_0356_),
    .B1(_0264_));
 sg13g2_o21ai_1 _1227_ (.B1(_0327_),
    .VDD(VPWR),
    .Y(_0357_),
    .VSS(VGND),
    .A1(net330),
    .A2(_0356_));
 sg13g2_a21oi_2 _1228_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_0261_),
    .Y(db[0]),
    .A2(_0357_),
    .A1(net334));
 sg13g2_o21ai_1 _1229_ (.B1(_0260_),
    .VDD(VPWR),
    .Y(_0358_),
    .VSS(VGND),
    .A1(net4),
    .A2(net334));
 sg13g2_nor2_1 _1230_ (.A(net4),
    .B(net359),
    .Y(_0359_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1231_ (.B1(net330),
    .VDD(VPWR),
    .Y(_0360_),
    .VSS(VGND),
    .A1(_0326_),
    .A2(_0359_));
 sg13g2_nand2_1 _1232_ (.Y(_0361_),
    .A(net392),
    .B(net406),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1233_ (.A(net392),
    .B(net405),
    .Y(_0362_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1234_ (.B(net406),
    .A(\rampc[1] ),
    .X(_0363_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1235_ (.Y(_0364_),
    .A(net356),
    .B(_0363_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1236_ (.Y(_0365_),
    .A(_0034_),
    .B(net364),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1237_ (.Y(_0366_),
    .A(_0364_),
    .B(_0365_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1238_ (.Y(_0367_),
    .A(_0364_),
    .B(_0365_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1239_ (.Y(_0368_),
    .A(_0351_),
    .B(_0367_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1240_ (.Y(_0369_),
    .A(net391),
    .B(net392),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1241_ (.Y(_0370_),
    .A(_0200_),
    .B(net364),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _1242_ (.A(\mode[2] ),
    .B(_0347_),
    .X(_0371_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1243_ (.Y(_0372_),
    .A(\mode[2] ),
    .B(_0347_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1244_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0369_),
    .A2(_0370_),
    .Y(_0373_),
    .B1(net341));
 sg13g2_o21ai_1 _1245_ (.B1(_0373_),
    .VDD(VPWR),
    .Y(_0374_),
    .VSS(VGND),
    .A1(_0369_),
    .A2(_0370_));
 sg13g2_nor2b_2 _1246_ (.A(net367),
    .B_N(_0335_),
    .Y(_0375_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _1247_ (.Y(_0376_),
    .B(_0335_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net367));
 sg13g2_a21o_1 _1248_ (.A2(_0375_),
    .A1(_0370_),
    .B1(net343),
    .X(_0377_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1249_ (.A(net356),
    .B(_0330_),
    .Y(_0378_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _1250_ (.A0(_0013_),
    .A1(_0023_),
    .S(net369),
    .X(_0379_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _1251_ (.A0(_0020_),
    .A1(_0021_),
    .S(net369),
    .X(_0380_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_2 _1252_ (.A0(_0380_),
    .A1(_0379_),
    .S(net368),
    .X(_0381_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _1253_ (.VSS(VGND),
    .VDD(VPWR),
    .B2(net371),
    .C1(_0378_),
    .B1(_0381_),
    .A1(_0022_),
    .Y(_0382_),
    .A2(_0331_));
 sg13g2_inv_1 _1254_ (.VDD(VPWR),
    .Y(_0383_),
    .A(_0382_),
    .VSS(VGND));
 sg13g2_a22oi_1 _1255_ (.Y(_0384_),
    .B1(_0383_),
    .B2(net325),
    .A2(_0377_),
    .A1(_0374_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1256_ (.B1(_0384_),
    .VDD(VPWR),
    .Y(_0385_),
    .VSS(VGND),
    .A1(net346),
    .A2(_0368_));
 sg13g2_nor2_2 _1257_ (.A(_0340_),
    .B(net351),
    .Y(_0386_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _1258_ (.Y(_0387_),
    .A(_0341_),
    .B(net349),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _1259_ (.VSS(VGND),
    .VDD(VPWR),
    .B2(_0382_),
    .C1(net361),
    .B1(_0387_),
    .A1(net348),
    .Y(_0388_),
    .A2(_0385_));
 sg13g2_nor2_1 _1260_ (.A(_0359_),
    .B(_0388_),
    .Y(_0389_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1261_ (.B1(_0360_),
    .VDD(VPWR),
    .Y(_0390_),
    .VSS(VGND),
    .A1(net330),
    .A2(_0389_));
 sg13g2_a21oi_2 _1262_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_0358_),
    .Y(db[1]),
    .A2(_0390_),
    .A1(net336));
 sg13g2_o21ai_1 _1263_ (.B1(_0260_),
    .VDD(VPWR),
    .Y(_0391_),
    .VSS(VGND),
    .A1(net5),
    .A2(net333));
 sg13g2_nor2_1 _1264_ (.A(net5),
    .B(net357),
    .Y(_0392_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1265_ (.B1(net329),
    .VDD(VPWR),
    .Y(_0393_),
    .VSS(VGND),
    .A1(_0326_),
    .A2(_0392_));
 sg13g2_mux4_1 _1266_ (.S0(net368),
    .A0(_0021_),
    .A1(_0023_),
    .A2(_0013_),
    .A3(_0015_),
    .S1(net369),
    .X(_0394_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _1267_ (.VDD(VPWR),
    .Y(_0395_),
    .A(_0394_),
    .VSS(VGND));
 sg13g2_nor2_1 _1268_ (.A(_0208_),
    .B(_0395_),
    .Y(_0396_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _1269_ (.VSS(VGND),
    .VDD(VPWR),
    .B2(_0024_),
    .C1(_0396_),
    .B1(_0331_),
    .A1(net327),
    .Y(_0397_),
    .A2(net363));
 sg13g2_and2_1 _1270_ (.A(net325),
    .B(_0397_),
    .X(_0398_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1271_ (.B1(_0366_),
    .VDD(VPWR),
    .Y(_0399_),
    .VSS(VGND),
    .A1(_0351_),
    .A2(_0367_));
 sg13g2_and2_1 _1272_ (.A(\rampc[2] ),
    .B(net403),
    .X(_0400_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1273_ (.B(net403),
    .A(\rampc[2] ),
    .X(_0401_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1274_ (.Y(_0402_),
    .A(_0303_),
    .B(_0401_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1275_ (.B1(_0361_),
    .VDD(VPWR),
    .Y(_0403_),
    .VSS(VGND),
    .A1(net355),
    .A2(_0362_));
 sg13g2_nor2b_1 _1276_ (.A(_0402_),
    .B_N(_0403_),
    .Y(_0404_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1277_ (.Y(_0405_),
    .A(_0402_),
    .B(_0403_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1278_ (.B(_0405_),
    .A(_0399_),
    .X(_0406_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1279_ (.Y(_0407_),
    .A(net406),
    .B(net355),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1280_ (.B1(net341),
    .VDD(VPWR),
    .Y(_0408_),
    .VSS(VGND),
    .A1(_0376_),
    .A2(_0407_));
 sg13g2_nand2_1 _1281_ (.Y(_0409_),
    .A(net392),
    .B(net408),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1282_ (.Y(_0410_),
    .A(net391),
    .B(net405),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1283_ (.Y(_0411_),
    .A(net391),
    .B(net405),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1284_ (.Y(_0412_),
    .A(_0409_),
    .B(_0411_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1285_ (.Y(_0413_),
    .A(net390),
    .B(net355),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1286_ (.Y(_0414_),
    .A(net389),
    .B(net355),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1287_ (.Y(_0415_),
    .A(net391),
    .B(net364),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1288_ (.B(_0415_),
    .A(_0414_),
    .X(_0416_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1289_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0412_),
    .A2(_0416_),
    .Y(_0417_),
    .B1(net339));
 sg13g2_o21ai_1 _1290_ (.B1(_0417_),
    .VDD(VPWR),
    .Y(_0418_),
    .VSS(VGND),
    .A1(_0412_),
    .A2(_0416_));
 sg13g2_a221oi_1 _1291_ (.VSS(VGND),
    .VDD(VPWR),
    .B2(_0418_),
    .C1(net354),
    .B1(_0408_),
    .A1(_0352_),
    .Y(_0419_),
    .A2(_0406_));
 sg13g2_o21ai_1 _1292_ (.B1(net347),
    .VDD(VPWR),
    .Y(_0420_),
    .VSS(VGND),
    .A1(_0398_),
    .A2(_0419_));
 sg13g2_o21ai_1 _1293_ (.B1(_0420_),
    .VDD(VPWR),
    .Y(_0421_),
    .VSS(VGND),
    .A1(_0386_),
    .A2(_0397_));
 sg13g2_a21oi_1 _1294_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net357),
    .A2(_0421_),
    .Y(_0422_),
    .B1(_0392_));
 sg13g2_o21ai_1 _1295_ (.B1(_0393_),
    .VDD(VPWR),
    .Y(_0423_),
    .VSS(VGND),
    .A1(net328),
    .A2(_0422_));
 sg13g2_a21oi_2 _1296_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_0391_),
    .Y(db[2]),
    .A2(_0423_),
    .A1(net332));
 sg13g2_o21ai_1 _1297_ (.B1(_0260_),
    .VDD(VPWR),
    .Y(_0424_),
    .VSS(VGND),
    .A1(net6),
    .A2(net333));
 sg13g2_nor2_1 _1298_ (.A(net6),
    .B(net357),
    .Y(_0425_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1299_ (.Y(_0426_),
    .A(_0199_),
    .B(net362),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1300_ (.B1(net329),
    .VDD(VPWR),
    .Y(_0427_),
    .VSS(VGND),
    .A1(_0326_),
    .A2(_0425_));
 sg13g2_nand2_1 _1301_ (.Y(_0428_),
    .A(net369),
    .B(_0026_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1302_ (.B1(_0428_),
    .VDD(VPWR),
    .Y(_0429_),
    .VSS(VGND),
    .A1(net369),
    .A2(_0207_));
 sg13g2_mux2_2 _1303_ (.A0(_0379_),
    .A1(_0429_),
    .S(net368),
    .X(_0430_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _1304_ (.Y(_0431_),
    .B1(_0430_),
    .B2(net370),
    .A2(_0331_),
    .A1(_0025_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1305_ (.B1(_0431_),
    .VDD(VPWR),
    .Y(_0432_),
    .VSS(VGND),
    .A1(net323),
    .A2(_0330_));
 sg13g2_a21oi_1 _1306_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0399_),
    .A2(_0405_),
    .Y(_0433_),
    .B1(_0404_));
 sg13g2_xor2_1 _1307_ (.B(net402),
    .A(net390),
    .X(_0434_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1308_ (.Y(_0435_),
    .B(_0434_),
    .A_N(net322),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1309_ (.Y(_0436_),
    .A(net322),
    .B(_0434_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _1310_ (.A2(_0401_),
    .A1(_0303_),
    .B1(_0400_),
    .X(_0437_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1311_ (.Y(_0438_),
    .A(_0436_),
    .B(_0437_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1312_ (.A(_0436_),
    .B(_0437_),
    .Y(_0439_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1313_ (.Y(_0440_),
    .A(_0436_),
    .B(_0437_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1314_ (.Y(_0441_),
    .A(_0433_),
    .B(_0440_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1315_ (.Y(_0442_),
    .A(_0202_),
    .B(net327),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1316_ (.B1(_0372_),
    .VDD(VPWR),
    .Y(_0443_),
    .VSS(VGND),
    .A1(_0376_),
    .A2(_0442_));
 sg13g2_o21ai_1 _1317_ (.B1(_0413_),
    .VDD(VPWR),
    .Y(_0444_),
    .VSS(VGND),
    .A1(_0414_),
    .A2(_0415_));
 sg13g2_xnor2_1 _1318_ (.Y(_0445_),
    .A(net387),
    .B(net327),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1319_ (.B(_0445_),
    .A(_0444_),
    .X(_0446_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1320_ (.A(_0197_),
    .B(_0202_),
    .Y(_0447_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1321_ (.B(net403),
    .A(net390),
    .X(_0448_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1322_ (.B1(_0410_),
    .VDD(VPWR),
    .Y(_0449_),
    .VSS(VGND),
    .A1(_0409_),
    .A2(_0411_));
 sg13g2_xnor2_1 _1323_ (.Y(_0450_),
    .A(_0448_),
    .B(_0449_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1324_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0446_),
    .A2(_0450_),
    .Y(_0451_),
    .B1(net339));
 sg13g2_o21ai_1 _1325_ (.B1(_0451_),
    .VDD(VPWR),
    .Y(_0452_),
    .VSS(VGND),
    .A1(_0446_),
    .A2(_0450_));
 sg13g2_a21oi_1 _1326_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0443_),
    .A2(_0452_),
    .Y(_0453_),
    .B1(net354));
 sg13g2_o21ai_1 _1327_ (.B1(_0453_),
    .VDD(VPWR),
    .Y(_0454_),
    .VSS(VGND),
    .A1(net346),
    .A2(_0441_));
 sg13g2_o21ai_1 _1328_ (.B1(_0454_),
    .VDD(VPWR),
    .Y(_0455_),
    .VSS(VGND),
    .A1(net324),
    .A2(_0432_));
 sg13g2_a22oi_1 _1329_ (.Y(_0456_),
    .B1(_0455_),
    .B2(net347),
    .A2(_0432_),
    .A1(_0387_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1330_ (.A(net361),
    .B(_0456_),
    .Y(_0457_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1331_ (.A(_0425_),
    .B(_0457_),
    .Y(_0458_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1332_ (.B1(_0427_),
    .VDD(VPWR),
    .Y(_0459_),
    .VSS(VGND),
    .A1(net329),
    .A2(_0458_));
 sg13g2_a21oi_2 _1333_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_0424_),
    .Y(db[3]),
    .A2(_0459_),
    .A1(net332));
 sg13g2_o21ai_1 _1334_ (.B1(_0260_),
    .VDD(VPWR),
    .Y(_0460_),
    .VSS(VGND),
    .A1(net7),
    .A2(net333));
 sg13g2_nor2_1 _1335_ (.A(net7),
    .B(net357),
    .Y(_0461_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1336_ (.B1(net329),
    .VDD(VPWR),
    .Y(_0462_),
    .VSS(VGND),
    .A1(_0326_),
    .A2(_0461_));
 sg13g2_mux4_1 _1337_ (.S0(\divider[1] ),
    .A0(_0023_),
    .A1(_0026_),
    .A2(_0015_),
    .A3(_0028_),
    .S1(\divider[0] ),
    .X(_0463_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _1338_ (.Y(_0464_),
    .B1(_0463_),
    .B2(net370),
    .A2(_0331_),
    .A1(_0027_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1339_ (.B1(_0464_),
    .VDD(VPWR),
    .Y(_0465_),
    .VSS(VGND),
    .A1(net321),
    .A2(_0330_));
 sg13g2_o21ai_1 _1340_ (.B1(_0438_),
    .VDD(VPWR),
    .Y(_0466_),
    .VSS(VGND),
    .A1(_0433_),
    .A2(_0439_));
 sg13g2_nand2_1 _1341_ (.Y(_0467_),
    .A(net388),
    .B(net400),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1342_ (.A(net388),
    .B(net400),
    .Y(_0468_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1343_ (.B(net400),
    .A(net388),
    .X(_0469_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1344_ (.Y(_0470_),
    .A(net320),
    .B(_0469_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1345_ (.B1(_0435_),
    .VDD(VPWR),
    .Y(_0471_),
    .VSS(VGND),
    .A1(_0197_),
    .A2(_0201_));
 sg13g2_and2_1 _1346_ (.A(_0470_),
    .B(_0471_),
    .X(_0472_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _1347_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0473_),
    .B(_0471_),
    .A(_0470_));
 sg13g2_nand2b_1 _1348_ (.Y(_0474_),
    .B(_0473_),
    .A_N(_0472_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1349_ (.Y(_0475_),
    .A(_0466_),
    .B(_0474_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1350_ (.Y(_0476_),
    .A(net401),
    .B(net323),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _1351_ (.VDD(VPWR),
    .Y(_0477_),
    .A(_0476_),
    .VSS(VGND));
 sg13g2_a21oi_1 _1352_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0375_),
    .A2(_0477_),
    .Y(_0478_),
    .B1(net343));
 sg13g2_a22oi_1 _1353_ (.Y(_0479_),
    .B1(_0444_),
    .B2(_0445_),
    .A2(_0304_),
    .A1(_0215_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1354_ (.Y(_0480_),
    .B(net323),
    .A_N(_0029_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _1355_ (.A(net322),
    .B_N(_0029_),
    .Y(_0481_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1356_ (.Y(_0482_),
    .A(_0029_),
    .B(net322),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1357_ (.Y(_0483_),
    .A(_0479_),
    .B(_0482_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1358_ (.Y(_0484_),
    .A(net388),
    .B(net401),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1359_ (.Y(_0485_),
    .A(net388),
    .B(net401),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1360_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0448_),
    .A2(_0449_),
    .Y(_0486_),
    .B1(_0447_));
 sg13g2_xnor2_1 _1361_ (.Y(_0487_),
    .A(_0485_),
    .B(_0486_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1362_ (.B1(net342),
    .VDD(VPWR),
    .Y(_0488_),
    .VSS(VGND),
    .A1(_0483_),
    .A2(_0487_));
 sg13g2_a21oi_1 _1363_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0483_),
    .A2(_0487_),
    .Y(_0489_),
    .B1(_0488_));
 sg13g2_o21ai_1 _1364_ (.B1(_0337_),
    .VDD(VPWR),
    .Y(_0490_),
    .VSS(VGND),
    .A1(_0478_),
    .A2(_0489_));
 sg13g2_a21o_1 _1365_ (.A2(_0475_),
    .A1(_0352_),
    .B1(_0490_),
    .X(_0491_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1366_ (.B1(_0491_),
    .VDD(VPWR),
    .Y(_0492_),
    .VSS(VGND),
    .A1(net324),
    .A2(_0465_));
 sg13g2_a22oi_1 _1367_ (.Y(_0493_),
    .B1(_0492_),
    .B2(net347),
    .A2(_0465_),
    .A1(_0387_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1368_ (.A(net361),
    .B(_0493_),
    .Y(_0494_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1369_ (.A(_0461_),
    .B(_0494_),
    .Y(_0495_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1370_ (.B1(_0462_),
    .VDD(VPWR),
    .Y(_0496_),
    .VSS(VGND),
    .A1(net328),
    .A2(_0495_));
 sg13g2_a21oi_2 _1371_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_0460_),
    .Y(db[4]),
    .A2(_0496_),
    .A1(net332));
 sg13g2_o21ai_1 _1372_ (.B1(_0260_),
    .VDD(VPWR),
    .Y(_0497_),
    .VSS(VGND),
    .A1(net8),
    .A2(net333));
 sg13g2_nor2_1 _1373_ (.A(net8),
    .B(net357),
    .Y(_0498_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1374_ (.B1(net328),
    .VDD(VPWR),
    .Y(_0499_),
    .VSS(VGND),
    .A1(_0326_),
    .A2(_0498_));
 sg13g2_nand2_1 _1375_ (.Y(_0500_),
    .A(net317),
    .B(_0329_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _1376_ (.A0(_0028_),
    .A1(_0014_),
    .S(net369),
    .X(_0501_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_2 _1377_ (.A0(_0429_),
    .A1(_0501_),
    .S(net368),
    .X(_0502_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _1378_ (.Y(_0503_),
    .B1(_0502_),
    .B2(net370),
    .A2(_0331_),
    .A1(_0029_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1379_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0500_),
    .A2(_0503_),
    .Y(_0504_),
    .B1(_0386_));
 sg13g2_nand3_1 _1380_ (.B(_0500_),
    .C(_0503_),
    .A(net326),
    .Y(_0505_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1381_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0466_),
    .A2(_0473_),
    .Y(_0506_),
    .B1(_0472_));
 sg13g2_and2_1 _1382_ (.A(net386),
    .B(net397),
    .X(_0507_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1383_ (.B(net397),
    .A(net386),
    .X(_0508_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1384_ (.B(_0508_),
    .A(net316),
    .X(_0509_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1385_ (.B1(_0467_),
    .VDD(VPWR),
    .Y(_0510_),
    .VSS(VGND),
    .A1(net320),
    .A2(_0468_));
 sg13g2_nand2_1 _1386_ (.Y(_0511_),
    .A(_0509_),
    .B(_0510_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1387_ (.Y(_0512_),
    .A(_0509_),
    .B(_0510_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1388_ (.Y(_0513_),
    .A(_0506_),
    .B(_0512_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1389_ (.B(net321),
    .A(net400),
    .X(_0514_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _1390_ (.A2(_0514_),
    .A1(_0375_),
    .B1(net343),
    .X(_0515_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1391_ (.B1(_0480_),
    .VDD(VPWR),
    .Y(_0516_),
    .VSS(VGND),
    .A1(_0479_),
    .A2(_0481_));
 sg13g2_xor2_1 _1392_ (.B(net320),
    .A(net384),
    .X(_0517_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1393_ (.Y(_0518_),
    .A(_0516_),
    .B(_0517_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _1394_ (.A(net386),
    .B(net400),
    .X(_0519_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1395_ (.B(net400),
    .A(net386),
    .X(_0520_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1396_ (.B1(_0484_),
    .VDD(VPWR),
    .Y(_0521_),
    .VSS(VGND),
    .A1(_0485_),
    .A2(_0486_));
 sg13g2_xor2_1 _1397_ (.B(_0521_),
    .A(_0520_),
    .X(_0522_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1398_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0518_),
    .A2(_0522_),
    .Y(_0523_),
    .B1(net340));
 sg13g2_o21ai_1 _1399_ (.B1(_0523_),
    .VDD(VPWR),
    .Y(_0524_),
    .VSS(VGND),
    .A1(_0518_),
    .A2(_0522_));
 sg13g2_a21oi_1 _1400_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0515_),
    .A2(_0524_),
    .Y(_0525_),
    .B1(net352));
 sg13g2_o21ai_1 _1401_ (.B1(_0525_),
    .VDD(VPWR),
    .Y(_0526_),
    .VSS(VGND),
    .A1(net344),
    .A2(_0513_));
 sg13g2_a21oi_1 _1402_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0505_),
    .A2(_0526_),
    .Y(_0527_),
    .B1(net350));
 sg13g2_o21ai_1 _1403_ (.B1(net360),
    .VDD(VPWR),
    .Y(_0528_),
    .VSS(VGND),
    .A1(_0504_),
    .A2(_0527_));
 sg13g2_nor2b_1 _1404_ (.A(_0498_),
    .B_N(_0528_),
    .Y(_0529_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1405_ (.B1(_0499_),
    .VDD(VPWR),
    .Y(_0530_),
    .VSS(VGND),
    .A1(net328),
    .A2(_0529_));
 sg13g2_a21oi_2 _1406_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_0497_),
    .Y(db[5]),
    .A2(_0530_),
    .A1(net332));
 sg13g2_o21ai_1 _1407_ (.B1(_0260_),
    .VDD(VPWR),
    .Y(_0531_),
    .VSS(VGND),
    .A1(net9),
    .A2(net336));
 sg13g2_nor2_1 _1408_ (.A(net9),
    .B(net360),
    .Y(_0532_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1409_ (.B1(_0263_),
    .VDD(VPWR),
    .Y(_0533_),
    .VSS(VGND),
    .A1(_0326_),
    .A2(_0532_));
 sg13g2_o21ai_1 _1410_ (.B1(_0511_),
    .VDD(VPWR),
    .Y(_0534_),
    .VSS(VGND),
    .A1(_0506_),
    .A2(_0512_));
 sg13g2_and2_1 _1411_ (.A(net384),
    .B(net395),
    .X(_0535_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1412_ (.B(net395),
    .A(\rampc[6] ),
    .X(_0536_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1413_ (.B(_0536_),
    .A(net318),
    .X(_0537_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1414_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net316),
    .A2(_0508_),
    .Y(_0538_),
    .B1(_0507_));
 sg13g2_nor2_1 _1415_ (.A(_0537_),
    .B(_0538_),
    .Y(_0539_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1416_ (.B(_0538_),
    .A(_0537_),
    .X(_0540_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1417_ (.A(_0534_),
    .B(_0540_),
    .Y(_0541_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1418_ (.Y(_0542_),
    .A(_0534_),
    .B(_0540_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1419_ (.A(net344),
    .B(_0541_),
    .Y(_0543_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1420_ (.Y(_0544_),
    .A(_0204_),
    .B(net317),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1421_ (.B1(net341),
    .VDD(VPWR),
    .Y(_0545_),
    .VSS(VGND),
    .A1(_0376_),
    .A2(_0544_));
 sg13g2_a22oi_1 _1422_ (.Y(_0546_),
    .B1(_0516_),
    .B2(_0517_),
    .A2(net320),
    .A1(_0216_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1423_ (.B(net316),
    .A(net382),
    .X(_0547_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1424_ (.Y(_0548_),
    .B(_0547_),
    .A_N(_0546_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1425_ (.B(_0547_),
    .A(_0546_),
    .X(_0549_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1426_ (.Y(_0550_),
    .A(\rampc[6] ),
    .B(net397),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _1427_ (.A2(_0521_),
    .A1(_0520_),
    .B1(_0519_),
    .X(_0551_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _1428_ (.A(_0550_),
    .B_N(_0551_),
    .Y(_0552_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1429_ (.Y(_0553_),
    .A(_0550_),
    .B(_0551_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1430_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0549_),
    .A2(_0553_),
    .Y(_0554_),
    .B1(net340));
 sg13g2_o21ai_1 _1431_ (.B1(_0554_),
    .VDD(VPWR),
    .Y(_0555_),
    .VSS(VGND),
    .A1(_0549_),
    .A2(_0553_));
 sg13g2_a221oi_1 _1432_ (.VSS(VGND),
    .VDD(VPWR),
    .B2(_0555_),
    .C1(net352),
    .B1(_0545_),
    .A1(_0542_),
    .Y(_0556_),
    .A2(_0543_));
 sg13g2_nor2_1 _1433_ (.A(net319),
    .B(_0330_),
    .Y(_0557_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _1434_ (.S0(\divider[0] ),
    .A0(_0026_),
    .A1(_0028_),
    .A2(_0014_),
    .A3(_0031_),
    .S1(net368),
    .X(_0558_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _1435_ (.VSS(VGND),
    .VDD(VPWR),
    .B2(net370),
    .C1(_0557_),
    .B1(_0558_),
    .A1(_0030_),
    .Y(_0559_),
    .A2(_0331_));
 sg13g2_nor2_1 _1436_ (.A(_0340_),
    .B(_0559_),
    .Y(_0560_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1437_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net324),
    .A2(_0559_),
    .Y(_0561_),
    .B1(_0560_));
 sg13g2_or3_1 _1438_ (.A(net351),
    .B(_0556_),
    .C(_0561_),
    .X(_0562_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1439_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net350),
    .A2(_0559_),
    .Y(_0563_),
    .B1(net362));
 sg13g2_a21oi_1 _1440_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0562_),
    .A2(_0563_),
    .Y(_0564_),
    .B1(_0532_));
 sg13g2_o21ai_1 _1441_ (.B1(_0533_),
    .VDD(VPWR),
    .Y(_0565_),
    .VSS(VGND),
    .A1(_0263_),
    .A2(_0564_));
 sg13g2_a21oi_2 _1442_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_0531_),
    .Y(b6),
    .A2(_0565_),
    .A1(net335));
 sg13g2_o21ai_1 _1443_ (.B1(_0260_),
    .VDD(VPWR),
    .Y(_0566_),
    .VSS(VGND),
    .A1(net10),
    .A2(net335));
 sg13g2_nor2_1 _1444_ (.A(net10),
    .B(net360),
    .Y(_0567_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1445_ (.B1(_0263_),
    .VDD(VPWR),
    .Y(_0568_),
    .VSS(VGND),
    .A1(_0326_),
    .A2(_0567_));
 sg13g2_xnor2_1 _1446_ (.Y(_0569_),
    .A(_0205_),
    .B(net318),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1447_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0375_),
    .A2(_0569_),
    .Y(_0570_),
    .B1(net343));
 sg13g2_o21ai_1 _1448_ (.B1(_0548_),
    .VDD(VPWR),
    .Y(_0571_),
    .VSS(VGND),
    .A1(net382),
    .A2(net316));
 sg13g2_xor2_1 _1449_ (.B(net319),
    .A(_0033_),
    .X(_0572_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1450_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\rampc[6] ),
    .A2(net397),
    .Y(_0573_),
    .B1(_0552_));
 sg13g2_xor2_1 _1451_ (.B(net395),
    .A(net383),
    .X(_0574_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1452_ (.Y(_0575_),
    .A(_0573_),
    .B(_0574_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1453_ (.Y(_0576_),
    .A(_0572_),
    .B(_0575_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1454_ (.Y(_0577_),
    .A(_0571_),
    .B(_0576_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1455_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net342),
    .A2(_0577_),
    .Y(_0578_),
    .B1(_0570_));
 sg13g2_a21oi_1 _1456_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0534_),
    .A2(_0540_),
    .Y(_0579_),
    .B1(_0539_));
 sg13g2_a21o_1 _1457_ (.A2(_0536_),
    .A1(_0319_),
    .B1(_0535_),
    .X(_0580_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1458_ (.Y(_0581_),
    .A(\rampc[7] ),
    .B(_0580_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1459_ (.Y(_0582_),
    .A(net393),
    .B(_0316_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1460_ (.Y(_0583_),
    .A(_0581_),
    .B(_0582_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1461_ (.Y(_0584_),
    .A(_0579_),
    .B(_0583_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _1462_ (.A0(_0578_),
    .A1(_0584_),
    .S(_0352_),
    .X(_0585_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1463_ (.A(_0316_),
    .B(_0330_),
    .Y(_0586_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _1464_ (.A(net369),
    .B_N(\h[9] ),
    .Y(_0587_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1465_ (.A(net368),
    .B(_0501_),
    .Y(_0588_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _1466_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_0588_),
    .Y(_0589_),
    .A2(_0587_),
    .A1(net368));
 sg13g2_a221oi_1 _1467_ (.VSS(VGND),
    .VDD(VPWR),
    .B2(net370),
    .C1(_0586_),
    .B1(_0589_),
    .A1(_0032_),
    .Y(_0590_),
    .A2(_0331_));
 sg13g2_nor2_1 _1468_ (.A(_0341_),
    .B(_0590_),
    .Y(_0591_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _1469_ (.VSS(VGND),
    .VDD(VPWR),
    .B2(net326),
    .C1(_0591_),
    .B1(_0590_),
    .A1(net367),
    .Y(_0592_),
    .A2(_0347_));
 sg13g2_o21ai_1 _1470_ (.B1(_0592_),
    .VDD(VPWR),
    .Y(_0593_),
    .VSS(VGND),
    .A1(net353),
    .A2(_0585_));
 sg13g2_a21oi_1 _1471_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net350),
    .A2(_0590_),
    .Y(_0594_),
    .B1(net362));
 sg13g2_a21oi_1 _1472_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0593_),
    .A2(_0594_),
    .Y(_0595_),
    .B1(_0567_));
 sg13g2_o21ai_1 _1473_ (.B1(_0568_),
    .VDD(VPWR),
    .Y(_0596_),
    .VSS(VGND),
    .A1(net331),
    .A2(_0595_));
 sg13g2_a21oi_2 _1474_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_0566_),
    .Y(b7),
    .A2(_0596_),
    .A1(net335));
 sg13g2_nor2_1 _1475_ (.A(_0208_),
    .B(net372),
    .Y(_0597_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _1476_ (.Y(_0598_),
    .B(net370),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net372));
 sg13g2_nor2_1 _1477_ (.A(net364),
    .B(_0332_),
    .Y(_0599_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _1478_ (.VSS(VGND),
    .VDD(VPWR),
    .B2(_0034_),
    .C1(_0599_),
    .B1(net337),
    .A1(net372),
    .Y(_0600_),
    .A2(_0328_));
 sg13g2_nand2b_1 _1479_ (.Y(_0601_),
    .B(net325),
    .A_N(_0600_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1480_ (.A(_0035_),
    .B(_0308_),
    .Y(_0602_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _1481_ (.Y(_0603_),
    .A(net345),
    .B(_0376_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1482_ (.A(_0328_),
    .B(_0603_),
    .Y(_0604_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _1483_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0605_),
    .B(_0604_),
    .A(_0377_));
 sg13g2_a22oi_1 _1484_ (.Y(_0606_),
    .B1(_0605_),
    .B2(_0374_),
    .A2(_0602_),
    .A1(_0352_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1485_ (.B1(_0601_),
    .VDD(VPWR),
    .Y(_0607_),
    .VSS(VGND),
    .A1(net354),
    .A2(_0606_));
 sg13g2_a221oi_1 _1486_ (.VSS(VGND),
    .VDD(VPWR),
    .B2(net347),
    .C1(net361),
    .B1(_0607_),
    .A1(_0387_),
    .Y(_0608_),
    .A2(_0600_));
 sg13g2_nor2_1 _1487_ (.A(_0264_),
    .B(_0608_),
    .Y(_0609_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1488_ (.B1(_0327_),
    .VDD(VPWR),
    .Y(_0610_),
    .VSS(VGND),
    .A1(net331),
    .A2(_0609_));
 sg13g2_a21oi_2 _1489_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_0261_),
    .Y(dg[0]),
    .A2(_0610_),
    .A1(net336));
 sg13g2_a22oi_1 _1490_ (.Y(_0611_),
    .B1(net337),
    .B2(_0022_),
    .A2(_0381_),
    .A1(net372),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1491_ (.B1(_0611_),
    .VDD(VPWR),
    .Y(_0612_),
    .VSS(VGND),
    .A1(net356),
    .A2(_0332_));
 sg13g2_nor2_1 _1492_ (.A(_0381_),
    .B(_0603_),
    .Y(_0613_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _1493_ (.A(net392),
    .B(net364),
    .X(_0614_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1494_ (.Y(_0615_),
    .A(_0024_),
    .B(net355),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1495_ (.Y(_0616_),
    .A(_0614_),
    .B(_0615_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1496_ (.Y(_0617_),
    .A(net391),
    .B(net408),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1497_ (.Y(_0618_),
    .A(net389),
    .B(net405),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1498_ (.A(net389),
    .B(net405),
    .Y(_0619_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1499_ (.B(net405),
    .A(net389),
    .X(_0620_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1500_ (.Y(_0621_),
    .A(_0617_),
    .B(_0620_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1501_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0616_),
    .A2(_0621_),
    .Y(_0622_),
    .B1(net339));
 sg13g2_o21ai_1 _1502_ (.B1(_0622_),
    .VDD(VPWR),
    .Y(_0623_),
    .VSS(VGND),
    .A1(_0616_),
    .A2(_0621_));
 sg13g2_o21ai_1 _1503_ (.B1(_0623_),
    .VDD(VPWR),
    .Y(_0624_),
    .VSS(VGND),
    .A1(_0408_),
    .A2(_0613_));
 sg13g2_nand3b_1 _1504_ (.B(net356),
    .C(_0352_),
    .Y(_0625_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_0020_));
 sg13g2_nand3_1 _1505_ (.B(_0624_),
    .C(_0625_),
    .A(_0337_),
    .Y(_0626_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1506_ (.B1(_0626_),
    .VDD(VPWR),
    .Y(_0627_),
    .VSS(VGND),
    .A1(net324),
    .A2(_0612_));
 sg13g2_a22oi_1 _1507_ (.Y(_0628_),
    .B1(_0627_),
    .B2(net348),
    .A2(_0612_),
    .A1(_0387_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1508_ (.A(net361),
    .B(_0628_),
    .Y(_0629_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1509_ (.A(_0359_),
    .B(_0629_),
    .Y(_0630_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1510_ (.B1(_0360_),
    .VDD(VPWR),
    .Y(_0631_),
    .VSS(VGND),
    .A1(net331),
    .A2(_0630_));
 sg13g2_a21oi_2 _1511_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_0358_),
    .Y(dg[1]),
    .A2(_0631_),
    .A1(net334));
 sg13g2_a22oi_1 _1512_ (.Y(_0632_),
    .B1(net337),
    .B2(_0024_),
    .A2(_0394_),
    .A1(net372),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1513_ (.B1(_0632_),
    .VDD(VPWR),
    .Y(_0633_),
    .VSS(VGND),
    .A1(_0304_),
    .A2(_0332_));
 sg13g2_nor2_1 _1514_ (.A(_0394_),
    .B(_0603_),
    .Y(_0634_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1515_ (.A(_0443_),
    .B(_0634_),
    .Y(_0635_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _1516_ (.Y(_0636_),
    .B1(_0614_),
    .B2(_0615_),
    .A2(net355),
    .A1(net391),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1517_ (.B(net327),
    .A(net390),
    .X(_0637_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1518_ (.Y(_0638_),
    .A(_0636_),
    .B(_0637_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _1519_ (.A(net387),
    .B(net403),
    .X(_0639_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _1520_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0640_),
    .B(net403),
    .A(net387));
 sg13g2_nand2b_1 _1521_ (.Y(_0641_),
    .B(_0640_),
    .A_N(_0639_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1522_ (.B1(_0618_),
    .VDD(VPWR),
    .Y(_0642_),
    .VSS(VGND),
    .A1(_0617_),
    .A2(_0619_));
 sg13g2_xnor2_1 _1523_ (.Y(_0643_),
    .A(_0641_),
    .B(_0642_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1524_ (.B1(net342),
    .VDD(VPWR),
    .Y(_0644_),
    .VSS(VGND),
    .A1(_0638_),
    .A2(_0643_));
 sg13g2_a21oi_1 _1525_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0638_),
    .A2(_0643_),
    .Y(_0645_),
    .B1(_0644_));
 sg13g2_nor3_1 _1526_ (.A(_0021_),
    .B(_0303_),
    .C(net345),
    .Y(_0646_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1527_ (.A(net352),
    .B(_0646_),
    .Y(_0647_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1528_ (.B1(_0647_),
    .VDD(VPWR),
    .Y(_0648_),
    .VSS(VGND),
    .A1(_0635_),
    .A2(_0645_));
 sg13g2_o21ai_1 _1529_ (.B1(_0648_),
    .VDD(VPWR),
    .Y(_0649_),
    .VSS(VGND),
    .A1(net324),
    .A2(_0633_));
 sg13g2_a22oi_1 _1530_ (.Y(_0650_),
    .B1(_0649_),
    .B2(net347),
    .A2(_0633_),
    .A1(_0387_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1531_ (.A(net361),
    .B(_0650_),
    .Y(_0651_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1532_ (.A(_0392_),
    .B(_0651_),
    .Y(_0652_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1533_ (.B1(_0393_),
    .VDD(VPWR),
    .Y(_0653_),
    .VSS(VGND),
    .A1(net328),
    .A2(_0652_));
 sg13g2_a21oi_1 _1534_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net332),
    .A2(_0653_),
    .Y(dg[2]),
    .B1(_0391_));
 sg13g2_a22oi_1 _1535_ (.Y(_0654_),
    .B1(net337),
    .B2(_0025_),
    .A2(_0430_),
    .A1(net372),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1536_ (.B1(_0654_),
    .VDD(VPWR),
    .Y(_0655_),
    .VSS(VGND),
    .A1(net323),
    .A2(_0332_));
 sg13g2_o21ai_1 _1537_ (.B1(_0478_),
    .VDD(VPWR),
    .Y(_0656_),
    .VSS(VGND),
    .A1(_0430_),
    .A2(_0603_));
 sg13g2_and2_1 _1538_ (.A(net385),
    .B(net401),
    .X(_0657_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1539_ (.B(net401),
    .A(net385),
    .X(_0658_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _1540_ (.A2(_0642_),
    .A1(_0640_),
    .B1(_0639_),
    .X(_0659_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1541_ (.B(_0659_),
    .A(_0658_),
    .X(_0660_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _1542_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0661_),
    .B(net327),
    .A(_0025_));
 sg13g2_o21ai_1 _1543_ (.B1(_0661_),
    .VDD(VPWR),
    .Y(_0662_),
    .VSS(VGND),
    .A1(_0636_),
    .A2(_0637_));
 sg13g2_and2_1 _1544_ (.A(_0215_),
    .B(net322),
    .X(_0663_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1545_ (.Y(_0664_),
    .A(_0027_),
    .B(net322),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1546_ (.Y(_0665_),
    .A(_0662_),
    .B(_0664_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1547_ (.Y(_0666_),
    .A(_0660_),
    .B(_0665_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1548_ (.B1(_0656_),
    .VDD(VPWR),
    .Y(_0667_),
    .VSS(VGND),
    .A1(_0372_),
    .A2(_0666_));
 sg13g2_nor2_1 _1549_ (.A(_0013_),
    .B(net344),
    .Y(_0668_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1550_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net323),
    .A2(_0668_),
    .Y(_0669_),
    .B1(net353));
 sg13g2_a21oi_1 _1551_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0340_),
    .A2(_0655_),
    .Y(_0670_),
    .B1(net351));
 sg13g2_o21ai_1 _1552_ (.B1(_0670_),
    .VDD(VPWR),
    .Y(_0671_),
    .VSS(VGND),
    .A1(net324),
    .A2(_0655_));
 sg13g2_a21oi_1 _1553_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0667_),
    .A2(_0669_),
    .Y(_0672_),
    .B1(_0671_));
 sg13g2_o21ai_1 _1554_ (.B1(net360),
    .VDD(VPWR),
    .Y(_0673_),
    .VSS(VGND),
    .A1(net349),
    .A2(_0655_));
 sg13g2_o21ai_1 _1555_ (.B1(_0426_),
    .VDD(VPWR),
    .Y(_0674_),
    .VSS(VGND),
    .A1(_0672_),
    .A2(_0673_));
 sg13g2_nand2b_1 _1556_ (.Y(_0675_),
    .B(_0674_),
    .A_N(net329),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1557_ (.Y(_0676_),
    .A(_0427_),
    .B(_0675_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _1558_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_0424_),
    .Y(dg[3]),
    .A2(_0676_),
    .A1(net332));
 sg13g2_nor2_1 _1559_ (.A(net321),
    .B(_0332_),
    .Y(_0677_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _1560_ (.VSS(VGND),
    .VDD(VPWR),
    .B2(_0027_),
    .C1(_0677_),
    .B1(net337),
    .A1(net373),
    .Y(_0678_),
    .A2(_0463_));
 sg13g2_or2_1 _1561_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0679_),
    .B(_0678_),
    .A(_0386_));
 sg13g2_nor2_1 _1562_ (.A(_0463_),
    .B(_0603_),
    .Y(_0680_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1563_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0662_),
    .A2(_0664_),
    .Y(_0681_),
    .B1(_0663_));
 sg13g2_xnor2_1 _1564_ (.Y(_0682_),
    .A(net386),
    .B(net320),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1565_ (.B(_0682_),
    .A(_0681_),
    .X(_0683_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1566_ (.Y(_0684_),
    .A(net384),
    .B(net400),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1567_ (.Y(_0685_),
    .A(net384),
    .B(net400),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1568_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0658_),
    .A2(_0659_),
    .Y(_0686_),
    .B1(_0657_));
 sg13g2_xnor2_1 _1569_ (.Y(_0687_),
    .A(_0685_),
    .B(_0686_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1570_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0683_),
    .A2(_0687_),
    .Y(_0688_),
    .B1(net339));
 sg13g2_o21ai_1 _1571_ (.B1(_0688_),
    .VDD(VPWR),
    .Y(_0689_),
    .VSS(VGND),
    .A1(_0683_),
    .A2(_0687_));
 sg13g2_o21ai_1 _1572_ (.B1(_0689_),
    .VDD(VPWR),
    .Y(_0690_),
    .VSS(VGND),
    .A1(_0515_),
    .A2(_0680_));
 sg13g2_nor2_1 _1573_ (.A(_0023_),
    .B(net344),
    .Y(_0691_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1574_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net321),
    .A2(_0691_),
    .Y(_0692_),
    .B1(net352));
 sg13g2_a22oi_1 _1575_ (.Y(_0693_),
    .B1(_0690_),
    .B2(_0692_),
    .A2(_0678_),
    .A1(net326),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1576_ (.B1(_0679_),
    .VDD(VPWR),
    .Y(_0694_),
    .VSS(VGND),
    .A1(net351),
    .A2(_0693_));
 sg13g2_a21oi_1 _1577_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net357),
    .A2(_0694_),
    .Y(_0695_),
    .B1(_0461_));
 sg13g2_o21ai_1 _1578_ (.B1(_0462_),
    .VDD(VPWR),
    .Y(_0696_),
    .VSS(VGND),
    .A1(net328),
    .A2(_0695_));
 sg13g2_a21oi_1 _1579_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net332),
    .A2(_0696_),
    .Y(dg[4]),
    .B1(_0460_));
 sg13g2_and2_1 _1580_ (.A(net373),
    .B(_0502_),
    .X(_0697_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _1581_ (.VSS(VGND),
    .VDD(VPWR),
    .B2(_0029_),
    .C1(_0697_),
    .B1(net338),
    .A1(net317),
    .Y(_0698_),
    .A2(_0331_));
 sg13g2_or2_1 _1582_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0699_),
    .B(_0698_),
    .A(_0386_));
 sg13g2_nor2_1 _1583_ (.A(_0502_),
    .B(_0603_),
    .Y(_0700_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1584_ (.Y(_0701_),
    .B(net320),
    .A_N(_0029_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1585_ (.B1(_0701_),
    .VDD(VPWR),
    .Y(_0702_),
    .VSS(VGND),
    .A1(_0681_),
    .A2(_0682_));
 sg13g2_nor2_1 _1586_ (.A(_0030_),
    .B(net316),
    .Y(_0703_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1587_ (.Y(_0704_),
    .A(_0216_),
    .B(net316),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1588_ (.Y(_0705_),
    .A(_0702_),
    .B(_0704_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _1589_ (.A(net383),
    .B(net397),
    .X(_0706_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1590_ (.B(net397),
    .A(net383),
    .X(_0707_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1591_ (.B1(_0684_),
    .VDD(VPWR),
    .Y(_0708_),
    .VSS(VGND),
    .A1(_0685_),
    .A2(_0686_));
 sg13g2_xor2_1 _1592_ (.B(_0708_),
    .A(_0707_),
    .X(_0709_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1593_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0705_),
    .A2(_0709_),
    .Y(_0710_),
    .B1(net340));
 sg13g2_o21ai_1 _1594_ (.B1(_0710_),
    .VDD(VPWR),
    .Y(_0711_),
    .VSS(VGND),
    .A1(_0705_),
    .A2(_0709_));
 sg13g2_o21ai_1 _1595_ (.B1(_0711_),
    .VDD(VPWR),
    .Y(_0712_),
    .VSS(VGND),
    .A1(_0545_),
    .A2(_0700_));
 sg13g2_nor3_1 _1596_ (.A(_0015_),
    .B(net317),
    .C(net344),
    .Y(_0713_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1597_ (.A(net352),
    .B(_0713_),
    .Y(_0714_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _1598_ (.Y(_0715_),
    .B1(_0712_),
    .B2(_0714_),
    .A2(_0698_),
    .A1(net326),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1599_ (.B1(_0699_),
    .VDD(VPWR),
    .Y(_0716_),
    .VSS(VGND),
    .A1(net350),
    .A2(_0715_));
 sg13g2_a21oi_1 _1600_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net357),
    .A2(_0716_),
    .Y(_0717_),
    .B1(_0498_));
 sg13g2_o21ai_1 _1601_ (.B1(_0499_),
    .VDD(VPWR),
    .Y(_0718_),
    .VSS(VGND),
    .A1(net328),
    .A2(_0717_));
 sg13g2_a21oi_1 _1602_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net332),
    .A2(_0718_),
    .Y(dg[5]),
    .B1(_0497_));
 sg13g2_o21ai_1 _1603_ (.B1(_0570_),
    .VDD(VPWR),
    .Y(_0719_),
    .VSS(VGND),
    .A1(_0558_),
    .A2(_0603_));
 sg13g2_nand2_1 _1604_ (.Y(_0720_),
    .A(\t[8] ),
    .B(net395),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1605_ (.A(\t[8] ),
    .B(net395),
    .Y(_0721_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1606_ (.Y(_0722_),
    .A(\t[8] ),
    .B(net395),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1607_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0707_),
    .A2(_0708_),
    .Y(_0723_),
    .B1(_0706_));
 sg13g2_xnor2_1 _1608_ (.Y(_0724_),
    .A(_0722_),
    .B(_0723_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _1609_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_0703_),
    .Y(_0725_),
    .A2(_0704_),
    .A1(_0702_));
 sg13g2_nand2b_1 _1610_ (.Y(_0726_),
    .B(net318),
    .A_N(net382),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _1611_ (.A(net318),
    .B_N(net382),
    .Y(_0727_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1612_ (.Y(_0728_),
    .A(net382),
    .B(net318),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1613_ (.Y(_0729_),
    .A(_0725_),
    .B(_0728_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1614_ (.Y(_0730_),
    .A(_0724_),
    .B(_0729_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1615_ (.B1(_0719_),
    .VDD(VPWR),
    .Y(_0731_),
    .VSS(VGND),
    .A1(net341),
    .A2(_0730_));
 sg13g2_nor2_1 _1616_ (.A(_0026_),
    .B(net345),
    .Y(_0732_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1617_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net318),
    .A2(_0732_),
    .Y(_0733_),
    .B1(net353));
 sg13g2_a22oi_1 _1618_ (.Y(_0734_),
    .B1(net338),
    .B2(_0030_),
    .A2(_0558_),
    .A1(net373),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1619_ (.B1(_0734_),
    .VDD(VPWR),
    .Y(_0735_),
    .VSS(VGND),
    .A1(net318),
    .A2(_0332_));
 sg13g2_o21ai_1 _1620_ (.B1(net349),
    .VDD(VPWR),
    .Y(_0736_),
    .VSS(VGND),
    .A1(_0344_),
    .A2(_0735_));
 sg13g2_a221oi_1 _1621_ (.VSS(VGND),
    .VDD(VPWR),
    .B2(_0340_),
    .C1(_0736_),
    .B1(_0735_),
    .A1(_0731_),
    .Y(_0737_),
    .A2(_0733_));
 sg13g2_o21ai_1 _1622_ (.B1(net360),
    .VDD(VPWR),
    .Y(_0738_),
    .VSS(VGND),
    .A1(net349),
    .A2(_0735_));
 sg13g2_nor2_1 _1623_ (.A(_0737_),
    .B(_0738_),
    .Y(_0739_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1624_ (.A(_0532_),
    .B(_0739_),
    .Y(_0740_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1625_ (.B1(_0533_),
    .VDD(VPWR),
    .Y(_0741_),
    .VSS(VGND),
    .A1(net331),
    .A2(_0740_));
 sg13g2_a21oi_2 _1626_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_0531_),
    .Y(g6),
    .A2(_0741_),
    .A1(net335));
 sg13g2_nor2_1 _1627_ (.A(_0316_),
    .B(_0332_),
    .Y(_0742_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _1628_ (.VSS(VGND),
    .VDD(VPWR),
    .B2(net382),
    .C1(_0742_),
    .B1(net338),
    .A1(net373),
    .Y(_0743_),
    .A2(_0589_));
 sg13g2_or2_1 _1629_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0744_),
    .B(_0743_),
    .A(_0386_));
 sg13g2_o21ai_1 _1630_ (.B1(net339),
    .VDD(VPWR),
    .Y(_0745_),
    .VSS(VGND),
    .A1(_0376_),
    .A2(_0582_));
 sg13g2_nor2_1 _1631_ (.A(_0589_),
    .B(_0603_),
    .Y(_0746_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _1632_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0747_),
    .B(_0746_),
    .A(_0745_));
 sg13g2_o21ai_1 _1633_ (.B1(_0726_),
    .VDD(VPWR),
    .Y(_0748_),
    .VSS(VGND),
    .A1(_0725_),
    .A2(_0727_));
 sg13g2_xnor2_1 _1634_ (.Y(_0749_),
    .A(_0033_),
    .B(_0316_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1635_ (.B1(_0720_),
    .VDD(VPWR),
    .Y(_0750_),
    .VSS(VGND),
    .A1(_0721_),
    .A2(_0723_));
 sg13g2_xnor2_1 _1636_ (.Y(_0751_),
    .A(\t[9] ),
    .B(net393),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1637_ (.Y(_0752_),
    .A(_0750_),
    .B(_0751_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1638_ (.Y(_0753_),
    .A(_0749_),
    .B(_0752_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _1639_ (.A(_0748_),
    .B(_0753_),
    .X(_0754_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1640_ (.B1(net342),
    .VDD(VPWR),
    .Y(_0755_),
    .VSS(VGND),
    .A1(_0748_),
    .A2(_0753_));
 sg13g2_o21ai_1 _1641_ (.B1(_0747_),
    .VDD(VPWR),
    .Y(_0756_),
    .VSS(VGND),
    .A1(_0754_),
    .A2(_0755_));
 sg13g2_nor2_1 _1642_ (.A(_0028_),
    .B(net344),
    .Y(_0757_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1643_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0316_),
    .A2(_0757_),
    .Y(_0758_),
    .B1(net352));
 sg13g2_a22oi_1 _1644_ (.Y(_0759_),
    .B1(_0756_),
    .B2(_0758_),
    .A2(_0743_),
    .A1(net326),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1645_ (.B1(_0744_),
    .VDD(VPWR),
    .Y(_0760_),
    .VSS(VGND),
    .A1(net350),
    .A2(_0759_));
 sg13g2_a21oi_1 _1646_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net360),
    .A2(_0760_),
    .Y(_0761_),
    .B1(_0567_));
 sg13g2_o21ai_1 _1647_ (.B1(_0568_),
    .VDD(VPWR),
    .Y(_0762_),
    .VSS(VGND),
    .A1(net331),
    .A2(_0761_));
 sg13g2_a21oi_2 _1648_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_0566_),
    .Y(g7),
    .A2(_0762_),
    .A1(net335));
 sg13g2_nor2_2 _1649_ (.A(net363),
    .B(net337),
    .Y(_0763_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1650_ (.A(net364),
    .B(_0598_),
    .Y(_0764_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _1651_ (.VSS(VGND),
    .VDD(VPWR),
    .B2(_0328_),
    .C1(_0764_),
    .B1(_0763_),
    .A1(_0034_),
    .Y(_0765_),
    .A2(net363));
 sg13g2_and2_1 _1652_ (.A(net325),
    .B(_0765_),
    .X(_0766_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1653_ (.Y(_0767_),
    .A(net390),
    .B(net364),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _1654_ (.VDD(VPWR),
    .Y(_0768_),
    .A(_0767_),
    .VSS(VGND));
 sg13g2_xnor2_1 _1655_ (.Y(_0769_),
    .A(_0027_),
    .B(net355),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1656_ (.Y(_0770_),
    .A(_0768_),
    .B(_0769_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1657_ (.Y(_0771_),
    .A(net389),
    .B(net408),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1658_ (.Y(_0772_),
    .A(net387),
    .B(net405),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1659_ (.Y(_0773_),
    .A(net387),
    .B(net405),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1660_ (.B(_0773_),
    .A(_0771_),
    .X(_0774_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1661_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0770_),
    .A2(_0774_),
    .Y(_0775_),
    .B1(net339));
 sg13g2_o21ai_1 _1662_ (.B1(_0775_),
    .VDD(VPWR),
    .Y(_0776_),
    .VSS(VGND),
    .A1(_0770_),
    .A2(_0774_));
 sg13g2_a221oi_1 _1663_ (.VSS(VGND),
    .VDD(VPWR),
    .B2(_0776_),
    .C1(net354),
    .B1(_0408_),
    .A1(_0352_),
    .Y(_0777_),
    .A2(_0370_));
 sg13g2_o21ai_1 _1664_ (.B1(net348),
    .VDD(VPWR),
    .Y(_0778_),
    .VSS(VGND),
    .A1(_0766_),
    .A2(_0777_));
 sg13g2_o21ai_1 _1665_ (.B1(_0778_),
    .VDD(VPWR),
    .Y(_0779_),
    .VSS(VGND),
    .A1(_0386_),
    .A2(_0765_));
 sg13g2_a21oi_1 _1666_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net359),
    .A2(_0779_),
    .Y(_0780_),
    .B1(_0264_));
 sg13g2_o21ai_1 _1667_ (.B1(_0327_),
    .VDD(VPWR),
    .Y(_0781_),
    .VSS(VGND),
    .A1(net330),
    .A2(_0780_));
 sg13g2_a21oi_1 _1668_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net334),
    .A2(_0781_),
    .Y(dr[0]),
    .B1(_0261_));
 sg13g2_a22oi_1 _1669_ (.Y(_0782_),
    .B1(_0381_),
    .B2(_0763_),
    .A2(net363),
    .A1(_0022_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1670_ (.B1(_0782_),
    .VDD(VPWR),
    .Y(_0783_),
    .VSS(VGND),
    .A1(net356),
    .A2(_0598_));
 sg13g2_a22oi_1 _1671_ (.Y(_0784_),
    .B1(_0768_),
    .B2(_0769_),
    .A2(net355),
    .A1(net387),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1672_ (.B(net327),
    .A(net385),
    .X(_0785_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1673_ (.B(_0785_),
    .A(_0784_),
    .X(_0786_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _1674_ (.A(net385),
    .B(net403),
    .X(_0787_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1675_ (.B(net403),
    .A(net385),
    .X(_0788_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1676_ (.B1(_0772_),
    .VDD(VPWR),
    .Y(_0789_),
    .VSS(VGND),
    .A1(_0771_),
    .A2(_0773_));
 sg13g2_xnor2_1 _1677_ (.Y(_0790_),
    .A(_0788_),
    .B(_0789_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1678_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0786_),
    .A2(_0790_),
    .Y(_0791_),
    .B1(net339));
 sg13g2_o21ai_1 _1679_ (.B1(_0791_),
    .VDD(VPWR),
    .Y(_0792_),
    .VSS(VGND),
    .A1(_0786_),
    .A2(_0790_));
 sg13g2_a21oi_1 _1680_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0443_),
    .A2(_0792_),
    .Y(_0793_),
    .B1(net354));
 sg13g2_o21ai_1 _1681_ (.B1(_0793_),
    .VDD(VPWR),
    .Y(_0794_),
    .VSS(VGND),
    .A1(net346),
    .A2(_0407_));
 sg13g2_o21ai_1 _1682_ (.B1(_0794_),
    .VDD(VPWR),
    .Y(_0795_),
    .VSS(VGND),
    .A1(net324),
    .A2(_0783_));
 sg13g2_a22oi_1 _1683_ (.Y(_0796_),
    .B1(_0795_),
    .B2(net348),
    .A2(_0783_),
    .A1(_0387_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _1684_ (.VDD(VPWR),
    .Y(_0797_),
    .A(_0796_),
    .VSS(VGND));
 sg13g2_a21oi_1 _1685_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net359),
    .A2(_0797_),
    .Y(_0798_),
    .B1(_0359_));
 sg13g2_o21ai_1 _1686_ (.B1(_0360_),
    .VDD(VPWR),
    .Y(_0799_),
    .VSS(VGND),
    .A1(net330),
    .A2(_0798_));
 sg13g2_a21oi_1 _1687_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net334),
    .A2(_0799_),
    .Y(dr[1]),
    .B1(_0358_));
 sg13g2_a22oi_1 _1688_ (.Y(_0800_),
    .B1(_0763_),
    .B2(_0395_),
    .A2(net337),
    .A1(_0304_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1689_ (.B1(_0800_),
    .VDD(VPWR),
    .Y(_0801_),
    .VSS(VGND),
    .A1(_0024_),
    .A2(_0330_));
 sg13g2_nand2_1 _1690_ (.Y(_0802_),
    .A(net325),
    .B(_0801_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1691_ (.Y(_0803_),
    .A(net384),
    .B(net401),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1692_ (.Y(_0804_),
    .A(net384),
    .B(net401),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1693_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0788_),
    .A2(_0789_),
    .Y(_0805_),
    .B1(_0787_));
 sg13g2_xnor2_1 _1694_ (.Y(_0806_),
    .A(_0804_),
    .B(_0805_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _1695_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0807_),
    .B(net327),
    .A(_0029_));
 sg13g2_o21ai_1 _1696_ (.B1(_0807_),
    .VDD(VPWR),
    .Y(_0808_),
    .VSS(VGND),
    .A1(_0784_),
    .A2(_0785_));
 sg13g2_and2_1 _1697_ (.A(_0216_),
    .B(net322),
    .X(_0809_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1698_ (.Y(_0810_),
    .A(_0030_),
    .B(net322),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1699_ (.B(_0810_),
    .A(_0808_),
    .X(_0811_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1700_ (.B1(net342),
    .VDD(VPWR),
    .Y(_0812_),
    .VSS(VGND),
    .A1(_0806_),
    .A2(_0811_));
 sg13g2_a21oi_1 _1701_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0806_),
    .A2(_0811_),
    .Y(_0813_),
    .B1(_0812_));
 sg13g2_nor2_1 _1702_ (.A(net346),
    .B(_0442_),
    .Y(_0814_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1703_ (.B1(_0337_),
    .VDD(VPWR),
    .Y(_0815_),
    .VSS(VGND),
    .A1(_0478_),
    .A2(_0813_));
 sg13g2_o21ai_1 _1704_ (.B1(_0802_),
    .VDD(VPWR),
    .Y(_0816_),
    .VSS(VGND),
    .A1(_0814_),
    .A2(_0815_));
 sg13g2_nand2_1 _1705_ (.Y(_0817_),
    .A(net347),
    .B(_0816_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1706_ (.B1(_0817_),
    .VDD(VPWR),
    .Y(_0818_),
    .VSS(VGND),
    .A1(_0386_),
    .A2(_0801_));
 sg13g2_a21oi_1 _1707_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net357),
    .A2(_0818_),
    .Y(_0819_),
    .B1(_0392_));
 sg13g2_o21ai_1 _1708_ (.B1(_0393_),
    .VDD(VPWR),
    .Y(_0820_),
    .VSS(VGND),
    .A1(net330),
    .A2(_0819_));
 sg13g2_a21oi_1 _1709_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net333),
    .A2(_0820_),
    .Y(dr[2]),
    .B1(_0391_));
 sg13g2_a21oi_2 _1710_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_0809_),
    .Y(_0821_),
    .A2(_0810_),
    .A1(_0808_));
 sg13g2_xnor2_1 _1711_ (.Y(_0822_),
    .A(\rampc[7] ),
    .B(net320),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1712_ (.Y(_0823_),
    .A(_0821_),
    .B(_0822_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _1713_ (.A(net383),
    .B(net399),
    .X(_0824_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1714_ (.B(net399),
    .A(net383),
    .X(_0825_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1715_ (.B1(_0803_),
    .VDD(VPWR),
    .Y(_0826_),
    .VSS(VGND),
    .A1(_0804_),
    .A2(_0805_));
 sg13g2_xor2_1 _1716_ (.B(_0826_),
    .A(_0825_),
    .X(_0827_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1717_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0823_),
    .A2(_0827_),
    .Y(_0828_),
    .B1(net340));
 sg13g2_o21ai_1 _1718_ (.B1(_0828_),
    .VDD(VPWR),
    .Y(_0829_),
    .VSS(VGND),
    .A1(_0823_),
    .A2(_0827_));
 sg13g2_nand2b_1 _1719_ (.Y(_0830_),
    .B(_0763_),
    .A_N(_0430_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1720_ (.B1(_0830_),
    .VDD(VPWR),
    .Y(_0831_),
    .VSS(VGND),
    .A1(_0025_),
    .A2(_0330_));
 sg13g2_a21oi_2 _1721_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_0831_),
    .Y(_0832_),
    .A2(net337),
    .A1(net323));
 sg13g2_a22oi_1 _1722_ (.Y(_0833_),
    .B1(_0832_),
    .B2(net325),
    .A2(_0829_),
    .A1(_0515_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1723_ (.B1(_0833_),
    .VDD(VPWR),
    .Y(_0834_),
    .VSS(VGND),
    .A1(net346),
    .A2(_0476_));
 sg13g2_o21ai_1 _1724_ (.B1(net358),
    .VDD(VPWR),
    .Y(_0835_),
    .VSS(VGND),
    .A1(_0386_),
    .A2(_0832_));
 sg13g2_a21oi_1 _1725_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net347),
    .A2(_0834_),
    .Y(_0836_),
    .B1(_0835_));
 sg13g2_nor2_1 _1726_ (.A(_0425_),
    .B(_0836_),
    .Y(_0837_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1727_ (.B1(_0427_),
    .VDD(VPWR),
    .Y(_0838_),
    .VSS(VGND),
    .A1(net329),
    .A2(_0837_));
 sg13g2_a21oi_1 _1728_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net333),
    .A2(_0838_),
    .Y(dr[3]),
    .B1(_0424_));
 sg13g2_nand2b_1 _1729_ (.Y(_0839_),
    .B(net320),
    .A_N(net382),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1730_ (.B1(_0839_),
    .VDD(VPWR),
    .Y(_0840_),
    .VSS(VGND),
    .A1(_0821_),
    .A2(_0822_));
 sg13g2_nor2_1 _1731_ (.A(_0033_),
    .B(net316),
    .Y(_0841_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1732_ (.B(net316),
    .A(_0033_),
    .X(_0842_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1733_ (.Y(_0843_),
    .A(_0840_),
    .B(_0842_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1734_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0825_),
    .A2(_0826_),
    .Y(_0844_),
    .B1(_0824_));
 sg13g2_nor2_1 _1735_ (.A(\t[8] ),
    .B(net398),
    .Y(_0845_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1736_ (.B(net397),
    .A(\t[8] ),
    .X(_0846_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1737_ (.Y(_0847_),
    .A(_0844_),
    .B(_0846_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1738_ (.Y(_0848_),
    .A(_0843_),
    .B(_0847_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1739_ (.B1(_0545_),
    .VDD(VPWR),
    .Y(_0849_),
    .VSS(VGND),
    .A1(net341),
    .A2(_0848_));
 sg13g2_a21oi_1 _1740_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0352_),
    .A2(_0514_),
    .Y(_0850_),
    .B1(net352));
 sg13g2_a22oi_1 _1741_ (.Y(_0851_),
    .B1(_0463_),
    .B2(_0763_),
    .A2(net363),
    .A1(_0027_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1742_ (.B1(_0851_),
    .VDD(VPWR),
    .Y(_0852_),
    .VSS(VGND),
    .A1(net321),
    .A2(_0598_));
 sg13g2_inv_1 _1743_ (.VDD(VPWR),
    .Y(_0853_),
    .A(_0852_),
    .VSS(VGND));
 sg13g2_o21ai_1 _1744_ (.B1(net349),
    .VDD(VPWR),
    .Y(_0854_),
    .VSS(VGND),
    .A1(_0344_),
    .A2(_0852_));
 sg13g2_a221oi_1 _1745_ (.VSS(VGND),
    .VDD(VPWR),
    .B2(_0340_),
    .C1(_0854_),
    .B1(_0852_),
    .A1(_0849_),
    .Y(_0855_),
    .A2(_0850_));
 sg13g2_a21oi_1 _1746_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net351),
    .A2(_0853_),
    .Y(_0856_),
    .B1(_0855_));
 sg13g2_a21oi_1 _1747_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net358),
    .A2(_0856_),
    .Y(_0857_),
    .B1(_0461_));
 sg13g2_o21ai_1 _1748_ (.B1(_0462_),
    .VDD(VPWR),
    .Y(_0858_),
    .VSS(VGND),
    .A1(net329),
    .A2(_0857_));
 sg13g2_a21oi_1 _1749_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net333),
    .A2(_0858_),
    .Y(dr[4]),
    .B1(_0460_));
 sg13g2_a21oi_2 _1750_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_0841_),
    .Y(_0859_),
    .A2(_0842_),
    .A1(_0840_));
 sg13g2_nor2b_1 _1751_ (.A(_0009_),
    .B_N(net319),
    .Y(_0860_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1752_ (.Y(_0861_),
    .A(_0009_),
    .B(net319),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1753_ (.Y(_0862_),
    .B(_0861_),
    .A_N(_0859_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1754_ (.B(_0861_),
    .A(_0859_),
    .X(_0863_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1755_ (.Y(_0864_),
    .A(\t[9] ),
    .B(net395),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _1756_ (.VSS(VGND),
    .VDD(VPWR),
    .B2(_0826_),
    .C1(_0824_),
    .B1(_0825_),
    .A1(\t[8] ),
    .Y(_0865_),
    .A2(net397));
 sg13g2_nor3_1 _1757_ (.A(_0845_),
    .B(_0864_),
    .C(_0865_),
    .Y(_0866_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1758_ (.B1(_0864_),
    .VDD(VPWR),
    .Y(_0867_),
    .VSS(VGND),
    .A1(_0845_),
    .A2(_0865_));
 sg13g2_nand2b_1 _1759_ (.Y(_0868_),
    .B(_0867_),
    .A_N(_0866_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1760_ (.Y(_0869_),
    .A(_0863_),
    .B(_0868_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1761_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net342),
    .A2(_0869_),
    .Y(_0870_),
    .B1(_0570_));
 sg13g2_o21ai_1 _1762_ (.B1(_0337_),
    .VDD(VPWR),
    .Y(_0871_),
    .VSS(VGND),
    .A1(net344),
    .A2(_0544_));
 sg13g2_nand2_1 _1763_ (.Y(_0872_),
    .A(net317),
    .B(net338),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _1764_ (.Y(_0873_),
    .B1(_0502_),
    .B2(_0763_),
    .A2(_0329_),
    .A1(_0029_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _1765_ (.Y(_0874_),
    .A(_0872_),
    .B(_0873_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1766_ (.B1(net349),
    .VDD(VPWR),
    .Y(_0875_),
    .VSS(VGND),
    .A1(_0344_),
    .A2(_0874_));
 sg13g2_a21oi_1 _1767_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0340_),
    .A2(_0874_),
    .Y(_0876_),
    .B1(_0875_));
 sg13g2_o21ai_1 _1768_ (.B1(_0876_),
    .VDD(VPWR),
    .Y(_0877_),
    .VSS(VGND),
    .A1(_0870_),
    .A2(_0871_));
 sg13g2_o21ai_1 _1769_ (.B1(net358),
    .VDD(VPWR),
    .Y(_0878_),
    .VSS(VGND),
    .A1(net347),
    .A2(_0874_));
 sg13g2_inv_1 _1770_ (.VDD(VPWR),
    .Y(_0879_),
    .A(_0878_),
    .VSS(VGND));
 sg13g2_a21oi_1 _1771_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0877_),
    .A2(_0879_),
    .Y(_0880_),
    .B1(_0498_));
 sg13g2_o21ai_1 _1772_ (.B1(_0499_),
    .VDD(VPWR),
    .Y(_0881_),
    .VSS(VGND),
    .A1(net328),
    .A2(_0880_));
 sg13g2_a21oi_1 _1773_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net333),
    .A2(_0881_),
    .Y(dr[5]),
    .B1(_0497_));
 sg13g2_nor3_1 _1774_ (.A(_0010_),
    .B(_0290_),
    .C(_0315_),
    .Y(_0882_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _1775_ (.A(_0010_),
    .B(_0290_),
    .C(_0315_),
    .X(_0883_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1776_ (.B1(_0010_),
    .VDD(VPWR),
    .Y(_0884_),
    .VSS(VGND),
    .A1(_0290_),
    .A2(_0315_));
 sg13g2_a21oi_1 _1777_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0883_),
    .A2(_0884_),
    .Y(_0885_),
    .B1(_0860_));
 sg13g2_nand3_1 _1778_ (.B(_0883_),
    .C(_0884_),
    .A(_0861_),
    .Y(_0886_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _1779_ (.B(_0883_),
    .C(_0884_),
    .A(_0860_),
    .Y(_0887_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1780_ (.B1(_0887_),
    .VDD(VPWR),
    .Y(_0888_),
    .VSS(VGND),
    .A1(_0859_),
    .A2(_0886_));
 sg13g2_a21oi_1 _1781_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0862_),
    .A2(_0885_),
    .Y(_0889_),
    .B1(_0888_));
 sg13g2_nand2_1 _1782_ (.Y(_0890_),
    .A(\t[10] ),
    .B(net394),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1783_ (.A(\t[10] ),
    .B(net394),
    .Y(_0891_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1784_ (.Y(_0892_),
    .A(\t[10] ),
    .B(net394),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1785_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\t[9] ),
    .A2(net395),
    .Y(_0893_),
    .B1(_0866_));
 sg13g2_xnor2_1 _1786_ (.Y(_0894_),
    .A(_0892_),
    .B(_0893_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1787_ (.Y(_0895_),
    .A(_0889_),
    .B(_0894_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1788_ (.B1(_0745_),
    .VDD(VPWR),
    .Y(_0896_),
    .VSS(VGND),
    .A1(net339),
    .A2(_0895_));
 sg13g2_a21oi_1 _1789_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0352_),
    .A2(_0569_),
    .Y(_0897_),
    .B1(net352));
 sg13g2_nor2_1 _1790_ (.A(net318),
    .B(_0598_),
    .Y(_0898_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _1791_ (.VSS(VGND),
    .VDD(VPWR),
    .B2(_0763_),
    .C1(_0898_),
    .B1(_0558_),
    .A1(_0030_),
    .Y(_0899_),
    .A2(net363));
 sg13g2_a21oi_1 _1792_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net325),
    .A2(_0899_),
    .Y(_0900_),
    .B1(net350));
 sg13g2_o21ai_1 _1793_ (.B1(_0900_),
    .VDD(VPWR),
    .Y(_0901_),
    .VSS(VGND),
    .A1(_0341_),
    .A2(_0899_));
 sg13g2_a21o_1 _1794_ (.A2(_0897_),
    .A1(_0896_),
    .B1(_0901_),
    .X(_0902_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1795_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net350),
    .A2(_0899_),
    .Y(_0903_),
    .B1(net362));
 sg13g2_a21oi_1 _1796_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0902_),
    .A2(_0903_),
    .Y(_0904_),
    .B1(_0532_));
 sg13g2_o21ai_1 _1797_ (.B1(_0533_),
    .VDD(VPWR),
    .Y(_0905_),
    .VSS(VGND),
    .A1(net331),
    .A2(_0904_));
 sg13g2_a21oi_2 _1798_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_0531_),
    .Y(r6),
    .A2(_0905_),
    .A1(net335));
 sg13g2_xor2_1 _1799_ (.B(_0295_),
    .A(\h[8] ),
    .X(_0906_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1800_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0375_),
    .A2(_0906_),
    .Y(_0907_),
    .B1(net342));
 sg13g2_o21ai_1 _1801_ (.B1(_0890_),
    .VDD(VPWR),
    .Y(_0908_),
    .VSS(VGND),
    .A1(_0891_),
    .A2(_0893_));
 sg13g2_xnor2_1 _1802_ (.Y(_0909_),
    .A(\t[11] ),
    .B(\h[8] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1803_ (.Y(_0910_),
    .A(_0908_),
    .B(_0909_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1804_ (.Y(_0911_),
    .A(\t[11] ),
    .B(_0295_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1805_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0860_),
    .A2(_0884_),
    .Y(_0912_),
    .B1(_0882_));
 sg13g2_o21ai_1 _1806_ (.B1(_0912_),
    .VDD(VPWR),
    .Y(_0913_),
    .VSS(VGND),
    .A1(_0859_),
    .A2(_0886_));
 sg13g2_xnor2_1 _1807_ (.Y(_0914_),
    .A(_0910_),
    .B(_0913_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1808_ (.Y(_0915_),
    .A(_0911_),
    .B(_0914_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1809_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net342),
    .A2(_0915_),
    .Y(_0916_),
    .B1(_0907_));
 sg13g2_o21ai_1 _1810_ (.B1(_0337_),
    .VDD(VPWR),
    .Y(_0917_),
    .VSS(VGND),
    .A1(net344),
    .A2(_0582_));
 sg13g2_nor2_1 _1811_ (.A(_0316_),
    .B(_0598_),
    .Y(_0918_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _1812_ (.VSS(VGND),
    .VDD(VPWR),
    .B2(_0763_),
    .C1(_0918_),
    .B1(_0589_),
    .A1(net382),
    .Y(_0919_),
    .A2(net363));
 sg13g2_nor2_1 _1813_ (.A(_0341_),
    .B(_0919_),
    .Y(_0920_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _1814_ (.VSS(VGND),
    .VDD(VPWR),
    .B2(net325),
    .C1(_0920_),
    .B1(_0919_),
    .A1(net367),
    .Y(_0921_),
    .A2(_0347_));
 sg13g2_o21ai_1 _1815_ (.B1(_0921_),
    .VDD(VPWR),
    .Y(_0922_),
    .VSS(VGND),
    .A1(_0916_),
    .A2(_0917_));
 sg13g2_a21oi_1 _1816_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net350),
    .A2(_0919_),
    .Y(_0923_),
    .B1(net362));
 sg13g2_a21oi_1 _1817_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0922_),
    .A2(_0923_),
    .Y(_0924_),
    .B1(_0567_));
 sg13g2_o21ai_1 _1818_ (.B1(_0568_),
    .VDD(VPWR),
    .Y(_0925_),
    .VSS(VGND),
    .A1(net331),
    .A2(_0924_));
 sg13g2_a21oi_2 _1819_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_0566_),
    .Y(r7),
    .A2(_0925_),
    .A1(net335));
 sg13g2_a21o_1 _1820_ (.A2(_0254_),
    .A1(_0246_),
    .B1(_0082_),
    .X(_0037_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _1821_ (.B(_0206_),
    .C(\h[9] ),
    .A(_0205_),
    .Y(_0926_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1822_ (.B1(net404),
    .VDD(VPWR),
    .Y(_0927_),
    .VSS(VGND),
    .A1(net365),
    .A2(_0926_));
 sg13g2_nand2_1 _1823_ (.Y(_0928_),
    .A(_0204_),
    .B(net399),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _1824_ (.A(_0013_),
    .B(_0014_),
    .C(_0310_),
    .D(_0928_),
    .Y(_0929_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _1825_ (.B(net396),
    .C(net393),
    .A(net365),
    .Y(_0930_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1826_ (.B1(_0202_),
    .VDD(VPWR),
    .Y(_0931_),
    .VSS(VGND),
    .A1(\h[9] ),
    .A2(_0930_));
 sg13g2_and3_2 _1827_ (.X(_0932_),
    .A(_0927_),
    .B(_0929_),
    .C(_0931_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _1828_ (.B(_0929_),
    .C(_0931_),
    .A(_0927_),
    .Y(_0933_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _1829_ (.A(net414),
    .B(_0932_),
    .Y(_0934_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _1830_ (.Y(_0935_),
    .A(net417),
    .B(_0933_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _1831_ (.A(net77),
    .B(_0934_),
    .X(_0039_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _1832_ (.A(_0222_),
    .B(net415),
    .C(_0309_),
    .Y(_0040_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1833_ (.Y(_0936_),
    .A(net403),
    .B(_0309_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1834_ (.A(_0935_),
    .B(_0936_),
    .Y(_0041_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1835_ (.A(net131),
    .B(_0310_),
    .Y(_0937_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1836_ (.Y(_0938_),
    .A(net402),
    .B(_0937_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1837_ (.A(_0935_),
    .B(net132),
    .Y(_0042_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1838_ (.Y(_0939_),
    .A(net117),
    .B(_0312_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1839_ (.A(_0935_),
    .B(_0939_),
    .Y(_0043_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1840_ (.Y(_0940_),
    .A(net398),
    .B(net399),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _1841_ (.A(_0312_),
    .B(_0940_),
    .Y(_0941_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1842_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net399),
    .A2(_0313_),
    .Y(_0942_),
    .B1(net398));
 sg13g2_nor3_1 _1843_ (.A(_0935_),
    .B(_0941_),
    .C(net129),
    .Y(_0044_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1844_ (.B1(_0934_),
    .VDD(VPWR),
    .Y(_0943_),
    .VSS(VGND),
    .A1(net396),
    .A2(_0941_));
 sg13g2_a21oi_1 _1845_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net396),
    .A2(_0941_),
    .Y(_0045_),
    .B1(_0943_));
 sg13g2_nor3_1 _1846_ (.A(_0026_),
    .B(_0312_),
    .C(_0940_),
    .Y(_0944_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1847_ (.Y(_0945_),
    .A(net394),
    .B(_0944_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1848_ (.A(_0935_),
    .B(net139),
    .Y(_0046_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _1849_ (.B(net393),
    .C(_0941_),
    .A(net396),
    .Y(_0946_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1850_ (.B(_0946_),
    .A(net137),
    .X(_0947_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1851_ (.A(_0935_),
    .B(_0947_),
    .Y(_0047_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1852_ (.A(net107),
    .B(_0946_),
    .Y(_0948_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1853_ (.Y(_0949_),
    .A(\h[9] ),
    .B(_0948_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1854_ (.A(_0935_),
    .B(net108),
    .Y(_0048_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _1855_ (.B(net378),
    .C(_0239_),
    .A(\v[3] ),
    .Y(_0950_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _1856_ (.A(net375),
    .B(\v[7] ),
    .C(net366),
    .D(_0950_),
    .Y(_0951_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1857_ (.A(net376),
    .B(_0951_),
    .Y(_0952_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _1858_ (.X(_0953_),
    .A(net379),
    .B(net381),
    .C(_0231_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _1859_ (.B(_0229_),
    .C(_0953_),
    .A(net366),
    .Y(_0954_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _1860_ (.A(net376),
    .B(_0954_),
    .X(_0955_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_2 _1861_ (.A(_0017_),
    .B(_0232_),
    .C(_0952_),
    .Y(_0956_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0955_));
 sg13g2_or4_1 _1862_ (.A(net375),
    .B(\v[7] ),
    .C(net376),
    .D(net366),
    .X(_0957_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _1863_ (.B(net366),
    .C(_0229_),
    .A(net376),
    .Y(_0958_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0953_));
 sg13g2_o21ai_1 _1864_ (.B1(_0958_),
    .VDD(VPWR),
    .Y(_0959_),
    .VSS(VGND),
    .A1(_0950_),
    .A2(_0957_));
 sg13g2_inv_1 _1865_ (.VDD(VPWR),
    .Y(_0960_),
    .A(_0959_),
    .VSS(VGND));
 sg13g2_nor3_1 _1866_ (.A(_0017_),
    .B(_0232_),
    .C(_0960_),
    .Y(_0961_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _1867_ (.A(_0933_),
    .B_N(_0961_),
    .Y(_0962_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1868_ (.A(\rampc[0] ),
    .B(_0962_),
    .Y(_0963_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _1869_ (.A(net87),
    .B_N(_0962_),
    .Y(_0964_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _1870_ (.A(net410),
    .B(_0963_),
    .C(_0964_),
    .Y(_0049_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1871_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net118),
    .A2(_0962_),
    .Y(_0965_),
    .B1(net392));
 sg13g2_and4_1 _1872_ (.A(net392),
    .B(\rampc[0] ),
    .C(_0932_),
    .D(_0956_),
    .X(_0966_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _1873_ (.X(_0967_),
    .A(net392),
    .B(\rampc[0] ),
    .C(_0962_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _1874_ (.A(net410),
    .B(net119),
    .C(_0966_),
    .Y(_0050_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1875_ (.A(net391),
    .B(_0966_),
    .Y(_0968_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _1876_ (.A(net391),
    .B(_0967_),
    .X(_0969_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _1877_ (.A(net411),
    .B(_0968_),
    .C(_0969_),
    .Y(_0051_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _1878_ (.A(net141),
    .B_N(_0967_),
    .Y(_0091_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1879_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net389),
    .A2(_0091_),
    .Y(_0092_),
    .B1(net411));
 sg13g2_o21ai_1 _1880_ (.B1(_0092_),
    .VDD(VPWR),
    .Y(_0093_),
    .VSS(VGND),
    .A1(net389),
    .A2(_0091_));
 sg13g2_inv_1 _1881_ (.VDD(VPWR),
    .Y(_0052_),
    .A(net142),
    .VSS(VGND));
 sg13g2_nand2_1 _1882_ (.Y(_0094_),
    .A(net389),
    .B(_0969_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1883_ (.B(_0094_),
    .A(net387),
    .X(_0095_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1884_ (.A(net411),
    .B(_0095_),
    .Y(_0053_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1885_ (.A(_0027_),
    .B(_0094_),
    .Y(_0096_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1886_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net385),
    .A2(_0096_),
    .Y(_0097_),
    .B1(net411));
 sg13g2_o21ai_1 _1887_ (.B1(_0097_),
    .VDD(VPWR),
    .Y(_0098_),
    .VSS(VGND),
    .A1(net385),
    .A2(_0096_));
 sg13g2_inv_1 _1888_ (.VDD(VPWR),
    .Y(_0054_),
    .A(_0098_),
    .VSS(VGND));
 sg13g2_and4_2 _1889_ (.A(net385),
    .B(net387),
    .C(net390),
    .D(_0969_),
    .X(_0099_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1890_ (.Y(_0100_),
    .A(net384),
    .B(_0099_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1891_ (.A(net411),
    .B(_0100_),
    .Y(_0055_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1892_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0216_),
    .A2(_0099_),
    .Y(_0101_),
    .B1(net383));
 sg13g2_and3_1 _1893_ (.X(_0102_),
    .A(net383),
    .B(_0216_),
    .C(_0099_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _1894_ (.A(net411),
    .B(_0101_),
    .C(_0102_),
    .Y(_0056_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _1895_ (.B(net384),
    .C(_0099_),
    .A(net383),
    .Y(_0103_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1896_ (.Y(_0104_),
    .A(_0196_),
    .B(_0103_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1897_ (.A(net415),
    .B(_0104_),
    .Y(_0057_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1898_ (.A(_0033_),
    .B(_0103_),
    .Y(_0105_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1899_ (.A(net113),
    .B(_0105_),
    .Y(_0106_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1900_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net113),
    .A2(_0105_),
    .Y(_0107_),
    .B1(net415));
 sg13g2_nor2b_1 _1901_ (.A(net114),
    .B_N(_0107_),
    .Y(_0058_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _1902_ (.A(_0195_),
    .B(_0196_),
    .C(_0103_),
    .X(_0108_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1903_ (.B(_0108_),
    .A(net115),
    .X(_0109_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1904_ (.A(net415),
    .B(_0109_),
    .Y(_0059_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1905_ (.A(_0010_),
    .B(_0108_),
    .Y(_0110_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1906_ (.A(net98),
    .B(_0110_),
    .Y(_0111_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1907_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net98),
    .A2(_0110_),
    .Y(_0112_),
    .B1(net415));
 sg13g2_nor2b_1 _1908_ (.A(net99),
    .B_N(_0112_),
    .Y(_0060_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1909_ (.B(net9),
    .A(\mode[2] ),
    .X(_0113_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1910_ (.B(net8),
    .A(\mode[1] ),
    .X(_0114_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1911_ (.B(net7),
    .A(\mode[0] ),
    .X(_0115_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _1912_ (.A(_0113_),
    .B(_0114_),
    .C(_0115_),
    .Y(_0116_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _1913_ (.A(_0228_),
    .B(net362),
    .C(_0116_),
    .Y(_0117_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1914_ (.A(net416),
    .B(_0117_),
    .Y(_0118_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _1915_ (.Y(_0119_),
    .A(net345),
    .B(net341),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _1916_ (.A(_0002_),
    .B(net414),
    .X(_0120_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _1917_ (.VSS(VGND),
    .VDD(VPWR),
    .B2(_0120_),
    .C1(net314),
    .B1(_0119_),
    .A1(net417),
    .Y(_0121_),
    .A2(_0115_));
 sg13g2_a21oi_1 _1918_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0214_),
    .A2(net314),
    .Y(_0061_),
    .B1(_0121_));
 sg13g2_and2_1 _1919_ (.A(_0003_),
    .B(net412),
    .X(_0122_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _1920_ (.VSS(VGND),
    .VDD(VPWR),
    .B2(_0122_),
    .C1(net315),
    .B1(_0119_),
    .A1(net418),
    .Y(_0123_),
    .A2(_0114_));
 sg13g2_a21oi_1 _1921_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0213_),
    .A2(net315),
    .Y(_0062_),
    .B1(_0123_));
 sg13g2_nand3_1 _1922_ (.B(net412),
    .C(_0119_),
    .A(net82),
    .Y(_0124_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1923_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net417),
    .A2(_0113_),
    .Y(_0125_),
    .B1(net314));
 sg13g2_a22oi_1 _1924_ (.Y(_0063_),
    .B1(_0124_),
    .B2(_0125_),
    .A2(net314),
    .A1(_0212_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _1925_ (.A(_0004_),
    .B(net414),
    .X(_0126_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _1926_ (.VSS(VGND),
    .VDD(VPWR),
    .B2(_0126_),
    .C1(net315),
    .B1(_0119_),
    .A1(net3),
    .Y(_0127_),
    .A2(net418));
 sg13g2_a21oi_1 _1927_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0211_),
    .A2(net315),
    .Y(_0064_),
    .B1(_0127_));
 sg13g2_nand2_1 _1928_ (.Y(_0128_),
    .A(\voffset[4] ),
    .B(net314),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _1929_ (.B(net417),
    .C(_0117_),
    .A(net4),
    .Y(_0129_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _1930_ (.B(_0128_),
    .C(_0129_),
    .A(_0124_),
    .Y(_0065_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _1931_ (.A(_0006_),
    .B(net412),
    .X(_0130_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _1932_ (.Y(_0131_),
    .B1(_0119_),
    .B2(_0130_),
    .A2(net418),
    .A1(net5),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1933_ (.Y(_0132_),
    .A(net78),
    .B(net314),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1934_ (.B1(_0132_),
    .VDD(VPWR),
    .Y(_0066_),
    .VSS(VGND),
    .A1(net314),
    .A2(_0131_));
 sg13g2_nand3_1 _1935_ (.B(net413),
    .C(_0119_),
    .A(_0007_),
    .Y(_0133_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1936_ (.B1(_0133_),
    .VDD(VPWR),
    .Y(_0134_),
    .VSS(VGND),
    .A1(_0199_),
    .A2(net413));
 sg13g2_mux2_1 _1937_ (.A0(_0134_),
    .A1(net94),
    .S(net315),
    .X(_0067_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _1938_ (.B(net413),
    .C(_0119_),
    .A(_0008_),
    .Y(_0135_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1939_ (.B1(_0135_),
    .VDD(VPWR),
    .Y(_0136_),
    .VSS(VGND),
    .A1(_0210_),
    .A2(net412));
 sg13g2_mux2_1 _1940_ (.A0(_0136_),
    .A1(net90),
    .S(net314),
    .X(_0068_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1941_ (.A(net402),
    .B(net404),
    .Y(_0137_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _1942_ (.B(net393),
    .C(_0305_),
    .A(_0205_),
    .Y(_0138_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0137_));
 sg13g2_nor4_1 _1943_ (.A(_0204_),
    .B(net399),
    .C(_0223_),
    .D(_0138_),
    .Y(_0139_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _1944_ (.Y(_0140_),
    .A(net365),
    .B(net417),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _1945_ (.B(net404),
    .C(net399),
    .A(net402),
    .Y(_0141_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1946_ (.A(_0218_),
    .B(_0141_),
    .Y(_0142_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1947_ (.Y(_0143_),
    .A(_0224_),
    .B(_0142_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1948_ (.A(_0139_),
    .B(_0140_),
    .Y(_0144_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _1949_ (.A(_0222_),
    .B(_0137_),
    .X(_0145_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _1950_ (.A(_0204_),
    .B(_0205_),
    .C(_0206_),
    .D(_0262_),
    .Y(_0146_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1951_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0145_),
    .A2(_0146_),
    .Y(_0147_),
    .B1(net414));
 sg13g2_nor4_1 _1952_ (.A(net398),
    .B(net396),
    .C(_0206_),
    .D(_0262_),
    .Y(_0148_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1953_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0145_),
    .A2(_0148_),
    .Y(_0149_),
    .B1(net365));
 sg13g2_a22oi_1 _1954_ (.Y(_0150_),
    .B1(_0147_),
    .B2(_0149_),
    .A2(_0144_),
    .A1(_0143_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1955_ (.A(net76),
    .B(_0150_),
    .Y(_0151_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1956_ (.Y(_0152_),
    .B(_0147_),
    .A_N(_0139_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1957_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0150_),
    .A2(_0152_),
    .Y(_0069_),
    .B1(_0151_));
 sg13g2_nor2_1 _1958_ (.A(_0933_),
    .B(_0961_),
    .Y(_0153_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1959_ (.B1(net417),
    .VDD(VPWR),
    .Y(_0154_),
    .VSS(VGND),
    .A1(net381),
    .A2(_0153_));
 sg13g2_a21oi_1 _1960_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net380),
    .A2(_0932_),
    .Y(_0070_),
    .B1(_0154_));
 sg13g2_a21oi_1 _1961_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net380),
    .A2(_0932_),
    .Y(_0155_),
    .B1(net379));
 sg13g2_and3_1 _1962_ (.X(_0156_),
    .A(net379),
    .B(net380),
    .C(_0932_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _1963_ (.A(net411),
    .B(_0155_),
    .C(_0156_),
    .Y(_0071_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _1964_ (.Y(_0157_),
    .B(net418),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_0962_));
 sg13g2_nand2_1 _1965_ (.Y(_0158_),
    .A(\v[2] ),
    .B(net380),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _1966_ (.B(net379),
    .C(net380),
    .A(net378),
    .Y(_0159_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1967_ (.Y(_0160_),
    .A(net378),
    .B(_0156_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1968_ (.A(_0157_),
    .B(_0160_),
    .Y(_0072_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1969_ (.Y(_0161_),
    .A(net127),
    .B(_0934_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _1970_ (.Y(_0162_),
    .A(net417),
    .B(_0153_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _1971_ (.VDD(VPWR),
    .Y(_0163_),
    .A(_0162_),
    .VSS(VGND));
 sg13g2_nor2_1 _1972_ (.A(_0194_),
    .B(_0159_),
    .Y(_0164_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1973_ (.Y(_0165_),
    .A(_0194_),
    .B(_0159_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1974_ (.B1(_0161_),
    .VDD(VPWR),
    .Y(_0073_),
    .VSS(VGND),
    .A1(_0162_),
    .A2(_0165_));
 sg13g2_a21oi_1 _1975_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0932_),
    .A2(_0164_),
    .Y(_0166_),
    .B1(net123));
 sg13g2_and3_1 _1976_ (.X(_0167_),
    .A(\v[4] ),
    .B(_0932_),
    .C(_0164_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1977_ (.Y(_0168_),
    .A(\v[4] ),
    .B(_0164_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _1978_ (.A(net414),
    .B(_0166_),
    .C(_0167_),
    .Y(_0074_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1979_ (.Y(_0169_),
    .A(net377),
    .B(_0934_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1980_ (.Y(_0170_),
    .A(net85),
    .B(_0168_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1981_ (.B1(_0169_),
    .VDD(VPWR),
    .Y(_0075_),
    .VSS(VGND),
    .A1(_0162_),
    .A2(_0170_));
 sg13g2_a21oi_1 _1982_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net376),
    .A2(_0167_),
    .Y(_0171_),
    .B1(net121));
 sg13g2_nor2b_1 _1983_ (.A(_0235_),
    .B_N(_0167_),
    .Y(_0172_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1984_ (.A(_0235_),
    .B(_0168_),
    .Y(_0173_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _1985_ (.A(net412),
    .B(net122),
    .C(_0172_),
    .Y(_0076_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1986_ (.Y(_0174_),
    .A(net124),
    .B(_0172_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1987_ (.A(_0157_),
    .B(_0174_),
    .Y(_0077_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1988_ (.Y(_0175_),
    .A(_0229_),
    .B(_0173_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _1989_ (.Y(_0176_),
    .B1(_0163_),
    .B2(_0175_),
    .A2(_0934_),
    .A1(net375),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1990_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net124),
    .A2(_0173_),
    .Y(_0177_),
    .B1(net375));
 sg13g2_nor2_1 _1991_ (.A(_0176_),
    .B(net125),
    .Y(_0078_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1992_ (.Y(_0178_),
    .A(net105),
    .B(_0934_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1993_ (.Y(_0179_),
    .A(_0017_),
    .B(_0175_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1994_ (.B1(_0178_),
    .VDD(VPWR),
    .Y(_0079_),
    .VSS(VGND),
    .A1(_0162_),
    .A2(_0179_));
 sg13g2_o21ai_1 _1995_ (.B1(net417),
    .VDD(VPWR),
    .Y(_0180_),
    .VSS(VGND),
    .A1(_0238_),
    .A2(_0950_));
 sg13g2_nor3_1 _1996_ (.A(_0194_),
    .B(net378),
    .C(net380),
    .Y(_0181_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _1997_ (.B(_0237_),
    .C(_0181_),
    .A(net379),
    .Y(_0182_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1998_ (.A(net365),
    .B(_0180_),
    .Y(_0183_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _1999_ (.A(\v[3] ),
    .B(net379),
    .C(_0230_),
    .D(_0158_),
    .Y(_0184_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2000_ (.A(net378),
    .B(_0230_),
    .Y(_0185_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _2001_ (.B(_0233_),
    .C(_0239_),
    .A(\v[3] ),
    .Y(_0186_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0185_));
 sg13g2_a21oi_1 _2002_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0233_),
    .A2(_0184_),
    .Y(_0187_),
    .B1(_0140_));
 sg13g2_a22oi_1 _2003_ (.Y(_0188_),
    .B1(_0186_),
    .B2(_0187_),
    .A2(_0183_),
    .A1(_0182_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2004_ (.A(net80),
    .B(_0188_),
    .Y(_0189_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2005_ (.Y(_0190_),
    .B(_0186_),
    .A_N(_0180_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2006_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0188_),
    .A2(_0190_),
    .Y(_0080_),
    .B1(_0189_));
 sg13g2_nor2_1 _2007_ (.A(_0249_),
    .B(_0253_),
    .Y(_0081_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2008_ (.A(net374),
    .B(net410),
    .Y(_0191_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2009_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0209_),
    .A2(net410),
    .Y(_0083_),
    .B1(_0191_));
 sg13g2_o21ai_1 _2010_ (.B1(_0247_),
    .VDD(VPWR),
    .Y(_0084_),
    .VSS(VGND),
    .A1(_0208_),
    .A2(net410));
 sg13g2_nand2_1 _2011_ (.Y(_0192_),
    .A(net89),
    .B(net418),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2012_ (.B1(_0192_),
    .VDD(VPWR),
    .Y(_0085_),
    .VSS(VGND),
    .A1(_0198_),
    .A2(net418));
 sg13g2_nand2_1 _2013_ (.Y(_0193_),
    .A(net81),
    .B(_0243_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2014_ (.B1(_0193_),
    .VDD(VPWR),
    .Y(_0086_),
    .VSS(VGND),
    .A1(_0199_),
    .A2(_0243_));
 sg13g2_mux2_1 _2015_ (.A0(net112),
    .A1(net7),
    .S(net410),
    .X(_0087_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2016_ (.A0(net120),
    .A1(net8),
    .S(net410),
    .X(_0088_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2017_ (.A0(net116),
    .A1(net9),
    .S(net416),
    .X(_0089_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2018_ (.B1(_0140_),
    .VDD(VPWR),
    .Y(_0090_),
    .VSS(VGND),
    .A1(_0210_),
    .A2(net418));
 sg13g2_dfrbp_1 _2019_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net26),
    .D(_0000_),
    .Q_N(_0998_),
    .Q(_0002_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbp_1 _2020_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net18),
    .D(net93),
    .Q_N(_0997_),
    .Q(_0003_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbp_1 _2021_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net58),
    .D(net110),
    .Q_N(_0996_),
    .Q(_0004_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbp_1 _2022_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net57),
    .D(_0037_),
    .Q_N(_0995_),
    .Q(_0006_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbp_1 _2023_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net56),
    .D(_0038_),
    .Q_N(_0994_),
    .Q(_0007_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbp_1 _2024_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net55),
    .D(_0039_),
    .Q_N(_0035_),
    .Q(\h[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbp_1 _2025_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net54),
    .D(_0040_),
    .Q_N(_0020_),
    .Q(\h[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbp_1 _2026_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net53),
    .D(_0041_),
    .Q_N(_0021_),
    .Q(\h[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbp_1 _2027_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net52),
    .D(_0042_),
    .Q_N(_0013_),
    .Q(\h[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbp_1 _2028_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net51),
    .D(_0043_),
    .Q_N(_0023_),
    .Q(\h[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbp_1 _2029_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net50),
    .D(_0044_),
    .Q_N(_0015_),
    .Q(\h[5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbp_1 _2030_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net49),
    .D(_0045_),
    .Q_N(_0026_),
    .Q(\h[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbp_1 _2031_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net48),
    .D(_0046_),
    .Q_N(_0028_),
    .Q(\h[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbp_1 _2032_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net47),
    .D(_0047_),
    .Q_N(_0014_),
    .Q(\h[8] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbp_1 _2033_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net46),
    .D(_0048_),
    .Q_N(_0031_),
    .Q(\h[9] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbp_1 _2034_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net45),
    .D(net88),
    .Q_N(_0034_),
    .Q(\rampc[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbp_1 _2035_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net43),
    .D(_0050_),
    .Q_N(_0022_),
    .Q(\rampc[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbp_1 _2036_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net41),
    .D(_0051_),
    .Q_N(_0024_),
    .Q(\rampc[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbp_1 _2037_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net39),
    .D(_0052_),
    .Q_N(_0025_),
    .Q(\rampc[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbp_1 _2038_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net37),
    .D(_0053_),
    .Q_N(_0027_),
    .Q(\rampc[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbp_1 _2039_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net35),
    .D(_0054_),
    .Q_N(_0029_),
    .Q(\rampc[5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbp_1 _2040_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net33),
    .D(_0055_),
    .Q_N(_0030_),
    .Q(\rampc[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbp_1 _2041_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net31),
    .D(_0056_),
    .Q_N(_0032_),
    .Q(\rampc[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbp_1 _2042_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net29),
    .D(_0057_),
    .Q_N(_0033_),
    .Q(\t[8] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbp_1 _2043_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net27),
    .D(_0058_),
    .Q_N(_0009_),
    .Q(\t[9] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbp_1 _2044_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net25),
    .D(_0059_),
    .Q_N(_0010_),
    .Q(\t[10] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbp_1 _2045_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net23),
    .D(net100),
    .Q_N(_0993_),
    .Q(\t[11] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbp_1 _2046_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net21),
    .D(net102),
    .Q_N(_0992_),
    .Q(\voffset[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbp_1 _2047_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net20),
    .D(net97),
    .Q_N(_0991_),
    .Q(\voffset[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbp_1 _2048_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net19),
    .D(_0063_),
    .Q_N(_0990_),
    .Q(\voffset[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbp_1 _2049_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net17),
    .D(net104),
    .Q_N(_0989_),
    .Q(\voffset[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbp_1 _2050_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net73),
    .D(net83),
    .Q_N(_0988_),
    .Q(\voffset[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbp_1 _2051_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net72),
    .D(net79),
    .Q_N(_0987_),
    .Q(\voffset[5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbp_1 _2052_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net71),
    .D(net95),
    .Q_N(_0986_),
    .Q(\voffset[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbp_1 _2053_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net70),
    .D(net91),
    .Q_N(_0985_),
    .Q(\voffset[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbp_1 _2054_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net69),
    .D(_0069_),
    .Q_N(hsync),
    .Q(\vga_sync.hsync ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbp_1 _2055_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net68),
    .D(_0070_),
    .Q_N(_0984_),
    .Q(\v[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbp_1 _2056_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net66),
    .D(_0071_),
    .Q_N(_0983_),
    .Q(\v[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbp_1 _2057_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net64),
    .D(_0072_),
    .Q_N(_0982_),
    .Q(\v[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbp_1 _2058_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net62),
    .D(_0073_),
    .Q_N(_0981_),
    .Q(\v[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbp_1 _2059_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net60),
    .D(_0074_),
    .Q_N(_0980_),
    .Q(\v[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbp_1 _2060_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net44),
    .D(net86),
    .Q_N(_0019_),
    .Q(\v[5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbp_1 _2061_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net40),
    .D(_0076_),
    .Q_N(_0979_),
    .Q(\v[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbp_1 _2062_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net36),
    .D(_0077_),
    .Q_N(_0978_),
    .Q(\v[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbp_1 _2063_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net32),
    .D(net126),
    .Q_N(_0977_),
    .Q(\v[8] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbp_1 _2064_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net28),
    .D(net106),
    .Q_N(_0017_),
    .Q(\v[9] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbp_1 _2065_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net24),
    .D(_0080_),
    .Q_N(_0976_),
    .Q(\vga_sync.vsync ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbp_1 _2066_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net22),
    .D(_0081_),
    .Q_N(_0975_),
    .Q(_0008_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbp_1 _2067_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net67),
    .D(_0082_),
    .Q_N(_0974_),
    .Q(_0005_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbp_1 _2068_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net65),
    .D(_0083_),
    .Q_N(_0973_),
    .Q(registered),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbp_1 _2069_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net63),
    .D(_0084_),
    .Q_N(_0018_),
    .Q(gate),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbp_1 _2070_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net61),
    .D(_0085_),
    .Q_N(_0011_),
    .Q(\divider[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbp_1 _2071_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net59),
    .D(_0086_),
    .Q_N(_0012_),
    .Q(\divider[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbp_1 _2072_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net42),
    .D(_0087_),
    .Q_N(_0972_),
    .Q(\mode[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbp_1 _2073_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net38),
    .D(_0088_),
    .Q_N(_0971_),
    .Q(\mode[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbp_1 _2074_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net34),
    .D(_0089_),
    .Q_N(_0016_),
    .Q(\mode[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbp_1 _2075_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net30),
    .D(_0090_),
    .Q_N(_0970_),
    .Q(\vga_sync.mode ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_tiehi _2020__18 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net18));
 sg13g2_tiehi _2048__19 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net19));
 sg13g2_tiehi _2047__20 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net20));
 sg13g2_tiehi _2046__21 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net21));
 sg13g2_tiehi _2066__22 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net22));
 sg13g2_tiehi _2045__23 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net23));
 sg13g2_tiehi _2065__24 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net24));
 sg13g2_tiehi _2044__25 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net25));
 sg13g2_tiehi _2019__26 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net26));
 sg13g2_tiehi _2043__27 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net27));
 sg13g2_tiehi _2064__28 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net28));
 sg13g2_tiehi _2042__29 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net29));
 sg13g2_tiehi _2075__30 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net30));
 sg13g2_tiehi _2041__31 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net31));
 sg13g2_tiehi _2063__32 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net32));
 sg13g2_tiehi _2040__33 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net33));
 sg13g2_tiehi _2074__34 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net34));
 sg13g2_tiehi _2039__35 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net35));
 sg13g2_tiehi _2062__36 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net36));
 sg13g2_tiehi _2038__37 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net37));
 sg13g2_tiehi _2073__38 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net38));
 sg13g2_tiehi _2037__39 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net39));
 sg13g2_tiehi _2061__40 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net40));
 sg13g2_tiehi _2036__41 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net41));
 sg13g2_tiehi _2072__42 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net42));
 sg13g2_tiehi _2035__43 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net43));
 sg13g2_tiehi _2060__44 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net44));
 sg13g2_tiehi _2034__45 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net45));
 sg13g2_tiehi _2033__46 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net46));
 sg13g2_tiehi _2032__47 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net47));
 sg13g2_tiehi _2031__48 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net48));
 sg13g2_tiehi _2030__49 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net49));
 sg13g2_tiehi _2029__50 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net50));
 sg13g2_tiehi _2028__51 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net51));
 sg13g2_tiehi _2027__52 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net52));
 sg13g2_tiehi _2026__53 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net53));
 sg13g2_tiehi _2025__54 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net54));
 sg13g2_tiehi _2024__55 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net55));
 sg13g2_tiehi _2023__56 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net56));
 sg13g2_tiehi _2022__57 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net57));
 sg13g2_tiehi _2021__58 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net58));
 sg13g2_tiehi _2071__59 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net59));
 sg13g2_tiehi _2059__60 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net60));
 sg13g2_tiehi _2070__61 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net61));
 sg13g2_tiehi _2058__62 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net62));
 sg13g2_tiehi _2069__63 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net63));
 sg13g2_tiehi _2057__64 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net64));
 sg13g2_tiehi _2068__65 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net65));
 sg13g2_tiehi _2056__66 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net66));
 sg13g2_tiehi _2067__67 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net67));
 sg13g2_tiehi _2055__68 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net68));
 sg13g2_tiehi _2054__69 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net69));
 sg13g2_tiehi _2053__70 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net70));
 sg13g2_tiehi _2052__71 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net71));
 sg13g2_tiehi _2051__72 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net72));
 sg13g2_tiehi _2050__73 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net73));
 sg13g2_tiehi controller_74 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net74));
 sg13g2_tiehi controller_75 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net75));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_tielo controller_12 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net12));
 sg13g2_tielo controller_13 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net13));
 sg13g2_tielo controller_14 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net14));
 sg13g2_tielo controller_15 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net15));
 sg13g2_tielo controller_16 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net16));
 sg13g2_tiehi _2049__17 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net17));
 sg13g2_buf_2 _2141_ (.A(b6),
    .X(db[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 _2142_ (.A(b7),
    .X(db[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 _2143_ (.A(g6),
    .X(dg[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 _2144_ (.A(g7),
    .X(dg[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _2145_ (.A(r6),
    .X(dr[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _2146_ (.A(r7),
    .X(dr[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout314 (.A(_0118_),
    .X(net314),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout315 (.A(_0118_),
    .X(net315),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout316 (.A(_0321_),
    .X(net316),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout317 (.A(_0321_),
    .X(net317),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout318 (.A(net319),
    .X(net318),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout319 (.A(_0318_),
    .X(net319),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_4 fanout320 (.X(net320),
    .A(_0322_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout321 (.A(_0322_),
    .X(net321),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout322 (.A(net323),
    .X(net322),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_4 fanout323 (.X(net323),
    .A(_0301_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout324 (.A(_0344_),
    .X(net324),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout325 (.A(_0343_),
    .X(net325),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout326 (.A(_0343_),
    .X(net326),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout327 (.A(_0303_),
    .X(net327),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout328 (.A(net329),
    .X(net328),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout329 (.A(net330),
    .X(net329),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout330 (.A(net331),
    .X(net330),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout331 (.A(_0263_),
    .X(net331),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_4 fanout332 (.X(net332),
    .A(net334),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout333 (.A(net334),
    .X(net333),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout334 (.A(net336),
    .X(net334),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_4 fanout335 (.X(net335),
    .A(net336),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout336 (.A(_0258_),
    .X(net336),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout337 (.A(_0597_),
    .X(net337),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout338 (.A(_0597_),
    .X(net338),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout339 (.A(net341),
    .X(net339),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout340 (.A(net341),
    .X(net340),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout341 (.A(_0372_),
    .X(net341),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout342 (.A(_0371_),
    .X(net342),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout343 (.A(_0371_),
    .X(net343),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout344 (.A(net345),
    .X(net344),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout345 (.A(net346),
    .X(net345),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout346 (.A(_0353_),
    .X(net346),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout347 (.A(net349),
    .X(net347),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout348 (.A(net349),
    .X(net348),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout349 (.A(_0349_),
    .X(net349),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout350 (.A(net351),
    .X(net350),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout351 (.A(_0348_),
    .X(net351),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout352 (.A(net354),
    .X(net352),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout353 (.A(net354),
    .X(net353),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout354 (.A(_0336_),
    .X(net354),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout355 (.A(net356),
    .X(net355),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout356 (.A(_0306_),
    .X(net356),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout357 (.A(net358),
    .X(net357),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout358 (.A(net359),
    .X(net358),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout359 (.A(net360),
    .X(net359),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout360 (.A(_0257_),
    .X(net360),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout361 (.A(_0256_),
    .X(net361),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout362 (.A(_0256_),
    .X(net362),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout363 (.A(_0329_),
    .X(net363),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_4 fanout364 (.X(net364),
    .A(_0307_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_4 fanout365 (.X(net365),
    .A(net146),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout366 (.A(\vga_sync.mode ),
    .X(net366),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout367 (.A(_0016_),
    .X(net367),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_4 fanout368 (.X(net368),
    .A(\divider[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout369 (.A(\divider[0] ),
    .X(net369),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_4 fanout370 (.X(net370),
    .A(net143),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout371 (.A(gate),
    .X(net371),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout372 (.A(net374),
    .X(net372),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout373 (.A(net374),
    .X(net373),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout374 (.A(net134),
    .X(net374),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout375 (.A(\v[8] ),
    .X(net375),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout376 (.A(\v[5] ),
    .X(net376),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout377 (.A(\v[5] ),
    .X(net377),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout378 (.A(net140),
    .X(net378),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout379 (.A(net135),
    .X(net379),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout380 (.A(net133),
    .X(net380),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout381 (.A(net133),
    .X(net381),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout382 (.A(_0032_),
    .X(net382),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout383 (.A(net148),
    .X(net383),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_4 fanout384 (.X(net384),
    .A(net151),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout385 (.A(net145),
    .X(net385),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout386 (.A(\rampc[5] ),
    .X(net386),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout387 (.A(net144),
    .X(net387),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout388 (.A(\rampc[4] ),
    .X(net388),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout389 (.A(\rampc[3] ),
    .X(net389),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout390 (.A(\rampc[3] ),
    .X(net390),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout391 (.A(net150),
    .X(net391),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout392 (.A(\rampc[1] ),
    .X(net392),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_4 fanout393 (.X(net393),
    .A(\h[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout394 (.A(net138),
    .X(net394),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_4 fanout395 (.X(net395),
    .A(\h[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout396 (.A(net130),
    .X(net396),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout397 (.A(net398),
    .X(net397),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout398 (.A(net128),
    .X(net398),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout399 (.A(\h[4] ),
    .X(net399),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_4 fanout400 (.X(net400),
    .A(\h[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_4 fanout401 (.X(net401),
    .A(net402),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout402 (.A(\h[3] ),
    .X(net402),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_4 fanout403 (.X(net403),
    .A(net136),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout404 (.A(\h[2] ),
    .X(net404),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout405 (.A(net406),
    .X(net405),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout406 (.A(net407),
    .X(net406),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout407 (.A(net147),
    .X(net407),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_4 fanout408 (.X(net408),
    .A(\h[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout409 (.A(\h[0] ),
    .X(net409),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout410 (.A(net411),
    .X(net410),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_4 fanout411 (.X(net411),
    .A(net416),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout412 (.A(net413),
    .X(net412),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout413 (.A(net414),
    .X(net413),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout414 (.A(net415),
    .X(net414),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout415 (.A(net416),
    .X(net415),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout416 (.A(_0244_),
    .X(net416),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_4 fanout417 (.X(net417),
    .A(net418),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_4 fanout418 (.X(net418),
    .A(_0243_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 input1 (.A(ena),
    .X(net1),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input2 (.A(rst_n),
    .X(net2),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 input3 (.A(ui_in[0]),
    .X(net3),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 input4 (.A(ui_in[1]),
    .X(net4),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 input5 (.A(ui_in[2]),
    .X(net5),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 input6 (.A(ui_in[3]),
    .X(net6),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 input7 (.A(ui_in[4]),
    .X(net7),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 input8 (.A(ui_in[5]),
    .X(net8),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 input9 (.A(ui_in[6]),
    .X(net9),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input10 (.A(ui_in[7]),
    .X(net10),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_tielo controller_11 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net11));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 clkload0 (.VDD(VPWR),
    .A(clknet_4_3_0_clk),
    .VSS(VGND));
 sg13g2_inv_1 clkload1 (.VDD(VPWR),
    .A(clknet_4_5_0_clk),
    .VSS(VGND));
 sg13g2_inv_1 clkload2 (.VDD(VPWR),
    .A(clknet_4_7_0_clk),
    .VSS(VGND));
 sg13g2_inv_1 clkload3 (.VDD(VPWR),
    .A(clknet_4_9_0_clk),
    .VSS(VGND));
 sg13g2_inv_1 clkload4 (.VDD(VPWR),
    .A(clknet_4_11_0_clk),
    .VSS(VGND));
 sg13g2_inv_1 clkload5 (.VDD(VPWR),
    .A(clknet_4_13_0_clk),
    .VSS(VGND));
 sg13g2_inv_1 clkload6 (.VDD(VPWR),
    .A(clknet_4_15_0_clk),
    .VSS(VGND));
 sg13g2_dlygate4sd3_1 hold1 (.A(\vga_sync.hsync ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0035_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold3 (.A(\voffset[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0066_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold5 (.A(\vga_sync.vsync ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold6 (.A(\divider[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0005_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0065_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold9 (.A(\voffset[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0019_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0075_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0034_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0049_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold14 (.A(\divider[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold15 (.A(\voffset[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0068_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0011_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0001_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold19 (.A(\voffset[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0067_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold21 (.A(\voffset[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0062_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold23 (.A(\t[11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0111_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0060_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold26 (.A(\voffset[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0061_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold28 (.A(\voffset[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0064_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold30 (.A(\v[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0079_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold32 (.A(_0014_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0949_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold34 (.A(_0012_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0036_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0018_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold37 (.A(\mode[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold38 (.A(\t[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0106_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold40 (.A(\t[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold41 (.A(\mode[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold42 (.A(_0023_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold43 (.A(\rampc[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold44 (.A(_0965_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold45 (.A(\mode[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold46 (.A(\v[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold47 (.A(_0171_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold48 (.A(\v[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold49 (.A(\v[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold50 (.A(_0177_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0078_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold52 (.A(\v[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold53 (.A(\h[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold54 (.A(_0942_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold55 (.A(\h[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold56 (.A(_0021_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold57 (.A(_0938_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold58 (.A(\v[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold59 (.A(registered),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold60 (.A(\v[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold61 (.A(\h[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold62 (.A(\h[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold63 (.A(\h[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold64 (.A(_0945_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold65 (.A(\v[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold66 (.A(_0024_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold67 (.A(_0093_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold68 (.A(gate),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold69 (.A(\rampc[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold70 (.A(\rampc[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold71 (.A(\vga_sync.mode ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold72 (.A(\h[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold73 (.A(\rampc[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold74 (.A(\t[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold75 (.A(\rampc[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold76 (.A(\rampc[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net151));
 sg13g2_decap_8 FILLER_0_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_178 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_41 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_13 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_15 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_58 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_78 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_29 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_86 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_12 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_37 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_178 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_27 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_107 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_65 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_20 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_58 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_50 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_27 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_34 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_48 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_12 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_23 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_29 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_37 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_31 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_23 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_66 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_80 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_38 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_107 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_15 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_36 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_22 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_36 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_38 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_59 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_17 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_19 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_59 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_86 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_92 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_26 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_62 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_19 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_38 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_178 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_9 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_86 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_320 (.VDD(VPWR),
    .VSS(VGND));
 assign uio_oe[0] = net74;
 assign uio_oe[1] = net75;
 assign uio_out2 = net11;
 assign uio_out3 = net12;
 assign uio_out4 = net13;
 assign uio_out5 = net14;
 assign uio_out6 = net15;
 assign uio_out7 = net16;
endmodule
