* NGSPICE file created from r2r_dac.ext - technology: ihp-sg13g2

.subckt rhigh a_0_1200# a_0_n86#
X0 a_0_1200# a_0_n86# rhigh l=6u w=1u
.ends

.subckt resistors B rhigh_0[0]/a_0_1200# rhigh_0[23]/a_0_n86# rhigh_0[11]/a_0_1200#
+ rhigh_0[21]/a_0_1200# rhigh_0[6]/a_0_n86# rhigh_0[1]/a_0_1200# rhigh_0[2]/a_0_n86#
+ rhigh_0[12]/a_0_1200# rhigh_0[18]/a_0_n86# rhigh_0[22]/a_0_1200# rhigh_0[2]/a_0_1200#
+ rhigh_0[14]/a_0_n86# rhigh_0[13]/a_0_1200# rhigh_0[10]/a_0_n86# rhigh_0[23]/a_0_1200#
+ rhigh_0[24]/a_0_n86# rhigh_0[3]/a_0_1200# rhigh_0[20]/a_0_n86# rhigh_0[14]/a_0_1200#
+ rhigh_0[7]/a_0_n86# rhigh_0[3]/a_0_n86# rhigh_0[24]/a_0_1200# rhigh_0[4]/a_0_1200#
+ rhigh_0[19]/a_0_n86# rhigh_0[15]/a_0_1200# rhigh_0[15]/a_0_n86# rhigh_0[5]/a_0_1200#
+ rhigh_0[11]/a_0_n86# rhigh_0[16]/a_0_1200# rhigh_0[21]/a_0_n86# rhigh_0[8]/a_0_n86#
+ rhigh_0[4]/a_0_n86# rhigh_0[6]/a_0_1200# rhigh_0[0]/a_0_n86# rhigh_0[17]/a_0_1200#
+ rhigh_0[18]/a_0_1200# rhigh_0[7]/a_0_1200# rhigh_0[16]/a_0_n86# rhigh_0[12]/a_0_n86#
+ rhigh_0[19]/a_0_1200# rhigh_0[8]/a_0_1200# rhigh_0[9]/a_0_n86# rhigh_0[22]/a_0_n86#
+ rhigh_0[5]/a_0_n86# rhigh_0[9]/a_0_1200# rhigh_0[1]/a_0_n86# rhigh_0[17]/a_0_n86#
+ rhigh_0[10]/a_0_1200# rhigh_0[13]/a_0_n86# rhigh_0[20]/a_0_1200#
Xrhigh_0[0] rhigh_0[0]/a_0_1200# rhigh_0[0]/a_0_n86# rhigh
Xrhigh_0[1] rhigh_0[1]/a_0_1200# rhigh_0[1]/a_0_n86# rhigh
Xrhigh_0[2] rhigh_0[2]/a_0_1200# rhigh_0[2]/a_0_n86# rhigh
Xrhigh_0[3] rhigh_0[3]/a_0_1200# rhigh_0[3]/a_0_n86# rhigh
Xrhigh_0[4] rhigh_0[4]/a_0_1200# rhigh_0[4]/a_0_n86# rhigh
Xrhigh_0[5] rhigh_0[5]/a_0_1200# rhigh_0[5]/a_0_n86# rhigh
Xrhigh_0[6] rhigh_0[6]/a_0_1200# rhigh_0[6]/a_0_n86# rhigh
Xrhigh_0[7] rhigh_0[7]/a_0_1200# rhigh_0[7]/a_0_n86# rhigh
Xrhigh_0[8] rhigh_0[8]/a_0_1200# rhigh_0[8]/a_0_n86# rhigh
Xrhigh_0[9] rhigh_0[9]/a_0_1200# rhigh_0[9]/a_0_n86# rhigh
Xrhigh_0[10] rhigh_0[10]/a_0_1200# rhigh_0[10]/a_0_n86# rhigh
Xrhigh_0[11] rhigh_0[11]/a_0_1200# rhigh_0[11]/a_0_n86# rhigh
Xrhigh_0[12] rhigh_0[12]/a_0_1200# rhigh_0[12]/a_0_n86# rhigh
Xrhigh_0[13] rhigh_0[13]/a_0_1200# rhigh_0[13]/a_0_n86# rhigh
Xrhigh_0[14] rhigh_0[14]/a_0_1200# rhigh_0[14]/a_0_n86# rhigh
Xrhigh_0[15] rhigh_0[15]/a_0_1200# rhigh_0[15]/a_0_n86# rhigh
Xrhigh_0[16] rhigh_0[16]/a_0_1200# rhigh_0[16]/a_0_n86# rhigh
Xrhigh_0[17] rhigh_0[17]/a_0_1200# rhigh_0[17]/a_0_n86# rhigh
Xrhigh_0[18] rhigh_0[18]/a_0_1200# rhigh_0[18]/a_0_n86# rhigh
Xrhigh_0[19] rhigh_0[19]/a_0_1200# rhigh_0[19]/a_0_n86# rhigh
Xrhigh_0[20] rhigh_0[20]/a_0_1200# rhigh_0[20]/a_0_n86# rhigh
Xrhigh_0[21] rhigh_0[21]/a_0_1200# rhigh_0[21]/a_0_n86# rhigh
Xrhigh_0[22] rhigh_0[22]/a_0_1200# rhigh_0[22]/a_0_n86# rhigh
Xrhigh_0[23] rhigh_0[23]/a_0_1200# rhigh_0[23]/a_0_n86# rhigh
Xrhigh_0[24] rhigh_0[24]/a_0_1200# rhigh_0[24]/a_0_n86# rhigh
.ends

.subckt r2r_dac GND IN[0] IN[1] IN[2] IN[3] IN[4] IN[5] IN[6] IN[7] OUT
Xresistors_0 GND m1_238_1630# m1_7044_332# m1_3186_1614# m1_6154_1622# m1_1716_324#
+ m1_238_1630# m1_538_330# IN[3] m1_5270_340# OUT m1_830_1624# m1_4080_334# m1_3186_1614#
+ m1_2308_316# OUT m1_7044_332# m1_830_1624# m1_5858_334# m1_4376_1620# m1_2308_316#
+ IN[0] IN[7] m1_1420_1618# m1_5858_334# m1_4376_1620# IN[4] m1_1420_1618# m1_3482_336#
+ m1_4976_1624# IN[6] m1_2308_316# m1_538_330# IN[1] GND m1_4976_1624# IN[5] m1_1420_1618#
+ m1_4080_334# m1_3482_336# m1_4976_1624# m1_2608_1626# IN[2] m1_5858_334# m1_1716_324#
+ m1_2608_1626# m1_538_330# m1_5270_340# m1_3186_1614# m1_4080_334# m1_6154_1622#
+ resistors
.ends

