magic
tech ihp-sg13g2
timestamp 1747537721
<< nwell >>
rect -24 175 312 417
<< pwell >>
rect 15 28 280 142
rect -13 -28 301 28
<< nmos >>
rect 66 57 79 129
rect 117 57 130 129
rect 169 57 182 129
rect 220 57 233 129
<< pmos >>
rect 66 206 79 318
rect 117 206 130 318
rect 169 206 182 318
rect 220 206 233 318
<< ndiff >>
rect 28 115 66 129
rect 28 99 37 115
rect 53 99 66 115
rect 28 81 66 99
rect 28 65 38 81
rect 54 65 66 81
rect 28 57 66 65
rect 79 80 117 129
rect 79 64 90 80
rect 106 64 117 80
rect 79 57 117 64
rect 130 116 169 129
rect 130 100 141 116
rect 157 100 169 116
rect 130 82 169 100
rect 130 66 141 82
rect 157 66 169 82
rect 130 57 169 66
rect 182 121 220 129
rect 182 105 193 121
rect 209 105 220 121
rect 182 57 220 105
rect 233 115 267 129
rect 233 99 244 115
rect 260 99 267 115
rect 233 81 267 99
rect 233 65 244 81
rect 260 65 267 81
rect 233 57 267 65
<< pdiff >>
rect 30 311 66 318
rect 30 295 37 311
rect 53 295 66 311
rect 30 270 66 295
rect 30 254 37 270
rect 53 254 66 270
rect 30 230 66 254
rect 30 214 37 230
rect 53 214 66 230
rect 30 206 66 214
rect 79 311 117 318
rect 79 295 90 311
rect 106 295 117 311
rect 79 271 117 295
rect 79 255 90 271
rect 106 255 117 271
rect 79 231 117 255
rect 79 215 90 231
rect 106 215 117 231
rect 79 206 117 215
rect 130 311 169 318
rect 130 295 141 311
rect 157 295 169 311
rect 130 206 169 295
rect 182 311 220 318
rect 182 295 193 311
rect 209 295 220 311
rect 182 271 220 295
rect 182 255 193 271
rect 209 255 220 271
rect 182 237 220 255
rect 182 221 193 237
rect 209 221 220 237
rect 182 206 220 221
rect 233 311 268 318
rect 233 295 244 311
rect 260 295 268 311
rect 233 271 268 295
rect 233 255 244 271
rect 260 255 268 271
rect 233 237 268 255
rect 233 221 244 237
rect 260 221 268 237
rect 233 206 268 221
<< ndiffc >>
rect 37 99 53 115
rect 38 65 54 81
rect 90 64 106 80
rect 141 100 157 116
rect 141 66 157 82
rect 193 105 209 121
rect 244 99 260 115
rect 244 65 260 81
<< pdiffc >>
rect 37 295 53 311
rect 37 254 53 270
rect 37 214 53 230
rect 90 295 106 311
rect 90 255 106 271
rect 90 215 106 231
rect 141 295 157 311
rect 193 295 209 311
rect 193 255 209 271
rect 193 221 209 237
rect 244 295 260 311
rect 244 255 260 271
rect 244 221 260 237
<< psubdiff >>
rect 0 8 288 15
rect 0 -8 16 8
rect 32 -8 64 8
rect 80 -8 112 8
rect 128 -8 160 8
rect 176 -8 208 8
rect 224 -8 256 8
rect 272 -8 288 8
rect 0 -15 288 -8
<< nsubdiff >>
rect 0 386 288 393
rect 0 370 16 386
rect 32 370 64 386
rect 80 370 112 386
rect 128 370 160 386
rect 176 370 208 386
rect 224 370 256 386
rect 272 370 288 386
rect 0 363 288 370
<< psubdiffcont >>
rect 16 -8 32 8
rect 64 -8 80 8
rect 112 -8 128 8
rect 160 -8 176 8
rect 208 -8 224 8
rect 256 -8 272 8
<< nsubdiffcont >>
rect 16 370 32 386
rect 64 370 80 386
rect 112 370 128 386
rect 160 370 176 386
rect 208 370 224 386
rect 256 370 272 386
<< poly >>
rect 66 318 79 336
rect 117 318 130 336
rect 169 318 182 336
rect 220 318 233 336
rect 66 187 79 206
rect 117 187 130 206
rect 66 180 130 187
rect 66 164 90 180
rect 106 164 130 180
rect 66 156 130 164
rect 66 129 79 156
rect 117 129 130 156
rect 169 199 182 206
rect 220 199 233 206
rect 169 192 233 199
rect 169 176 193 192
rect 209 176 233 192
rect 169 168 233 176
rect 169 129 182 168
rect 220 129 233 168
rect 66 39 79 57
rect 117 39 130 57
rect 169 39 182 57
rect 220 39 233 57
<< polycont >>
rect 90 164 106 180
rect 193 176 209 192
<< metal1 >>
rect 0 386 288 400
rect 0 370 16 386
rect 32 370 64 386
rect 80 370 112 386
rect 128 370 160 386
rect 176 370 208 386
rect 224 370 256 386
rect 272 370 288 386
rect 0 356 288 370
rect 32 311 58 356
rect 32 295 37 311
rect 53 295 58 311
rect 32 270 58 295
rect 32 254 37 270
rect 53 254 58 270
rect 32 230 58 254
rect 32 214 37 230
rect 53 214 58 230
rect 84 311 110 318
rect 84 295 90 311
rect 106 295 110 311
rect 84 271 110 295
rect 135 311 161 356
rect 135 295 141 311
rect 157 295 161 311
rect 135 290 161 295
rect 189 311 215 318
rect 189 295 193 311
rect 209 295 215 311
rect 84 255 90 271
rect 106 255 110 271
rect 84 236 110 255
rect 189 271 215 295
rect 189 255 193 271
rect 209 255 215 271
rect 189 237 215 255
rect 189 236 193 237
rect 84 231 193 236
rect 84 215 90 231
rect 106 221 193 231
rect 209 221 215 237
rect 106 216 215 221
rect 239 311 265 356
rect 239 295 244 311
rect 260 295 265 311
rect 239 271 265 295
rect 239 255 244 271
rect 260 255 265 271
rect 239 237 265 255
rect 239 221 244 237
rect 260 221 265 237
rect 239 216 265 221
rect 106 215 162 216
rect 84 214 162 215
rect 32 212 58 214
rect 82 180 115 192
rect 82 164 90 180
rect 106 164 115 180
rect 82 139 115 164
rect 138 155 162 214
rect 181 192 264 198
rect 181 176 193 192
rect 209 176 264 192
rect 181 173 264 176
rect 138 139 214 155
rect 237 144 264 173
rect 188 121 214 139
rect 32 116 162 120
rect 32 115 141 116
rect 32 99 37 115
rect 53 103 141 115
rect 53 99 58 103
rect 32 81 58 99
rect 135 100 141 103
rect 157 100 162 116
rect 188 105 193 121
rect 209 105 214 121
rect 188 100 214 105
rect 237 115 265 120
rect 32 65 38 81
rect 54 65 58 81
rect 32 50 58 65
rect 85 80 111 85
rect 85 64 90 80
rect 106 64 111 80
rect 85 22 111 64
rect 135 82 162 100
rect 135 66 141 82
rect 157 76 162 82
rect 237 99 244 115
rect 260 99 265 115
rect 237 81 265 99
rect 237 76 244 81
rect 157 66 244 76
rect 135 65 244 66
rect 260 65 265 81
rect 135 53 265 65
rect 0 8 288 22
rect 0 -8 16 8
rect 32 -8 64 8
rect 80 -8 112 8
rect 128 -8 160 8
rect 176 -8 208 8
rect 224 -8 256 8
rect 272 -8 288 8
rect 0 -22 288 -8
<< labels >>
flabel metal1 s 138 139 162 236 0 FreeSans 200 0 0 0 Y
port 2 nsew
flabel metal1 s 0 356 288 400 0 FreeSans 200 0 0 0 VDD
port 3 nsew
flabel metal1 s 181 173 264 198 0 FreeSans 200 0 0 0 A
port 4 nsew
flabel metal1 s 0 -22 288 22 0 FreeSans 200 0 0 0 VSS
port 5 nsew
flabel metal1 s 82 139 115 192 0 FreeSans 200 0 0 0 B
port 6 nsew
<< properties >>
string FIXED_BBOX 0 0 288 378
string GDS_END 183608
string GDS_FILE ../gds/controller.gds
string GDS_START 178738
<< end >>
