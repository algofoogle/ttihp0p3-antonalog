magic
tech ihp-sg13g2
magscale 1 2
timestamp 1747537721
<< nwell >>
rect -48 350 720 834
<< pwell >>
rect 181 284 665 314
rect 159 56 665 284
rect -26 -56 698 56
<< nmos >>
rect 253 140 279 288
rect 366 160 392 288
rect 468 160 494 288
rect 545 160 571 288
<< pmos >>
rect 124 412 150 636
rect 332 436 358 636
rect 443 436 469 636
rect 545 436 571 636
<< ndiff >>
rect 207 258 253 288
rect 185 219 253 258
rect 185 187 199 219
rect 231 187 253 219
rect 185 140 253 187
rect 279 188 366 288
rect 279 156 301 188
rect 333 160 366 188
rect 392 208 468 288
rect 392 176 414 208
rect 446 176 468 208
rect 392 160 468 176
rect 494 160 545 288
rect 571 271 639 288
rect 571 239 593 271
rect 625 239 639 271
rect 571 160 639 239
rect 333 156 352 160
rect 279 140 352 156
<< pdiff >>
rect 56 619 124 636
rect 56 587 70 619
rect 102 587 124 619
rect 56 540 124 587
rect 56 508 70 540
rect 102 508 124 540
rect 56 462 124 508
rect 56 430 70 462
rect 102 430 124 462
rect 56 412 124 430
rect 150 619 218 636
rect 150 587 172 619
rect 204 587 218 619
rect 150 540 218 587
rect 150 508 172 540
rect 204 508 218 540
rect 150 462 218 508
rect 150 430 172 462
rect 204 430 218 462
rect 262 622 332 636
rect 262 590 277 622
rect 309 590 332 622
rect 262 553 332 590
rect 262 521 277 553
rect 309 521 332 553
rect 262 483 332 521
rect 262 451 277 483
rect 309 451 332 483
rect 262 436 332 451
rect 358 622 443 636
rect 358 590 381 622
rect 413 590 443 622
rect 358 553 443 590
rect 358 521 381 553
rect 413 521 443 553
rect 358 483 443 521
rect 358 451 381 483
rect 413 451 443 483
rect 358 436 443 451
rect 469 622 545 636
rect 469 590 491 622
rect 523 590 545 622
rect 469 551 545 590
rect 469 519 491 551
rect 523 519 545 551
rect 469 436 545 519
rect 571 622 639 636
rect 571 590 593 622
rect 625 590 639 622
rect 571 552 639 590
rect 571 520 593 552
rect 625 520 639 552
rect 571 483 639 520
rect 571 451 593 483
rect 625 451 639 483
rect 571 436 639 451
rect 150 412 218 430
<< ndiffc >>
rect 199 187 231 219
rect 301 156 333 188
rect 414 176 446 208
rect 593 239 625 271
<< pdiffc >>
rect 70 587 102 619
rect 70 508 102 540
rect 70 430 102 462
rect 172 587 204 619
rect 172 508 204 540
rect 172 430 204 462
rect 277 590 309 622
rect 277 521 309 553
rect 277 451 309 483
rect 381 590 413 622
rect 381 521 413 553
rect 381 451 413 483
rect 491 590 523 622
rect 491 519 523 551
rect 593 590 625 622
rect 593 520 625 552
rect 593 451 625 483
<< psubdiff >>
rect 0 16 672 30
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 608 16
rect 640 -16 672 16
rect 0 -30 672 -16
<< nsubdiff >>
rect 0 772 672 786
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 608 772
rect 640 740 672 772
rect 0 726 672 740
<< psubdiffcont >>
rect 32 -16 64 16
rect 128 -16 160 16
rect 224 -16 256 16
rect 320 -16 352 16
rect 416 -16 448 16
rect 512 -16 544 16
rect 608 -16 640 16
<< nsubdiffcont >>
rect 32 740 64 772
rect 128 740 160 772
rect 224 740 256 772
rect 320 740 352 772
rect 416 740 448 772
rect 512 740 544 772
rect 608 740 640 772
<< poly >>
rect 124 636 150 672
rect 332 636 358 672
rect 443 636 469 672
rect 545 636 571 672
rect 332 421 358 436
rect 124 374 150 412
rect 332 383 401 421
rect 115 357 185 374
rect 115 325 136 357
rect 168 353 185 357
rect 168 325 279 353
rect 332 351 352 383
rect 384 351 401 383
rect 332 334 401 351
rect 443 400 469 436
rect 443 383 509 400
rect 443 351 460 383
rect 492 351 509 383
rect 443 334 509 351
rect 115 323 279 325
rect 115 308 185 323
rect 253 288 279 323
rect 366 288 392 334
rect 468 288 494 334
rect 545 288 571 436
rect 253 104 279 140
rect 366 124 392 160
rect 468 124 494 160
rect 545 140 571 160
rect 545 123 629 140
rect 545 91 580 123
rect 612 91 629 123
rect 545 74 629 91
<< polycont >>
rect 136 325 168 357
rect 352 351 384 383
rect 460 351 492 383
rect 580 91 612 123
<< metal1 >>
rect 0 772 672 800
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 608 772
rect 640 740 672 772
rect 0 712 672 740
rect 41 619 112 621
rect 41 587 70 619
rect 102 587 112 619
rect 41 540 112 587
rect 41 508 70 540
rect 102 508 112 540
rect 41 462 112 508
rect 41 430 70 462
rect 102 430 112 462
rect 41 419 112 430
rect 162 619 214 712
rect 162 587 172 619
rect 204 587 214 619
rect 162 540 214 587
rect 162 508 172 540
rect 204 508 214 540
rect 162 462 214 508
rect 162 430 172 462
rect 204 430 214 462
rect 162 428 214 430
rect 267 622 319 625
rect 267 590 277 622
rect 309 590 319 622
rect 267 553 319 590
rect 267 521 277 553
rect 309 521 319 553
rect 267 483 319 521
rect 267 451 277 483
rect 309 451 319 483
rect 267 434 319 451
rect 371 622 423 625
rect 371 590 381 622
rect 413 590 423 622
rect 371 553 423 590
rect 371 521 381 553
rect 413 521 423 553
rect 371 483 423 521
rect 481 622 533 712
rect 481 590 491 622
rect 523 590 533 622
rect 481 551 533 590
rect 481 519 491 551
rect 523 519 533 551
rect 481 517 533 519
rect 583 622 635 625
rect 583 590 593 622
rect 625 590 635 622
rect 583 552 635 590
rect 583 520 593 552
rect 625 520 635 552
rect 371 451 381 483
rect 413 481 423 483
rect 583 483 635 520
rect 583 481 593 483
rect 413 451 593 481
rect 625 451 635 483
rect 371 442 635 451
rect 41 229 89 419
rect 267 374 315 434
rect 125 357 315 374
rect 125 325 136 357
rect 168 325 315 357
rect 125 308 315 325
rect 351 383 401 400
rect 351 351 352 383
rect 384 351 401 383
rect 351 314 401 351
rect 443 383 509 400
rect 443 351 460 383
rect 492 351 509 383
rect 443 313 509 351
rect 283 277 315 308
rect 283 244 454 277
rect 584 271 633 282
rect 584 262 593 271
rect 41 219 245 229
rect 41 187 199 219
rect 231 187 245 219
rect 404 208 454 244
rect 41 177 245 187
rect 291 188 343 193
rect 291 156 301 188
rect 333 156 343 188
rect 404 176 414 208
rect 446 176 454 208
rect 404 165 454 176
rect 491 239 593 262
rect 625 239 633 271
rect 491 229 633 239
rect 291 44 343 156
rect 491 44 523 229
rect 562 123 643 193
rect 562 91 580 123
rect 612 91 643 123
rect 562 81 643 91
rect 0 16 672 44
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 608 16
rect 640 -16 672 16
rect 0 -44 672 -16
<< labels >>
flabel metal1 s 351 314 401 400 0 FreeSans 400 0 0 0 B1
port 2 nsew
flabel metal1 s 57 419 112 621 0 FreeSans 400 0 0 0 X
port 3 nsew
flabel metal1 s 0 712 672 800 0 FreeSans 400 0 0 0 VDD
port 4 nsew
flabel metal1 s 0 -44 672 44 0 FreeSans 400 0 0 0 VSS
port 5 nsew
flabel metal1 s 443 313 509 400 0 FreeSans 400 0 0 0 A1
port 6 nsew
flabel metal1 s 562 81 643 193 0 FreeSans 400 0 0 0 A2
port 7 nsew
<< properties >>
string FIXED_BBOX 0 0 672 756
string GDS_END 89618
string GDS_FILE ../gds/controller.gds
string GDS_START 84462
<< end >>
