magic
tech ihp-sg13g2
magscale 1 2
timestamp 1746869612
<< metal1 >>
rect 576 27992 31392 28016
rect 576 27952 4352 27992
rect 4720 27952 12126 27992
rect 12494 27952 19900 27992
rect 20268 27952 27674 27992
rect 28042 27952 31392 27992
rect 576 27928 31392 27952
rect 843 27824 885 27833
rect 843 27784 844 27824
rect 884 27784 885 27824
rect 843 27775 885 27784
rect 1611 27824 1653 27833
rect 1611 27784 1612 27824
rect 1652 27784 1653 27824
rect 1611 27775 1653 27784
rect 17739 27824 17781 27833
rect 17739 27784 17740 27824
rect 17780 27784 17781 27824
rect 17739 27775 17781 27784
rect 17979 27824 18021 27833
rect 17979 27784 17980 27824
rect 18020 27784 18021 27824
rect 17979 27775 18021 27784
rect 30298 27824 30356 27825
rect 30298 27784 30307 27824
rect 30347 27784 30356 27824
rect 30298 27783 30356 27784
rect 1899 27740 1941 27749
rect 1899 27700 1900 27740
rect 1940 27700 1941 27740
rect 1899 27691 1941 27700
rect 3706 27740 3764 27741
rect 3706 27700 3715 27740
rect 3755 27700 3764 27740
rect 3706 27699 3764 27700
rect 4570 27740 4628 27741
rect 4570 27700 4579 27740
rect 4619 27700 4628 27740
rect 4570 27699 4628 27700
rect 12154 27740 12212 27741
rect 12154 27700 12163 27740
rect 12203 27700 12212 27740
rect 12154 27699 12212 27700
rect 14458 27740 14516 27741
rect 14458 27700 14467 27740
rect 14507 27700 14516 27740
rect 14458 27699 14516 27700
rect 1803 27656 1845 27665
rect 1803 27616 1804 27656
rect 1844 27616 1845 27656
rect 1803 27607 1845 27616
rect 1978 27656 2036 27657
rect 1978 27616 1987 27656
rect 2027 27616 2036 27656
rect 1978 27615 2036 27616
rect 2194 27656 2236 27665
rect 2194 27616 2195 27656
rect 2235 27616 2236 27656
rect 2194 27607 2236 27616
rect 2362 27656 2420 27657
rect 2362 27616 2371 27656
rect 2411 27616 2420 27656
rect 2362 27615 2420 27616
rect 2950 27656 2992 27665
rect 2950 27616 2951 27656
rect 2991 27616 2992 27656
rect 2950 27607 2992 27616
rect 3130 27656 3188 27657
rect 3130 27616 3139 27656
rect 3179 27616 3188 27656
rect 3130 27615 3188 27616
rect 4395 27656 4437 27665
rect 4395 27616 4396 27656
rect 4436 27616 4437 27656
rect 4395 27607 4437 27616
rect 4954 27656 5012 27657
rect 4954 27616 4963 27656
rect 5003 27616 5012 27656
rect 4954 27615 5012 27616
rect 7450 27656 7508 27657
rect 7450 27616 7459 27656
rect 7499 27616 7508 27656
rect 7450 27615 7508 27616
rect 9946 27656 10004 27657
rect 9946 27616 9955 27656
rect 9995 27616 10004 27656
rect 9946 27615 10004 27616
rect 14074 27656 14132 27657
rect 14074 27616 14083 27656
rect 14123 27616 14132 27656
rect 14074 27615 14132 27616
rect 15418 27656 15476 27657
rect 15418 27616 15427 27656
rect 15467 27616 15476 27656
rect 15418 27615 15476 27616
rect 17533 27656 17575 27665
rect 18123 27656 18165 27665
rect 17533 27616 17534 27656
rect 17574 27616 17575 27656
rect 17533 27607 17575 27616
rect 17835 27647 17877 27656
rect 17835 27607 17836 27647
rect 17876 27607 17877 27647
rect 18123 27616 18124 27656
rect 18164 27616 18165 27656
rect 18123 27607 18165 27616
rect 18315 27656 18357 27665
rect 18315 27616 18316 27656
rect 18356 27616 18357 27656
rect 18315 27607 18357 27616
rect 19546 27656 19604 27657
rect 19546 27616 19555 27656
rect 19595 27616 19604 27656
rect 19546 27615 19604 27616
rect 22330 27656 22388 27657
rect 22330 27616 22339 27656
rect 22379 27616 22388 27656
rect 22330 27615 22388 27616
rect 26362 27656 26420 27657
rect 26362 27616 26371 27656
rect 26411 27616 26420 27656
rect 26362 27615 26420 27616
rect 26746 27656 26804 27657
rect 26746 27616 26755 27656
rect 26795 27616 26804 27656
rect 26746 27615 26804 27616
rect 27322 27656 27380 27657
rect 27322 27616 27331 27656
rect 27371 27616 27380 27656
rect 27322 27615 27380 27616
rect 30123 27656 30165 27665
rect 30123 27616 30124 27656
rect 30164 27616 30165 27656
rect 30123 27607 30165 27616
rect 30459 27656 30501 27665
rect 30459 27616 30460 27656
rect 30500 27616 30501 27656
rect 30459 27607 30501 27616
rect 30603 27656 30645 27665
rect 30603 27616 30604 27656
rect 30644 27616 30645 27656
rect 30603 27607 30645 27616
rect 30786 27647 30832 27656
rect 30786 27607 30787 27647
rect 30827 27607 30832 27647
rect 17835 27598 17877 27607
rect 30786 27598 30832 27607
rect 7083 27572 7125 27581
rect 7083 27532 7084 27572
rect 7124 27532 7125 27572
rect 7083 27523 7125 27532
rect 9579 27572 9621 27581
rect 9579 27532 9580 27572
rect 9620 27532 9621 27572
rect 9579 27523 9621 27532
rect 15051 27572 15093 27581
rect 15051 27532 15052 27572
rect 15092 27532 15093 27572
rect 15051 27523 15093 27532
rect 18987 27572 19029 27581
rect 18987 27532 18988 27572
rect 19028 27532 19029 27572
rect 18987 27523 19029 27532
rect 19179 27572 19221 27581
rect 19179 27532 19180 27572
rect 19220 27532 19221 27572
rect 19179 27523 19221 27532
rect 21963 27572 22005 27581
rect 21963 27532 21964 27572
rect 22004 27532 22005 27572
rect 21963 27523 22005 27532
rect 26955 27572 26997 27581
rect 26955 27532 26956 27572
rect 26996 27532 26997 27572
rect 26955 27523 26997 27532
rect 30939 27572 30981 27581
rect 30939 27532 30940 27572
rect 30980 27532 30981 27572
rect 30939 27523 30981 27532
rect 1227 27488 1269 27497
rect 1227 27448 1228 27488
rect 1268 27448 1269 27488
rect 1227 27439 1269 27448
rect 2362 27488 2420 27489
rect 2362 27448 2371 27488
rect 2411 27448 2420 27488
rect 2362 27447 2420 27448
rect 2763 27488 2805 27497
rect 2763 27448 2764 27488
rect 2804 27448 2805 27488
rect 2763 27439 2805 27448
rect 3531 27488 3573 27497
rect 3531 27448 3532 27488
rect 3572 27448 3573 27488
rect 3531 27439 3573 27448
rect 14859 27488 14901 27497
rect 14859 27448 14860 27488
rect 14900 27448 14901 27488
rect 14859 27439 14901 27448
rect 17355 27488 17397 27497
rect 17355 27448 17356 27488
rect 17396 27448 17397 27488
rect 17355 27439 17397 27448
rect 3130 27404 3188 27405
rect 3130 27364 3139 27404
rect 3179 27364 3188 27404
rect 3130 27363 3188 27364
rect 6891 27404 6933 27413
rect 6891 27364 6892 27404
rect 6932 27364 6933 27404
rect 6891 27355 6933 27364
rect 9387 27404 9429 27413
rect 9387 27364 9388 27404
rect 9428 27364 9429 27404
rect 9387 27355 9429 27364
rect 11883 27404 11925 27413
rect 11883 27364 11884 27404
rect 11924 27364 11925 27404
rect 11883 27355 11925 27364
rect 17530 27404 17588 27405
rect 17530 27364 17539 27404
rect 17579 27364 17588 27404
rect 17530 27363 17588 27364
rect 21483 27404 21525 27413
rect 21483 27364 21484 27404
rect 21524 27364 21525 27404
rect 21483 27355 21525 27364
rect 24267 27404 24309 27413
rect 24267 27364 24268 27404
rect 24308 27364 24309 27404
rect 24267 27355 24309 27364
rect 24459 27404 24501 27413
rect 24459 27364 24460 27404
rect 24500 27364 24501 27404
rect 24459 27355 24501 27364
rect 29259 27404 29301 27413
rect 29259 27364 29260 27404
rect 29300 27364 29301 27404
rect 29259 27355 29301 27364
rect 29451 27404 29493 27413
rect 29451 27364 29452 27404
rect 29492 27364 29493 27404
rect 29451 27355 29493 27364
rect 576 27236 31392 27260
rect 576 27196 3112 27236
rect 3480 27196 10886 27236
rect 11254 27196 18660 27236
rect 19028 27196 26434 27236
rect 26802 27196 31392 27236
rect 576 27172 31392 27196
rect 2091 27068 2133 27077
rect 2091 27028 2092 27068
rect 2132 27028 2133 27068
rect 2091 27019 2133 27028
rect 2650 27068 2708 27069
rect 2650 27028 2659 27068
rect 2699 27028 2708 27068
rect 2650 27027 2708 27028
rect 6682 27068 6740 27069
rect 6682 27028 6691 27068
rect 6731 27028 6740 27068
rect 6682 27027 6740 27028
rect 7930 27068 7988 27069
rect 7930 27028 7939 27068
rect 7979 27028 7988 27068
rect 7930 27027 7988 27028
rect 9850 27068 9908 27069
rect 9850 27028 9859 27068
rect 9899 27028 9908 27068
rect 9850 27027 9908 27028
rect 12075 27068 12117 27077
rect 12075 27028 12076 27068
rect 12116 27028 12117 27068
rect 12075 27019 12117 27028
rect 14955 27068 14997 27077
rect 14955 27028 14956 27068
rect 14996 27028 14997 27068
rect 14955 27019 14997 27028
rect 19179 27068 19221 27077
rect 19179 27028 19180 27068
rect 19220 27028 19221 27068
rect 19179 27019 19221 27028
rect 22923 27068 22965 27077
rect 22923 27028 22924 27068
rect 22964 27028 22965 27068
rect 22923 27019 22965 27028
rect 26379 27068 26421 27077
rect 26379 27028 26380 27068
rect 26420 27028 26421 27068
rect 26379 27019 26421 27028
rect 28299 27068 28341 27077
rect 28299 27028 28300 27068
rect 28340 27028 28341 27068
rect 28299 27019 28341 27028
rect 1131 26984 1173 26993
rect 1131 26944 1132 26984
rect 1172 26944 1173 26984
rect 1131 26935 1173 26944
rect 6507 26984 6549 26993
rect 6507 26944 6508 26984
rect 6548 26944 6549 26984
rect 6507 26935 6549 26944
rect 11115 26984 11157 26993
rect 11115 26944 11116 26984
rect 11156 26944 11157 26984
rect 11115 26935 11157 26944
rect 12747 26984 12789 26993
rect 12747 26944 12748 26984
rect 12788 26944 12789 26984
rect 12747 26935 12789 26944
rect 13419 26984 13461 26993
rect 13419 26944 13420 26984
rect 13460 26944 13461 26984
rect 13419 26935 13461 26944
rect 15627 26984 15669 26993
rect 15627 26944 15628 26984
rect 15668 26944 15669 26984
rect 15627 26935 15669 26944
rect 3226 26900 3284 26901
rect 3226 26860 3235 26900
rect 3275 26860 3284 26900
rect 3226 26859 3284 26860
rect 7755 26900 7797 26909
rect 7755 26860 7756 26900
rect 7796 26860 7797 26900
rect 6975 26849 7017 26858
rect 7755 26851 7797 26860
rect 13515 26900 13557 26909
rect 13515 26860 13516 26900
rect 13556 26860 13557 26900
rect 13515 26851 13557 26860
rect 20602 26900 20660 26901
rect 20602 26860 20611 26900
rect 20651 26860 20660 26900
rect 20602 26859 20660 26860
rect 2091 26816 2133 26825
rect 2091 26776 2092 26816
rect 2132 26776 2133 26816
rect 2091 26767 2133 26776
rect 2283 26816 2325 26825
rect 2283 26776 2284 26816
rect 2324 26776 2325 26816
rect 2283 26767 2325 26776
rect 2475 26816 2517 26825
rect 2475 26776 2476 26816
rect 2516 26776 2517 26816
rect 2475 26767 2517 26776
rect 2650 26816 2708 26817
rect 2650 26776 2659 26816
rect 2699 26776 2708 26816
rect 2650 26775 2708 26776
rect 4762 26816 4820 26817
rect 4762 26776 4771 26816
rect 4811 26776 4820 26816
rect 4762 26775 4820 26776
rect 5146 26816 5204 26817
rect 5146 26776 5155 26816
rect 5195 26776 5204 26816
rect 5146 26775 5204 26776
rect 5547 26816 5589 26825
rect 5547 26776 5548 26816
rect 5588 26776 5589 26816
rect 5547 26767 5589 26776
rect 5635 26816 5693 26817
rect 5635 26776 5644 26816
rect 5684 26776 5693 26816
rect 5635 26775 5693 26776
rect 5883 26816 5925 26825
rect 5883 26776 5884 26816
rect 5924 26776 5925 26816
rect 6975 26809 6976 26849
rect 7016 26809 7017 26849
rect 6975 26800 7017 26809
rect 7066 26816 7124 26817
rect 5883 26767 5925 26776
rect 7066 26776 7075 26816
rect 7115 26776 7124 26816
rect 7066 26775 7124 26776
rect 8139 26816 8181 26825
rect 8139 26776 8140 26816
rect 8180 26776 8181 26816
rect 8139 26767 8181 26776
rect 8227 26816 8285 26817
rect 8227 26776 8236 26816
rect 8276 26776 8285 26816
rect 8227 26775 8285 26776
rect 8619 26816 8661 26825
rect 8619 26776 8620 26816
rect 8660 26776 8661 26816
rect 8619 26767 8661 26776
rect 8707 26816 8765 26817
rect 8707 26776 8716 26816
rect 8756 26776 8765 26816
rect 8707 26775 8765 26776
rect 8907 26816 8949 26825
rect 8907 26776 8908 26816
rect 8948 26776 8949 26816
rect 8907 26767 8949 26776
rect 10147 26816 10205 26817
rect 10147 26776 10156 26816
rect 10196 26776 10205 26816
rect 10147 26775 10205 26776
rect 10443 26816 10485 26825
rect 10443 26776 10444 26816
rect 10484 26776 10485 26816
rect 10443 26767 10485 26776
rect 10923 26816 10965 26825
rect 10923 26776 10924 26816
rect 10964 26776 10965 26816
rect 10923 26767 10965 26776
rect 11403 26816 11445 26825
rect 11403 26776 11404 26816
rect 11444 26776 11445 26816
rect 11403 26767 11445 26776
rect 11787 26816 11829 26825
rect 11787 26776 11788 26816
rect 11828 26776 11829 26816
rect 11787 26767 11829 26776
rect 11901 26816 11959 26817
rect 11901 26776 11910 26816
rect 11950 26776 11959 26816
rect 11901 26775 11959 26776
rect 12028 26816 12086 26817
rect 12028 26776 12037 26816
rect 12077 26776 12086 26816
rect 12028 26775 12086 26776
rect 12250 26816 12308 26817
rect 12250 26776 12259 26816
rect 12299 26776 12308 26816
rect 12250 26775 12308 26776
rect 12939 26816 12981 26825
rect 12939 26776 12940 26816
rect 12980 26776 12981 26816
rect 12939 26767 12981 26776
rect 13188 26816 13246 26817
rect 13188 26776 13197 26816
rect 13237 26776 13246 26816
rect 13188 26775 13246 26776
rect 13344 26816 13386 26825
rect 13344 26776 13345 26816
rect 13385 26776 13386 26816
rect 13344 26767 13386 26776
rect 13642 26816 13700 26817
rect 13642 26776 13651 26816
rect 13691 26776 13700 26816
rect 13642 26775 13700 26776
rect 13803 26816 13845 26825
rect 13803 26776 13804 26816
rect 13844 26776 13845 26816
rect 13803 26767 13845 26776
rect 14746 26816 14804 26817
rect 14746 26776 14755 26816
rect 14795 26776 14804 26816
rect 14746 26775 14804 26776
rect 15819 26816 15861 26825
rect 15819 26776 15820 26816
rect 15860 26776 15861 26816
rect 15819 26767 15861 26776
rect 17050 26816 17108 26817
rect 17050 26776 17059 26816
rect 17099 26776 17108 26816
rect 17050 26775 17108 26776
rect 19467 26816 19509 26825
rect 19851 26816 19893 26825
rect 19467 26776 19468 26816
rect 19508 26776 19509 26816
rect 19467 26767 19509 26776
rect 19563 26807 19605 26816
rect 19563 26767 19564 26807
rect 19604 26767 19605 26807
rect 19851 26776 19852 26816
rect 19892 26776 19893 26816
rect 19851 26767 19893 26776
rect 20331 26816 20373 26825
rect 20331 26776 20332 26816
rect 20372 26776 20373 26816
rect 20331 26767 20373 26776
rect 21291 26816 21333 26825
rect 21291 26776 21292 26816
rect 21332 26776 21333 26816
rect 21291 26767 21333 26776
rect 21526 26816 21568 26825
rect 21526 26776 21527 26816
rect 21567 26776 21568 26816
rect 21526 26767 21568 26776
rect 21658 26816 21716 26817
rect 21658 26776 21667 26816
rect 21707 26776 21716 26816
rect 21658 26775 21716 26776
rect 21771 26816 21813 26825
rect 21771 26776 21772 26816
rect 21812 26776 21813 26816
rect 21771 26767 21813 26776
rect 22731 26816 22773 26825
rect 22731 26776 22732 26816
rect 22772 26776 22773 26816
rect 22731 26767 22773 26776
rect 23595 26816 23637 26825
rect 23595 26776 23596 26816
rect 23636 26776 23637 26816
rect 23595 26767 23637 26776
rect 24459 26816 24501 26825
rect 24459 26776 24460 26816
rect 24500 26776 24501 26816
rect 24459 26767 24501 26776
rect 25323 26816 25365 26825
rect 25323 26776 25324 26816
rect 25364 26776 25365 26816
rect 25323 26767 25365 26776
rect 26187 26816 26229 26825
rect 26187 26776 26188 26816
rect 26228 26776 26229 26816
rect 26187 26767 26229 26776
rect 27051 26816 27093 26825
rect 27051 26776 27052 26816
rect 27092 26776 27093 26816
rect 27051 26767 27093 26776
rect 27915 26816 27957 26825
rect 27915 26776 27916 26816
rect 27956 26776 27957 26816
rect 27915 26767 27957 26776
rect 30202 26816 30260 26817
rect 30202 26776 30211 26816
rect 30251 26776 30260 26816
rect 30202 26775 30260 26776
rect 30891 26816 30933 26825
rect 30891 26776 30892 26816
rect 30932 26776 30933 26816
rect 30891 26767 30933 26776
rect 19563 26758 19605 26767
rect 5341 26732 5383 26741
rect 5341 26692 5342 26732
rect 5382 26692 5383 26732
rect 5341 26683 5383 26692
rect 7933 26732 7975 26741
rect 7933 26692 7934 26732
rect 7974 26692 7975 26732
rect 7933 26683 7975 26692
rect 8413 26732 8455 26741
rect 8413 26692 8414 26732
rect 8454 26692 8455 26732
rect 8413 26683 8455 26692
rect 9853 26732 9895 26741
rect 9853 26692 9854 26732
rect 9894 26692 9895 26732
rect 9853 26683 9895 26692
rect 12569 26732 12611 26741
rect 12569 26692 12570 26732
rect 12610 26692 12611 26732
rect 12569 26683 12611 26692
rect 15034 26732 15092 26733
rect 15034 26692 15043 26732
rect 15083 26692 15092 26732
rect 15034 26691 15092 26692
rect 16491 26732 16533 26741
rect 16491 26692 16492 26732
rect 16532 26692 16533 26732
rect 16491 26683 16533 26692
rect 16666 26732 16724 26733
rect 16666 26692 16675 26732
rect 16715 26692 16724 26732
rect 16666 26691 16724 26692
rect 21850 26732 21908 26733
rect 21850 26692 21859 26732
rect 21899 26692 21908 26732
rect 21850 26691 21908 26692
rect 25498 26732 25556 26733
rect 25498 26692 25507 26732
rect 25547 26692 25556 26732
rect 25498 26691 25556 26692
rect 30586 26732 30644 26733
rect 30586 26692 30595 26732
rect 30635 26692 30644 26732
rect 30586 26691 30644 26692
rect 1515 26648 1557 26657
rect 1515 26608 1516 26648
rect 1556 26608 1557 26648
rect 1515 26599 1557 26608
rect 1899 26648 1941 26657
rect 1899 26608 1900 26648
rect 1940 26608 1941 26648
rect 1899 26599 1941 26608
rect 2859 26648 2901 26657
rect 2859 26608 2860 26648
rect 2900 26608 2901 26648
rect 2859 26599 2901 26608
rect 5434 26648 5492 26649
rect 5434 26608 5443 26648
rect 5483 26608 5492 26648
rect 5434 26607 5492 26608
rect 7515 26648 7557 26657
rect 7515 26608 7516 26648
rect 7556 26608 7557 26648
rect 7210 26606 7268 26607
rect 7210 26566 7219 26606
rect 7259 26566 7268 26606
rect 7515 26599 7557 26608
rect 8139 26648 8181 26657
rect 8139 26608 8140 26648
rect 8180 26608 8181 26648
rect 8139 26599 8181 26608
rect 8506 26648 8564 26649
rect 8506 26608 8515 26648
rect 8555 26608 8564 26648
rect 8506 26607 8564 26608
rect 9579 26648 9621 26657
rect 9579 26608 9580 26648
rect 9620 26608 9621 26648
rect 9579 26599 9621 26608
rect 10059 26648 10101 26657
rect 10059 26608 10060 26648
rect 10100 26608 10101 26648
rect 10059 26599 10101 26608
rect 10330 26648 10388 26649
rect 10330 26608 10339 26648
rect 10379 26608 10388 26648
rect 10330 26607 10388 26608
rect 10635 26648 10677 26657
rect 10635 26608 10636 26648
rect 10676 26608 10677 26648
rect 10635 26599 10677 26608
rect 10810 26648 10868 26649
rect 10810 26608 10819 26648
rect 10859 26608 10868 26648
rect 10810 26607 10868 26608
rect 11290 26648 11348 26649
rect 11290 26608 11299 26648
rect 11339 26608 11348 26648
rect 11290 26607 11348 26608
rect 11595 26648 11637 26657
rect 11595 26608 11596 26648
rect 11636 26608 11637 26648
rect 11595 26599 11637 26608
rect 12346 26648 12404 26649
rect 12346 26608 12355 26648
rect 12395 26608 12404 26648
rect 12346 26607 12404 26608
rect 12459 26648 12501 26657
rect 12459 26608 12460 26648
rect 12500 26608 12501 26648
rect 12459 26599 12501 26608
rect 12987 26648 13029 26657
rect 12987 26608 12988 26648
rect 13028 26608 13029 26648
rect 12987 26599 13029 26608
rect 14475 26648 14517 26657
rect 14475 26608 14476 26648
rect 14516 26608 14517 26648
rect 14475 26599 14517 26608
rect 18987 26648 19029 26657
rect 18987 26608 18988 26648
rect 19028 26608 19029 26648
rect 18987 26599 19029 26608
rect 20139 26648 20181 26657
rect 20139 26608 20140 26648
rect 20180 26608 20181 26648
rect 20139 26599 20181 26608
rect 20410 26648 20468 26649
rect 20410 26608 20419 26648
rect 20459 26608 20468 26648
rect 20410 26607 20468 26608
rect 22059 26648 22101 26657
rect 22059 26608 22060 26648
rect 22100 26608 22101 26648
rect 22059 26599 22101 26608
rect 23787 26648 23829 26657
rect 23787 26608 23788 26648
rect 23828 26608 23829 26648
rect 23787 26599 23829 26608
rect 24651 26648 24693 26657
rect 24651 26608 24652 26648
rect 24692 26608 24693 26648
rect 24651 26599 24693 26608
rect 27243 26648 27285 26657
rect 27243 26608 27244 26648
rect 27284 26608 27285 26648
rect 27243 26599 27285 26608
rect 28299 26648 28341 26657
rect 28299 26608 28300 26648
rect 28340 26608 28341 26648
rect 28299 26599 28341 26608
rect 30778 26648 30836 26649
rect 30778 26608 30787 26648
rect 30827 26608 30836 26648
rect 30778 26607 30836 26608
rect 31083 26648 31125 26657
rect 31083 26608 31084 26648
rect 31124 26608 31125 26648
rect 31083 26599 31125 26608
rect 7210 26565 7268 26566
rect 576 26480 31392 26504
rect 576 26440 4352 26480
rect 4720 26440 12126 26480
rect 12494 26440 19900 26480
rect 20268 26440 27674 26480
rect 28042 26440 31392 26480
rect 576 26416 31392 26440
rect 18010 26354 18068 26355
rect 2667 26312 2709 26321
rect 2667 26272 2668 26312
rect 2708 26272 2709 26312
rect 2667 26263 2709 26272
rect 5019 26312 5061 26321
rect 5019 26272 5020 26312
rect 5060 26272 5061 26312
rect 5019 26263 5061 26272
rect 8811 26312 8853 26321
rect 8811 26272 8812 26312
rect 8852 26272 8853 26312
rect 8811 26263 8853 26272
rect 11307 26312 11349 26321
rect 11307 26272 11308 26312
rect 11348 26272 11349 26312
rect 11307 26263 11349 26272
rect 12171 26312 12213 26321
rect 12171 26272 12172 26312
rect 12212 26272 12213 26312
rect 12171 26263 12213 26272
rect 12730 26312 12788 26313
rect 12730 26272 12739 26312
rect 12779 26272 12788 26312
rect 12730 26271 12788 26272
rect 13498 26312 13556 26313
rect 13498 26272 13507 26312
rect 13547 26272 13556 26312
rect 13498 26271 13556 26272
rect 13611 26312 13653 26321
rect 13611 26272 13612 26312
rect 13652 26272 13653 26312
rect 13611 26263 13653 26272
rect 16347 26312 16389 26321
rect 18010 26314 18019 26354
rect 18059 26314 18068 26354
rect 18010 26313 18068 26314
rect 16347 26272 16348 26312
rect 16388 26272 16389 26312
rect 18891 26312 18933 26321
rect 16347 26263 16389 26272
rect 18135 26270 18177 26279
rect 3003 26228 3045 26237
rect 3003 26188 3004 26228
rect 3044 26188 3045 26228
rect 3003 26179 3045 26188
rect 4011 26228 4053 26237
rect 4011 26188 4012 26228
rect 4052 26188 4053 26228
rect 4011 26179 4053 26188
rect 4683 26228 4725 26237
rect 18135 26230 18136 26270
rect 18176 26230 18177 26270
rect 18891 26272 18892 26312
rect 18932 26272 18933 26312
rect 18891 26263 18933 26272
rect 20506 26312 20564 26313
rect 20506 26272 20515 26312
rect 20555 26272 20564 26312
rect 20506 26271 20564 26272
rect 25179 26312 25221 26321
rect 25179 26272 25180 26312
rect 25220 26272 25221 26312
rect 25179 26263 25221 26272
rect 25498 26312 25556 26313
rect 25498 26272 25507 26312
rect 25547 26272 25556 26312
rect 25498 26271 25556 26272
rect 27051 26312 27093 26321
rect 27051 26272 27052 26312
rect 27092 26272 27093 26312
rect 27051 26263 27093 26272
rect 27819 26312 27861 26321
rect 27819 26272 27820 26312
rect 27860 26272 27861 26312
rect 27819 26263 27861 26272
rect 31275 26312 31317 26321
rect 31275 26272 31276 26312
rect 31316 26272 31317 26312
rect 31275 26263 31317 26272
rect 4683 26188 4684 26228
rect 4724 26188 4725 26228
rect 4683 26179 4725 26188
rect 6490 26228 6548 26229
rect 6490 26188 6499 26228
rect 6539 26188 6548 26228
rect 6490 26187 6548 26188
rect 8986 26228 9044 26229
rect 8986 26188 8995 26228
rect 9035 26188 9044 26228
rect 8986 26187 9044 26188
rect 13882 26228 13940 26229
rect 13882 26188 13891 26228
rect 13931 26188 13940 26228
rect 18135 26221 18177 26230
rect 22042 26228 22100 26229
rect 13882 26187 13940 26188
rect 18055 26186 18097 26195
rect 22042 26188 22051 26228
rect 22091 26188 22100 26228
rect 22042 26187 22100 26188
rect 26427 26228 26469 26237
rect 26427 26188 26428 26228
rect 26468 26188 26469 26228
rect 2091 26144 2133 26153
rect 2091 26104 2092 26144
rect 2132 26104 2133 26144
rect 2091 26095 2133 26104
rect 2266 26144 2324 26145
rect 3339 26144 3381 26153
rect 2266 26104 2275 26144
rect 2315 26104 2324 26144
rect 2266 26103 2324 26104
rect 2850 26135 2896 26144
rect 2850 26095 2851 26135
rect 2891 26095 2896 26135
rect 3339 26104 3340 26144
rect 3380 26104 3381 26144
rect 3339 26095 3381 26104
rect 4299 26144 4341 26153
rect 4299 26104 4300 26144
rect 4340 26104 4341 26144
rect 4299 26095 4341 26104
rect 4570 26144 4628 26145
rect 4570 26104 4579 26144
rect 4619 26104 4628 26144
rect 4570 26103 4628 26104
rect 5163 26144 5205 26153
rect 5163 26104 5164 26144
rect 5204 26104 5205 26144
rect 5163 26095 5205 26104
rect 6874 26144 6932 26145
rect 6874 26104 6883 26144
rect 6923 26104 6932 26144
rect 6874 26103 6932 26104
rect 9370 26144 9428 26145
rect 9370 26104 9379 26144
rect 9419 26104 9428 26144
rect 9370 26103 9428 26104
rect 11499 26144 11541 26153
rect 11499 26104 11500 26144
rect 11540 26104 11541 26144
rect 6346 26102 6404 26103
rect 2850 26086 2896 26095
rect 843 26060 885 26069
rect 6346 26062 6355 26102
rect 6395 26062 6404 26102
rect 11499 26095 11541 26104
rect 12459 26144 12501 26153
rect 12459 26104 12460 26144
rect 12500 26104 12501 26144
rect 12459 26095 12501 26104
rect 12667 26144 12725 26145
rect 12667 26104 12676 26144
rect 12716 26104 12725 26144
rect 12667 26103 12725 26104
rect 12848 26144 12890 26153
rect 12848 26104 12849 26144
rect 12889 26104 12890 26144
rect 12848 26095 12890 26104
rect 12952 26144 13010 26145
rect 12952 26104 12961 26144
rect 13001 26104 13010 26144
rect 13210 26144 13268 26145
rect 12952 26103 13010 26104
rect 13083 26133 13125 26142
rect 13083 26093 13084 26133
rect 13124 26093 13125 26133
rect 13210 26104 13219 26144
rect 13259 26104 13268 26144
rect 13210 26103 13268 26104
rect 13400 26144 13458 26145
rect 13400 26104 13409 26144
rect 13449 26104 13458 26144
rect 13400 26103 13458 26104
rect 13721 26144 13763 26153
rect 13721 26104 13722 26144
rect 13762 26104 13763 26144
rect 13721 26095 13763 26104
rect 14266 26144 14324 26145
rect 14266 26104 14275 26144
rect 14315 26104 14324 26144
rect 14266 26103 14324 26104
rect 16491 26144 16533 26153
rect 16491 26104 16492 26144
rect 16532 26104 16533 26144
rect 16491 26095 16533 26104
rect 16666 26144 16724 26145
rect 16666 26104 16675 26144
rect 16715 26104 16724 26144
rect 16666 26103 16724 26104
rect 17355 26144 17397 26153
rect 17355 26104 17356 26144
rect 17396 26104 17397 26144
rect 18055 26146 18056 26186
rect 18096 26146 18097 26186
rect 26427 26179 26469 26188
rect 18055 26137 18097 26146
rect 18346 26144 18404 26145
rect 17355 26095 17397 26104
rect 18346 26104 18355 26144
rect 18395 26104 18404 26144
rect 18346 26103 18404 26104
rect 18502 26144 18544 26153
rect 18502 26104 18503 26144
rect 18543 26104 18544 26144
rect 18502 26095 18544 26104
rect 18699 26144 18741 26153
rect 18699 26104 18700 26144
rect 18740 26104 18741 26144
rect 18699 26095 18741 26104
rect 19563 26144 19605 26153
rect 19563 26104 19564 26144
rect 19604 26104 19605 26144
rect 19563 26095 19605 26104
rect 19755 26144 19797 26153
rect 19755 26104 19756 26144
rect 19796 26104 19797 26144
rect 19755 26095 19797 26104
rect 20043 26144 20085 26153
rect 20043 26104 20044 26144
rect 20084 26104 20085 26144
rect 20043 26095 20085 26104
rect 20667 26144 20709 26153
rect 20667 26104 20668 26144
rect 20708 26104 20709 26144
rect 20667 26095 20709 26104
rect 20811 26144 20853 26153
rect 20811 26104 20812 26144
rect 20852 26104 20853 26144
rect 20811 26095 20853 26104
rect 21370 26144 21428 26145
rect 21370 26104 21379 26144
rect 21419 26104 21428 26144
rect 21370 26103 21428 26104
rect 22426 26144 22484 26145
rect 22426 26104 22435 26144
rect 22475 26104 22484 26144
rect 22426 26103 22484 26104
rect 24555 26144 24597 26153
rect 24555 26104 24556 26144
rect 24596 26104 24597 26144
rect 24555 26095 24597 26104
rect 24730 26144 24788 26145
rect 24730 26104 24739 26144
rect 24779 26104 24788 26144
rect 24730 26103 24788 26104
rect 24843 26144 24885 26153
rect 25803 26144 25845 26153
rect 26763 26144 26805 26153
rect 24843 26104 24844 26144
rect 24884 26104 24885 26144
rect 24843 26095 24885 26104
rect 25026 26135 25072 26144
rect 25026 26095 25027 26135
rect 25067 26095 25072 26135
rect 25803 26104 25804 26144
rect 25844 26104 25845 26144
rect 25803 26095 25845 26104
rect 26274 26135 26320 26144
rect 26274 26095 26275 26135
rect 26315 26095 26320 26135
rect 26763 26104 26764 26144
rect 26804 26104 26805 26144
rect 27339 26144 27381 26153
rect 26763 26095 26805 26104
rect 26891 26120 26933 26129
rect 13083 26084 13125 26093
rect 25026 26086 25072 26095
rect 26274 26086 26320 26095
rect 26891 26080 26892 26120
rect 26932 26080 26933 26120
rect 27339 26104 27340 26144
rect 27380 26104 27381 26144
rect 27339 26095 27381 26104
rect 27723 26144 27765 26153
rect 27723 26104 27724 26144
rect 27764 26104 27765 26144
rect 27723 26095 27765 26104
rect 28779 26144 28821 26153
rect 28779 26104 28780 26144
rect 28820 26104 28821 26144
rect 28779 26095 28821 26104
rect 29338 26144 29396 26145
rect 29338 26104 29347 26144
rect 29387 26104 29396 26144
rect 29338 26103 29396 26104
rect 26891 26071 26933 26080
rect 6346 26061 6404 26062
rect 843 26020 844 26060
rect 884 26020 885 26060
rect 843 26011 885 26020
rect 6154 26060 6212 26061
rect 6154 26020 6163 26060
rect 6203 26020 6212 26060
rect 6154 26019 6212 26020
rect 18219 26060 18261 26069
rect 18219 26020 18220 26060
rect 18260 26020 18261 26060
rect 18219 26011 18261 26020
rect 25713 26060 25755 26069
rect 25713 26020 25714 26060
rect 25754 26020 25755 26060
rect 25713 26011 25755 26020
rect 28971 26060 29013 26069
rect 28971 26020 28972 26060
rect 29012 26020 29013 26060
rect 28971 26011 29013 26020
rect 603 25976 645 25985
rect 603 25936 604 25976
rect 644 25936 645 25976
rect 603 25927 645 25936
rect 1515 25976 1557 25985
rect 1515 25936 1516 25976
rect 1556 25936 1557 25976
rect 1515 25927 1557 25936
rect 1899 25976 1941 25985
rect 1899 25936 1900 25976
rect 1940 25936 1941 25976
rect 1899 25927 1941 25936
rect 2266 25976 2324 25977
rect 2266 25936 2275 25976
rect 2315 25936 2324 25976
rect 2266 25935 2324 25936
rect 16203 25976 16245 25985
rect 16203 25936 16204 25976
rect 16244 25936 16245 25976
rect 16203 25927 16245 25936
rect 17547 25976 17589 25985
rect 17547 25936 17548 25976
rect 17588 25936 17589 25976
rect 17547 25927 17589 25936
rect 18603 25976 18645 25985
rect 18603 25936 18604 25976
rect 18644 25936 18645 25976
rect 18603 25927 18645 25936
rect 20379 25976 20421 25985
rect 20379 25936 20380 25976
rect 20420 25936 20421 25976
rect 20379 25927 20421 25936
rect 24363 25976 24405 25985
rect 24363 25936 24364 25976
rect 24404 25936 24405 25976
rect 24363 25927 24405 25936
rect 24843 25976 24885 25985
rect 24843 25936 24844 25976
rect 24884 25936 24885 25976
rect 24843 25927 24885 25936
rect 28107 25976 28149 25985
rect 28107 25936 28108 25976
rect 28148 25936 28149 25976
rect 28107 25927 28149 25936
rect 5835 25892 5877 25901
rect 5835 25852 5836 25892
rect 5876 25852 5877 25892
rect 5835 25843 5877 25852
rect 21771 25892 21813 25901
rect 21771 25852 21772 25892
rect 21812 25852 21813 25892
rect 21771 25843 21813 25852
rect 576 25724 31392 25748
rect 576 25684 3112 25724
rect 3480 25684 10886 25724
rect 11254 25684 18660 25724
rect 19028 25684 26434 25724
rect 26802 25684 31392 25724
rect 576 25660 31392 25684
rect 5547 25556 5589 25565
rect 5547 25516 5548 25556
rect 5588 25516 5589 25556
rect 5547 25507 5589 25516
rect 7834 25556 7892 25557
rect 7834 25516 7843 25556
rect 7883 25516 7892 25556
rect 7834 25515 7892 25516
rect 8859 25556 8901 25565
rect 8859 25516 8860 25556
rect 8900 25516 8901 25556
rect 8859 25507 8901 25516
rect 21082 25556 21140 25557
rect 21082 25516 21091 25556
rect 21131 25516 21140 25556
rect 21082 25515 21140 25516
rect 26859 25556 26901 25565
rect 26859 25516 26860 25556
rect 26900 25516 26901 25556
rect 26859 25507 26901 25516
rect 28107 25556 28149 25565
rect 28107 25516 28108 25556
rect 28148 25516 28149 25556
rect 28107 25507 28149 25516
rect 1611 25472 1653 25481
rect 1611 25432 1612 25472
rect 1652 25432 1653 25472
rect 1611 25423 1653 25432
rect 2379 25472 2421 25481
rect 9195 25472 9237 25481
rect 2379 25432 2380 25472
rect 2420 25432 2421 25472
rect 2379 25423 2421 25432
rect 7611 25463 7653 25472
rect 7611 25423 7612 25463
rect 7652 25423 7653 25463
rect 9195 25432 9196 25472
rect 9236 25432 9237 25472
rect 9195 25423 9237 25432
rect 10779 25472 10821 25481
rect 10779 25432 10780 25472
rect 10820 25432 10821 25472
rect 10779 25423 10821 25432
rect 11595 25472 11637 25481
rect 11595 25432 11596 25472
rect 11636 25432 11637 25472
rect 11595 25423 11637 25432
rect 14187 25472 14229 25481
rect 14187 25432 14188 25472
rect 14228 25432 14229 25472
rect 14187 25423 14229 25432
rect 14763 25472 14805 25481
rect 14763 25432 14764 25472
rect 14804 25432 14805 25472
rect 14763 25423 14805 25432
rect 18699 25472 18741 25481
rect 18699 25432 18700 25472
rect 18740 25432 18741 25472
rect 18699 25423 18741 25432
rect 25227 25472 25269 25481
rect 26379 25472 26421 25481
rect 25227 25432 25228 25472
rect 25268 25432 25269 25472
rect 25227 25423 25269 25432
rect 25675 25463 25717 25472
rect 25675 25423 25676 25463
rect 25716 25423 25717 25463
rect 26379 25432 26380 25472
rect 26420 25432 26421 25472
rect 26379 25423 26421 25432
rect 30987 25472 31029 25481
rect 30987 25432 30988 25472
rect 31028 25432 31029 25472
rect 30987 25423 31029 25432
rect 7611 25414 7653 25423
rect 25675 25414 25717 25423
rect 651 25388 693 25397
rect 651 25348 652 25388
rect 692 25348 693 25388
rect 651 25339 693 25348
rect 1227 25388 1269 25397
rect 1227 25348 1228 25388
rect 1268 25348 1269 25388
rect 1227 25339 1269 25348
rect 2650 25388 2708 25389
rect 2650 25348 2659 25388
rect 2699 25348 2708 25388
rect 2650 25347 2708 25348
rect 3051 25388 3093 25397
rect 3051 25348 3052 25388
rect 3092 25348 3093 25388
rect 3051 25339 3093 25348
rect 8619 25388 8661 25397
rect 8619 25348 8620 25388
rect 8660 25348 8661 25388
rect 8619 25339 8661 25348
rect 9579 25388 9621 25397
rect 9579 25348 9580 25388
rect 9620 25348 9621 25388
rect 9579 25339 9621 25348
rect 13851 25388 13893 25397
rect 13851 25348 13852 25388
rect 13892 25348 13893 25388
rect 13851 25339 13893 25348
rect 14667 25388 14709 25397
rect 14667 25348 14668 25388
rect 14708 25348 14709 25388
rect 14667 25339 14709 25348
rect 16395 25388 16437 25397
rect 16395 25348 16396 25388
rect 16436 25348 16437 25388
rect 16395 25339 16437 25348
rect 25323 25388 25365 25397
rect 25323 25348 25324 25388
rect 25364 25348 25365 25388
rect 25323 25339 25365 25348
rect 27339 25388 27381 25397
rect 27339 25348 27340 25388
rect 27380 25348 27381 25388
rect 27339 25339 27381 25348
rect 12304 25315 12346 25324
rect 1803 25304 1845 25313
rect 1803 25264 1804 25304
rect 1844 25264 1845 25304
rect 1803 25255 1845 25264
rect 1995 25304 2037 25313
rect 1995 25264 1996 25304
rect 2036 25264 2037 25304
rect 1995 25255 2037 25264
rect 2518 25304 2560 25313
rect 2518 25264 2519 25304
rect 2559 25264 2560 25304
rect 2518 25255 2560 25264
rect 2748 25304 2806 25305
rect 2748 25264 2757 25304
rect 2797 25264 2806 25304
rect 2748 25263 2806 25264
rect 3418 25304 3476 25305
rect 6219 25304 6261 25313
rect 3418 25264 3427 25304
rect 3467 25264 3476 25304
rect 3418 25263 3476 25264
rect 5931 25295 5973 25304
rect 5931 25255 5932 25295
rect 5972 25255 5973 25295
rect 6219 25264 6220 25304
rect 6260 25264 6261 25304
rect 6219 25255 6261 25264
rect 6507 25304 6549 25313
rect 6507 25264 6508 25304
rect 6548 25264 6549 25304
rect 6507 25255 6549 25264
rect 6891 25304 6933 25313
rect 6891 25264 6892 25304
rect 6932 25264 6933 25304
rect 6891 25255 6933 25264
rect 7275 25304 7317 25313
rect 7275 25264 7276 25304
rect 7316 25264 7317 25304
rect 7275 25255 7317 25264
rect 7642 25304 7700 25305
rect 7642 25264 7651 25304
rect 7691 25264 7700 25304
rect 7642 25263 7700 25264
rect 8335 25304 8393 25305
rect 8335 25264 8344 25304
rect 8384 25264 8393 25304
rect 8335 25263 8393 25264
rect 9946 25304 10004 25305
rect 9946 25264 9955 25304
rect 9995 25264 10004 25304
rect 9946 25263 10004 25264
rect 10347 25304 10389 25313
rect 10347 25264 10348 25304
rect 10388 25264 10389 25304
rect 10347 25255 10389 25264
rect 10635 25304 10677 25313
rect 10635 25264 10636 25304
rect 10676 25264 10677 25304
rect 10635 25255 10677 25264
rect 10858 25304 10916 25305
rect 10858 25264 10867 25304
rect 10907 25264 10916 25304
rect 10858 25263 10916 25264
rect 11403 25304 11445 25313
rect 11403 25264 11404 25304
rect 11444 25264 11445 25304
rect 11403 25255 11445 25264
rect 11518 25304 11560 25313
rect 11518 25264 11519 25304
rect 11559 25264 11560 25304
rect 11518 25255 11560 25264
rect 11691 25304 11733 25313
rect 11691 25264 11692 25304
rect 11732 25264 11733 25304
rect 11691 25255 11733 25264
rect 11911 25304 11969 25305
rect 11911 25264 11920 25304
rect 11960 25264 11969 25304
rect 11911 25263 11969 25264
rect 12058 25304 12116 25305
rect 12058 25264 12067 25304
rect 12107 25264 12116 25304
rect 12058 25263 12116 25264
rect 12183 25304 12225 25313
rect 12183 25264 12184 25304
rect 12224 25264 12225 25304
rect 12304 25275 12305 25315
rect 12345 25275 12346 25315
rect 12304 25266 12346 25275
rect 12442 25304 12500 25305
rect 12183 25255 12225 25264
rect 12442 25264 12451 25304
rect 12491 25264 12500 25304
rect 12442 25263 12500 25264
rect 12744 25304 12786 25313
rect 12744 25264 12745 25304
rect 12785 25264 12786 25304
rect 12744 25255 12786 25264
rect 12861 25304 12919 25305
rect 12861 25264 12870 25304
rect 12910 25264 12919 25304
rect 12861 25263 12919 25264
rect 12987 25304 13029 25313
rect 12987 25264 12988 25304
rect 13028 25264 13029 25304
rect 12987 25255 13029 25264
rect 13207 25304 13265 25305
rect 13207 25264 13216 25304
rect 13256 25264 13265 25304
rect 13207 25263 13265 25264
rect 13657 25304 13715 25305
rect 13657 25264 13666 25304
rect 13706 25264 13715 25304
rect 13657 25263 13715 25264
rect 14523 25304 14565 25313
rect 14523 25264 14524 25304
rect 14564 25264 14565 25304
rect 14523 25255 14565 25264
rect 14838 25304 14880 25313
rect 14838 25264 14839 25304
rect 14879 25264 14880 25304
rect 14838 25255 14880 25264
rect 14986 25304 15044 25305
rect 14986 25264 14995 25304
rect 15035 25264 15044 25304
rect 14986 25263 15044 25264
rect 15819 25304 15861 25313
rect 15819 25264 15820 25304
rect 15860 25264 15861 25304
rect 15819 25255 15861 25264
rect 15994 25304 16036 25313
rect 15994 25264 15995 25304
rect 16035 25264 16036 25304
rect 15994 25255 16036 25264
rect 16203 25304 16245 25313
rect 16203 25264 16204 25304
rect 16244 25264 16245 25304
rect 16203 25255 16245 25264
rect 16762 25304 16820 25305
rect 16762 25264 16771 25304
rect 16811 25264 16820 25304
rect 16762 25263 16820 25264
rect 18987 25304 19029 25313
rect 18987 25264 18988 25304
rect 19028 25264 19029 25304
rect 18987 25255 19029 25264
rect 19851 25304 19893 25313
rect 19851 25264 19852 25304
rect 19892 25264 19893 25304
rect 19851 25255 19893 25264
rect 20139 25304 20181 25313
rect 20139 25264 20140 25304
rect 20180 25264 20181 25304
rect 20139 25255 20181 25264
rect 20554 25304 20612 25305
rect 20554 25264 20563 25304
rect 20603 25264 20612 25304
rect 20554 25263 20612 25264
rect 21379 25304 21437 25305
rect 21379 25264 21388 25304
rect 21428 25264 21437 25304
rect 21379 25263 21437 25264
rect 21946 25304 22004 25305
rect 21946 25264 21955 25304
rect 21995 25264 22004 25304
rect 21946 25263 22004 25264
rect 24747 25304 24789 25313
rect 24747 25264 24748 25304
rect 24788 25264 24789 25304
rect 24747 25255 24789 25264
rect 24987 25304 25029 25313
rect 24987 25264 24988 25304
rect 25028 25264 25029 25304
rect 25444 25304 25486 25313
rect 24987 25255 25029 25264
rect 25159 25262 25201 25271
rect 5931 25246 5973 25255
rect 891 25220 933 25229
rect 891 25180 892 25220
rect 932 25180 933 25220
rect 891 25171 933 25180
rect 5835 25220 5877 25229
rect 5835 25180 5836 25220
rect 5876 25180 5877 25220
rect 5835 25171 5877 25180
rect 8170 25220 8228 25221
rect 8170 25180 8179 25220
rect 8219 25180 8228 25220
rect 8170 25179 8228 25180
rect 9339 25220 9381 25229
rect 9339 25180 9340 25220
rect 9380 25180 9381 25220
rect 9339 25171 9381 25180
rect 12442 25220 12500 25221
rect 12442 25180 12451 25220
rect 12491 25180 12500 25220
rect 12442 25179 12500 25180
rect 21085 25220 21127 25229
rect 25159 25222 25160 25262
rect 25200 25222 25201 25262
rect 25444 25264 25445 25304
rect 25485 25264 25486 25304
rect 25444 25255 25486 25264
rect 25690 25304 25748 25305
rect 25690 25264 25699 25304
rect 25739 25264 25748 25304
rect 25690 25263 25748 25264
rect 26091 25304 26133 25313
rect 26091 25264 26092 25304
rect 26132 25264 26133 25304
rect 26091 25255 26133 25264
rect 26266 25304 26324 25305
rect 26266 25264 26275 25304
rect 26315 25264 26324 25304
rect 26266 25263 26324 25264
rect 26379 25304 26421 25313
rect 26379 25264 26380 25304
rect 26420 25264 26421 25304
rect 26379 25255 26421 25264
rect 26554 25304 26612 25305
rect 26554 25264 26563 25304
rect 26603 25264 26612 25304
rect 26554 25263 26612 25264
rect 26998 25304 27040 25313
rect 26998 25264 26999 25304
rect 27039 25264 27040 25304
rect 26998 25255 27040 25264
rect 27130 25304 27188 25305
rect 27130 25264 27139 25304
rect 27179 25264 27188 25304
rect 27130 25263 27188 25264
rect 27243 25304 27285 25313
rect 27243 25264 27244 25304
rect 27284 25264 27285 25304
rect 27243 25255 27285 25264
rect 27514 25304 27572 25305
rect 27514 25264 27523 25304
rect 27563 25264 27572 25304
rect 27514 25263 27572 25264
rect 28779 25304 28821 25313
rect 28779 25264 28780 25304
rect 28820 25264 28821 25304
rect 28779 25255 28821 25264
rect 29643 25304 29685 25313
rect 29643 25264 29644 25304
rect 29684 25264 29685 25304
rect 29643 25255 29685 25264
rect 30507 25304 30549 25313
rect 30507 25264 30508 25304
rect 30548 25264 30549 25304
rect 30507 25255 30549 25264
rect 30795 25304 30837 25313
rect 30795 25264 30796 25304
rect 30836 25264 30837 25304
rect 30795 25255 30837 25264
rect 21085 25180 21086 25220
rect 21126 25180 21127 25220
rect 21085 25171 21127 25180
rect 21562 25220 21620 25221
rect 21562 25180 21571 25220
rect 21611 25180 21620 25220
rect 25159 25213 25201 25222
rect 26667 25220 26709 25229
rect 21562 25179 21620 25180
rect 26667 25180 26668 25220
rect 26708 25180 26709 25220
rect 26667 25171 26709 25180
rect 26870 25220 26912 25229
rect 26870 25180 26871 25220
rect 26911 25180 26912 25220
rect 26870 25171 26912 25180
rect 27830 25220 27872 25229
rect 27830 25180 27831 25220
rect 27871 25180 27872 25220
rect 27830 25171 27872 25180
rect 28954 25220 29012 25221
rect 28954 25180 28963 25220
rect 29003 25180 29012 25220
rect 28954 25179 29012 25180
rect 987 25136 1029 25145
rect 987 25096 988 25136
rect 1028 25096 1029 25136
rect 987 25087 1029 25096
rect 1978 25136 2036 25137
rect 1978 25096 1987 25136
rect 2027 25096 2036 25136
rect 1978 25095 2036 25096
rect 2842 25136 2900 25137
rect 2842 25096 2851 25136
rect 2891 25096 2900 25136
rect 2842 25095 2900 25096
rect 5355 25136 5397 25145
rect 5355 25096 5356 25136
rect 5396 25096 5397 25136
rect 5355 25087 5397 25096
rect 6987 25136 7029 25145
rect 6987 25096 6988 25136
rect 7028 25096 7029 25136
rect 6987 25087 7029 25096
rect 7834 25136 7892 25137
rect 7834 25096 7843 25136
rect 7883 25096 7892 25136
rect 7834 25095 7892 25096
rect 11067 25136 11109 25145
rect 11067 25096 11068 25136
rect 11108 25096 11109 25136
rect 11067 25087 11109 25096
rect 13035 25136 13077 25145
rect 13035 25096 13036 25136
rect 13076 25096 13077 25136
rect 13035 25087 13077 25096
rect 13371 25136 13413 25145
rect 13371 25096 13372 25136
rect 13412 25096 13413 25136
rect 13371 25087 13413 25096
rect 15147 25136 15189 25145
rect 15147 25096 15148 25136
rect 15188 25096 15189 25136
rect 15147 25087 15189 25096
rect 16186 25136 16244 25137
rect 16186 25096 16195 25136
rect 16235 25096 16244 25136
rect 16186 25095 16244 25096
rect 19659 25136 19701 25145
rect 19659 25096 19660 25136
rect 19700 25096 19701 25136
rect 19659 25087 19701 25096
rect 20331 25136 20373 25145
rect 20331 25096 20332 25136
rect 20372 25096 20373 25136
rect 20331 25087 20373 25096
rect 20763 25136 20805 25145
rect 20763 25096 20764 25136
rect 20804 25096 20805 25136
rect 20763 25087 20805 25096
rect 21291 25136 21333 25145
rect 21291 25096 21292 25136
rect 21332 25096 21333 25136
rect 21291 25087 21333 25096
rect 23883 25136 23925 25145
rect 23883 25096 23884 25136
rect 23924 25096 23925 25136
rect 23883 25087 23925 25096
rect 24075 25136 24117 25145
rect 24075 25096 24076 25136
rect 24116 25096 24117 25136
rect 24075 25087 24117 25096
rect 25882 25136 25940 25137
rect 25882 25096 25891 25136
rect 25931 25096 25940 25136
rect 25882 25095 25940 25096
rect 27610 25136 27668 25137
rect 27610 25096 27619 25136
rect 27659 25096 27668 25136
rect 27610 25095 27668 25096
rect 27723 25136 27765 25145
rect 27723 25096 27724 25136
rect 27764 25096 27765 25136
rect 27723 25087 27765 25096
rect 29835 25136 29877 25145
rect 29835 25096 29836 25136
rect 29876 25096 29877 25136
rect 29835 25087 29877 25096
rect 30682 25136 30740 25137
rect 30682 25096 30691 25136
rect 30731 25096 30740 25136
rect 30682 25095 30740 25096
rect 576 24968 31392 24992
rect 576 24928 4352 24968
rect 4720 24928 12126 24968
rect 12494 24928 19900 24968
rect 20268 24928 27674 24968
rect 28042 24928 31392 24968
rect 576 24904 31392 24928
rect 1707 24800 1749 24809
rect 1707 24760 1708 24800
rect 1748 24760 1749 24800
rect 1707 24751 1749 24760
rect 13690 24800 13748 24801
rect 13690 24760 13699 24800
rect 13739 24760 13748 24800
rect 13690 24759 13748 24760
rect 17451 24800 17493 24809
rect 17451 24760 17452 24800
rect 17492 24760 17493 24800
rect 17451 24751 17493 24760
rect 19834 24800 19892 24801
rect 19834 24760 19843 24800
rect 19883 24760 19892 24800
rect 19834 24759 19892 24760
rect 20506 24800 20564 24801
rect 20506 24760 20515 24800
rect 20555 24760 20564 24800
rect 20506 24759 20564 24760
rect 22155 24800 22197 24809
rect 22155 24760 22156 24800
rect 22196 24760 22197 24800
rect 22155 24751 22197 24760
rect 22539 24800 22581 24809
rect 22539 24760 22540 24800
rect 22580 24760 22581 24800
rect 22539 24751 22581 24760
rect 23098 24800 23156 24801
rect 23098 24760 23107 24800
rect 23147 24760 23156 24800
rect 23098 24759 23156 24760
rect 23722 24800 23780 24801
rect 23722 24760 23731 24800
rect 23771 24760 23780 24800
rect 23722 24759 23780 24760
rect 24459 24800 24501 24809
rect 24459 24760 24460 24800
rect 24500 24760 24501 24800
rect 24459 24751 24501 24760
rect 25210 24800 25268 24801
rect 25210 24760 25219 24800
rect 25259 24760 25268 24800
rect 25210 24759 25268 24760
rect 26571 24800 26613 24809
rect 26571 24760 26572 24800
rect 26612 24760 26613 24800
rect 26571 24751 26613 24760
rect 31275 24800 31317 24809
rect 31275 24760 31276 24800
rect 31316 24760 31317 24800
rect 31275 24751 31317 24760
rect 1882 24716 1940 24717
rect 1882 24676 1891 24716
rect 1931 24676 1940 24716
rect 1882 24675 1940 24676
rect 6106 24716 6164 24717
rect 6106 24676 6115 24716
rect 6155 24676 6164 24716
rect 6106 24675 6164 24676
rect 8410 24716 8468 24717
rect 8410 24676 8419 24716
rect 8459 24676 8468 24716
rect 8410 24675 8468 24676
rect 9195 24716 9237 24725
rect 15130 24716 15188 24717
rect 9195 24676 9196 24716
rect 9236 24676 9237 24716
rect 9195 24667 9237 24676
rect 13506 24707 13552 24716
rect 13506 24667 13507 24707
rect 13547 24667 13552 24707
rect 15130 24676 15139 24716
rect 15179 24676 15188 24716
rect 15130 24675 15188 24676
rect 27613 24716 27655 24725
rect 27613 24676 27614 24716
rect 27654 24676 27655 24716
rect 27613 24667 27655 24676
rect 27819 24716 27861 24725
rect 27819 24676 27820 24716
rect 27860 24676 27861 24716
rect 27819 24667 27861 24676
rect 13506 24658 13552 24667
rect 2266 24632 2324 24633
rect 2266 24592 2275 24632
rect 2315 24592 2324 24632
rect 2266 24591 2324 24592
rect 4395 24632 4437 24641
rect 4395 24592 4396 24632
rect 4436 24592 4437 24632
rect 4395 24583 4437 24592
rect 8026 24632 8084 24633
rect 8026 24592 8035 24632
rect 8075 24592 8084 24632
rect 8026 24591 8084 24592
rect 8701 24632 8743 24641
rect 8701 24592 8702 24632
rect 8742 24592 8743 24632
rect 8701 24583 8743 24592
rect 8907 24632 8949 24641
rect 9291 24632 9333 24641
rect 8907 24592 8908 24632
rect 8948 24592 8949 24632
rect 8907 24583 8949 24592
rect 9003 24623 9045 24632
rect 9003 24583 9004 24623
rect 9044 24583 9045 24623
rect 9291 24592 9292 24632
rect 9332 24592 9333 24632
rect 9291 24583 9333 24592
rect 9508 24632 9550 24641
rect 9508 24592 9509 24632
rect 9549 24592 9550 24632
rect 9508 24583 9550 24592
rect 10234 24632 10292 24633
rect 10234 24592 10243 24632
rect 10283 24592 10292 24632
rect 10234 24591 10292 24592
rect 12363 24632 12405 24641
rect 12363 24592 12364 24632
rect 12404 24592 12405 24632
rect 12363 24583 12405 24592
rect 13210 24632 13268 24633
rect 13590 24632 13648 24633
rect 13210 24592 13219 24632
rect 13259 24592 13268 24632
rect 13210 24591 13268 24592
rect 13323 24623 13365 24632
rect 13323 24583 13324 24623
rect 13364 24583 13365 24623
rect 13590 24592 13599 24632
rect 13639 24592 13648 24632
rect 13590 24591 13648 24592
rect 13771 24632 13829 24633
rect 14667 24632 14709 24641
rect 13771 24592 13780 24632
rect 13820 24592 13829 24632
rect 13771 24591 13829 24592
rect 14178 24623 14224 24632
rect 9003 24574 9045 24583
rect 13323 24574 13365 24583
rect 14178 24583 14179 24623
rect 14219 24583 14224 24623
rect 14667 24592 14668 24632
rect 14708 24592 14709 24632
rect 14667 24583 14709 24592
rect 14781 24632 14839 24633
rect 14781 24592 14790 24632
rect 14830 24592 14839 24632
rect 14781 24591 14839 24592
rect 14908 24632 14966 24633
rect 14908 24592 14917 24632
rect 14957 24592 14966 24632
rect 14908 24591 14966 24592
rect 15514 24632 15572 24633
rect 15514 24592 15523 24632
rect 15563 24592 15572 24632
rect 15514 24591 15572 24592
rect 18123 24632 18165 24641
rect 18123 24592 18124 24632
rect 18164 24592 18165 24632
rect 18123 24583 18165 24592
rect 18315 24632 18357 24641
rect 19275 24632 19317 24641
rect 18315 24592 18316 24632
rect 18356 24592 18357 24632
rect 18315 24583 18357 24592
rect 18498 24623 18544 24632
rect 18498 24583 18499 24623
rect 18539 24583 18544 24623
rect 19275 24592 19276 24632
rect 19316 24592 19317 24632
rect 19275 24583 19317 24592
rect 19492 24632 19534 24641
rect 19492 24592 19493 24632
rect 19533 24592 19534 24632
rect 19492 24583 19534 24592
rect 19947 24632 19989 24641
rect 19947 24592 19948 24632
rect 19988 24592 19989 24632
rect 19947 24583 19989 24592
rect 20331 24632 20373 24641
rect 20331 24592 20332 24632
rect 20372 24592 20373 24632
rect 20331 24583 20373 24592
rect 20619 24632 20661 24641
rect 20619 24592 20620 24632
rect 20660 24592 20661 24632
rect 20619 24583 20661 24592
rect 21295 24632 21353 24633
rect 21295 24592 21304 24632
rect 21344 24592 21353 24632
rect 21295 24591 21353 24592
rect 21483 24632 21525 24641
rect 21483 24592 21484 24632
rect 21524 24592 21525 24632
rect 21483 24583 21525 24592
rect 22333 24632 22375 24641
rect 22333 24592 22334 24632
rect 22374 24592 22375 24632
rect 22333 24583 22375 24592
rect 22539 24632 22581 24641
rect 22774 24632 22816 24641
rect 22539 24592 22540 24632
rect 22580 24592 22581 24632
rect 22539 24583 22581 24592
rect 22635 24623 22677 24632
rect 22635 24583 22636 24623
rect 22676 24583 22677 24623
rect 22774 24592 22775 24632
rect 22815 24592 22816 24632
rect 22774 24583 22816 24592
rect 22906 24632 22964 24633
rect 22906 24592 22915 24632
rect 22955 24592 22964 24632
rect 22906 24591 22964 24592
rect 23019 24632 23061 24641
rect 23019 24592 23020 24632
rect 23060 24592 23061 24632
rect 23019 24583 23061 24592
rect 23403 24632 23445 24641
rect 23403 24592 23404 24632
rect 23444 24592 23445 24632
rect 23403 24583 23445 24592
rect 23887 24632 23945 24633
rect 23887 24592 23896 24632
rect 23936 24592 23945 24632
rect 23887 24591 23945 24592
rect 24075 24632 24117 24641
rect 24075 24592 24076 24632
rect 24116 24592 24117 24632
rect 24075 24583 24117 24592
rect 24189 24632 24247 24633
rect 24651 24632 24693 24641
rect 24189 24592 24198 24632
rect 24238 24592 24247 24632
rect 24189 24591 24247 24592
rect 24414 24623 24456 24632
rect 24307 24590 24365 24591
rect 14178 24574 14224 24583
rect 18498 24574 18544 24583
rect 22635 24574 22677 24583
rect 1323 24548 1365 24557
rect 1323 24508 1324 24548
rect 1364 24508 1365 24548
rect 1323 24499 1365 24508
rect 9410 24548 9452 24557
rect 9410 24508 9411 24548
rect 9451 24508 9452 24548
rect 9410 24499 9452 24508
rect 9867 24548 9909 24557
rect 9867 24508 9868 24548
rect 9908 24508 9909 24548
rect 9867 24499 9909 24508
rect 11787 24548 11829 24557
rect 11787 24508 11788 24548
rect 11828 24508 11829 24548
rect 11787 24499 11829 24508
rect 14331 24548 14373 24557
rect 14331 24508 14332 24548
rect 14372 24508 14373 24548
rect 14331 24499 14373 24508
rect 18651 24548 18693 24557
rect 18651 24508 18652 24548
rect 18692 24508 18693 24548
rect 18651 24499 18693 24508
rect 19179 24548 19221 24557
rect 19179 24508 19180 24548
rect 19220 24508 19221 24548
rect 19179 24499 19221 24508
rect 19394 24548 19436 24557
rect 19394 24508 19395 24548
rect 19435 24508 19436 24548
rect 19394 24499 19436 24508
rect 21130 24548 21188 24549
rect 21130 24508 21139 24548
rect 21179 24508 21188 24548
rect 21130 24507 21188 24508
rect 23259 24548 23301 24557
rect 24307 24550 24316 24590
rect 24356 24550 24365 24590
rect 24414 24583 24415 24623
rect 24455 24583 24456 24623
rect 24651 24592 24652 24632
rect 24692 24592 24693 24632
rect 24651 24583 24693 24592
rect 24886 24632 24928 24641
rect 24886 24592 24887 24632
rect 24927 24592 24928 24632
rect 24886 24583 24928 24592
rect 25131 24632 25173 24641
rect 25899 24632 25941 24641
rect 25131 24592 25132 24632
rect 25172 24592 25173 24632
rect 25131 24583 25173 24592
rect 25410 24623 25456 24632
rect 25410 24583 25411 24623
rect 25451 24583 25456 24623
rect 25899 24592 25900 24632
rect 25940 24592 25941 24632
rect 25899 24583 25941 24592
rect 26016 24632 26074 24633
rect 26016 24592 26025 24632
rect 26065 24592 26074 24632
rect 26016 24591 26074 24592
rect 26187 24632 26229 24641
rect 26187 24592 26188 24632
rect 26228 24592 26229 24632
rect 26187 24583 26229 24592
rect 26368 24632 26410 24641
rect 26907 24632 26949 24641
rect 26368 24592 26369 24632
rect 26409 24592 26410 24632
rect 26368 24583 26410 24592
rect 26667 24623 26709 24632
rect 26667 24583 26668 24623
rect 26708 24583 26709 24623
rect 26907 24592 26908 24632
rect 26948 24592 26949 24632
rect 26907 24583 26949 24592
rect 27137 24632 27179 24641
rect 27137 24592 27138 24632
rect 27178 24592 27179 24632
rect 27137 24583 27179 24592
rect 27322 24632 27380 24633
rect 27322 24592 27331 24632
rect 27371 24592 27380 24632
rect 27322 24591 27380 24592
rect 27435 24632 27477 24641
rect 28107 24632 28149 24641
rect 27435 24592 27436 24632
rect 27476 24592 27477 24632
rect 27435 24583 27477 24592
rect 27915 24623 27957 24632
rect 27915 24583 27916 24623
rect 27956 24583 27957 24623
rect 28107 24592 28108 24632
rect 28148 24592 28149 24632
rect 28107 24583 28149 24592
rect 29338 24632 29396 24633
rect 29338 24592 29347 24632
rect 29387 24592 29396 24632
rect 29338 24591 29396 24592
rect 24414 24574 24456 24583
rect 25410 24574 25456 24583
rect 26667 24574 26709 24583
rect 27915 24574 27957 24583
rect 24307 24549 24365 24550
rect 23259 24508 23260 24548
rect 23300 24508 23301 24548
rect 23259 24499 23301 24508
rect 24795 24548 24837 24557
rect 24795 24508 24796 24548
rect 24836 24508 24837 24548
rect 24795 24499 24837 24508
rect 25018 24548 25076 24549
rect 25018 24508 25027 24548
rect 25067 24508 25076 24548
rect 25018 24507 25076 24508
rect 25563 24548 25605 24557
rect 25563 24508 25564 24548
rect 25604 24508 25605 24548
rect 25563 24499 25605 24508
rect 28971 24548 29013 24557
rect 28971 24508 28972 24548
rect 29012 24508 29013 24548
rect 28971 24499 29013 24508
rect 939 24464 981 24473
rect 939 24424 940 24464
rect 980 24424 981 24464
rect 939 24415 981 24424
rect 4203 24464 4245 24473
rect 4203 24424 4204 24464
rect 4244 24424 4245 24464
rect 4203 24415 4245 24424
rect 5547 24464 5589 24473
rect 5547 24424 5548 24464
rect 5588 24424 5589 24464
rect 5547 24415 5589 24424
rect 5931 24464 5973 24473
rect 5931 24424 5932 24464
rect 5972 24424 5973 24464
rect 5931 24415 5973 24424
rect 13035 24464 13077 24473
rect 13035 24424 13036 24464
rect 13076 24424 13077 24464
rect 13035 24415 13077 24424
rect 14955 24464 14997 24473
rect 14955 24424 14956 24464
rect 14996 24424 14997 24464
rect 14955 24415 14997 24424
rect 17643 24464 17685 24473
rect 17643 24424 17644 24464
rect 17684 24424 17685 24464
rect 17643 24415 17685 24424
rect 20811 24464 20853 24473
rect 20811 24424 20812 24464
rect 20852 24424 20853 24464
rect 20811 24415 20853 24424
rect 26091 24464 26133 24473
rect 26091 24424 26092 24464
rect 26132 24424 26133 24464
rect 26091 24415 26133 24424
rect 26811 24464 26853 24473
rect 26811 24424 26812 24464
rect 26852 24424 26853 24464
rect 26811 24415 26853 24424
rect 27435 24464 27477 24473
rect 27435 24424 27436 24464
rect 27476 24424 27477 24464
rect 27435 24415 27477 24424
rect 1083 24380 1125 24389
rect 1083 24340 1084 24380
rect 1124 24340 1125 24380
rect 1083 24331 1125 24340
rect 5067 24380 5109 24389
rect 5067 24340 5068 24380
rect 5108 24340 5109 24380
rect 5067 24331 5109 24340
rect 6507 24380 6549 24389
rect 6507 24340 6508 24380
rect 6548 24340 6549 24380
rect 6507 24331 6549 24340
rect 8698 24380 8756 24381
rect 8698 24340 8707 24380
rect 8747 24340 8756 24380
rect 8698 24339 8756 24340
rect 12171 24380 12213 24389
rect 12171 24340 12172 24380
rect 12212 24340 12213 24380
rect 12171 24331 12213 24340
rect 18219 24380 18261 24389
rect 18219 24340 18220 24380
rect 18260 24340 18261 24380
rect 18219 24331 18261 24340
rect 22330 24380 22388 24381
rect 22330 24340 22339 24380
rect 22379 24340 22388 24380
rect 22330 24339 22388 24340
rect 26362 24380 26420 24381
rect 26362 24340 26371 24380
rect 26411 24340 26420 24380
rect 26362 24339 26420 24340
rect 27610 24380 27668 24381
rect 27610 24340 27619 24380
rect 27659 24340 27668 24380
rect 27610 24339 27668 24340
rect 28779 24380 28821 24389
rect 28779 24340 28780 24380
rect 28820 24340 28821 24380
rect 28779 24331 28821 24340
rect 576 24212 31392 24236
rect 576 24172 3112 24212
rect 3480 24172 10886 24212
rect 11254 24172 18660 24212
rect 19028 24172 26434 24212
rect 26802 24172 31392 24212
rect 576 24148 31392 24172
rect 1035 24044 1077 24053
rect 1035 24004 1036 24044
rect 1076 24004 1077 24044
rect 1035 23995 1077 24004
rect 4587 24044 4629 24053
rect 4587 24004 4588 24044
rect 4628 24004 4629 24044
rect 4587 23995 4629 24004
rect 6171 24044 6213 24053
rect 6171 24004 6172 24044
rect 6212 24004 6213 24044
rect 6171 23995 6213 24004
rect 10810 24044 10868 24045
rect 10810 24004 10819 24044
rect 10859 24004 10868 24044
rect 10810 24003 10868 24004
rect 16875 24044 16917 24053
rect 16875 24004 16876 24044
rect 16916 24004 16917 24044
rect 16875 23995 16917 24004
rect 24363 24044 24405 24053
rect 24363 24004 24364 24044
rect 24404 24004 24405 24044
rect 24363 23995 24405 24004
rect 25467 24044 25509 24053
rect 25467 24004 25468 24044
rect 25508 24004 25509 24044
rect 25467 23995 25509 24004
rect 28107 24044 28149 24053
rect 28107 24004 28108 24044
rect 28148 24004 28149 24044
rect 28107 23995 28149 24004
rect 12651 23960 12693 23969
rect 12651 23920 12652 23960
rect 12692 23920 12693 23960
rect 12651 23911 12693 23920
rect 14667 23960 14709 23969
rect 14667 23920 14668 23960
rect 14708 23920 14709 23960
rect 14667 23911 14709 23920
rect 19515 23960 19557 23969
rect 19515 23920 19516 23960
rect 19556 23920 19557 23960
rect 19515 23911 19557 23920
rect 24490 23960 24548 23961
rect 24490 23920 24499 23960
rect 24539 23920 24548 23960
rect 24490 23919 24548 23920
rect 27243 23960 27285 23969
rect 27243 23920 27244 23960
rect 27284 23920 27285 23960
rect 27243 23911 27285 23920
rect 9291 23876 9333 23885
rect 9291 23836 9292 23876
rect 9332 23836 9333 23876
rect 9291 23827 9333 23836
rect 9627 23876 9669 23885
rect 9627 23836 9628 23876
rect 9668 23836 9669 23876
rect 9627 23827 9669 23836
rect 10443 23876 10485 23885
rect 10443 23836 10444 23876
rect 10484 23836 10485 23876
rect 10443 23827 10485 23836
rect 14955 23876 14997 23885
rect 14955 23836 14956 23876
rect 14996 23836 14997 23876
rect 14955 23827 14997 23836
rect 18394 23876 18452 23877
rect 18394 23836 18403 23876
rect 18443 23836 18452 23876
rect 18394 23835 18452 23836
rect 23595 23876 23637 23885
rect 23595 23836 23596 23876
rect 23636 23836 23637 23876
rect 23595 23827 23637 23836
rect 28971 23876 29013 23885
rect 28971 23836 28972 23876
rect 29012 23836 29013 23876
rect 28971 23827 29013 23836
rect 2554 23792 2612 23793
rect 2554 23752 2563 23792
rect 2603 23752 2612 23792
rect 2554 23751 2612 23752
rect 4107 23792 4149 23801
rect 4107 23752 4108 23792
rect 4148 23752 4149 23792
rect 4107 23743 4149 23752
rect 4395 23792 4437 23801
rect 5259 23792 5301 23801
rect 4395 23752 4396 23792
rect 4436 23752 4437 23792
rect 4395 23743 4437 23752
rect 4971 23783 5013 23792
rect 4971 23743 4972 23783
rect 5012 23743 5013 23783
rect 5259 23752 5260 23792
rect 5300 23752 5301 23792
rect 5259 23743 5301 23752
rect 5547 23792 5589 23801
rect 5547 23752 5548 23792
rect 5588 23752 5589 23792
rect 5547 23743 5589 23752
rect 5931 23792 5973 23801
rect 5931 23752 5932 23792
rect 5972 23752 5973 23792
rect 5931 23743 5973 23752
rect 6637 23792 6695 23793
rect 6637 23752 6646 23792
rect 6686 23752 6695 23792
rect 6637 23751 6695 23752
rect 6970 23792 7028 23793
rect 6970 23752 6979 23792
rect 7019 23752 7028 23792
rect 6970 23751 7028 23752
rect 7659 23792 7701 23801
rect 7659 23752 7660 23792
rect 7700 23752 7701 23792
rect 7659 23743 7701 23752
rect 8715 23792 8757 23801
rect 8715 23752 8716 23792
rect 8756 23752 8757 23792
rect 8715 23743 8757 23752
rect 8803 23792 8861 23793
rect 8803 23752 8812 23792
rect 8852 23752 8861 23792
rect 8803 23751 8861 23752
rect 8962 23792 9020 23793
rect 8962 23752 8971 23792
rect 9011 23752 9020 23792
rect 8962 23751 9020 23752
rect 9082 23792 9140 23793
rect 9082 23752 9091 23792
rect 9131 23752 9140 23792
rect 9082 23751 9140 23752
rect 9195 23792 9237 23801
rect 9195 23752 9196 23792
rect 9236 23752 9237 23792
rect 9195 23743 9237 23752
rect 9483 23792 9525 23801
rect 9483 23752 9484 23792
rect 9524 23752 9525 23792
rect 9483 23743 9525 23752
rect 9771 23792 9813 23801
rect 9771 23752 9772 23792
rect 9812 23752 9813 23792
rect 9771 23743 9813 23752
rect 9963 23792 10005 23801
rect 9963 23752 9964 23792
rect 10004 23752 10005 23792
rect 9963 23743 10005 23752
rect 10102 23792 10144 23801
rect 10102 23752 10103 23792
rect 10143 23752 10144 23792
rect 10102 23743 10144 23752
rect 10234 23792 10292 23793
rect 10234 23752 10243 23792
rect 10283 23752 10292 23792
rect 10234 23751 10292 23752
rect 10347 23792 10389 23801
rect 10347 23752 10348 23792
rect 10388 23752 10389 23792
rect 10347 23743 10389 23752
rect 10630 23792 10672 23801
rect 10630 23752 10631 23792
rect 10671 23752 10672 23792
rect 10630 23743 10672 23752
rect 10810 23792 10868 23793
rect 10810 23752 10819 23792
rect 10859 23752 10868 23792
rect 10810 23751 10868 23752
rect 10999 23792 11057 23793
rect 10999 23752 11008 23792
rect 11048 23752 11057 23792
rect 10999 23751 11057 23752
rect 11163 23792 11205 23801
rect 11163 23752 11164 23792
rect 11204 23752 11205 23792
rect 11163 23743 11205 23752
rect 12363 23792 12405 23801
rect 12363 23752 12364 23792
rect 12404 23752 12405 23792
rect 12363 23743 12405 23752
rect 12651 23792 12693 23801
rect 12651 23752 12652 23792
rect 12692 23752 12693 23792
rect 12651 23743 12693 23752
rect 12766 23792 12808 23801
rect 12766 23752 12767 23792
rect 12807 23752 12808 23792
rect 12766 23743 12808 23752
rect 12939 23792 12981 23801
rect 12939 23752 12940 23792
rect 12980 23752 12981 23792
rect 12939 23743 12981 23752
rect 13131 23792 13173 23801
rect 13131 23752 13132 23792
rect 13172 23752 13173 23792
rect 13131 23743 13173 23752
rect 13515 23792 13557 23801
rect 13515 23752 13516 23792
rect 13556 23752 13557 23792
rect 13515 23743 13557 23752
rect 13995 23792 14037 23801
rect 13995 23752 13996 23792
rect 14036 23752 14037 23792
rect 13995 23743 14037 23752
rect 14266 23792 14324 23793
rect 14266 23752 14275 23792
rect 14315 23752 14324 23792
rect 14266 23751 14324 23752
rect 15322 23792 15380 23793
rect 15322 23752 15331 23792
rect 15371 23752 15380 23792
rect 15322 23751 15380 23752
rect 18123 23792 18165 23801
rect 18123 23752 18124 23792
rect 18164 23752 18165 23792
rect 18123 23743 18165 23752
rect 18795 23792 18837 23801
rect 18795 23752 18796 23792
rect 18836 23752 18837 23792
rect 18795 23743 18837 23752
rect 19018 23792 19076 23793
rect 19018 23752 19027 23792
rect 19067 23752 19076 23792
rect 19018 23751 19076 23752
rect 19659 23792 19701 23801
rect 19659 23752 19660 23792
rect 19700 23752 19701 23792
rect 19659 23743 19701 23752
rect 20026 23792 20084 23793
rect 20026 23752 20035 23792
rect 20075 23752 20084 23792
rect 20026 23751 20084 23752
rect 20139 23792 20181 23801
rect 20139 23752 20140 23792
rect 20180 23752 20181 23792
rect 20139 23743 20181 23752
rect 20763 23792 20805 23801
rect 20763 23752 20764 23792
rect 20804 23752 20805 23792
rect 20763 23743 20805 23752
rect 20907 23792 20949 23801
rect 20907 23752 20908 23792
rect 20948 23752 20949 23792
rect 20907 23743 20949 23752
rect 21723 23792 21765 23801
rect 21723 23752 21724 23792
rect 21764 23752 21765 23792
rect 21723 23743 21765 23752
rect 21867 23792 21909 23801
rect 21867 23752 21868 23792
rect 21908 23752 21909 23792
rect 21867 23743 21909 23752
rect 22330 23792 22388 23793
rect 22330 23752 22339 23792
rect 22379 23752 22388 23792
rect 22330 23751 22388 23752
rect 22448 23792 22506 23793
rect 22448 23752 22457 23792
rect 22497 23752 22506 23792
rect 22448 23751 22506 23752
rect 22616 23792 22658 23801
rect 22616 23752 22617 23792
rect 22657 23752 22658 23792
rect 22616 23743 22658 23752
rect 22714 23792 22772 23793
rect 22714 23752 22723 23792
rect 22763 23752 22772 23792
rect 22714 23751 22772 23752
rect 22848 23792 22906 23793
rect 22848 23752 22857 23792
rect 22897 23752 22906 23792
rect 22848 23751 22906 23752
rect 23407 23792 23465 23793
rect 23407 23752 23416 23792
rect 23456 23752 23465 23792
rect 23407 23751 23465 23752
rect 23691 23792 23733 23801
rect 23691 23752 23692 23792
rect 23732 23752 23733 23792
rect 23691 23743 23733 23752
rect 23810 23792 23852 23801
rect 23810 23752 23811 23792
rect 23851 23752 23852 23792
rect 23810 23743 23852 23752
rect 23931 23792 23973 23801
rect 23931 23752 23932 23792
rect 23972 23752 23973 23792
rect 23931 23743 23973 23752
rect 24058 23792 24116 23793
rect 24058 23752 24067 23792
rect 24107 23752 24116 23792
rect 24058 23751 24116 23752
rect 24699 23792 24757 23793
rect 24699 23752 24708 23792
rect 24748 23752 24757 23792
rect 24699 23751 24757 23752
rect 24843 23792 24885 23801
rect 24843 23752 24844 23792
rect 24884 23752 24885 23792
rect 24843 23743 24885 23752
rect 25078 23792 25120 23801
rect 25323 23792 25365 23801
rect 25078 23752 25079 23792
rect 25119 23752 25120 23792
rect 25078 23743 25120 23752
rect 25218 23783 25264 23792
rect 25218 23743 25219 23783
rect 25259 23743 25264 23783
rect 25323 23752 25324 23792
rect 25364 23752 25365 23792
rect 25323 23743 25365 23752
rect 25611 23792 25653 23801
rect 25611 23752 25612 23792
rect 25652 23752 25653 23792
rect 25611 23743 25653 23752
rect 25846 23792 25888 23801
rect 26091 23792 26133 23801
rect 25846 23752 25847 23792
rect 25887 23752 25888 23792
rect 25846 23743 25888 23752
rect 25986 23783 26032 23792
rect 25986 23743 25987 23783
rect 26027 23743 26032 23783
rect 26091 23752 26092 23792
rect 26132 23752 26133 23792
rect 26091 23743 26133 23752
rect 26458 23792 26516 23793
rect 26458 23752 26467 23792
rect 26507 23752 26516 23792
rect 26458 23751 26516 23752
rect 26774 23792 26816 23801
rect 26774 23752 26775 23792
rect 26815 23752 26816 23792
rect 26774 23743 26816 23752
rect 26938 23792 26996 23793
rect 26938 23752 26947 23792
rect 26987 23752 26996 23792
rect 26938 23751 26996 23752
rect 27243 23792 27285 23801
rect 27243 23752 27244 23792
rect 27284 23752 27285 23792
rect 27243 23743 27285 23752
rect 27627 23792 27669 23801
rect 27627 23752 27628 23792
rect 27668 23752 27669 23792
rect 27627 23743 27669 23752
rect 27771 23792 27813 23801
rect 27771 23752 27772 23792
rect 27812 23752 27813 23792
rect 27771 23743 27813 23752
rect 28779 23792 28821 23801
rect 28779 23752 28780 23792
rect 28820 23752 28821 23792
rect 28779 23743 28821 23752
rect 29338 23792 29396 23793
rect 29338 23752 29347 23792
rect 29387 23752 29396 23792
rect 29338 23751 29396 23752
rect 4971 23734 5013 23743
rect 25218 23734 25264 23743
rect 25986 23734 26032 23743
rect 634 23708 692 23709
rect 634 23668 643 23708
rect 683 23668 692 23708
rect 634 23667 692 23668
rect 2938 23708 2996 23709
rect 2938 23668 2947 23708
rect 2987 23668 2996 23708
rect 2938 23667 2996 23668
rect 3418 23708 3476 23709
rect 3418 23668 3427 23708
rect 3467 23668 3476 23708
rect 3418 23667 3476 23668
rect 4875 23708 4917 23717
rect 4875 23668 4876 23708
rect 4916 23668 4917 23708
rect 4875 23659 4917 23668
rect 6442 23708 6500 23709
rect 6442 23668 6451 23708
rect 6491 23668 6500 23708
rect 6442 23667 6500 23668
rect 7289 23708 7331 23717
rect 7289 23668 7290 23708
rect 7330 23668 7331 23708
rect 7289 23659 7331 23668
rect 8509 23708 8551 23717
rect 8509 23668 8510 23708
rect 8550 23668 8551 23708
rect 8509 23659 8551 23668
rect 14379 23708 14421 23717
rect 14379 23668 14380 23708
rect 14420 23668 14421 23708
rect 14379 23659 14421 23668
rect 17434 23708 17492 23709
rect 17434 23668 17443 23708
rect 17483 23668 17492 23708
rect 17434 23667 17492 23668
rect 19227 23708 19269 23717
rect 19227 23668 19228 23708
rect 19268 23668 19269 23708
rect 19227 23659 19269 23668
rect 23242 23708 23300 23709
rect 23242 23668 23251 23708
rect 23291 23668 23300 23708
rect 23242 23667 23300 23668
rect 24377 23708 24419 23717
rect 24377 23668 24378 23708
rect 24418 23668 24419 23708
rect 24377 23659 24419 23668
rect 27418 23708 27476 23709
rect 27418 23668 27427 23708
rect 27467 23668 27476 23708
rect 27418 23667 27476 23668
rect 4251 23624 4293 23633
rect 4251 23584 4252 23624
rect 4292 23584 4293 23624
rect 4251 23575 4293 23584
rect 7066 23624 7124 23625
rect 7066 23584 7075 23624
rect 7115 23584 7124 23624
rect 7066 23583 7124 23584
rect 7179 23624 7221 23633
rect 7179 23584 7180 23624
rect 7220 23584 7221 23624
rect 7179 23575 7221 23584
rect 8331 23624 8373 23633
rect 8331 23584 8332 23624
rect 8372 23584 8373 23624
rect 8331 23575 8373 23584
rect 8602 23624 8660 23625
rect 8602 23584 8611 23624
rect 8651 23584 8660 23624
rect 8602 23583 8660 23584
rect 9946 23624 10004 23625
rect 9946 23584 9955 23624
rect 9995 23584 10004 23624
rect 9946 23583 10004 23584
rect 11691 23624 11733 23633
rect 11691 23584 11692 23624
rect 11732 23584 11733 23624
rect 11691 23575 11733 23584
rect 13611 23624 13653 23633
rect 13611 23584 13612 23624
rect 13652 23584 13653 23624
rect 13611 23575 13653 23584
rect 17259 23624 17301 23633
rect 17259 23584 17260 23624
rect 17300 23584 17301 23624
rect 17259 23575 17301 23584
rect 20427 23624 20469 23633
rect 20427 23584 20428 23624
rect 20468 23584 20469 23624
rect 20427 23575 20469 23584
rect 20602 23624 20660 23625
rect 20602 23584 20611 23624
rect 20651 23584 20660 23624
rect 20602 23583 20660 23584
rect 21562 23624 21620 23625
rect 21562 23584 21571 23624
rect 21611 23584 21620 23624
rect 21562 23583 21620 23584
rect 22810 23624 22868 23625
rect 22810 23584 22819 23624
rect 22859 23584 22868 23624
rect 22810 23583 22868 23584
rect 24154 23624 24212 23625
rect 24154 23584 24163 23624
rect 24203 23584 24212 23624
rect 24154 23583 24212 23584
rect 25035 23624 25077 23633
rect 25035 23584 25036 23624
rect 25076 23584 25077 23624
rect 25035 23575 25077 23584
rect 25803 23624 25845 23633
rect 25803 23584 25804 23624
rect 25844 23584 25845 23624
rect 25803 23575 25845 23584
rect 26554 23624 26612 23625
rect 26554 23584 26563 23624
rect 26603 23584 26612 23624
rect 26554 23583 26612 23584
rect 26667 23624 26709 23633
rect 26667 23584 26668 23624
rect 26708 23584 26709 23624
rect 26667 23575 26709 23584
rect 27723 23624 27765 23633
rect 27723 23584 27724 23624
rect 27764 23584 27765 23624
rect 27723 23575 27765 23584
rect 31275 23624 31317 23633
rect 31275 23584 31276 23624
rect 31316 23584 31317 23624
rect 31275 23575 31317 23584
rect 576 23456 31392 23480
rect 576 23416 4352 23456
rect 4720 23416 12126 23456
rect 12494 23416 19900 23456
rect 20268 23416 27674 23456
rect 28042 23416 31392 23456
rect 576 23392 31392 23416
rect 1690 23288 1748 23289
rect 1690 23248 1699 23288
rect 1739 23248 1748 23288
rect 1690 23247 1748 23248
rect 3562 23288 3620 23289
rect 3562 23248 3571 23288
rect 3611 23248 3620 23288
rect 3562 23247 3620 23248
rect 3994 23288 4052 23289
rect 3994 23248 4003 23288
rect 4043 23248 4052 23288
rect 3994 23247 4052 23248
rect 4107 23288 4149 23297
rect 4107 23248 4108 23288
rect 4148 23248 4149 23288
rect 4107 23239 4149 23248
rect 4779 23288 4821 23297
rect 4779 23248 4780 23288
rect 4820 23248 4821 23288
rect 4779 23239 4821 23248
rect 5067 23288 5109 23297
rect 5067 23248 5068 23288
rect 5108 23248 5109 23288
rect 5067 23239 5109 23248
rect 5626 23288 5684 23289
rect 5626 23248 5635 23288
rect 5675 23248 5684 23288
rect 5626 23247 5684 23248
rect 11482 23288 11540 23289
rect 11482 23248 11491 23288
rect 11531 23248 11540 23288
rect 11482 23247 11540 23248
rect 12891 23288 12933 23297
rect 12891 23248 12892 23288
rect 12932 23248 12933 23288
rect 12891 23239 12933 23248
rect 15034 23288 15092 23289
rect 15034 23248 15043 23288
rect 15083 23248 15092 23288
rect 15034 23247 15092 23248
rect 18202 23288 18260 23289
rect 18202 23248 18211 23288
rect 18251 23248 18260 23288
rect 18202 23247 18260 23248
rect 18507 23288 18549 23297
rect 18507 23248 18508 23288
rect 18548 23248 18549 23288
rect 18507 23239 18549 23248
rect 19179 23288 19221 23297
rect 19179 23248 19180 23288
rect 19220 23248 19221 23288
rect 19179 23239 19221 23248
rect 20410 23288 20468 23289
rect 20410 23248 20419 23288
rect 20459 23248 20468 23288
rect 20410 23247 20468 23248
rect 20523 23288 20565 23297
rect 20523 23248 20524 23288
rect 20564 23248 20565 23288
rect 20523 23239 20565 23248
rect 21610 23288 21668 23289
rect 21610 23248 21619 23288
rect 21659 23248 21668 23288
rect 21610 23247 21668 23248
rect 28491 23288 28533 23297
rect 28491 23248 28492 23288
rect 28532 23248 28533 23288
rect 28491 23239 28533 23248
rect 2170 23204 2228 23205
rect 2170 23164 2179 23204
rect 2219 23164 2228 23204
rect 2170 23163 2228 23164
rect 2283 23204 2325 23213
rect 2283 23164 2284 23204
rect 2324 23164 2325 23204
rect 2283 23155 2325 23164
rect 3243 23204 3285 23213
rect 3243 23164 3244 23204
rect 3284 23164 3285 23204
rect 3243 23155 3285 23164
rect 4666 23204 4724 23205
rect 4666 23164 4675 23204
rect 4715 23164 4724 23204
rect 4666 23163 4724 23164
rect 5533 23204 5575 23213
rect 5533 23164 5534 23204
rect 5574 23164 5575 23204
rect 5533 23155 5575 23164
rect 6106 23204 6164 23205
rect 6106 23164 6115 23204
rect 6155 23164 6164 23204
rect 6106 23163 6164 23164
rect 10731 23204 10773 23213
rect 10731 23164 10732 23204
rect 10772 23164 10773 23204
rect 10731 23155 10773 23164
rect 15339 23204 15381 23213
rect 15339 23164 15340 23204
rect 15380 23164 15381 23204
rect 15339 23155 15381 23164
rect 16666 23204 16724 23205
rect 16666 23164 16675 23204
rect 16715 23164 16724 23204
rect 16666 23163 16724 23164
rect 17931 23204 17973 23213
rect 17931 23164 17932 23204
rect 17972 23164 17973 23204
rect 17931 23155 17973 23164
rect 19978 23204 20036 23205
rect 19978 23164 19987 23204
rect 20027 23164 20036 23204
rect 19978 23163 20036 23164
rect 20633 23204 20675 23213
rect 20633 23164 20634 23204
rect 20674 23164 20675 23204
rect 20633 23155 20675 23164
rect 20955 23204 20997 23213
rect 20955 23164 20956 23204
rect 20996 23164 20997 23204
rect 20955 23155 20997 23164
rect 25131 23204 25173 23213
rect 26955 23204 26997 23213
rect 25131 23164 25132 23204
rect 25172 23164 25173 23204
rect 25131 23155 25173 23164
rect 25794 23195 25840 23204
rect 25794 23155 25795 23195
rect 25835 23155 25840 23195
rect 26955 23164 26956 23204
rect 26996 23164 26997 23204
rect 26955 23155 26997 23164
rect 25794 23146 25840 23155
rect 843 23120 885 23129
rect 843 23080 844 23120
rect 884 23080 885 23120
rect 843 23071 885 23080
rect 1018 23120 1076 23121
rect 1018 23080 1027 23120
rect 1067 23080 1076 23120
rect 1018 23079 1076 23080
rect 1227 23120 1269 23129
rect 1227 23080 1228 23120
rect 1268 23080 1269 23120
rect 1227 23071 1269 23080
rect 1402 23120 1460 23121
rect 1402 23080 1411 23120
rect 1451 23080 1460 23120
rect 1402 23079 1460 23080
rect 1594 23120 1652 23121
rect 1594 23080 1603 23120
rect 1643 23080 1652 23120
rect 1594 23079 1652 23080
rect 1913 23120 1955 23129
rect 1913 23080 1914 23120
rect 1954 23080 1955 23120
rect 1913 23071 1955 23080
rect 2080 23120 2122 23129
rect 2571 23120 2613 23129
rect 2080 23080 2081 23120
rect 2121 23080 2122 23120
rect 2080 23071 2122 23080
rect 2379 23111 2421 23120
rect 2379 23071 2380 23111
rect 2420 23071 2421 23111
rect 2571 23080 2572 23120
rect 2612 23080 2613 23120
rect 2571 23071 2613 23080
rect 3727 23120 3785 23121
rect 3727 23080 3736 23120
rect 3776 23080 3785 23120
rect 3727 23079 3785 23080
rect 3904 23120 3946 23129
rect 4573 23120 4615 23129
rect 5163 23120 5205 23129
rect 3904 23080 3905 23120
rect 3945 23080 3946 23120
rect 3904 23071 3946 23080
rect 4203 23111 4245 23120
rect 4203 23071 4204 23111
rect 4244 23071 4245 23111
rect 4573 23080 4574 23120
rect 4614 23080 4615 23120
rect 4573 23071 4615 23080
rect 4875 23111 4917 23120
rect 4875 23071 4876 23111
rect 4916 23071 4917 23111
rect 5163 23080 5164 23120
rect 5204 23080 5205 23120
rect 5163 23071 5205 23080
rect 5392 23120 5450 23121
rect 5392 23080 5401 23120
rect 5441 23080 5450 23120
rect 5392 23079 5450 23080
rect 5739 23120 5781 23129
rect 7083 23120 7125 23129
rect 5739 23080 5740 23120
rect 5780 23080 5781 23120
rect 5739 23071 5781 23080
rect 5835 23111 5877 23120
rect 5835 23071 5836 23111
rect 5876 23071 5877 23111
rect 7083 23080 7084 23120
rect 7124 23080 7125 23120
rect 7083 23071 7125 23080
rect 7467 23120 7509 23129
rect 7467 23080 7468 23120
rect 7508 23080 7509 23120
rect 7467 23071 7509 23080
rect 8331 23120 8373 23129
rect 8331 23080 8332 23120
rect 8372 23080 8373 23120
rect 8331 23071 8373 23080
rect 8506 23120 8564 23121
rect 8506 23080 8515 23120
rect 8555 23080 8564 23120
rect 8506 23079 8564 23080
rect 9771 23120 9813 23129
rect 9771 23080 9772 23120
rect 9812 23080 9813 23120
rect 9771 23071 9813 23080
rect 10347 23120 10389 23129
rect 10347 23080 10348 23120
rect 10388 23080 10389 23120
rect 10347 23071 10389 23080
rect 10576 23120 10634 23121
rect 10576 23080 10585 23120
rect 10625 23080 10634 23120
rect 10576 23079 10634 23080
rect 10827 23120 10869 23129
rect 10827 23080 10828 23120
rect 10868 23080 10869 23120
rect 10827 23071 10869 23080
rect 11044 23120 11086 23129
rect 11044 23080 11045 23120
rect 11085 23080 11086 23120
rect 11044 23071 11086 23080
rect 11163 23120 11205 23129
rect 11163 23080 11164 23120
rect 11204 23080 11205 23120
rect 11163 23071 11205 23080
rect 11290 23120 11348 23121
rect 11290 23080 11299 23120
rect 11339 23080 11348 23120
rect 11290 23079 11348 23080
rect 11403 23120 11445 23129
rect 11403 23080 11404 23120
rect 11444 23080 11445 23120
rect 11403 23071 11445 23080
rect 11883 23120 11925 23129
rect 11883 23080 11884 23120
rect 11924 23080 11925 23120
rect 11883 23071 11925 23080
rect 12112 23120 12170 23121
rect 12112 23080 12121 23120
rect 12161 23080 12170 23120
rect 12112 23079 12170 23080
rect 12363 23120 12405 23129
rect 12363 23080 12364 23120
rect 12404 23080 12405 23120
rect 12363 23071 12405 23080
rect 12555 23120 12597 23129
rect 12555 23080 12556 23120
rect 12596 23080 12597 23120
rect 12555 23071 12597 23080
rect 12747 23120 12789 23129
rect 12747 23080 12748 23120
rect 12788 23080 12789 23120
rect 12747 23071 12789 23080
rect 13419 23120 13461 23129
rect 13419 23080 13420 23120
rect 13460 23080 13461 23120
rect 13419 23071 13461 23080
rect 13611 23120 13653 23129
rect 13611 23080 13612 23120
rect 13652 23080 13653 23120
rect 13611 23071 13653 23080
rect 13803 23120 13845 23129
rect 13803 23080 13804 23120
rect 13844 23080 13845 23120
rect 13803 23071 13845 23080
rect 13978 23120 14036 23121
rect 13978 23080 13987 23120
rect 14027 23080 14036 23120
rect 13978 23079 14036 23080
rect 14283 23120 14325 23129
rect 14283 23080 14284 23120
rect 14324 23080 14325 23120
rect 14283 23071 14325 23080
rect 14512 23120 14570 23121
rect 14512 23080 14521 23120
rect 14561 23080 14570 23120
rect 14512 23079 14570 23080
rect 14859 23115 14901 23124
rect 14859 23075 14860 23115
rect 14900 23075 14901 23115
rect 15046 23120 15104 23121
rect 15046 23080 15055 23120
rect 15095 23080 15104 23120
rect 15046 23079 15104 23080
rect 15243 23120 15285 23129
rect 15243 23080 15244 23120
rect 15284 23080 15285 23120
rect 2379 23062 2421 23071
rect 4203 23062 4245 23071
rect 4875 23062 4917 23071
rect 5835 23062 5877 23071
rect 14859 23066 14901 23075
rect 15243 23071 15285 23080
rect 15435 23120 15477 23129
rect 15435 23080 15436 23120
rect 15476 23080 15477 23120
rect 15435 23071 15477 23080
rect 17451 23120 17493 23129
rect 17451 23080 17452 23120
rect 17492 23080 17493 23120
rect 17451 23071 17493 23080
rect 17835 23120 17877 23129
rect 17835 23080 17836 23120
rect 17876 23080 17877 23120
rect 17835 23071 17877 23080
rect 18027 23120 18069 23129
rect 18027 23080 18028 23120
rect 18068 23080 18069 23120
rect 18027 23071 18069 23080
rect 18315 23120 18357 23129
rect 18315 23080 18316 23120
rect 18356 23080 18357 23120
rect 18315 23071 18357 23080
rect 19179 23120 19221 23129
rect 19179 23080 19180 23120
rect 19220 23080 19221 23120
rect 19179 23071 19221 23080
rect 19371 23120 19413 23129
rect 19371 23080 19372 23120
rect 19412 23080 19413 23120
rect 19371 23071 19413 23080
rect 20143 23120 20201 23121
rect 20143 23080 20152 23120
rect 20192 23080 20201 23120
rect 20143 23079 20201 23080
rect 20314 23120 20372 23121
rect 20314 23080 20323 23120
rect 20363 23080 20372 23120
rect 20314 23079 20372 23080
rect 20811 23120 20853 23129
rect 21466 23120 21524 23121
rect 20811 23080 20812 23120
rect 20852 23080 20853 23120
rect 20811 23071 20853 23080
rect 21375 23111 21417 23120
rect 21375 23071 21376 23111
rect 21416 23071 21417 23111
rect 21466 23080 21475 23120
rect 21515 23080 21524 23120
rect 21466 23079 21524 23080
rect 21771 23120 21813 23129
rect 21771 23080 21772 23120
rect 21812 23080 21813 23120
rect 21771 23071 21813 23080
rect 21963 23120 22005 23129
rect 21963 23080 21964 23120
rect 22004 23080 22005 23120
rect 21963 23071 22005 23080
rect 22522 23120 22580 23121
rect 22522 23080 22531 23120
rect 22571 23080 22580 23120
rect 22522 23079 22580 23080
rect 24826 23120 24884 23121
rect 24826 23080 24835 23120
rect 24875 23080 24884 23120
rect 24826 23079 24884 23080
rect 25498 23120 25556 23121
rect 25882 23120 25940 23121
rect 25498 23080 25507 23120
rect 25547 23080 25556 23120
rect 25498 23079 25556 23080
rect 25611 23111 25653 23120
rect 25611 23071 25612 23111
rect 25652 23071 25653 23111
rect 25882 23080 25891 23120
rect 25931 23080 25940 23120
rect 25882 23079 25940 23080
rect 26059 23120 26117 23121
rect 26059 23080 26068 23120
rect 26108 23080 26117 23120
rect 26059 23079 26117 23080
rect 26458 23120 26516 23121
rect 26458 23080 26467 23120
rect 26507 23080 26516 23120
rect 26458 23079 26516 23080
rect 26650 23120 26708 23121
rect 26650 23080 26659 23120
rect 26699 23080 26708 23120
rect 26650 23079 26708 23080
rect 26763 23120 26805 23129
rect 26763 23080 26764 23120
rect 26804 23080 26805 23120
rect 27202 23120 27260 23121
rect 26763 23071 26805 23080
rect 27068 23105 27110 23114
rect 21375 23062 21417 23071
rect 25611 23062 25653 23071
rect 27068 23065 27069 23105
rect 27109 23065 27110 23105
rect 27202 23080 27211 23120
rect 27251 23080 27260 23120
rect 27202 23079 27260 23080
rect 27435 23120 27477 23129
rect 27435 23080 27436 23120
rect 27476 23080 27477 23120
rect 27435 23071 27477 23080
rect 28044 23120 28102 23121
rect 28044 23080 28053 23120
rect 28093 23080 28102 23120
rect 28044 23079 28102 23080
rect 28203 23120 28245 23129
rect 28203 23080 28204 23120
rect 28244 23080 28245 23120
rect 29355 23120 29397 23129
rect 28203 23071 28245 23080
rect 28337 23088 28395 23089
rect 27068 23056 27110 23065
rect 28337 23048 28346 23088
rect 28386 23048 28395 23088
rect 29355 23080 29356 23120
rect 29396 23080 29397 23120
rect 29355 23071 29397 23080
rect 29547 23120 29589 23129
rect 29547 23080 29548 23120
rect 29588 23080 29589 23120
rect 29547 23071 29589 23080
rect 30394 23120 30452 23121
rect 30394 23080 30403 23120
rect 30443 23080 30452 23120
rect 30394 23079 30452 23080
rect 31083 23120 31125 23129
rect 31083 23080 31084 23120
rect 31124 23080 31125 23120
rect 31083 23071 31125 23080
rect 28337 23047 28395 23048
rect 5067 23036 5109 23045
rect 5067 22996 5068 23036
rect 5108 22996 5109 23036
rect 5067 22987 5109 22996
rect 5282 23036 5324 23045
rect 5282 22996 5283 23036
rect 5323 22996 5324 23036
rect 5282 22987 5324 22996
rect 10251 23036 10293 23045
rect 10251 22996 10252 23036
rect 10292 22996 10293 23036
rect 10251 22987 10293 22996
rect 10466 23036 10508 23045
rect 10466 22996 10467 23036
rect 10507 22996 10508 23036
rect 10466 22987 10508 22996
rect 10946 23036 10988 23045
rect 10946 22996 10947 23036
rect 10987 22996 10988 23036
rect 10946 22987 10988 22996
rect 11787 23036 11829 23045
rect 13227 23036 13269 23045
rect 11787 22996 11788 23036
rect 11828 22996 11829 23036
rect 11787 22987 11829 22996
rect 12018 23027 12064 23036
rect 12018 22987 12019 23027
rect 12059 22987 12064 23027
rect 13227 22996 13228 23036
rect 13268 22996 13269 23036
rect 13227 22987 13269 22996
rect 14187 23036 14229 23045
rect 14187 22996 14188 23036
rect 14228 22996 14229 23036
rect 14187 22987 14229 22996
rect 14402 23036 14444 23045
rect 14402 22996 14403 23036
rect 14443 22996 14444 23036
rect 14402 22987 14444 22996
rect 22155 23036 22197 23045
rect 22155 22996 22156 23036
rect 22196 22996 22197 23036
rect 22155 22987 22197 22996
rect 24651 23036 24693 23045
rect 24651 22996 24652 23036
rect 24692 22996 24693 23036
rect 24651 22987 24693 22996
rect 25227 23036 25269 23045
rect 25227 22996 25228 23036
rect 25268 22996 25269 23036
rect 25227 22987 25269 22996
rect 27322 23036 27380 23037
rect 27322 22996 27331 23036
rect 27371 22996 27380 23036
rect 27322 22995 27380 22996
rect 27531 23036 27573 23045
rect 27531 22996 27532 23036
rect 27572 22996 27573 23036
rect 27531 22987 27573 22996
rect 27850 23036 27908 23037
rect 27850 22996 27859 23036
rect 27899 22996 27908 23036
rect 27850 22995 27908 22996
rect 12018 22978 12064 22987
rect 1018 22952 1076 22953
rect 1018 22912 1027 22952
rect 1067 22912 1076 22952
rect 1018 22911 1076 22912
rect 1402 22952 1460 22953
rect 1402 22912 1411 22952
rect 1451 22912 1460 22952
rect 1402 22911 1460 22912
rect 8506 22952 8564 22953
rect 8506 22912 8515 22952
rect 8555 22912 8564 22952
rect 8506 22911 8564 22912
rect 8986 22952 9044 22953
rect 8986 22912 8995 22952
rect 9035 22912 9044 22952
rect 8986 22911 9044 22912
rect 13978 22952 14036 22953
rect 13978 22912 13987 22952
rect 14027 22912 14036 22952
rect 13978 22911 14036 22912
rect 15819 22952 15861 22961
rect 15819 22912 15820 22952
rect 15860 22912 15861 22952
rect 15819 22903 15861 22912
rect 16011 22952 16053 22961
rect 16011 22912 16012 22952
rect 16052 22912 16053 22952
rect 16011 22903 16053 22912
rect 18699 22952 18741 22961
rect 18699 22912 18700 22952
rect 18740 22912 18741 22952
rect 18699 22903 18741 22912
rect 21771 22952 21813 22961
rect 21771 22912 21772 22952
rect 21812 22912 21813 22952
rect 21771 22903 21813 22912
rect 24459 22952 24501 22961
rect 24459 22912 24460 22952
rect 24500 22912 24501 22952
rect 24459 22903 24501 22912
rect 1899 22868 1941 22877
rect 1899 22828 1900 22868
rect 1940 22828 1941 22868
rect 1899 22819 1941 22828
rect 8139 22868 8181 22877
rect 8139 22828 8140 22868
rect 8180 22828 8181 22868
rect 8139 22819 8181 22828
rect 12459 22868 12501 22877
rect 12459 22828 12460 22868
rect 12500 22828 12501 22868
rect 12459 22819 12501 22828
rect 12987 22868 13029 22877
rect 12987 22828 12988 22868
rect 13028 22828 13029 22868
rect 12987 22819 13029 22828
rect 13419 22868 13461 22877
rect 13419 22828 13420 22868
rect 13460 22828 13461 22868
rect 13419 22819 13461 22828
rect 21082 22868 21140 22869
rect 21082 22828 21091 22868
rect 21131 22828 21140 22868
rect 21082 22827 21140 22828
rect 25498 22868 25556 22869
rect 25498 22828 25507 22868
rect 25547 22828 25556 22868
rect 25498 22827 25556 22828
rect 28683 22868 28725 22877
rect 28683 22828 28684 22868
rect 28724 22828 28725 22868
rect 28683 22819 28725 22828
rect 30219 22868 30261 22877
rect 30219 22828 30220 22868
rect 30260 22828 30261 22868
rect 30219 22819 30261 22828
rect 576 22700 31392 22724
rect 576 22660 3112 22700
rect 3480 22660 10886 22700
rect 11254 22660 18660 22700
rect 19028 22660 26434 22700
rect 26802 22660 31392 22700
rect 576 22636 31392 22660
rect 6010 22532 6068 22533
rect 6010 22492 6019 22532
rect 6059 22492 6068 22532
rect 6010 22491 6068 22492
rect 7258 22532 7316 22533
rect 7258 22492 7267 22532
rect 7307 22492 7316 22532
rect 7258 22491 7316 22492
rect 10635 22532 10677 22541
rect 10635 22492 10636 22532
rect 10676 22492 10677 22532
rect 10635 22483 10677 22492
rect 11403 22532 11445 22541
rect 11403 22492 11404 22532
rect 11444 22492 11445 22532
rect 11403 22483 11445 22492
rect 11691 22532 11733 22541
rect 11691 22492 11692 22532
rect 11732 22492 11733 22532
rect 11691 22483 11733 22492
rect 14554 22532 14612 22533
rect 14554 22492 14563 22532
rect 14603 22492 14612 22532
rect 14554 22491 14612 22492
rect 20314 22532 20372 22533
rect 20314 22492 20323 22532
rect 20363 22492 20372 22532
rect 20314 22491 20372 22492
rect 21178 22532 21236 22533
rect 21178 22492 21187 22532
rect 21227 22492 21236 22532
rect 21178 22491 21236 22492
rect 21946 22532 22004 22533
rect 21946 22492 21955 22532
rect 21995 22492 22004 22532
rect 21946 22491 22004 22492
rect 23962 22532 24020 22533
rect 23962 22492 23971 22532
rect 24011 22492 24020 22532
rect 23962 22491 24020 22492
rect 25899 22532 25941 22541
rect 25899 22492 25900 22532
rect 25940 22492 25941 22532
rect 25899 22483 25941 22492
rect 27147 22532 27189 22541
rect 27147 22492 27148 22532
rect 27188 22492 27189 22532
rect 27147 22483 27189 22492
rect 27723 22532 27765 22541
rect 27723 22492 27724 22532
rect 27764 22492 27765 22532
rect 27723 22483 27765 22492
rect 8986 22448 9044 22449
rect 8986 22408 8995 22448
rect 9035 22408 9044 22448
rect 8986 22407 9044 22408
rect 16474 22448 16532 22449
rect 16474 22408 16483 22448
rect 16523 22408 16532 22448
rect 16474 22407 16532 22408
rect 17739 22448 17781 22457
rect 17739 22408 17740 22448
rect 17780 22408 17781 22448
rect 17739 22399 17781 22408
rect 18891 22448 18933 22457
rect 18891 22408 18892 22448
rect 18932 22408 18933 22448
rect 18891 22399 18933 22408
rect 19258 22448 19316 22449
rect 19258 22408 19267 22448
rect 19307 22408 19316 22448
rect 19258 22407 19316 22408
rect 24267 22448 24309 22457
rect 24267 22408 24268 22448
rect 24308 22408 24309 22448
rect 24267 22399 24309 22408
rect 29355 22448 29397 22457
rect 29355 22408 29356 22448
rect 29396 22408 29397 22448
rect 29355 22399 29397 22408
rect 2379 22364 2421 22373
rect 3754 22364 3812 22365
rect 2379 22324 2380 22364
rect 2420 22324 2421 22364
rect 2379 22315 2421 22324
rect 2610 22355 2656 22364
rect 2610 22315 2611 22355
rect 2651 22315 2656 22355
rect 3754 22324 3763 22364
rect 3803 22324 3812 22364
rect 3754 22323 3812 22324
rect 4107 22364 4149 22373
rect 5355 22364 5397 22373
rect 4107 22324 4108 22364
rect 4148 22324 4149 22364
rect 4107 22315 4149 22324
rect 4338 22355 4384 22364
rect 4338 22315 4339 22355
rect 4379 22315 4384 22355
rect 5355 22324 5356 22364
rect 5396 22324 5397 22364
rect 5355 22315 5397 22324
rect 5835 22364 5877 22373
rect 5835 22324 5836 22364
rect 5876 22324 5877 22364
rect 6795 22364 6837 22373
rect 5835 22315 5877 22324
rect 6459 22322 6501 22331
rect 2610 22306 2656 22315
rect 4338 22306 4384 22315
rect 6305 22313 6363 22314
rect 1707 22280 1749 22289
rect 1707 22240 1708 22280
rect 1748 22240 1749 22280
rect 1707 22231 1749 22240
rect 1882 22280 1940 22281
rect 1882 22240 1891 22280
rect 1931 22240 1940 22280
rect 1882 22239 1940 22240
rect 2198 22280 2240 22289
rect 2198 22240 2199 22280
rect 2239 22240 2240 22280
rect 2198 22231 2240 22240
rect 2475 22280 2517 22289
rect 2475 22240 2476 22280
rect 2516 22240 2517 22280
rect 2475 22231 2517 22240
rect 2704 22280 2762 22281
rect 2704 22240 2713 22280
rect 2753 22240 2762 22280
rect 2704 22239 2762 22240
rect 3291 22280 3349 22281
rect 3291 22240 3300 22280
rect 3340 22240 3349 22280
rect 3291 22239 3349 22240
rect 3435 22280 3477 22289
rect 3435 22240 3436 22280
rect 3476 22240 3477 22280
rect 3435 22231 3477 22240
rect 3919 22280 3977 22281
rect 3919 22240 3928 22280
rect 3968 22240 3977 22280
rect 3919 22239 3977 22240
rect 4203 22280 4245 22289
rect 4203 22240 4204 22280
rect 4244 22240 4245 22280
rect 4203 22231 4245 22240
rect 4432 22280 4490 22281
rect 4432 22240 4441 22280
rect 4481 22240 4490 22280
rect 4432 22239 4490 22240
rect 4779 22280 4821 22289
rect 4779 22240 4780 22280
rect 4820 22240 4821 22280
rect 4779 22231 4821 22240
rect 4971 22280 5013 22289
rect 4971 22240 4972 22280
rect 5012 22240 5013 22280
rect 4971 22231 5013 22240
rect 5494 22280 5536 22289
rect 5494 22240 5495 22280
rect 5535 22240 5536 22280
rect 5494 22231 5536 22240
rect 5626 22280 5684 22281
rect 5626 22240 5635 22280
rect 5675 22240 5684 22280
rect 5626 22239 5684 22240
rect 5739 22280 5781 22289
rect 5739 22240 5740 22280
rect 5780 22240 5781 22280
rect 6305 22273 6314 22313
rect 6354 22273 6363 22313
rect 6459 22282 6460 22322
rect 6500 22282 6501 22322
rect 6795 22324 6796 22364
rect 6836 22324 6837 22364
rect 6795 22315 6837 22324
rect 7834 22364 7892 22365
rect 7834 22324 7843 22364
rect 7883 22324 7892 22364
rect 7834 22323 7892 22324
rect 13690 22364 13748 22365
rect 13690 22324 13699 22364
rect 13739 22324 13748 22364
rect 13690 22323 13748 22324
rect 18442 22364 18500 22365
rect 18442 22324 18451 22364
rect 18491 22324 18500 22364
rect 18442 22323 18500 22324
rect 18987 22364 19029 22373
rect 18987 22324 18988 22364
rect 19028 22324 19029 22364
rect 11211 22313 11253 22322
rect 18987 22315 19029 22324
rect 19162 22364 19220 22365
rect 19162 22324 19171 22364
rect 19211 22324 19220 22364
rect 19162 22323 19220 22324
rect 19738 22364 19796 22365
rect 19738 22324 19747 22364
rect 19787 22324 19796 22364
rect 19738 22323 19796 22324
rect 20337 22364 20379 22373
rect 20337 22324 20338 22364
rect 20378 22324 20379 22364
rect 20337 22315 20379 22324
rect 22714 22364 22772 22365
rect 22714 22324 22723 22364
rect 22763 22324 22772 22364
rect 22714 22323 22772 22324
rect 25498 22364 25556 22365
rect 25498 22324 25507 22364
rect 25547 22324 25556 22364
rect 25498 22323 25556 22324
rect 27825 22364 27867 22373
rect 27825 22324 27826 22364
rect 27866 22324 27867 22364
rect 26506 22322 26564 22323
rect 6459 22273 6501 22282
rect 6586 22280 6644 22281
rect 6305 22272 6363 22273
rect 5739 22231 5781 22240
rect 6586 22240 6595 22280
rect 6635 22240 6644 22280
rect 6586 22239 6644 22240
rect 6699 22280 6741 22289
rect 6699 22240 6700 22280
rect 6740 22240 6741 22280
rect 6699 22231 6741 22240
rect 7264 22280 7306 22289
rect 7264 22240 7265 22280
rect 7305 22240 7306 22280
rect 7264 22231 7306 22240
rect 7555 22280 7613 22281
rect 7555 22240 7564 22280
rect 7604 22240 7613 22280
rect 7555 22239 7613 22240
rect 7702 22280 7744 22289
rect 7702 22240 7703 22280
rect 7743 22240 7744 22280
rect 7702 22231 7744 22240
rect 7947 22280 7989 22289
rect 7947 22240 7948 22280
rect 7988 22240 7989 22280
rect 7947 22231 7989 22240
rect 8515 22280 8573 22281
rect 8515 22240 8524 22280
rect 8564 22240 8573 22280
rect 8515 22239 8573 22240
rect 9658 22280 9716 22281
rect 9658 22240 9667 22280
rect 9707 22240 9716 22280
rect 9658 22239 9716 22240
rect 9963 22280 10005 22289
rect 9963 22240 9964 22280
rect 10004 22240 10005 22280
rect 9963 22231 10005 22240
rect 10153 22280 10195 22289
rect 10153 22240 10154 22280
rect 10194 22240 10195 22280
rect 10153 22231 10195 22240
rect 10445 22280 10487 22289
rect 10445 22240 10446 22280
rect 10486 22240 10487 22280
rect 10445 22231 10487 22240
rect 10827 22280 10869 22289
rect 10827 22240 10828 22280
rect 10868 22240 10869 22280
rect 10827 22231 10869 22240
rect 10980 22280 11038 22281
rect 10980 22240 10989 22280
rect 11029 22240 11038 22280
rect 10980 22239 11038 22240
rect 11098 22280 11156 22281
rect 11098 22240 11107 22280
rect 11147 22240 11156 22280
rect 11211 22273 11212 22313
rect 11252 22273 11253 22313
rect 22239 22313 22281 22322
rect 11211 22264 11253 22273
rect 11595 22280 11637 22289
rect 11098 22239 11156 22240
rect 11595 22240 11596 22280
rect 11636 22240 11637 22280
rect 11595 22231 11637 22240
rect 11787 22280 11829 22289
rect 11787 22240 11788 22280
rect 11828 22240 11829 22280
rect 11787 22231 11829 22240
rect 12271 22280 12329 22281
rect 12271 22240 12280 22280
rect 12320 22240 12329 22280
rect 12271 22239 12329 22240
rect 13323 22280 13365 22289
rect 13323 22240 13324 22280
rect 13364 22240 13365 22280
rect 13323 22231 13365 22240
rect 13803 22280 13845 22289
rect 13803 22240 13804 22280
rect 13844 22240 13845 22280
rect 13803 22231 13845 22240
rect 13995 22280 14037 22289
rect 13995 22240 13996 22280
rect 14036 22240 14037 22280
rect 13995 22231 14037 22240
rect 15147 22280 15189 22289
rect 15147 22240 15148 22280
rect 15188 22240 15189 22280
rect 15147 22231 15189 22240
rect 15723 22280 15765 22289
rect 15723 22240 15724 22280
rect 15764 22240 15765 22280
rect 15723 22231 15765 22240
rect 15811 22280 15869 22281
rect 15811 22240 15820 22280
rect 15860 22240 15869 22280
rect 15811 22239 15869 22240
rect 17067 22280 17109 22289
rect 17067 22240 17068 22280
rect 17108 22240 17109 22280
rect 17067 22231 17109 22240
rect 18027 22280 18069 22289
rect 18027 22240 18028 22280
rect 18068 22240 18069 22280
rect 18027 22231 18069 22240
rect 18146 22280 18188 22289
rect 18146 22240 18147 22280
rect 18187 22240 18188 22280
rect 18146 22231 18188 22240
rect 18256 22280 18314 22281
rect 18256 22240 18265 22280
rect 18305 22240 18314 22280
rect 18256 22239 18314 22240
rect 18586 22280 18644 22281
rect 18586 22240 18595 22280
rect 18635 22240 18644 22280
rect 18586 22239 18644 22240
rect 19546 22280 19604 22281
rect 19546 22240 19555 22280
rect 19595 22240 19604 22280
rect 19546 22239 19604 22240
rect 20427 22280 20469 22289
rect 20427 22240 20428 22280
rect 20468 22240 20469 22280
rect 20427 22231 20469 22240
rect 21180 22280 21222 22289
rect 21180 22240 21181 22280
rect 21221 22240 21222 22280
rect 21180 22231 21222 22240
rect 21291 22280 21333 22289
rect 21291 22240 21292 22280
rect 21332 22240 21333 22280
rect 22239 22273 22240 22313
rect 22280 22273 22281 22313
rect 22239 22264 22281 22273
rect 22330 22280 22388 22281
rect 21291 22231 21333 22240
rect 22330 22240 22339 22280
rect 22379 22240 22388 22280
rect 22330 22239 22388 22240
rect 22594 22280 22652 22281
rect 22594 22240 22603 22280
rect 22643 22240 22652 22280
rect 22594 22239 22652 22240
rect 22827 22280 22869 22289
rect 22827 22240 22828 22280
rect 22868 22240 22869 22280
rect 22827 22231 22869 22240
rect 23098 22280 23140 22289
rect 23098 22240 23099 22280
rect 23139 22240 23140 22280
rect 23098 22231 23140 22240
rect 23307 22280 23349 22289
rect 23307 22240 23308 22280
rect 23348 22240 23349 22280
rect 23307 22231 23349 22240
rect 23674 22280 23732 22281
rect 23674 22240 23683 22280
rect 23723 22240 23732 22280
rect 23674 22239 23732 22240
rect 23787 22280 23829 22289
rect 23787 22240 23788 22280
rect 23828 22240 23829 22280
rect 23787 22231 23829 22240
rect 24267 22280 24309 22289
rect 24267 22240 24268 22280
rect 24308 22240 24309 22280
rect 24267 22231 24309 22240
rect 24457 22280 24499 22289
rect 24457 22240 24458 22280
rect 24498 22240 24499 22280
rect 24457 22231 24499 22240
rect 24641 22280 24683 22289
rect 24641 22240 24642 22280
rect 24682 22240 24683 22280
rect 24641 22231 24683 22240
rect 24826 22280 24884 22281
rect 24826 22240 24835 22280
rect 24875 22240 24884 22280
rect 24826 22239 24884 22240
rect 24939 22280 24981 22289
rect 24939 22240 24940 22280
rect 24980 22240 24981 22280
rect 24939 22231 24981 22240
rect 25378 22280 25436 22281
rect 25378 22240 25387 22280
rect 25427 22240 25436 22280
rect 25378 22239 25436 22240
rect 25611 22280 25653 22289
rect 25611 22240 25612 22280
rect 25652 22240 25653 22280
rect 25611 22231 25653 22240
rect 25942 22280 25984 22289
rect 25942 22240 25943 22280
rect 25983 22240 25984 22280
rect 25942 22231 25984 22240
rect 26038 22280 26096 22281
rect 26038 22240 26047 22280
rect 26087 22240 26096 22280
rect 26038 22239 26096 22240
rect 26187 22280 26229 22289
rect 26187 22240 26188 22280
rect 26228 22240 26229 22280
rect 26187 22231 26229 22240
rect 26376 22280 26418 22289
rect 26506 22282 26515 22322
rect 26555 22282 26564 22322
rect 27825 22315 27867 22324
rect 31258 22364 31316 22365
rect 31258 22324 31267 22364
rect 31307 22324 31316 22364
rect 31258 22323 31316 22324
rect 26506 22281 26564 22282
rect 26376 22240 26377 22280
rect 26417 22240 26418 22280
rect 26376 22231 26418 22240
rect 26620 22280 26678 22281
rect 26620 22240 26629 22280
rect 26669 22240 26678 22280
rect 26620 22239 26678 22240
rect 26842 22280 26900 22281
rect 26842 22240 26851 22280
rect 26891 22240 26900 22280
rect 26842 22239 26900 22240
rect 27147 22280 27189 22289
rect 27147 22240 27148 22280
rect 27188 22240 27189 22280
rect 27147 22231 27189 22240
rect 27435 22280 27477 22289
rect 27435 22240 27436 22280
rect 27476 22240 27477 22280
rect 27435 22231 27477 22240
rect 27915 22280 27957 22289
rect 27915 22240 27916 22280
rect 27956 22240 27957 22280
rect 27915 22231 27957 22240
rect 28687 22280 28745 22281
rect 28687 22240 28696 22280
rect 28736 22240 28745 22280
rect 28687 22239 28745 22240
rect 30874 22280 30932 22281
rect 30874 22240 30883 22280
rect 30923 22240 30932 22280
rect 30874 22239 30932 22240
rect 730 22196 788 22197
rect 730 22156 739 22196
rect 779 22156 788 22196
rect 730 22155 788 22156
rect 2091 22196 2133 22205
rect 2091 22156 2092 22196
rect 2132 22156 2133 22196
rect 2091 22147 2133 22156
rect 4875 22196 4917 22205
rect 4875 22156 4876 22196
rect 4916 22156 4917 22196
rect 4875 22147 4917 22156
rect 6016 22196 6058 22205
rect 6016 22156 6017 22196
rect 6057 22156 6058 22196
rect 6016 22147 6058 22156
rect 7467 22196 7509 22205
rect 7467 22156 7468 22196
rect 7508 22156 7509 22196
rect 7467 22147 7509 22156
rect 8221 22196 8263 22205
rect 8221 22156 8222 22196
rect 8262 22156 8263 22196
rect 8221 22147 8263 22156
rect 8427 22196 8469 22205
rect 8427 22156 8428 22196
rect 8468 22156 8469 22196
rect 8427 22147 8469 22156
rect 15517 22196 15559 22205
rect 15517 22156 15518 22196
rect 15558 22156 15559 22196
rect 15517 22147 15559 22156
rect 23211 22196 23253 22205
rect 23211 22156 23212 22196
rect 23252 22156 23253 22196
rect 23211 22147 23253 22156
rect 24730 22196 24788 22197
rect 24730 22156 24739 22196
rect 24779 22156 24788 22196
rect 24730 22155 24788 22156
rect 28522 22196 28580 22197
rect 28522 22156 28531 22196
rect 28571 22156 28580 22196
rect 28522 22155 28580 22156
rect 1978 22112 2036 22113
rect 1978 22072 1987 22112
rect 2027 22072 2036 22112
rect 1978 22071 2036 22072
rect 3130 22112 3188 22113
rect 3130 22072 3139 22112
rect 3179 22072 3188 22112
rect 3130 22071 3188 22072
rect 5115 22112 5157 22121
rect 5115 22072 5116 22112
rect 5156 22072 5157 22112
rect 5115 22063 5157 22072
rect 6219 22112 6261 22121
rect 6219 22072 6220 22112
rect 6260 22072 6261 22112
rect 6219 22063 6261 22072
rect 8026 22112 8084 22113
rect 8026 22072 8035 22112
rect 8075 22072 8084 22112
rect 8026 22071 8084 22072
rect 8314 22112 8372 22113
rect 8314 22072 8323 22112
rect 8363 22072 8372 22112
rect 8314 22071 8372 22072
rect 10059 22112 10101 22121
rect 10059 22072 10060 22112
rect 10100 22072 10101 22112
rect 10059 22063 10101 22072
rect 10330 22112 10388 22113
rect 10330 22072 10339 22112
rect 10379 22072 10388 22112
rect 10330 22071 10388 22072
rect 12106 22112 12164 22113
rect 12106 22072 12115 22112
rect 12155 22072 12164 22112
rect 12106 22071 12164 22072
rect 12730 22112 12788 22113
rect 12730 22072 12739 22112
rect 12779 22072 12788 22112
rect 12730 22071 12788 22072
rect 15610 22112 15668 22113
rect 15610 22072 15619 22112
rect 15659 22072 15668 22112
rect 15610 22071 15668 22072
rect 17931 22112 17973 22121
rect 17931 22072 17932 22112
rect 17972 22072 17973 22112
rect 17931 22063 17973 22072
rect 20122 22112 20180 22113
rect 20122 22072 20131 22112
rect 20171 22072 20180 22112
rect 20122 22071 20180 22072
rect 22450 22112 22508 22113
rect 22450 22072 22459 22112
rect 22499 22072 22508 22112
rect 22450 22071 22508 22072
rect 22906 22112 22964 22113
rect 22906 22072 22915 22112
rect 22955 22072 22964 22112
rect 22906 22071 22964 22072
rect 25690 22112 25748 22113
rect 25690 22072 25699 22112
rect 25739 22072 25748 22112
rect 25690 22071 25748 22072
rect 26667 22112 26709 22121
rect 26667 22072 26668 22112
rect 26708 22072 26709 22112
rect 26667 22063 26709 22072
rect 28971 22112 29013 22121
rect 28971 22072 28972 22112
rect 29012 22072 29013 22112
rect 28971 22063 29013 22072
rect 576 21944 31392 21968
rect 576 21904 4352 21944
rect 4720 21904 12126 21944
rect 12494 21904 19900 21944
rect 20268 21904 27674 21944
rect 28042 21904 31392 21944
rect 576 21880 31392 21904
rect 1306 21776 1364 21777
rect 1306 21736 1315 21776
rect 1355 21736 1364 21776
rect 1306 21735 1364 21736
rect 3531 21776 3573 21785
rect 3531 21736 3532 21776
rect 3572 21736 3573 21776
rect 3531 21727 3573 21736
rect 5338 21776 5396 21777
rect 5338 21736 5347 21776
rect 5387 21736 5396 21776
rect 5338 21735 5396 21736
rect 5914 21776 5972 21777
rect 5914 21736 5923 21776
rect 5963 21736 5972 21776
rect 5914 21735 5972 21736
rect 6315 21776 6357 21785
rect 6315 21736 6316 21776
rect 6356 21736 6357 21776
rect 6315 21727 6357 21736
rect 6874 21776 6932 21777
rect 6874 21736 6883 21776
rect 6923 21736 6932 21776
rect 6874 21735 6932 21736
rect 7371 21776 7413 21785
rect 7371 21736 7372 21776
rect 7412 21736 7413 21776
rect 7371 21727 7413 21736
rect 8619 21776 8661 21785
rect 8619 21736 8620 21776
rect 8660 21736 8661 21776
rect 8619 21727 8661 21736
rect 9754 21776 9812 21777
rect 9754 21736 9763 21776
rect 9803 21736 9812 21776
rect 9754 21735 9812 21736
rect 10426 21776 10484 21777
rect 10426 21736 10435 21776
rect 10475 21736 10484 21776
rect 10426 21735 10484 21736
rect 10714 21776 10772 21777
rect 10714 21736 10723 21776
rect 10763 21736 10772 21776
rect 10714 21735 10772 21736
rect 11194 21776 11252 21777
rect 11194 21736 11203 21776
rect 11243 21736 11252 21776
rect 11194 21735 11252 21736
rect 13594 21776 13652 21777
rect 13594 21736 13603 21776
rect 13643 21736 13652 21776
rect 13594 21735 13652 21736
rect 15898 21776 15956 21777
rect 15898 21736 15907 21776
rect 15947 21736 15956 21776
rect 15898 21735 15956 21736
rect 22155 21776 22197 21785
rect 22155 21736 22156 21776
rect 22196 21736 22197 21776
rect 22155 21727 22197 21736
rect 23595 21776 23637 21785
rect 23595 21736 23596 21776
rect 23636 21736 23637 21776
rect 23595 21727 23637 21736
rect 24171 21776 24213 21785
rect 24171 21736 24172 21776
rect 24212 21736 24213 21776
rect 24171 21727 24213 21736
rect 25563 21776 25605 21785
rect 25563 21736 25564 21776
rect 25604 21736 25605 21776
rect 25563 21727 25605 21736
rect 26379 21776 26421 21785
rect 26379 21736 26380 21776
rect 26420 21736 26421 21776
rect 26379 21727 26421 21736
rect 27250 21776 27308 21777
rect 27250 21736 27259 21776
rect 27299 21736 27308 21776
rect 27250 21735 27308 21736
rect 27579 21776 27621 21785
rect 27579 21736 27580 21776
rect 27620 21736 27621 21776
rect 27579 21727 27621 21736
rect 28635 21776 28677 21785
rect 28635 21736 28636 21776
rect 28676 21736 28677 21776
rect 28635 21727 28677 21736
rect 2845 21692 2887 21701
rect 2845 21652 2846 21692
rect 2886 21652 2887 21692
rect 2845 21643 2887 21652
rect 3638 21692 3680 21701
rect 3638 21652 3639 21692
rect 3679 21652 3680 21692
rect 3638 21643 3680 21652
rect 4762 21692 4820 21693
rect 4762 21652 4771 21692
rect 4811 21652 4820 21692
rect 4762 21651 4820 21652
rect 6027 21692 6069 21701
rect 6027 21652 6028 21692
rect 6068 21652 6069 21692
rect 6027 21643 6069 21652
rect 6781 21692 6823 21701
rect 6781 21652 6782 21692
rect 6822 21652 6823 21692
rect 6781 21643 6823 21652
rect 7851 21692 7893 21701
rect 7851 21652 7852 21692
rect 7892 21652 7893 21692
rect 7851 21643 7893 21652
rect 8091 21692 8133 21701
rect 8091 21652 8092 21692
rect 8132 21652 8133 21692
rect 8091 21643 8133 21652
rect 9387 21692 9429 21701
rect 9387 21652 9388 21692
rect 9428 21652 9429 21692
rect 9387 21643 9429 21652
rect 10937 21692 10979 21701
rect 10937 21652 10938 21692
rect 10978 21652 10979 21692
rect 10937 21643 10979 21652
rect 11417 21692 11459 21701
rect 11417 21652 11418 21692
rect 11458 21652 11459 21692
rect 11417 21643 11459 21652
rect 11739 21692 11781 21701
rect 11739 21652 11740 21692
rect 11780 21652 11781 21692
rect 11739 21643 11781 21652
rect 14763 21692 14805 21701
rect 14763 21652 14764 21692
rect 14804 21652 14805 21692
rect 14763 21643 14805 21652
rect 16714 21692 16772 21693
rect 16714 21652 16723 21692
rect 16763 21652 16772 21692
rect 16714 21651 16772 21652
rect 18298 21692 18356 21693
rect 18298 21652 18307 21692
rect 18347 21652 18356 21692
rect 18298 21651 18356 21652
rect 26283 21692 26325 21701
rect 26283 21652 26284 21692
rect 26324 21652 26325 21692
rect 26283 21643 26325 21652
rect 27997 21692 28039 21701
rect 27997 21652 27998 21692
rect 28038 21652 28039 21692
rect 27997 21643 28039 21652
rect 28954 21692 29012 21693
rect 28954 21652 28963 21692
rect 29003 21652 29012 21692
rect 28954 21651 29012 21652
rect 1131 21608 1173 21617
rect 1131 21568 1132 21608
rect 1172 21568 1173 21608
rect 1131 21559 1173 21568
rect 1318 21608 1376 21609
rect 1318 21568 1327 21608
rect 1367 21568 1376 21608
rect 1318 21567 1376 21568
rect 1515 21608 1557 21617
rect 1515 21568 1516 21608
rect 1556 21568 1557 21608
rect 1515 21559 1557 21568
rect 1620 21608 1662 21617
rect 1620 21568 1621 21608
rect 1661 21568 1662 21608
rect 1620 21559 1662 21568
rect 1842 21608 1884 21617
rect 1842 21568 1843 21608
rect 1883 21568 1884 21608
rect 1842 21559 1884 21568
rect 2043 21608 2085 21617
rect 2043 21568 2044 21608
rect 2084 21568 2085 21608
rect 2043 21559 2085 21568
rect 3051 21608 3093 21617
rect 3322 21608 3380 21609
rect 3051 21568 3052 21608
rect 3092 21568 3093 21608
rect 3051 21559 3093 21568
rect 3147 21599 3189 21608
rect 3147 21559 3148 21599
rect 3188 21559 3189 21599
rect 3322 21568 3331 21608
rect 3371 21568 3380 21608
rect 3322 21567 3380 21568
rect 3435 21608 3477 21617
rect 4438 21608 4480 21617
rect 3435 21568 3436 21608
rect 3476 21568 3477 21608
rect 3435 21559 3477 21568
rect 4002 21599 4048 21608
rect 4002 21559 4003 21599
rect 4043 21559 4048 21599
rect 4438 21568 4439 21608
rect 4479 21568 4480 21608
rect 4438 21559 4480 21568
rect 4683 21608 4725 21617
rect 4683 21568 4684 21608
rect 4724 21568 4725 21608
rect 4683 21559 4725 21568
rect 5499 21608 5541 21617
rect 5499 21568 5500 21608
rect 5540 21568 5541 21608
rect 5499 21559 5541 21568
rect 5643 21608 5685 21617
rect 5643 21568 5644 21608
rect 5684 21568 5685 21608
rect 5643 21559 5685 21568
rect 5821 21608 5863 21617
rect 6411 21608 6453 21617
rect 5821 21568 5822 21608
rect 5862 21568 5863 21608
rect 5821 21559 5863 21568
rect 6123 21599 6165 21608
rect 6123 21559 6124 21599
rect 6164 21559 6165 21599
rect 6411 21568 6412 21608
rect 6452 21568 6453 21608
rect 6411 21559 6453 21568
rect 6628 21608 6670 21617
rect 6628 21568 6629 21608
rect 6669 21568 6670 21608
rect 6628 21559 6670 21568
rect 6987 21608 7029 21617
rect 7371 21608 7413 21617
rect 6987 21568 6988 21608
rect 7028 21568 7029 21608
rect 6987 21559 7029 21568
rect 7083 21599 7125 21608
rect 7083 21559 7084 21599
rect 7124 21559 7125 21599
rect 7371 21568 7372 21608
rect 7412 21568 7413 21608
rect 7371 21559 7413 21568
rect 7563 21608 7605 21617
rect 7563 21568 7564 21608
rect 7604 21568 7605 21608
rect 7563 21559 7605 21568
rect 7755 21608 7797 21617
rect 7755 21568 7756 21608
rect 7796 21568 7797 21608
rect 7755 21559 7797 21568
rect 7947 21608 7989 21617
rect 7947 21568 7948 21608
rect 7988 21568 7989 21608
rect 7947 21559 7989 21568
rect 8283 21608 8325 21617
rect 8283 21568 8284 21608
rect 8324 21568 8325 21608
rect 8283 21559 8325 21568
rect 8427 21608 8469 21617
rect 8427 21568 8428 21608
rect 8468 21568 8469 21608
rect 8427 21559 8469 21568
rect 8715 21608 8757 21617
rect 8715 21568 8716 21608
rect 8756 21568 8757 21608
rect 8715 21559 8757 21568
rect 8944 21608 9002 21609
rect 8944 21568 8953 21608
rect 8993 21568 9002 21608
rect 8944 21567 9002 21568
rect 9291 21608 9333 21617
rect 9291 21568 9292 21608
rect 9332 21568 9333 21608
rect 9291 21559 9333 21568
rect 9483 21608 9525 21617
rect 9483 21568 9484 21608
rect 9524 21568 9525 21608
rect 9483 21559 9525 21568
rect 9658 21608 9716 21609
rect 9658 21568 9667 21608
rect 9707 21568 9716 21608
rect 9658 21567 9716 21568
rect 9974 21608 10016 21617
rect 9974 21568 9975 21608
rect 10015 21568 10016 21608
rect 9974 21559 10016 21568
rect 10130 21608 10172 21617
rect 10130 21568 10131 21608
rect 10171 21568 10172 21608
rect 10130 21559 10172 21568
rect 10347 21608 10389 21617
rect 10347 21568 10348 21608
rect 10388 21568 10389 21608
rect 10347 21559 10389 21568
rect 10618 21608 10676 21609
rect 10618 21568 10627 21608
rect 10667 21568 10676 21608
rect 10618 21567 10676 21568
rect 11098 21608 11156 21609
rect 12202 21608 12260 21609
rect 11098 21568 11107 21608
rect 11147 21568 11156 21608
rect 11098 21567 11156 21568
rect 11586 21599 11632 21608
rect 11586 21559 11587 21599
rect 11627 21559 11632 21599
rect 12202 21568 12211 21608
rect 12251 21568 12260 21608
rect 12202 21567 12260 21568
rect 12634 21608 12692 21609
rect 12634 21568 12643 21608
rect 12683 21568 12692 21608
rect 12634 21567 12692 21568
rect 13515 21608 13557 21617
rect 13515 21568 13516 21608
rect 13556 21568 13557 21608
rect 3147 21550 3189 21559
rect 4002 21550 4048 21559
rect 6123 21550 6165 21559
rect 7083 21550 7125 21559
rect 11586 21550 11632 21559
rect 12394 21566 12452 21567
rect 843 21524 885 21533
rect 4155 21524 4197 21533
rect 843 21484 844 21524
rect 884 21484 885 21524
rect 843 21475 885 21484
rect 1746 21515 1792 21524
rect 1746 21475 1747 21515
rect 1787 21475 1792 21515
rect 4155 21484 4156 21524
rect 4196 21484 4197 21524
rect 4155 21475 4197 21484
rect 4570 21524 4628 21525
rect 4570 21484 4579 21524
rect 4619 21484 4628 21524
rect 4570 21483 4628 21484
rect 4971 21524 5013 21533
rect 4971 21484 4972 21524
rect 5012 21484 5013 21524
rect 4971 21475 5013 21484
rect 6530 21524 6572 21533
rect 6530 21484 6531 21524
rect 6571 21484 6572 21524
rect 6530 21475 6572 21484
rect 8834 21524 8876 21533
rect 12394 21526 12403 21566
rect 12443 21526 12452 21566
rect 13515 21559 13557 21568
rect 13750 21608 13792 21617
rect 13750 21568 13751 21608
rect 13791 21568 13792 21608
rect 13750 21559 13792 21568
rect 13995 21608 14037 21617
rect 13995 21568 13996 21608
rect 14036 21568 14037 21608
rect 13995 21559 14037 21568
rect 14458 21608 14516 21609
rect 14458 21568 14467 21608
rect 14507 21568 14516 21608
rect 14458 21567 14516 21568
rect 15051 21608 15093 21617
rect 15051 21568 15052 21608
rect 15092 21568 15093 21608
rect 15532 21608 15574 21617
rect 15051 21559 15093 21568
rect 15291 21566 15333 21575
rect 12394 21525 12452 21526
rect 8834 21484 8835 21524
rect 8875 21484 8876 21524
rect 8834 21475 8876 21484
rect 10234 21524 10292 21525
rect 10234 21484 10243 21524
rect 10283 21484 10292 21524
rect 10234 21483 10292 21484
rect 13882 21524 13940 21525
rect 13882 21484 13891 21524
rect 13931 21484 13940 21524
rect 13882 21483 13940 21484
rect 14091 21524 14133 21533
rect 14091 21484 14092 21524
rect 14132 21484 14133 21524
rect 14091 21475 14133 21484
rect 14283 21524 14325 21533
rect 14283 21484 14284 21524
rect 14324 21484 14325 21524
rect 14283 21475 14325 21484
rect 14859 21524 14901 21533
rect 14859 21484 14860 21524
rect 14900 21484 14901 21524
rect 15291 21526 15292 21566
rect 15332 21526 15333 21566
rect 15532 21568 15533 21608
rect 15573 21568 15574 21608
rect 15532 21559 15574 21568
rect 16186 21608 16244 21609
rect 16186 21568 16195 21608
rect 16235 21568 16244 21608
rect 16186 21567 16244 21568
rect 16879 21608 16937 21609
rect 16879 21568 16888 21608
rect 16928 21568 16937 21608
rect 16879 21567 16937 21568
rect 17067 21608 17109 21617
rect 17067 21568 17068 21608
rect 17108 21568 17109 21608
rect 17067 21559 17109 21568
rect 17259 21608 17301 21617
rect 17259 21568 17260 21608
rect 17300 21568 17301 21608
rect 17259 21559 17301 21568
rect 18586 21608 18644 21609
rect 18586 21568 18595 21608
rect 18635 21568 18644 21608
rect 18586 21567 18644 21568
rect 18987 21608 19029 21617
rect 18987 21568 18988 21608
rect 19028 21568 19029 21608
rect 18987 21559 19029 21568
rect 19179 21608 19221 21617
rect 19179 21568 19180 21608
rect 19220 21568 19221 21608
rect 19179 21559 19221 21568
rect 19755 21608 19797 21617
rect 19755 21568 19756 21608
rect 19796 21568 19797 21608
rect 19755 21559 19797 21568
rect 19984 21608 20042 21609
rect 19984 21568 19993 21608
rect 20033 21568 20042 21608
rect 19984 21567 20042 21568
rect 20331 21608 20373 21617
rect 20331 21568 20332 21608
rect 20372 21568 20373 21608
rect 20331 21559 20373 21568
rect 20715 21608 20757 21617
rect 20715 21568 20716 21608
rect 20756 21568 20757 21608
rect 20715 21559 20757 21568
rect 21099 21608 21141 21617
rect 21099 21568 21100 21608
rect 21140 21568 21141 21608
rect 21099 21559 21141 21568
rect 21483 21608 21525 21617
rect 21483 21568 21484 21608
rect 21524 21568 21525 21608
rect 21483 21559 21525 21568
rect 21670 21608 21712 21617
rect 21670 21568 21671 21608
rect 21711 21568 21712 21608
rect 21670 21559 21712 21568
rect 21867 21608 21909 21617
rect 21867 21568 21868 21608
rect 21908 21568 21909 21608
rect 21867 21559 21909 21568
rect 22059 21608 22101 21617
rect 22059 21568 22060 21608
rect 22100 21568 22101 21608
rect 22059 21559 22101 21568
rect 22234 21608 22292 21609
rect 22234 21568 22243 21608
rect 22283 21568 22292 21608
rect 22234 21567 22292 21568
rect 22714 21608 22772 21609
rect 22714 21568 22723 21608
rect 22763 21568 22772 21608
rect 22714 21567 22772 21568
rect 22827 21608 22869 21617
rect 22827 21568 22828 21608
rect 22868 21568 22869 21608
rect 22827 21559 22869 21568
rect 23403 21608 23445 21617
rect 23403 21568 23404 21608
rect 23444 21568 23445 21608
rect 23403 21559 23445 21568
rect 23595 21608 23637 21617
rect 23595 21568 23596 21608
rect 23636 21568 23637 21608
rect 23595 21559 23637 21568
rect 24154 21608 24212 21609
rect 24154 21568 24163 21608
rect 24203 21568 24212 21608
rect 24154 21567 24212 21568
rect 24267 21608 24309 21617
rect 24267 21568 24268 21608
rect 24308 21568 24309 21608
rect 24267 21559 24309 21568
rect 24598 21608 24640 21617
rect 24598 21568 24599 21608
rect 24639 21568 24640 21608
rect 24598 21559 24640 21568
rect 24843 21608 24885 21617
rect 24843 21568 24844 21608
rect 24884 21568 24885 21608
rect 24843 21559 24885 21568
rect 25130 21608 25172 21617
rect 25130 21568 25131 21608
rect 25171 21568 25172 21608
rect 25130 21559 25172 21568
rect 25306 21608 25364 21609
rect 25306 21568 25315 21608
rect 25355 21568 25364 21608
rect 25306 21567 25364 21568
rect 25419 21608 25461 21617
rect 25419 21568 25420 21608
rect 25460 21568 25461 21608
rect 25419 21559 25461 21568
rect 25707 21608 25749 21617
rect 26475 21608 26517 21617
rect 27130 21608 27188 21609
rect 28203 21608 28245 21617
rect 29338 21608 29396 21609
rect 25707 21568 25708 21608
rect 25748 21568 25749 21608
rect 25707 21559 25749 21568
rect 26178 21599 26224 21608
rect 26178 21559 26179 21599
rect 26219 21559 26224 21599
rect 26475 21568 26476 21608
rect 26516 21568 26517 21608
rect 26475 21559 26517 21568
rect 27047 21599 27089 21608
rect 27047 21559 27048 21599
rect 27088 21559 27089 21599
rect 27130 21568 27139 21608
rect 27179 21568 27188 21608
rect 27130 21567 27188 21568
rect 27426 21599 27472 21608
rect 26178 21550 26224 21559
rect 27047 21550 27089 21559
rect 27426 21559 27427 21599
rect 27467 21559 27472 21599
rect 28203 21568 28204 21608
rect 28244 21568 28245 21608
rect 28203 21559 28245 21568
rect 28299 21599 28341 21608
rect 28299 21559 28300 21599
rect 28340 21559 28341 21599
rect 27426 21550 27472 21559
rect 28299 21550 28341 21559
rect 28482 21599 28528 21608
rect 28482 21559 28483 21599
rect 28523 21559 28528 21599
rect 29338 21568 29347 21608
rect 29387 21568 29396 21608
rect 29338 21567 29396 21568
rect 28482 21550 28528 21559
rect 15291 21517 15333 21526
rect 15418 21524 15476 21525
rect 14859 21475 14901 21484
rect 15418 21484 15427 21524
rect 15467 21484 15476 21524
rect 15418 21483 15476 21484
rect 15627 21524 15669 21533
rect 15627 21484 15628 21524
rect 15668 21484 15669 21524
rect 15627 21475 15669 21484
rect 15802 21524 15860 21525
rect 15802 21484 15811 21524
rect 15851 21484 15860 21524
rect 15802 21483 15860 21484
rect 16378 21524 16436 21525
rect 16378 21484 16387 21524
rect 16427 21484 16436 21524
rect 16378 21483 16436 21484
rect 18202 21524 18260 21525
rect 18202 21484 18211 21524
rect 18251 21484 18260 21524
rect 18202 21483 18260 21484
rect 18778 21524 18836 21525
rect 18778 21484 18787 21524
rect 18827 21484 18836 21524
rect 18778 21483 18836 21484
rect 19659 21524 19701 21533
rect 24730 21524 24788 21525
rect 19659 21484 19660 21524
rect 19700 21484 19701 21524
rect 19659 21475 19701 21484
rect 19890 21515 19936 21524
rect 19890 21475 19891 21515
rect 19931 21475 19936 21515
rect 24730 21484 24739 21524
rect 24779 21484 24788 21524
rect 24730 21483 24788 21484
rect 24939 21524 24981 21533
rect 24939 21484 24940 21524
rect 24980 21484 24981 21524
rect 24939 21475 24981 21484
rect 1746 21466 1792 21475
rect 19890 21466 19936 21475
rect 5211 21440 5253 21449
rect 5211 21400 5212 21440
rect 5252 21400 5253 21440
rect 5211 21391 5253 21400
rect 12843 21440 12885 21449
rect 12843 21400 12844 21440
rect 12884 21400 12885 21440
rect 12843 21391 12885 21400
rect 17643 21440 17685 21449
rect 17643 21400 17644 21440
rect 17684 21400 17685 21440
rect 17643 21391 17685 21400
rect 18027 21440 18069 21449
rect 18027 21400 18028 21440
rect 18068 21400 18069 21440
rect 18027 21391 18069 21400
rect 20091 21440 20133 21449
rect 20091 21400 20092 21440
rect 20132 21400 20133 21440
rect 20091 21391 20133 21400
rect 20859 21440 20901 21449
rect 20859 21400 20860 21440
rect 20900 21400 20901 21440
rect 20859 21391 20901 21400
rect 23386 21440 23444 21441
rect 23386 21400 23395 21440
rect 23435 21400 23444 21440
rect 23386 21399 23444 21400
rect 25419 21440 25461 21449
rect 25419 21400 25420 21440
rect 25460 21400 25461 21440
rect 25419 21391 25461 21400
rect 603 21356 645 21365
rect 603 21316 604 21356
rect 644 21316 645 21356
rect 603 21307 645 21316
rect 2667 21356 2709 21365
rect 2667 21316 2668 21356
rect 2708 21316 2709 21356
rect 2667 21307 2709 21316
rect 2842 21356 2900 21357
rect 2842 21316 2851 21356
rect 2891 21316 2900 21356
rect 2842 21315 2900 21316
rect 7851 21356 7893 21365
rect 7851 21316 7852 21356
rect 7892 21316 7893 21356
rect 7851 21307 7893 21316
rect 9963 21356 10005 21365
rect 9963 21316 9964 21356
rect 10004 21316 10005 21356
rect 9963 21307 10005 21316
rect 10923 21356 10965 21365
rect 10923 21316 10924 21356
rect 10964 21316 10965 21356
rect 10923 21307 10965 21316
rect 11403 21356 11445 21365
rect 11403 21316 11404 21356
rect 11444 21316 11445 21356
rect 11403 21307 11445 21316
rect 13035 21356 13077 21365
rect 13035 21316 13036 21356
rect 13076 21316 13077 21356
rect 13035 21307 13077 21316
rect 13323 21356 13365 21365
rect 13323 21316 13324 21356
rect 13364 21316 13365 21356
rect 13323 21307 13365 21316
rect 15195 21356 15237 21365
rect 15195 21316 15196 21356
rect 15236 21316 15237 21356
rect 15195 21307 15237 21316
rect 17163 21356 17205 21365
rect 17163 21316 17164 21356
rect 17204 21316 17205 21356
rect 17163 21307 17205 21316
rect 18987 21356 19029 21365
rect 18987 21316 18988 21356
rect 19028 21316 19029 21356
rect 18987 21307 19029 21316
rect 21771 21356 21813 21365
rect 21771 21316 21772 21356
rect 21812 21316 21813 21356
rect 21771 21307 21813 21316
rect 23002 21356 23060 21357
rect 23002 21316 23011 21356
rect 23051 21316 23060 21356
rect 23002 21315 23060 21316
rect 24459 21356 24501 21365
rect 24459 21316 24460 21356
rect 24500 21316 24501 21356
rect 24459 21307 24501 21316
rect 25995 21356 26037 21365
rect 25995 21316 25996 21356
rect 26036 21316 26037 21356
rect 25995 21307 26037 21316
rect 26746 21356 26804 21357
rect 26746 21316 26755 21356
rect 26795 21316 26804 21356
rect 26746 21315 26804 21316
rect 27994 21356 28052 21357
rect 27994 21316 28003 21356
rect 28043 21316 28052 21356
rect 27994 21315 28052 21316
rect 31275 21356 31317 21365
rect 31275 21316 31276 21356
rect 31316 21316 31317 21356
rect 31275 21307 31317 21316
rect 576 21188 31392 21212
rect 576 21148 3112 21188
rect 3480 21148 10886 21188
rect 11254 21148 18660 21188
rect 19028 21148 26434 21188
rect 26802 21148 31392 21188
rect 576 21124 31392 21148
rect 603 21020 645 21029
rect 603 20980 604 21020
rect 644 20980 645 21020
rect 603 20971 645 20980
rect 1227 21020 1269 21029
rect 1227 20980 1228 21020
rect 1268 20980 1269 21020
rect 1227 20971 1269 20980
rect 3531 21020 3573 21029
rect 3531 20980 3532 21020
rect 3572 20980 3573 21020
rect 3531 20971 3573 20980
rect 4954 21020 5012 21021
rect 4954 20980 4963 21020
rect 5003 20980 5012 21020
rect 4954 20979 5012 20980
rect 7371 21020 7413 21029
rect 7371 20980 7372 21020
rect 7412 20980 7413 21020
rect 7371 20971 7413 20980
rect 7947 21020 7989 21029
rect 7947 20980 7948 21020
rect 7988 20980 7989 21020
rect 7947 20971 7989 20980
rect 9051 21020 9093 21029
rect 9051 20980 9052 21020
rect 9092 20980 9093 21020
rect 9051 20971 9093 20980
rect 13083 21020 13125 21029
rect 13083 20980 13084 21020
rect 13124 20980 13125 21020
rect 13083 20971 13125 20980
rect 14362 21020 14420 21021
rect 14362 20980 14371 21020
rect 14411 20980 14420 21020
rect 14362 20979 14420 20980
rect 15627 21020 15669 21029
rect 15627 20980 15628 21020
rect 15668 20980 15669 21020
rect 15627 20971 15669 20980
rect 17146 21020 17204 21021
rect 17146 20980 17155 21020
rect 17195 20980 17204 21020
rect 17146 20979 17204 20980
rect 20506 21020 20564 21021
rect 20506 20980 20515 21020
rect 20555 20980 20564 21020
rect 20506 20979 20564 20980
rect 21291 21020 21333 21029
rect 21291 20980 21292 21020
rect 21332 20980 21333 21020
rect 21291 20971 21333 20980
rect 24442 21020 24500 21021
rect 24442 20980 24451 21020
rect 24491 20980 24500 21020
rect 24442 20979 24500 20980
rect 25803 21020 25845 21029
rect 25803 20980 25804 21020
rect 25844 20980 25845 21020
rect 25803 20971 25845 20980
rect 26379 21020 26421 21029
rect 26379 20980 26380 21020
rect 26420 20980 26421 21020
rect 26379 20971 26421 20980
rect 27706 21020 27764 21021
rect 27706 20980 27715 21020
rect 27755 20980 27764 21020
rect 27706 20979 27764 20980
rect 29835 21020 29877 21029
rect 29835 20980 29836 21020
rect 29876 20980 29877 21020
rect 29835 20971 29877 20980
rect 21867 20936 21909 20945
rect 21867 20896 21868 20936
rect 21908 20896 21909 20936
rect 21867 20887 21909 20896
rect 843 20852 885 20861
rect 843 20812 844 20852
rect 884 20812 885 20852
rect 843 20803 885 20812
rect 3915 20852 3957 20861
rect 5163 20852 5205 20861
rect 3915 20812 3916 20852
rect 3956 20812 3957 20852
rect 3915 20803 3957 20812
rect 4338 20843 4384 20852
rect 4338 20803 4339 20843
rect 4379 20803 4384 20843
rect 5163 20812 5164 20852
rect 5204 20812 5205 20852
rect 5163 20803 5205 20812
rect 6843 20852 6885 20861
rect 6843 20812 6844 20852
rect 6884 20812 6885 20852
rect 6843 20803 6885 20812
rect 7083 20852 7125 20861
rect 7083 20812 7084 20852
rect 7124 20812 7125 20852
rect 7083 20803 7125 20812
rect 8139 20852 8181 20861
rect 8139 20812 8140 20852
rect 8180 20812 8181 20852
rect 8139 20803 8181 20812
rect 8354 20852 8396 20861
rect 8354 20812 8355 20852
rect 8395 20812 8396 20852
rect 8354 20803 8396 20812
rect 8619 20852 8661 20861
rect 8619 20812 8620 20852
rect 8660 20812 8661 20852
rect 8619 20803 8661 20812
rect 9291 20852 9333 20861
rect 9291 20812 9292 20852
rect 9332 20812 9333 20852
rect 9291 20803 9333 20812
rect 14938 20852 14996 20853
rect 14938 20812 14947 20852
rect 14987 20812 14996 20852
rect 14938 20811 14996 20812
rect 19258 20852 19316 20853
rect 19258 20812 19267 20852
rect 19307 20812 19316 20852
rect 19258 20811 19316 20812
rect 19467 20852 19509 20861
rect 19467 20812 19468 20852
rect 19508 20812 19509 20852
rect 11050 20810 11108 20811
rect 4338 20794 4384 20803
rect 1131 20768 1173 20777
rect 1131 20728 1132 20768
rect 1172 20728 1173 20768
rect 1131 20719 1173 20728
rect 1323 20768 1365 20777
rect 1323 20728 1324 20768
rect 1364 20728 1365 20768
rect 1323 20719 1365 20728
rect 1515 20768 1557 20777
rect 1515 20728 1516 20768
rect 1556 20728 1557 20768
rect 1515 20719 1557 20728
rect 1707 20773 1749 20782
rect 1707 20733 1708 20773
rect 1748 20733 1749 20773
rect 1707 20724 1749 20733
rect 1899 20768 1941 20777
rect 1899 20728 1900 20768
rect 1940 20728 1941 20768
rect 1899 20719 1941 20728
rect 2091 20768 2133 20777
rect 2091 20728 2092 20768
rect 2132 20728 2133 20768
rect 2091 20719 2133 20728
rect 2565 20768 2623 20769
rect 2565 20728 2574 20768
rect 2614 20728 2623 20768
rect 2565 20727 2623 20728
rect 3082 20768 3140 20769
rect 3082 20728 3091 20768
rect 3131 20728 3140 20768
rect 3082 20727 3140 20728
rect 3226 20768 3284 20769
rect 3226 20728 3235 20768
rect 3275 20728 3284 20768
rect 3226 20727 3284 20728
rect 4203 20768 4245 20777
rect 4203 20728 4204 20768
rect 4244 20728 4245 20768
rect 4203 20719 4245 20728
rect 4432 20768 4490 20769
rect 4432 20728 4441 20768
rect 4481 20728 4490 20768
rect 4432 20727 4490 20728
rect 4779 20768 4821 20777
rect 4779 20728 4780 20768
rect 4820 20728 4821 20768
rect 4779 20719 4821 20728
rect 4954 20768 5012 20769
rect 4954 20728 4963 20768
rect 5003 20728 5012 20768
rect 4954 20727 5012 20728
rect 5259 20768 5301 20777
rect 5259 20728 5260 20768
rect 5300 20728 5301 20768
rect 5259 20719 5301 20728
rect 5378 20768 5420 20777
rect 5378 20728 5379 20768
rect 5419 20728 5420 20768
rect 5378 20719 5420 20728
rect 5488 20768 5546 20769
rect 5488 20728 5497 20768
rect 5537 20728 5546 20768
rect 5488 20727 5546 20728
rect 5643 20768 5685 20777
rect 5643 20728 5644 20768
rect 5684 20728 5685 20768
rect 5643 20719 5685 20728
rect 5818 20768 5876 20769
rect 5818 20728 5827 20768
rect 5867 20728 5876 20768
rect 5818 20727 5876 20728
rect 6028 20768 6070 20777
rect 6028 20728 6029 20768
rect 6069 20728 6070 20768
rect 6028 20719 6070 20728
rect 6217 20768 6259 20777
rect 6217 20728 6218 20768
rect 6258 20728 6259 20768
rect 6217 20719 6259 20728
rect 6411 20768 6453 20777
rect 6411 20728 6412 20768
rect 6452 20728 6453 20768
rect 6411 20719 6453 20728
rect 6603 20768 6645 20777
rect 6603 20728 6604 20768
rect 6644 20728 6645 20768
rect 6603 20719 6645 20728
rect 7275 20768 7317 20777
rect 7275 20728 7276 20768
rect 7316 20728 7317 20768
rect 7275 20719 7317 20728
rect 7466 20768 7508 20777
rect 7466 20728 7467 20768
rect 7507 20728 7508 20768
rect 7466 20719 7508 20728
rect 7642 20768 7700 20769
rect 7642 20728 7651 20768
rect 7691 20728 7700 20768
rect 7642 20727 7700 20728
rect 8235 20768 8277 20777
rect 8235 20728 8236 20768
rect 8276 20728 8277 20768
rect 8235 20719 8277 20728
rect 8464 20768 8522 20769
rect 8464 20728 8473 20768
rect 8513 20728 8522 20768
rect 8464 20727 8522 20728
rect 8715 20768 8757 20777
rect 8944 20768 9002 20769
rect 8715 20728 8716 20768
rect 8756 20728 8757 20768
rect 8715 20719 8757 20728
rect 8850 20759 8896 20768
rect 8850 20719 8851 20759
rect 8891 20719 8896 20759
rect 8944 20728 8953 20768
rect 8993 20728 9002 20768
rect 8944 20727 9002 20728
rect 9579 20768 9621 20777
rect 11050 20770 11059 20810
rect 11099 20770 11108 20810
rect 19467 20803 19509 20812
rect 19947 20852 19989 20861
rect 19947 20812 19948 20852
rect 19988 20812 19989 20852
rect 19947 20803 19989 20812
rect 24730 20852 24788 20853
rect 24730 20812 24739 20852
rect 24779 20812 24788 20852
rect 24730 20811 24788 20812
rect 25306 20852 25364 20853
rect 25306 20812 25315 20852
rect 25355 20812 25364 20852
rect 25306 20811 25364 20812
rect 28954 20852 29012 20853
rect 28954 20812 28963 20852
rect 29003 20812 29012 20852
rect 28954 20811 29012 20812
rect 11050 20769 11108 20770
rect 9579 20728 9580 20768
rect 9620 20728 9621 20768
rect 9579 20719 9621 20728
rect 9754 20768 9812 20769
rect 9754 20728 9763 20768
rect 9803 20728 9812 20768
rect 9754 20727 9812 20728
rect 10243 20768 10301 20769
rect 10243 20728 10252 20768
rect 10292 20728 10301 20768
rect 10243 20727 10301 20728
rect 11533 20768 11591 20769
rect 11533 20728 11542 20768
rect 11582 20728 11591 20768
rect 11533 20727 11591 20728
rect 11674 20768 11732 20769
rect 11674 20728 11683 20768
rect 11723 20728 11732 20768
rect 11674 20727 11732 20728
rect 12363 20768 12405 20777
rect 12363 20728 12364 20768
rect 12404 20728 12405 20768
rect 12363 20719 12405 20728
rect 12651 20768 12693 20777
rect 12651 20728 12652 20768
rect 12692 20728 12693 20768
rect 12651 20719 12693 20728
rect 12843 20768 12885 20777
rect 12843 20728 12844 20768
rect 12884 20728 12885 20768
rect 12843 20719 12885 20728
rect 13227 20768 13269 20777
rect 13227 20728 13228 20768
rect 13268 20728 13269 20768
rect 13227 20719 13269 20728
rect 13741 20768 13799 20769
rect 13741 20728 13750 20768
rect 13790 20728 13799 20768
rect 13741 20727 13799 20728
rect 14043 20768 14101 20769
rect 14043 20728 14052 20768
rect 14092 20728 14101 20768
rect 14043 20727 14101 20728
rect 14187 20768 14229 20777
rect 14187 20728 14188 20768
rect 14228 20728 14229 20768
rect 14187 20719 14229 20728
rect 14571 20768 14613 20777
rect 14571 20728 14572 20768
rect 14612 20728 14613 20768
rect 14571 20719 14613 20728
rect 14659 20768 14717 20769
rect 14659 20728 14668 20768
rect 14708 20728 14717 20768
rect 14659 20727 14717 20728
rect 14818 20768 14876 20769
rect 14818 20728 14827 20768
rect 14867 20728 14876 20768
rect 14818 20727 14876 20728
rect 15051 20768 15093 20777
rect 15051 20728 15052 20768
rect 15092 20728 15093 20768
rect 15051 20719 15093 20728
rect 15322 20768 15380 20769
rect 15322 20728 15331 20768
rect 15371 20728 15380 20768
rect 15322 20727 15380 20728
rect 16141 20768 16199 20769
rect 16141 20728 16150 20768
rect 16190 20728 16199 20768
rect 16141 20727 16199 20728
rect 16779 20768 16821 20777
rect 17355 20768 17397 20777
rect 16779 20728 16780 20768
rect 16820 20728 16821 20768
rect 16779 20719 16821 20728
rect 17058 20759 17104 20768
rect 17058 20719 17059 20759
rect 17099 20719 17104 20759
rect 17355 20728 17356 20768
rect 17396 20728 17397 20768
rect 17355 20719 17397 20728
rect 17686 20768 17728 20777
rect 17686 20728 17687 20768
rect 17727 20728 17728 20768
rect 17686 20719 17728 20728
rect 17818 20768 17876 20769
rect 17818 20728 17827 20768
rect 17867 20728 17876 20768
rect 17818 20727 17876 20728
rect 17931 20768 17973 20777
rect 17931 20728 17932 20768
rect 17972 20728 17973 20768
rect 17931 20719 17973 20728
rect 18202 20768 18260 20769
rect 18202 20728 18211 20768
rect 18251 20728 18260 20768
rect 18202 20727 18260 20728
rect 18521 20768 18563 20777
rect 18521 20728 18522 20768
rect 18562 20728 18563 20768
rect 18521 20719 18563 20728
rect 18699 20768 18741 20777
rect 18699 20728 18700 20768
rect 18740 20728 18741 20768
rect 18699 20719 18741 20728
rect 18838 20768 18880 20777
rect 18838 20728 18839 20768
rect 18879 20728 18880 20768
rect 18838 20719 18880 20728
rect 19126 20768 19168 20777
rect 19126 20728 19127 20768
rect 19167 20728 19168 20768
rect 19126 20719 19168 20728
rect 19352 20768 19394 20777
rect 19352 20728 19353 20768
rect 19393 20728 19394 20768
rect 19352 20719 19394 20728
rect 19606 20768 19648 20777
rect 19606 20728 19607 20768
rect 19647 20728 19648 20768
rect 19606 20719 19648 20728
rect 19738 20768 19796 20769
rect 19738 20728 19747 20768
rect 19787 20728 19796 20768
rect 19738 20727 19796 20728
rect 19851 20768 19893 20777
rect 19851 20728 19852 20768
rect 19892 20728 19893 20768
rect 19851 20719 19893 20728
rect 20907 20768 20949 20777
rect 20907 20728 20908 20768
rect 20948 20728 20949 20768
rect 20907 20719 20949 20728
rect 21291 20768 21333 20777
rect 21291 20728 21292 20768
rect 21332 20728 21333 20768
rect 21291 20719 21333 20728
rect 21483 20768 21525 20777
rect 21483 20728 21484 20768
rect 21524 20728 21525 20768
rect 21483 20719 21525 20728
rect 22155 20768 22197 20777
rect 22155 20728 22156 20768
rect 22196 20728 22197 20768
rect 22155 20719 22197 20728
rect 23098 20768 23156 20769
rect 23098 20728 23107 20768
rect 23147 20728 23156 20768
rect 23098 20727 23156 20728
rect 24154 20768 24212 20769
rect 24154 20728 24163 20768
rect 24203 20728 24212 20768
rect 24154 20727 24212 20728
rect 24261 20768 24319 20769
rect 24261 20728 24270 20768
rect 24310 20728 24319 20768
rect 24261 20727 24319 20728
rect 25114 20768 25172 20769
rect 25114 20728 25123 20768
rect 25163 20728 25172 20768
rect 25114 20727 25172 20728
rect 25611 20768 25653 20777
rect 25611 20728 25612 20768
rect 25652 20728 25653 20768
rect 25611 20719 25653 20728
rect 26091 20768 26133 20777
rect 26091 20728 26092 20768
rect 26132 20728 26133 20768
rect 26091 20719 26133 20728
rect 26266 20768 26324 20769
rect 26266 20728 26275 20768
rect 26315 20728 26324 20768
rect 26266 20727 26324 20728
rect 26379 20768 26421 20777
rect 26379 20728 26380 20768
rect 26420 20728 26421 20768
rect 26379 20719 26421 20728
rect 26650 20768 26708 20769
rect 26650 20728 26659 20768
rect 26699 20728 26708 20768
rect 26650 20727 26708 20728
rect 26966 20768 27008 20777
rect 26966 20728 26967 20768
rect 27007 20728 27008 20768
rect 26966 20719 27008 20728
rect 27147 20768 27189 20777
rect 27147 20728 27148 20768
rect 27188 20728 27189 20768
rect 27147 20719 27189 20728
rect 27281 20768 27339 20769
rect 27915 20768 27957 20777
rect 27281 20728 27290 20768
rect 27330 20728 27339 20768
rect 27281 20727 27339 20728
rect 27618 20759 27664 20768
rect 27618 20719 27619 20759
rect 27659 20719 27664 20759
rect 27915 20728 27916 20768
rect 27956 20728 27957 20768
rect 27915 20719 27957 20728
rect 28378 20768 28436 20769
rect 28378 20728 28387 20768
rect 28427 20728 28436 20768
rect 28378 20727 28436 20728
rect 28491 20768 28533 20777
rect 28491 20728 28492 20768
rect 28532 20728 28533 20768
rect 28491 20719 28533 20728
rect 29643 20768 29685 20777
rect 29643 20728 29644 20768
rect 29684 20728 29685 20768
rect 29643 20719 29685 20728
rect 30507 20768 30549 20777
rect 30507 20728 30508 20768
rect 30548 20728 30549 20768
rect 30507 20719 30549 20728
rect 30891 20768 30933 20777
rect 30891 20728 30892 20768
rect 30932 20728 30933 20768
rect 30891 20719 30933 20728
rect 31179 20768 31221 20777
rect 31179 20728 31180 20768
rect 31220 20728 31221 20768
rect 31179 20719 31221 20728
rect 8850 20710 8896 20719
rect 17058 20710 17104 20719
rect 27618 20710 27664 20719
rect 1611 20684 1653 20693
rect 1611 20644 1612 20684
rect 1652 20644 1653 20684
rect 1611 20635 1653 20644
rect 2272 20684 2314 20693
rect 2272 20644 2273 20684
rect 2313 20644 2314 20684
rect 2272 20635 2314 20644
rect 3542 20684 3584 20693
rect 3542 20644 3543 20684
rect 3583 20644 3584 20684
rect 3542 20635 3584 20644
rect 4107 20684 4149 20693
rect 4107 20644 4108 20684
rect 4148 20644 4149 20684
rect 4107 20635 4149 20644
rect 6123 20684 6165 20693
rect 6123 20644 6124 20684
rect 6164 20644 6165 20684
rect 6123 20635 6165 20644
rect 7755 20684 7797 20693
rect 7755 20644 7756 20684
rect 7796 20644 7797 20684
rect 7755 20635 7797 20644
rect 7961 20684 8003 20693
rect 7961 20644 7962 20684
rect 8002 20644 8003 20684
rect 7961 20635 8003 20644
rect 9675 20684 9717 20693
rect 9675 20644 9676 20684
rect 9716 20644 9717 20684
rect 9675 20635 9717 20644
rect 9949 20684 9991 20693
rect 9949 20644 9950 20684
rect 9990 20644 9991 20684
rect 9949 20635 9991 20644
rect 12939 20684 12981 20693
rect 12939 20644 12940 20684
rect 12980 20644 12981 20684
rect 12939 20635 12981 20644
rect 14365 20684 14407 20693
rect 14365 20644 14366 20684
rect 14406 20644 14407 20684
rect 14365 20635 14407 20644
rect 15641 20684 15683 20693
rect 15641 20644 15642 20684
rect 15682 20644 15683 20684
rect 15641 20635 15683 20644
rect 16570 20684 16628 20685
rect 16570 20644 16579 20684
rect 16619 20644 16628 20684
rect 16570 20643 16628 20644
rect 18411 20684 18453 20693
rect 18411 20644 18412 20684
rect 18452 20644 18453 20684
rect 18411 20635 18453 20644
rect 23290 20684 23348 20685
rect 23290 20644 23299 20684
rect 23339 20644 23348 20684
rect 23290 20643 23348 20644
rect 27723 20684 27765 20693
rect 27723 20644 27724 20684
rect 27764 20644 27765 20684
rect 27723 20635 27765 20644
rect 30682 20684 30740 20685
rect 30682 20644 30691 20684
rect 30731 20644 30740 20684
rect 30682 20643 30740 20644
rect 1995 20600 2037 20609
rect 1995 20560 1996 20600
rect 2036 20560 2037 20600
rect 1995 20551 2037 20560
rect 2362 20600 2420 20601
rect 2362 20560 2371 20600
rect 2411 20560 2420 20600
rect 2362 20559 2420 20560
rect 2475 20600 2517 20609
rect 2475 20560 2476 20600
rect 2516 20560 2517 20600
rect 2475 20551 2517 20560
rect 2890 20600 2948 20601
rect 2890 20560 2899 20600
rect 2939 20560 2948 20600
rect 2890 20559 2948 20560
rect 3322 20600 3380 20601
rect 3322 20560 3331 20600
rect 3371 20560 3380 20600
rect 3322 20559 3380 20560
rect 3675 20600 3717 20609
rect 3675 20560 3676 20600
rect 3716 20560 3717 20600
rect 3675 20551 3717 20560
rect 5739 20600 5781 20609
rect 5739 20560 5740 20600
rect 5780 20560 5781 20600
rect 5739 20551 5781 20560
rect 6411 20600 6453 20609
rect 6411 20560 6412 20600
rect 6452 20560 6453 20600
rect 6411 20551 6453 20560
rect 10042 20600 10100 20601
rect 10042 20560 10051 20600
rect 10091 20560 10100 20600
rect 10042 20559 10100 20560
rect 10155 20600 10197 20609
rect 10155 20560 10156 20600
rect 10196 20560 10197 20600
rect 10155 20551 10197 20560
rect 10858 20600 10916 20601
rect 10858 20560 10867 20600
rect 10907 20560 10916 20600
rect 10858 20559 10916 20560
rect 11338 20600 11396 20601
rect 11338 20560 11347 20600
rect 11387 20560 11396 20600
rect 11338 20559 11396 20560
rect 13546 20600 13604 20601
rect 13546 20560 13555 20600
rect 13595 20560 13604 20600
rect 13546 20559 13604 20560
rect 13882 20600 13940 20601
rect 13882 20560 13891 20600
rect 13931 20560 13940 20600
rect 13882 20559 13940 20560
rect 15130 20600 15188 20601
rect 15130 20560 15139 20600
rect 15179 20560 15188 20600
rect 15130 20559 15188 20560
rect 15418 20600 15476 20601
rect 15418 20560 15427 20600
rect 15467 20560 15476 20600
rect 15418 20559 15476 20560
rect 15946 20600 16004 20601
rect 15946 20560 15955 20600
rect 15995 20560 16004 20600
rect 15946 20559 16004 20560
rect 18010 20600 18068 20601
rect 18010 20560 18019 20600
rect 18059 20560 18068 20600
rect 18010 20559 18068 20560
rect 18298 20600 18356 20601
rect 18298 20560 18307 20600
rect 18347 20560 18356 20600
rect 18298 20559 18356 20560
rect 18987 20600 19029 20609
rect 18987 20560 18988 20600
rect 19028 20560 19029 20600
rect 18987 20551 19029 20560
rect 20715 20600 20757 20609
rect 20715 20560 20716 20600
rect 20756 20560 20757 20600
rect 20715 20551 20757 20560
rect 22827 20600 22869 20609
rect 22827 20560 22828 20600
rect 22868 20560 22869 20600
rect 22827 20551 22869 20560
rect 24826 20600 24884 20601
rect 24826 20560 24835 20600
rect 24875 20560 24884 20600
rect 24826 20559 24884 20560
rect 25498 20600 25556 20601
rect 25498 20560 25507 20600
rect 25547 20560 25556 20600
rect 25498 20559 25556 20560
rect 25786 20600 25844 20601
rect 25786 20560 25795 20600
rect 25835 20560 25844 20600
rect 25786 20559 25844 20560
rect 26746 20600 26804 20601
rect 26746 20560 26755 20600
rect 26795 20560 26804 20600
rect 26746 20559 26804 20560
rect 26859 20600 26901 20609
rect 26859 20560 26860 20600
rect 26900 20560 26901 20600
rect 26859 20551 26901 20560
rect 27435 20600 27477 20609
rect 27435 20560 27436 20600
rect 27476 20560 27477 20600
rect 27435 20551 27477 20560
rect 28779 20600 28821 20609
rect 28779 20560 28780 20600
rect 28820 20560 28821 20600
rect 28779 20551 28821 20560
rect 30970 20600 31028 20601
rect 30970 20560 30979 20600
rect 31019 20560 31028 20600
rect 30970 20559 31028 20560
rect 576 20432 31392 20456
rect 576 20392 4352 20432
rect 4720 20392 12126 20432
rect 12494 20392 19900 20432
rect 20268 20392 27674 20432
rect 28042 20392 31392 20432
rect 576 20368 31392 20392
rect 2667 20264 2709 20273
rect 2667 20224 2668 20264
rect 2708 20224 2709 20264
rect 2667 20215 2709 20224
rect 3226 20264 3284 20265
rect 3226 20224 3235 20264
rect 3275 20224 3284 20264
rect 3226 20223 3284 20224
rect 5355 20264 5397 20273
rect 5355 20224 5356 20264
rect 5396 20224 5397 20264
rect 5355 20215 5397 20224
rect 6202 20264 6260 20265
rect 6202 20224 6211 20264
rect 6251 20224 6260 20264
rect 6202 20223 6260 20224
rect 6315 20264 6357 20273
rect 6315 20224 6316 20264
rect 6356 20224 6357 20264
rect 6315 20215 6357 20224
rect 7371 20264 7413 20273
rect 7371 20224 7372 20264
rect 7412 20224 7413 20264
rect 7371 20215 7413 20224
rect 8763 20264 8805 20273
rect 8763 20224 8764 20264
rect 8804 20224 8805 20264
rect 8763 20215 8805 20224
rect 11691 20264 11733 20273
rect 11691 20224 11692 20264
rect 11732 20224 11733 20264
rect 11691 20215 11733 20224
rect 12739 20264 12797 20265
rect 12739 20224 12748 20264
rect 12788 20224 12797 20264
rect 12739 20223 12797 20224
rect 12922 20264 12980 20265
rect 12922 20224 12931 20264
rect 12971 20224 12980 20264
rect 12922 20223 12980 20224
rect 13131 20264 13173 20273
rect 13131 20224 13132 20264
rect 13172 20224 13173 20264
rect 13131 20215 13173 20224
rect 14170 20264 14228 20265
rect 14170 20224 14179 20264
rect 14219 20224 14228 20264
rect 14170 20223 14228 20224
rect 14842 20264 14900 20265
rect 14842 20224 14851 20264
rect 14891 20224 14900 20264
rect 14842 20223 14900 20224
rect 14955 20264 14997 20273
rect 14955 20224 14956 20264
rect 14996 20224 14997 20264
rect 14955 20215 14997 20224
rect 16203 20264 16245 20273
rect 16203 20224 16204 20264
rect 16244 20224 16245 20264
rect 16203 20215 16245 20224
rect 16570 20264 16628 20265
rect 16570 20224 16579 20264
rect 16619 20224 16628 20264
rect 16570 20223 16628 20224
rect 17259 20264 17301 20273
rect 17259 20224 17260 20264
rect 17300 20224 17301 20264
rect 17259 20215 17301 20224
rect 18682 20264 18740 20265
rect 18682 20224 18691 20264
rect 18731 20224 18740 20264
rect 18682 20223 18740 20224
rect 18795 20264 18837 20273
rect 18795 20224 18796 20264
rect 18836 20224 18837 20264
rect 18795 20215 18837 20224
rect 19258 20264 19316 20265
rect 19258 20224 19267 20264
rect 19307 20224 19316 20264
rect 19258 20223 19316 20224
rect 19707 20264 19749 20273
rect 19707 20224 19708 20264
rect 19748 20224 19749 20264
rect 19707 20215 19749 20224
rect 24970 20264 25028 20265
rect 24970 20224 24979 20264
rect 25019 20224 25028 20264
rect 24970 20223 25028 20224
rect 28971 20264 29013 20273
rect 28971 20224 28972 20264
rect 29012 20224 29013 20264
rect 28971 20215 29013 20224
rect 4059 20180 4101 20189
rect 4059 20140 4060 20180
rect 4100 20140 4101 20180
rect 4059 20131 4101 20140
rect 4672 20180 4714 20189
rect 4672 20140 4673 20180
rect 4713 20140 4714 20180
rect 4672 20131 4714 20140
rect 4875 20180 4917 20189
rect 4875 20140 4876 20180
rect 4916 20140 4917 20180
rect 4875 20131 4917 20140
rect 13786 20180 13844 20181
rect 13786 20140 13795 20180
rect 13835 20140 13844 20180
rect 13786 20139 13844 20140
rect 17163 20180 17205 20189
rect 17163 20140 17164 20180
rect 17204 20140 17205 20180
rect 17163 20131 17205 20140
rect 17846 20180 17888 20189
rect 17846 20140 17847 20180
rect 17887 20140 17888 20180
rect 17846 20131 17888 20140
rect 20602 20180 20660 20181
rect 20602 20140 20611 20180
rect 20651 20140 20660 20180
rect 20602 20139 20660 20140
rect 24747 20180 24789 20189
rect 24747 20140 24748 20180
rect 24788 20140 24789 20180
rect 24747 20131 24789 20140
rect 25899 20180 25941 20189
rect 25899 20140 25900 20180
rect 25940 20140 25941 20180
rect 25899 20131 25941 20140
rect 27819 20180 27861 20189
rect 27819 20140 27820 20180
rect 27860 20140 27861 20180
rect 27819 20131 27861 20140
rect 28779 20180 28821 20189
rect 28779 20140 28780 20180
rect 28820 20140 28821 20180
rect 28779 20131 28821 20140
rect 31258 20180 31316 20181
rect 31258 20140 31267 20180
rect 31307 20140 31316 20180
rect 31258 20139 31316 20140
rect 1707 20096 1749 20105
rect 1707 20056 1708 20096
rect 1748 20056 1749 20096
rect 1707 20047 1749 20056
rect 2134 20096 2176 20105
rect 2134 20056 2135 20096
rect 2175 20056 2176 20096
rect 2134 20047 2176 20056
rect 2379 20096 2421 20105
rect 2379 20056 2380 20096
rect 2420 20056 2421 20096
rect 2379 20047 2421 20056
rect 2763 20096 2805 20105
rect 2763 20056 2764 20096
rect 2804 20056 2805 20096
rect 2763 20047 2805 20056
rect 2992 20096 3050 20097
rect 2992 20056 3001 20096
rect 3041 20056 3050 20096
rect 2992 20055 3050 20056
rect 3387 20096 3429 20105
rect 3387 20056 3388 20096
rect 3428 20056 3429 20096
rect 3387 20047 3429 20056
rect 3531 20096 3573 20105
rect 5152 20096 5194 20105
rect 5739 20096 5781 20105
rect 3531 20056 3532 20096
rect 3572 20056 3573 20096
rect 3531 20047 3573 20056
rect 4971 20087 5013 20096
rect 4971 20047 4972 20087
rect 5012 20047 5013 20087
rect 5152 20056 5153 20096
rect 5193 20056 5194 20096
rect 5152 20047 5194 20056
rect 5451 20087 5493 20096
rect 5451 20047 5452 20087
rect 5492 20047 5493 20087
rect 5739 20056 5740 20096
rect 5780 20056 5781 20096
rect 5739 20047 5781 20056
rect 5968 20096 6026 20097
rect 5968 20056 5977 20096
rect 6017 20056 6026 20096
rect 5968 20055 6026 20056
rect 6112 20096 6154 20105
rect 6603 20096 6645 20105
rect 6112 20056 6113 20096
rect 6153 20056 6154 20096
rect 6112 20047 6154 20056
rect 6411 20087 6453 20096
rect 6411 20047 6412 20087
rect 6452 20047 6453 20087
rect 6603 20056 6604 20096
rect 6644 20056 6645 20096
rect 6603 20047 6645 20056
rect 6708 20096 6750 20105
rect 6708 20056 6709 20096
rect 6749 20056 6750 20096
rect 6708 20047 6750 20056
rect 6930 20096 6972 20105
rect 6930 20056 6931 20096
rect 6971 20056 6972 20096
rect 6930 20047 6972 20056
rect 7083 20096 7125 20105
rect 7083 20056 7084 20096
rect 7124 20056 7125 20096
rect 7083 20047 7125 20056
rect 7217 20096 7275 20097
rect 7217 20056 7226 20096
rect 7266 20056 7275 20096
rect 7217 20055 7275 20056
rect 7755 20096 7797 20105
rect 9387 20096 9429 20105
rect 7755 20056 7756 20096
rect 7796 20056 7797 20096
rect 7755 20047 7797 20056
rect 8130 20087 8176 20096
rect 8130 20047 8131 20087
rect 8171 20047 8176 20087
rect 4971 20038 5013 20047
rect 5451 20038 5493 20047
rect 6411 20038 6453 20047
rect 8130 20038 8176 20047
rect 8610 20087 8656 20096
rect 8610 20047 8611 20087
rect 8651 20047 8656 20087
rect 9387 20056 9388 20096
rect 9428 20056 9429 20096
rect 9387 20047 9429 20056
rect 9754 20096 9812 20097
rect 9754 20056 9763 20096
rect 9803 20056 9812 20096
rect 9754 20055 9812 20056
rect 12346 20096 12404 20097
rect 12346 20056 12355 20096
rect 12395 20056 12404 20096
rect 12346 20055 12404 20056
rect 13306 20096 13364 20097
rect 13306 20056 13315 20096
rect 13355 20056 13364 20096
rect 13306 20055 13364 20056
rect 13707 20096 13749 20105
rect 13707 20056 13708 20096
rect 13748 20056 13749 20096
rect 13707 20047 13749 20056
rect 13899 20096 13941 20105
rect 13899 20056 13900 20096
rect 13940 20056 13941 20096
rect 13899 20047 13941 20056
rect 14283 20096 14325 20105
rect 14283 20056 14284 20096
rect 14324 20056 14325 20096
rect 14283 20047 14325 20056
rect 14749 20096 14791 20105
rect 15339 20096 15381 20105
rect 14749 20056 14750 20096
rect 14790 20056 14791 20096
rect 14749 20047 14791 20056
rect 15051 20087 15093 20096
rect 15051 20047 15052 20087
rect 15092 20047 15093 20087
rect 15339 20056 15340 20096
rect 15380 20056 15381 20096
rect 15339 20047 15381 20056
rect 15531 20096 15573 20105
rect 15531 20056 15532 20096
rect 15572 20056 15573 20096
rect 15531 20047 15573 20056
rect 15723 20096 15765 20105
rect 15723 20056 15724 20096
rect 15764 20056 15765 20096
rect 15723 20047 15765 20056
rect 15915 20096 15957 20105
rect 15915 20056 15916 20096
rect 15956 20056 15957 20096
rect 15915 20047 15957 20056
rect 16107 20096 16149 20105
rect 16107 20056 16108 20096
rect 16148 20056 16149 20096
rect 16107 20047 16149 20056
rect 16299 20096 16341 20105
rect 16299 20056 16300 20096
rect 16340 20056 16341 20096
rect 16299 20047 16341 20056
rect 16683 20096 16725 20105
rect 16683 20056 16684 20096
rect 16724 20056 16725 20096
rect 16683 20047 16725 20056
rect 17050 20096 17108 20097
rect 17050 20056 17059 20096
rect 17099 20056 17108 20096
rect 17050 20055 17108 20056
rect 17366 20096 17408 20105
rect 17366 20056 17367 20096
rect 17407 20056 17408 20096
rect 17366 20047 17408 20056
rect 17530 20096 17588 20097
rect 17530 20056 17539 20096
rect 17579 20056 17588 20096
rect 17530 20055 17588 20056
rect 17643 20096 17685 20105
rect 17643 20056 17644 20096
rect 17684 20056 17685 20096
rect 17643 20047 17685 20056
rect 18106 20096 18164 20097
rect 18106 20056 18115 20096
rect 18155 20056 18164 20096
rect 18106 20055 18164 20056
rect 18219 20096 18261 20105
rect 18219 20056 18220 20096
rect 18260 20056 18261 20096
rect 18219 20047 18261 20056
rect 18422 20096 18464 20105
rect 18422 20056 18423 20096
rect 18463 20056 18464 20096
rect 18422 20047 18464 20056
rect 18586 20096 18644 20097
rect 18586 20056 18595 20096
rect 18635 20056 18644 20096
rect 18586 20055 18644 20056
rect 18902 20096 18944 20105
rect 18902 20056 18903 20096
rect 18943 20056 18944 20096
rect 18902 20047 18944 20056
rect 19083 20096 19125 20105
rect 19083 20056 19084 20096
rect 19124 20056 19125 20096
rect 19083 20047 19125 20056
rect 19275 20096 19317 20105
rect 19275 20056 19276 20096
rect 19316 20056 19317 20096
rect 19275 20047 19317 20056
rect 19519 20096 19577 20097
rect 19519 20056 19528 20096
rect 19568 20056 19577 20096
rect 19519 20055 19577 20056
rect 20218 20096 20276 20097
rect 20218 20056 20227 20096
rect 20267 20056 20276 20096
rect 20218 20055 20276 20056
rect 22522 20096 22580 20097
rect 22522 20056 22531 20096
rect 22571 20056 22580 20096
rect 22522 20055 22580 20056
rect 23403 20096 23445 20105
rect 23403 20056 23404 20096
rect 23444 20056 23445 20096
rect 23403 20047 23445 20056
rect 23524 20096 23582 20097
rect 23524 20056 23533 20096
rect 23573 20056 23582 20096
rect 23524 20055 23582 20056
rect 23787 20096 23829 20105
rect 23787 20056 23788 20096
rect 23828 20056 23829 20096
rect 23787 20047 23829 20056
rect 24442 20096 24500 20097
rect 24442 20056 24451 20096
rect 24491 20056 24500 20096
rect 24442 20055 24500 20056
rect 25114 20096 25172 20097
rect 25995 20096 26037 20105
rect 25114 20056 25123 20096
rect 25163 20056 25172 20096
rect 25114 20055 25172 20056
rect 25227 20087 25269 20096
rect 25227 20047 25228 20087
rect 25268 20047 25269 20087
rect 25995 20056 25996 20096
rect 26036 20056 26037 20096
rect 25995 20047 26037 20056
rect 26224 20096 26282 20097
rect 26224 20056 26233 20096
rect 26273 20056 26282 20096
rect 26224 20055 26282 20056
rect 26701 20096 26759 20097
rect 26701 20056 26710 20096
rect 26750 20056 26759 20096
rect 26701 20055 26759 20056
rect 27136 20096 27178 20105
rect 27136 20056 27137 20096
rect 27177 20056 27178 20096
rect 27136 20047 27178 20056
rect 27243 20096 27285 20105
rect 27243 20056 27244 20096
rect 27284 20056 27285 20096
rect 27243 20047 27285 20056
rect 27610 20096 27668 20097
rect 27610 20056 27619 20096
rect 27659 20056 27668 20096
rect 27610 20055 27668 20056
rect 27911 20096 27953 20105
rect 27911 20056 27912 20096
rect 27952 20056 27953 20096
rect 27911 20047 27953 20056
rect 28155 20096 28197 20105
rect 28155 20056 28156 20096
rect 28196 20056 28197 20096
rect 28155 20047 28197 20056
rect 30874 20096 30932 20097
rect 30874 20056 30883 20096
rect 30923 20056 30932 20096
rect 30874 20055 30932 20056
rect 8610 20038 8656 20047
rect 15051 20038 15093 20047
rect 25227 20038 25269 20047
rect 2266 20012 2324 20013
rect 2266 19972 2275 20012
rect 2315 19972 2324 20012
rect 2266 19971 2324 19972
rect 2475 20012 2517 20021
rect 3915 20012 3957 20021
rect 2475 19972 2476 20012
rect 2516 19972 2517 20012
rect 2475 19963 2517 19972
rect 2898 20003 2944 20012
rect 2898 19963 2899 20003
rect 2939 19963 2944 20003
rect 3915 19972 3916 20012
rect 3956 19972 3957 20012
rect 3915 19963 3957 19972
rect 4299 20012 4341 20021
rect 4299 19972 4300 20012
rect 4340 19972 4341 20012
rect 4299 19963 4341 19972
rect 5643 20012 5685 20021
rect 8283 20012 8325 20021
rect 5643 19972 5644 20012
rect 5684 19972 5685 20012
rect 5643 19963 5685 19972
rect 5874 20003 5920 20012
rect 5874 19963 5875 20003
rect 5915 19963 5920 20003
rect 2898 19954 2944 19963
rect 5874 19954 5920 19963
rect 6834 20003 6880 20012
rect 6834 19963 6835 20003
rect 6875 19963 6880 20003
rect 8283 19972 8284 20012
rect 8324 19972 8325 20012
rect 8283 19963 8325 19972
rect 12538 20012 12596 20013
rect 12538 19972 12547 20012
rect 12587 19972 12596 20012
rect 12538 19971 12596 19972
rect 22906 20012 22964 20013
rect 22906 19972 22915 20012
rect 22955 19972 22964 20012
rect 22906 19971 22964 19972
rect 24267 20012 24309 20021
rect 24267 19972 24268 20012
rect 24308 19972 24309 20012
rect 24267 19963 24309 19972
rect 24843 20012 24885 20021
rect 24843 19972 24844 20012
rect 24884 19972 24885 20012
rect 24843 19963 24885 19972
rect 26114 20012 26156 20021
rect 26114 19972 26115 20012
rect 26155 19972 26156 20012
rect 26114 19963 26156 19972
rect 26506 20012 26564 20013
rect 26506 19972 26515 20012
rect 26555 19972 26564 20012
rect 26506 19971 26564 19972
rect 6834 19954 6880 19963
rect 11883 19928 11925 19937
rect 11883 19888 11884 19928
rect 11924 19888 11925 19928
rect 11883 19879 11925 19888
rect 14475 19928 14517 19937
rect 14475 19888 14476 19928
rect 14516 19888 14517 19928
rect 14475 19879 14517 19888
rect 20271 19928 20313 19937
rect 20271 19888 20272 19928
rect 20312 19888 20313 19928
rect 20271 19879 20313 19888
rect 23115 19928 23157 19937
rect 23115 19888 23116 19928
rect 23156 19888 23157 19928
rect 23115 19879 23157 19888
rect 922 19844 980 19845
rect 922 19804 931 19844
rect 971 19804 980 19844
rect 922 19803 980 19804
rect 3675 19844 3717 19853
rect 3675 19804 3676 19844
rect 3716 19804 3717 19844
rect 3675 19795 3717 19804
rect 4666 19844 4724 19845
rect 4666 19804 4675 19844
rect 4715 19804 4724 19844
rect 4666 19803 4724 19804
rect 5146 19844 5204 19845
rect 5146 19804 5155 19844
rect 5195 19804 5204 19844
rect 5146 19803 5204 19804
rect 7851 19844 7893 19853
rect 7851 19804 7852 19844
rect 7892 19804 7893 19844
rect 7851 19795 7893 19804
rect 15435 19844 15477 19853
rect 15435 19804 15436 19844
rect 15476 19804 15477 19844
rect 15435 19795 15477 19804
rect 15723 19844 15765 19853
rect 15723 19804 15724 19844
rect 15764 19804 15765 19844
rect 15723 19795 15765 19804
rect 16875 19844 16917 19853
rect 16875 19804 16876 19844
rect 16916 19804 16917 19844
rect 16875 19795 16917 19804
rect 17835 19844 17877 19853
rect 17835 19804 17836 19844
rect 17876 19804 17877 19844
rect 17835 19795 17877 19804
rect 18411 19844 18453 19853
rect 18411 19804 18412 19844
rect 18452 19804 18453 19844
rect 18411 19795 18453 19804
rect 20043 19844 20085 19853
rect 20043 19804 20044 19844
rect 20084 19804 20085 19844
rect 20043 19795 20085 19804
rect 21003 19844 21045 19853
rect 21003 19804 21004 19844
rect 21044 19804 21045 19844
rect 21003 19795 21045 19804
rect 25515 19844 25557 19853
rect 25515 19804 25516 19844
rect 25556 19804 25557 19844
rect 25515 19795 25557 19804
rect 27243 19844 27285 19853
rect 27243 19804 27244 19844
rect 27284 19804 27285 19844
rect 27243 19795 27285 19804
rect 576 19676 31392 19700
rect 576 19636 3112 19676
rect 3480 19636 10886 19676
rect 11254 19636 18660 19676
rect 19028 19636 26434 19676
rect 26802 19636 31392 19676
rect 576 19612 31392 19636
rect 2170 19508 2228 19509
rect 2170 19468 2179 19508
rect 2219 19468 2228 19508
rect 2170 19467 2228 19468
rect 3723 19508 3765 19517
rect 3723 19468 3724 19508
rect 3764 19468 3765 19508
rect 3723 19459 3765 19468
rect 4378 19508 4436 19509
rect 4378 19468 4387 19508
rect 4427 19468 4436 19508
rect 4378 19467 4436 19468
rect 5914 19508 5972 19509
rect 5914 19468 5923 19508
rect 5963 19468 5972 19508
rect 5914 19467 5972 19468
rect 6874 19508 6932 19509
rect 6874 19468 6883 19508
rect 6923 19468 6932 19508
rect 6874 19467 6932 19468
rect 9579 19508 9621 19517
rect 9579 19468 9580 19508
rect 9620 19468 9621 19508
rect 9579 19459 9621 19468
rect 11002 19508 11060 19509
rect 11002 19468 11011 19508
rect 11051 19468 11060 19508
rect 11002 19467 11060 19468
rect 13467 19508 13509 19517
rect 13467 19468 13468 19508
rect 13508 19468 13509 19508
rect 13467 19459 13509 19468
rect 14571 19508 14613 19517
rect 14571 19468 14572 19508
rect 14612 19468 14613 19508
rect 14571 19459 14613 19468
rect 16491 19508 16533 19517
rect 16491 19468 16492 19508
rect 16532 19468 16533 19508
rect 16491 19459 16533 19468
rect 18411 19508 18453 19517
rect 18411 19468 18412 19508
rect 18452 19468 18453 19508
rect 18411 19459 18453 19468
rect 19450 19508 19508 19509
rect 19450 19468 19459 19508
rect 19499 19468 19508 19508
rect 19450 19467 19508 19468
rect 22443 19508 22485 19517
rect 22443 19468 22444 19508
rect 22484 19468 22485 19508
rect 22443 19459 22485 19468
rect 23115 19508 23157 19517
rect 23115 19468 23116 19508
rect 23156 19468 23157 19508
rect 23115 19459 23157 19468
rect 31275 19508 31317 19517
rect 31275 19468 31276 19508
rect 31316 19468 31317 19508
rect 31275 19459 31317 19468
rect 1611 19424 1653 19433
rect 1611 19384 1612 19424
rect 1652 19384 1653 19424
rect 1611 19375 1653 19384
rect 12939 19424 12981 19433
rect 12939 19384 12940 19424
rect 12980 19384 12981 19424
rect 12939 19375 12981 19384
rect 843 19340 885 19349
rect 843 19300 844 19340
rect 884 19300 885 19340
rect 843 19291 885 19300
rect 5451 19340 5493 19349
rect 5451 19300 5452 19340
rect 5492 19300 5493 19340
rect 5451 19291 5493 19300
rect 5666 19340 5708 19349
rect 5666 19300 5667 19340
rect 5707 19300 5708 19340
rect 5666 19291 5708 19300
rect 6699 19340 6741 19349
rect 6699 19300 6700 19340
rect 6740 19300 6741 19340
rect 6699 19291 6741 19300
rect 7755 19340 7797 19349
rect 7755 19300 7756 19340
rect 7796 19300 7797 19340
rect 7755 19291 7797 19300
rect 9771 19340 9813 19349
rect 9771 19300 9772 19340
rect 9812 19300 9813 19340
rect 7169 19289 7227 19290
rect 1803 19256 1845 19265
rect 1803 19216 1804 19256
rect 1844 19216 1845 19256
rect 1803 19207 1845 19216
rect 1995 19256 2037 19265
rect 1995 19216 1996 19256
rect 2036 19216 2037 19256
rect 1995 19207 2037 19216
rect 2176 19256 2218 19265
rect 2176 19216 2177 19256
rect 2217 19216 2218 19256
rect 2176 19207 2218 19216
rect 2467 19256 2525 19257
rect 2467 19216 2476 19256
rect 2516 19216 2525 19256
rect 2467 19215 2525 19216
rect 2938 19256 2996 19257
rect 2938 19216 2947 19256
rect 2987 19216 2996 19256
rect 2938 19215 2996 19216
rect 3051 19256 3093 19265
rect 3051 19216 3052 19256
rect 3092 19216 3093 19256
rect 3051 19207 3093 19216
rect 3418 19256 3476 19257
rect 3418 19216 3427 19256
rect 3467 19216 3476 19256
rect 3418 19215 3476 19216
rect 3737 19256 3779 19265
rect 3737 19216 3738 19256
rect 3778 19216 3779 19256
rect 3737 19207 3779 19216
rect 4011 19256 4053 19265
rect 4011 19216 4012 19256
rect 4052 19216 4053 19256
rect 4011 19207 4053 19216
rect 4130 19256 4172 19265
rect 4130 19216 4131 19256
rect 4171 19216 4172 19256
rect 4130 19207 4172 19216
rect 4240 19256 4298 19257
rect 4240 19216 4249 19256
rect 4289 19216 4298 19256
rect 4240 19215 4298 19216
rect 4381 19256 4423 19265
rect 4381 19216 4382 19256
rect 4422 19216 4423 19256
rect 4381 19207 4423 19216
rect 4675 19256 4733 19257
rect 4675 19216 4684 19256
rect 4724 19216 4733 19256
rect 4675 19215 4733 19216
rect 5067 19256 5109 19265
rect 5067 19216 5068 19256
rect 5108 19216 5109 19256
rect 5067 19207 5109 19216
rect 5259 19256 5301 19265
rect 5259 19216 5260 19256
rect 5300 19216 5301 19256
rect 5259 19207 5301 19216
rect 5547 19256 5589 19265
rect 5547 19216 5548 19256
rect 5588 19216 5589 19256
rect 5547 19207 5589 19216
rect 5776 19256 5834 19257
rect 5776 19216 5785 19256
rect 5825 19216 5834 19256
rect 5776 19215 5834 19216
rect 5920 19256 5962 19265
rect 5920 19216 5921 19256
rect 5961 19216 5962 19256
rect 5920 19207 5962 19216
rect 6211 19256 6269 19257
rect 6211 19216 6220 19256
rect 6260 19216 6269 19256
rect 6211 19215 6269 19216
rect 6358 19256 6400 19265
rect 6358 19216 6359 19256
rect 6399 19216 6400 19256
rect 6358 19207 6400 19216
rect 6490 19256 6548 19257
rect 6490 19216 6499 19256
rect 6539 19216 6548 19256
rect 6490 19215 6548 19216
rect 6603 19256 6645 19265
rect 6603 19216 6604 19256
rect 6644 19216 6645 19256
rect 6603 19207 6645 19216
rect 6880 19256 6922 19265
rect 6880 19216 6881 19256
rect 6921 19216 6922 19256
rect 7169 19249 7178 19289
rect 7218 19249 7227 19289
rect 9303 19289 9345 19298
rect 9771 19291 9813 19300
rect 10443 19340 10485 19349
rect 10443 19300 10444 19340
rect 10484 19300 10485 19340
rect 10443 19291 10485 19300
rect 13227 19340 13269 19349
rect 13227 19300 13228 19340
rect 13268 19300 13269 19340
rect 13227 19291 13269 19300
rect 15938 19340 15980 19349
rect 15938 19300 15939 19340
rect 15979 19300 15980 19340
rect 18699 19340 18741 19349
rect 15938 19291 15980 19300
rect 16059 19298 16101 19307
rect 18699 19300 18700 19340
rect 18740 19300 18741 19340
rect 7169 19248 7227 19249
rect 7851 19256 7893 19265
rect 6880 19207 6922 19216
rect 7851 19216 7852 19256
rect 7892 19216 7893 19256
rect 7851 19207 7893 19216
rect 7970 19256 8012 19265
rect 7970 19216 7971 19256
rect 8011 19216 8012 19256
rect 7970 19207 8012 19216
rect 8080 19256 8138 19257
rect 8080 19216 8089 19256
rect 8129 19216 8138 19256
rect 8080 19215 8138 19216
rect 8715 19256 8757 19265
rect 8715 19216 8716 19256
rect 8756 19216 8757 19256
rect 8715 19207 8757 19216
rect 8907 19256 8949 19265
rect 8907 19216 8908 19256
rect 8948 19216 8949 19256
rect 8907 19207 8949 19216
rect 9178 19256 9236 19257
rect 9178 19216 9187 19256
rect 9227 19216 9236 19256
rect 9303 19249 9304 19289
rect 9344 19249 9345 19289
rect 9303 19240 9345 19249
rect 9867 19256 9909 19265
rect 9178 19215 9236 19216
rect 9867 19216 9868 19256
rect 9908 19216 9909 19256
rect 9867 19207 9909 19216
rect 9986 19256 10028 19265
rect 9986 19216 9987 19256
rect 10027 19216 10028 19256
rect 9986 19207 10028 19216
rect 10098 19256 10140 19265
rect 10098 19216 10099 19256
rect 10139 19216 10140 19256
rect 10098 19207 10140 19216
rect 11299 19256 11357 19257
rect 11299 19216 11308 19256
rect 11348 19216 11357 19256
rect 11299 19215 11357 19216
rect 11671 19256 11729 19257
rect 12939 19256 12981 19265
rect 11671 19216 11680 19256
rect 11720 19216 11729 19256
rect 11671 19215 11729 19216
rect 12642 19247 12688 19256
rect 12642 19207 12643 19247
rect 12683 19207 12688 19247
rect 12939 19216 12940 19256
rect 12980 19216 12981 19256
rect 12939 19207 12981 19216
rect 13903 19256 13961 19257
rect 13903 19216 13912 19256
rect 13952 19216 13961 19256
rect 13903 19215 13961 19216
rect 14074 19256 14132 19257
rect 14074 19216 14083 19256
rect 14123 19216 14132 19256
rect 14074 19215 14132 19216
rect 14393 19256 14435 19265
rect 14393 19216 14394 19256
rect 14434 19216 14435 19256
rect 14393 19207 14435 19216
rect 14763 19256 14805 19265
rect 14763 19216 14764 19256
rect 14804 19216 14805 19256
rect 14763 19207 14805 19216
rect 14882 19256 14924 19265
rect 14882 19216 14883 19256
rect 14923 19216 14924 19256
rect 14882 19207 14924 19216
rect 15051 19256 15093 19265
rect 15051 19216 15052 19256
rect 15092 19216 15093 19256
rect 15051 19207 15093 19216
rect 15190 19256 15232 19265
rect 15190 19216 15191 19256
rect 15231 19216 15232 19256
rect 15190 19207 15232 19216
rect 15322 19256 15380 19257
rect 15322 19216 15331 19256
rect 15371 19216 15380 19256
rect 15322 19215 15380 19216
rect 15435 19256 15477 19265
rect 15435 19216 15436 19256
rect 15476 19216 15477 19256
rect 15435 19207 15477 19216
rect 15819 19256 15861 19265
rect 15819 19216 15820 19256
rect 15860 19216 15861 19256
rect 16059 19258 16060 19298
rect 16100 19258 16101 19298
rect 18135 19289 18177 19298
rect 18699 19291 18741 19300
rect 19738 19340 19796 19341
rect 19738 19300 19747 19340
rect 19787 19300 19796 19340
rect 19738 19299 19796 19300
rect 21867 19340 21909 19349
rect 21867 19300 21868 19340
rect 21908 19300 21909 19340
rect 21867 19291 21909 19300
rect 24038 19340 24096 19341
rect 24038 19300 24047 19340
rect 24087 19300 24096 19340
rect 24038 19299 24096 19300
rect 26571 19340 26613 19349
rect 26571 19300 26572 19340
rect 26612 19300 26613 19340
rect 26571 19291 26613 19300
rect 27051 19340 27093 19349
rect 27051 19300 27052 19340
rect 27092 19300 27093 19340
rect 27051 19291 27093 19300
rect 27266 19340 27308 19349
rect 27266 19300 27267 19340
rect 27307 19300 27308 19340
rect 27266 19291 27308 19300
rect 16059 19249 16101 19258
rect 16299 19256 16341 19265
rect 15819 19207 15861 19216
rect 16299 19216 16300 19256
rect 16340 19216 16341 19256
rect 16299 19207 16341 19216
rect 16975 19256 17033 19257
rect 16975 19216 16984 19256
rect 17024 19216 17033 19256
rect 16975 19215 17033 19216
rect 17163 19256 17205 19265
rect 17163 19216 17164 19256
rect 17204 19216 17205 19256
rect 17163 19207 17205 19216
rect 17302 19256 17344 19265
rect 17302 19216 17303 19256
rect 17343 19216 17344 19256
rect 17302 19207 17344 19216
rect 18010 19256 18068 19257
rect 18010 19216 18019 19256
rect 18059 19216 18068 19256
rect 18135 19249 18136 19289
rect 18176 19249 18177 19289
rect 18135 19240 18177 19249
rect 18603 19256 18645 19265
rect 18010 19215 18068 19216
rect 18603 19216 18604 19256
rect 18644 19216 18645 19256
rect 18603 19207 18645 19216
rect 18795 19256 18837 19265
rect 18795 19216 18796 19256
rect 18836 19216 18837 19256
rect 18795 19207 18837 19216
rect 19275 19256 19317 19265
rect 19275 19216 19276 19256
rect 19316 19216 19317 19256
rect 19275 19207 19317 19216
rect 19444 19256 19486 19265
rect 19444 19216 19445 19256
rect 19485 19216 19486 19256
rect 19444 19207 19486 19216
rect 19606 19256 19648 19265
rect 19606 19216 19607 19256
rect 19647 19216 19648 19256
rect 19606 19207 19648 19216
rect 19851 19256 19893 19265
rect 19851 19216 19852 19256
rect 19892 19216 19893 19256
rect 19851 19207 19893 19216
rect 20394 19256 20452 19257
rect 20394 19216 20403 19256
rect 20443 19216 20452 19256
rect 20394 19215 20452 19216
rect 20794 19256 20852 19257
rect 20794 19216 20803 19256
rect 20843 19216 20852 19256
rect 20794 19215 20852 19216
rect 20986 19256 21044 19257
rect 20986 19216 20995 19256
rect 21035 19216 21044 19256
rect 20986 19215 21044 19216
rect 21291 19256 21333 19265
rect 21291 19216 21292 19256
rect 21332 19216 21333 19256
rect 21291 19207 21333 19216
rect 21483 19256 21525 19265
rect 21483 19216 21484 19256
rect 21524 19216 21525 19256
rect 21483 19207 21525 19216
rect 21771 19256 21813 19265
rect 21771 19216 21772 19256
rect 21812 19216 21813 19256
rect 21771 19207 21813 19216
rect 21963 19256 22005 19265
rect 21963 19216 21964 19256
rect 22004 19216 22005 19256
rect 21963 19207 22005 19216
rect 22138 19256 22196 19257
rect 22138 19216 22147 19256
rect 22187 19216 22196 19256
rect 22138 19215 22196 19216
rect 22618 19256 22676 19257
rect 22618 19216 22627 19256
rect 22667 19216 22676 19256
rect 22618 19215 22676 19216
rect 22923 19256 22965 19265
rect 22923 19216 22924 19256
rect 22964 19216 22965 19256
rect 22923 19207 22965 19216
rect 23115 19256 23157 19265
rect 23115 19216 23116 19256
rect 23156 19216 23157 19256
rect 23115 19207 23157 19216
rect 23232 19256 23290 19257
rect 23232 19216 23241 19256
rect 23281 19216 23290 19256
rect 23232 19215 23290 19216
rect 23403 19256 23445 19265
rect 23403 19216 23404 19256
rect 23444 19216 23445 19256
rect 23403 19207 23445 19216
rect 23936 19256 23994 19257
rect 23936 19216 23945 19256
rect 23985 19216 23994 19256
rect 23936 19215 23994 19216
rect 24154 19256 24212 19257
rect 24154 19216 24163 19256
rect 24203 19216 24212 19256
rect 24154 19215 24212 19216
rect 24267 19256 24309 19265
rect 24267 19216 24268 19256
rect 24308 19216 24309 19256
rect 24267 19207 24309 19216
rect 24651 19256 24693 19265
rect 24651 19216 24652 19256
rect 24692 19216 24693 19256
rect 24651 19207 24693 19216
rect 24826 19256 24884 19257
rect 24826 19216 24835 19256
rect 24875 19216 24884 19256
rect 24826 19215 24884 19216
rect 25323 19256 25365 19265
rect 25323 19216 25324 19256
rect 25364 19216 25365 19256
rect 25323 19207 25365 19216
rect 25611 19256 25653 19265
rect 25611 19216 25612 19256
rect 25652 19216 25653 19256
rect 25611 19207 25653 19216
rect 25995 19256 26037 19265
rect 25995 19216 25996 19256
rect 26036 19216 26037 19256
rect 25995 19207 26037 19216
rect 26650 19256 26708 19257
rect 26650 19216 26659 19256
rect 26699 19216 26708 19256
rect 26650 19215 26708 19216
rect 27147 19256 27189 19265
rect 27147 19216 27148 19256
rect 27188 19216 27189 19256
rect 27147 19207 27189 19216
rect 27376 19256 27434 19257
rect 27376 19216 27385 19256
rect 27425 19216 27434 19256
rect 27376 19215 27434 19216
rect 27623 19256 27665 19265
rect 27623 19216 27624 19256
rect 27664 19216 27665 19256
rect 27623 19207 27665 19216
rect 27819 19256 27861 19265
rect 27819 19216 27820 19256
rect 27860 19216 27861 19256
rect 27819 19207 27861 19216
rect 28107 19256 28149 19265
rect 28107 19216 28108 19256
rect 28148 19216 28149 19256
rect 28107 19207 28149 19216
rect 29338 19256 29396 19257
rect 29338 19216 29347 19256
rect 29387 19216 29396 19256
rect 29338 19215 29396 19216
rect 12642 19198 12688 19207
rect 3257 19172 3299 19181
rect 3257 19132 3258 19172
rect 3298 19132 3299 19172
rect 3257 19123 3299 19132
rect 11005 19172 11047 19181
rect 11005 19132 11006 19172
rect 11046 19132 11047 19172
rect 11005 19123 11047 19132
rect 15514 19172 15572 19173
rect 15514 19132 15523 19172
rect 15563 19132 15572 19172
rect 15514 19131 15572 19132
rect 21387 19172 21429 19181
rect 21387 19132 21388 19172
rect 21428 19132 21429 19172
rect 21387 19123 21429 19132
rect 22457 19172 22499 19181
rect 22457 19132 22458 19172
rect 22498 19132 22499 19172
rect 22457 19123 22499 19132
rect 24747 19172 24789 19181
rect 24747 19132 24748 19172
rect 24788 19132 24789 19172
rect 24747 19123 24789 19132
rect 28954 19172 29012 19173
rect 28954 19132 28963 19172
rect 29003 19132 29012 19172
rect 28954 19131 29012 19132
rect 603 19088 645 19097
rect 603 19048 604 19088
rect 644 19048 645 19088
rect 603 19039 645 19048
rect 1803 19088 1845 19097
rect 1803 19048 1804 19088
rect 1844 19048 1845 19088
rect 1803 19039 1845 19048
rect 2379 19088 2421 19097
rect 2379 19048 2380 19088
rect 2420 19048 2421 19088
rect 2379 19039 2421 19048
rect 3147 19088 3189 19097
rect 3147 19048 3148 19088
rect 3188 19048 3189 19088
rect 3147 19039 3189 19048
rect 3514 19088 3572 19089
rect 3514 19048 3523 19088
rect 3563 19048 3572 19088
rect 3514 19047 3572 19048
rect 3915 19088 3957 19097
rect 3915 19048 3916 19088
rect 3956 19048 3957 19088
rect 3915 19039 3957 19048
rect 4587 19088 4629 19097
rect 4587 19048 4588 19088
rect 4628 19048 4629 19088
rect 4587 19039 4629 19048
rect 5242 19088 5300 19089
rect 5242 19048 5251 19088
rect 5291 19048 5300 19088
rect 5242 19047 5300 19048
rect 6123 19088 6165 19097
rect 6123 19048 6124 19088
rect 6164 19048 6165 19088
rect 6123 19039 6165 19048
rect 7083 19088 7125 19097
rect 7083 19048 7084 19088
rect 7124 19048 7125 19088
rect 7083 19039 7125 19048
rect 8715 19088 8757 19097
rect 8715 19048 8716 19088
rect 8756 19048 8757 19088
rect 8715 19039 8757 19048
rect 9034 19088 9092 19089
rect 9034 19048 9043 19088
rect 9083 19048 9092 19088
rect 9034 19047 9092 19048
rect 10203 19088 10245 19097
rect 10203 19048 10204 19088
rect 10244 19048 10245 19088
rect 10203 19039 10245 19048
rect 11211 19088 11253 19097
rect 11211 19048 11212 19088
rect 11252 19048 11253 19088
rect 11211 19039 11253 19048
rect 11835 19088 11877 19097
rect 11835 19048 11836 19088
rect 11876 19048 11877 19088
rect 11835 19039 11877 19048
rect 13738 19088 13796 19089
rect 13738 19048 13747 19088
rect 13787 19048 13796 19088
rect 13738 19047 13796 19048
rect 14170 19088 14228 19089
rect 14170 19048 14179 19088
rect 14219 19048 14228 19088
rect 14170 19047 14228 19048
rect 14283 19088 14325 19097
rect 14283 19048 14284 19088
rect 14324 19048 14325 19088
rect 14283 19039 14325 19048
rect 15723 19088 15765 19097
rect 15723 19048 15724 19088
rect 15764 19048 15765 19088
rect 15723 19039 15765 19048
rect 16186 19088 16244 19089
rect 16186 19048 16195 19088
rect 16235 19048 16244 19088
rect 16186 19047 16244 19048
rect 16810 19088 16868 19089
rect 16810 19048 16819 19088
rect 16859 19048 16868 19088
rect 16810 19047 16868 19048
rect 17451 19088 17493 19097
rect 19930 19088 19988 19089
rect 17451 19048 17452 19088
rect 17492 19048 17493 19088
rect 17451 19039 17493 19048
rect 17922 19079 17968 19088
rect 17922 19039 17923 19079
rect 17963 19039 17968 19079
rect 19930 19048 19939 19088
rect 19979 19048 19988 19088
rect 19930 19047 19988 19048
rect 20506 19088 20564 19089
rect 20506 19048 20515 19088
rect 20555 19048 20564 19088
rect 20506 19047 20564 19048
rect 22234 19088 22292 19089
rect 22234 19048 22243 19088
rect 22283 19048 22292 19088
rect 22234 19047 22292 19048
rect 22827 19088 22869 19097
rect 22827 19048 22828 19088
rect 22868 19048 22869 19088
rect 22827 19039 22869 19048
rect 23979 19088 24021 19097
rect 23979 19048 23980 19088
rect 24020 19048 24021 19088
rect 23979 19039 24021 19048
rect 25114 19088 25172 19089
rect 25114 19048 25123 19088
rect 25163 19048 25172 19088
rect 25114 19047 25172 19048
rect 25803 19088 25845 19097
rect 25803 19048 25804 19088
rect 25844 19048 25845 19088
rect 25803 19039 25845 19048
rect 26074 19088 26132 19089
rect 27627 19088 27669 19097
rect 26074 19048 26083 19088
rect 26123 19048 26132 19088
rect 26074 19047 26132 19048
rect 26282 19079 26324 19088
rect 26282 19039 26283 19079
rect 26323 19039 26324 19079
rect 27627 19048 27628 19088
rect 27668 19048 27669 19088
rect 27627 19039 27669 19048
rect 28779 19088 28821 19097
rect 28779 19048 28780 19088
rect 28820 19048 28821 19088
rect 28779 19039 28821 19048
rect 17922 19030 17968 19039
rect 26282 19030 26324 19039
rect 576 18920 31392 18944
rect 576 18880 4352 18920
rect 4720 18880 12126 18920
rect 12494 18880 19900 18920
rect 20268 18880 27674 18920
rect 28042 18880 31392 18920
rect 576 18856 31392 18880
rect 747 18752 789 18761
rect 747 18712 748 18752
rect 788 18712 789 18752
rect 747 18703 789 18712
rect 5259 18752 5301 18761
rect 5259 18712 5260 18752
rect 5300 18712 5301 18752
rect 5259 18703 5301 18712
rect 6490 18752 6548 18753
rect 6490 18712 6499 18752
rect 6539 18712 6548 18752
rect 6490 18711 6548 18712
rect 6874 18752 6932 18753
rect 6874 18712 6883 18752
rect 6923 18712 6932 18752
rect 6874 18711 6932 18712
rect 7642 18752 7700 18753
rect 7642 18712 7651 18752
rect 7691 18712 7700 18752
rect 7642 18711 7700 18712
rect 8122 18752 8180 18753
rect 8122 18712 8131 18752
rect 8171 18712 8180 18752
rect 8122 18711 8180 18712
rect 9178 18752 9236 18753
rect 9178 18712 9187 18752
rect 9227 18712 9236 18752
rect 9178 18711 9236 18712
rect 9514 18752 9572 18753
rect 9514 18712 9523 18752
rect 9563 18712 9572 18752
rect 9514 18711 9572 18712
rect 10731 18752 10773 18761
rect 10731 18712 10732 18752
rect 10772 18712 10773 18752
rect 10731 18703 10773 18712
rect 12154 18752 12212 18753
rect 12154 18712 12163 18752
rect 12203 18712 12212 18752
rect 12154 18711 12212 18712
rect 13786 18752 13844 18753
rect 13786 18712 13795 18752
rect 13835 18712 13844 18752
rect 13786 18711 13844 18712
rect 15514 18752 15572 18753
rect 15514 18712 15523 18752
rect 15563 18712 15572 18752
rect 15514 18711 15572 18712
rect 17338 18752 17396 18753
rect 17338 18712 17347 18752
rect 17387 18712 17396 18752
rect 17338 18711 17396 18712
rect 20218 18752 20276 18753
rect 20218 18712 20227 18752
rect 20267 18712 20276 18752
rect 20218 18711 20276 18712
rect 20907 18752 20949 18761
rect 20907 18712 20908 18752
rect 20948 18712 20949 18752
rect 20907 18703 20949 18712
rect 21195 18752 21237 18761
rect 21195 18712 21196 18752
rect 21236 18712 21237 18752
rect 21195 18703 21237 18712
rect 23019 18752 23061 18761
rect 23019 18712 23020 18752
rect 23060 18712 23061 18752
rect 23019 18703 23061 18712
rect 24267 18752 24309 18761
rect 24267 18712 24268 18752
rect 24308 18712 24309 18752
rect 24267 18703 24309 18712
rect 25690 18752 25748 18753
rect 25690 18712 25699 18752
rect 25739 18712 25748 18752
rect 25690 18711 25748 18712
rect 10635 18668 10677 18677
rect 10635 18628 10636 18668
rect 10676 18628 10677 18668
rect 10635 18619 10677 18628
rect 10841 18668 10883 18677
rect 10841 18628 10842 18668
rect 10882 18628 10883 18668
rect 10841 18619 10883 18628
rect 11019 18668 11061 18677
rect 11019 18628 11020 18668
rect 11060 18628 11061 18668
rect 11019 18619 11061 18628
rect 14650 18668 14708 18669
rect 14650 18628 14659 18668
rect 14699 18628 14708 18668
rect 14650 18627 14708 18628
rect 17245 18668 17287 18677
rect 17245 18628 17246 18668
rect 17286 18628 17287 18668
rect 17245 18619 17287 18628
rect 18795 18668 18837 18677
rect 18795 18628 18796 18668
rect 18836 18628 18837 18668
rect 18795 18619 18837 18628
rect 19563 18668 19605 18677
rect 21850 18668 21908 18669
rect 19563 18628 19564 18668
rect 19604 18628 19605 18668
rect 19563 18619 19605 18628
rect 20130 18659 20176 18668
rect 20130 18619 20131 18659
rect 20171 18619 20176 18659
rect 21850 18628 21859 18668
rect 21899 18628 21908 18668
rect 21850 18627 21908 18628
rect 22443 18668 22485 18677
rect 22443 18628 22444 18668
rect 22484 18628 22485 18668
rect 22443 18619 22485 18628
rect 30411 18668 30453 18677
rect 30411 18628 30412 18668
rect 30452 18628 30453 18668
rect 30411 18619 30453 18628
rect 20130 18610 20176 18619
rect 2650 18584 2708 18585
rect 2650 18544 2659 18584
rect 2699 18544 2708 18584
rect 2650 18543 2708 18544
rect 3915 18584 3957 18593
rect 3915 18544 3916 18584
rect 3956 18544 3957 18584
rect 3915 18535 3957 18544
rect 4203 18584 4245 18593
rect 4203 18544 4204 18584
rect 4244 18544 4245 18584
rect 4203 18535 4245 18544
rect 4432 18584 4490 18585
rect 4432 18544 4441 18584
rect 4481 18544 4490 18584
rect 4432 18543 4490 18544
rect 4971 18584 5013 18593
rect 4971 18544 4972 18584
rect 5012 18544 5013 18584
rect 4971 18535 5013 18544
rect 5098 18584 5156 18585
rect 5098 18544 5107 18584
rect 5147 18544 5156 18584
rect 5098 18543 5156 18544
rect 5739 18584 5781 18593
rect 5739 18544 5740 18584
rect 5780 18544 5781 18584
rect 5739 18535 5781 18544
rect 5914 18584 5972 18585
rect 5914 18544 5923 18584
rect 5963 18544 5972 18584
rect 5914 18543 5972 18544
rect 6139 18584 6197 18585
rect 6139 18544 6148 18584
rect 6188 18544 6197 18584
rect 6139 18543 6197 18544
rect 6298 18584 6356 18585
rect 6298 18544 6307 18584
rect 6347 18544 6356 18584
rect 6298 18543 6356 18544
rect 6423 18584 6465 18593
rect 6423 18544 6424 18584
rect 6464 18544 6465 18584
rect 6682 18584 6740 18585
rect 6423 18535 6465 18544
rect 6582 18573 6640 18574
rect 6582 18533 6591 18573
rect 6631 18533 6640 18573
rect 6682 18544 6691 18584
rect 6731 18544 6740 18584
rect 6682 18543 6740 18544
rect 6987 18584 7029 18593
rect 6987 18544 6988 18584
rect 7028 18544 7029 18584
rect 7561 18584 7603 18593
rect 6987 18535 7029 18544
rect 7323 18542 7365 18551
rect 6582 18532 6640 18533
rect 3034 18500 3092 18501
rect 3034 18460 3043 18500
rect 3083 18460 3092 18500
rect 3034 18459 3092 18460
rect 4107 18500 4149 18509
rect 7323 18502 7324 18542
rect 7364 18502 7365 18542
rect 7561 18544 7562 18584
rect 7602 18544 7603 18584
rect 7561 18535 7603 18544
rect 7798 18584 7840 18593
rect 7798 18544 7799 18584
rect 7839 18544 7840 18584
rect 7798 18535 7840 18544
rect 8043 18584 8085 18593
rect 8043 18544 8044 18584
rect 8084 18544 8085 18584
rect 8043 18535 8085 18544
rect 8278 18584 8320 18593
rect 8278 18544 8279 18584
rect 8319 18544 8320 18584
rect 8278 18535 8320 18544
rect 8523 18584 8565 18593
rect 8523 18544 8524 18584
rect 8564 18544 8565 18584
rect 8523 18535 8565 18544
rect 8866 18584 8924 18585
rect 8866 18544 8875 18584
rect 8915 18544 8924 18584
rect 8866 18543 8924 18544
rect 9099 18584 9141 18593
rect 9099 18544 9100 18584
rect 9140 18544 9141 18584
rect 9099 18535 9141 18544
rect 9709 18584 9767 18585
rect 9709 18544 9718 18584
rect 9758 18544 9767 18584
rect 9709 18543 9767 18544
rect 10522 18584 10580 18585
rect 10522 18544 10531 18584
rect 10571 18544 10580 18584
rect 10522 18543 10580 18544
rect 11115 18584 11157 18593
rect 11115 18544 11116 18584
rect 11156 18544 11157 18584
rect 10378 18542 10436 18543
rect 4107 18460 4108 18500
rect 4148 18460 4149 18500
rect 4107 18451 4149 18460
rect 4338 18491 4384 18500
rect 7323 18493 7365 18502
rect 7450 18500 7508 18501
rect 4338 18451 4339 18491
rect 4379 18451 4384 18491
rect 7450 18460 7459 18500
rect 7499 18460 7508 18500
rect 7450 18459 7508 18460
rect 7930 18500 7988 18501
rect 7930 18460 7939 18500
rect 7979 18460 7988 18500
rect 7930 18459 7988 18460
rect 8410 18500 8468 18501
rect 8410 18460 8419 18500
rect 8459 18460 8468 18500
rect 8410 18459 8468 18460
rect 8619 18500 8661 18509
rect 10378 18502 10387 18542
rect 10427 18502 10436 18542
rect 11115 18535 11157 18544
rect 11344 18584 11402 18585
rect 11344 18544 11353 18584
rect 11393 18544 11402 18584
rect 11344 18543 11402 18544
rect 11821 18584 11879 18585
rect 11821 18544 11830 18584
rect 11870 18544 11879 18584
rect 11821 18543 11879 18544
rect 12267 18584 12309 18593
rect 12267 18544 12268 18584
rect 12308 18544 12309 18584
rect 12267 18535 12309 18544
rect 12607 18584 12665 18585
rect 12607 18544 12616 18584
rect 12656 18544 12665 18584
rect 12607 18543 12665 18544
rect 13450 18584 13508 18585
rect 13450 18544 13459 18584
rect 13499 18544 13508 18584
rect 13450 18543 13508 18544
rect 13645 18584 13703 18585
rect 13645 18544 13654 18584
rect 13694 18544 13703 18584
rect 13645 18543 13703 18544
rect 13947 18584 14005 18585
rect 13947 18544 13956 18584
rect 13996 18544 14005 18584
rect 13947 18543 14005 18544
rect 14091 18584 14133 18593
rect 14091 18544 14092 18584
rect 14132 18544 14133 18584
rect 14091 18535 14133 18544
rect 14326 18584 14368 18593
rect 14326 18544 14327 18584
rect 14367 18544 14368 18584
rect 14326 18535 14368 18544
rect 14458 18584 14516 18585
rect 14458 18544 14467 18584
rect 14507 18544 14516 18584
rect 14458 18543 14516 18544
rect 14571 18584 14613 18593
rect 14571 18544 14572 18584
rect 14612 18544 14613 18584
rect 14571 18535 14613 18544
rect 14806 18584 14848 18593
rect 14806 18544 14807 18584
rect 14847 18544 14848 18584
rect 14806 18535 14848 18544
rect 15051 18584 15093 18593
rect 15051 18544 15052 18584
rect 15092 18544 15093 18584
rect 15051 18535 15093 18544
rect 15339 18584 15381 18593
rect 15339 18544 15340 18584
rect 15380 18544 15381 18584
rect 15339 18535 15381 18544
rect 15531 18584 15573 18593
rect 15531 18544 15532 18584
rect 15572 18544 15573 18584
rect 15531 18535 15573 18544
rect 15906 18584 15948 18593
rect 15906 18544 15907 18584
rect 15947 18544 15948 18584
rect 15906 18535 15948 18544
rect 16011 18584 16053 18593
rect 16011 18544 16012 18584
rect 16052 18544 16053 18584
rect 16011 18535 16053 18544
rect 16203 18584 16245 18593
rect 16203 18544 16204 18584
rect 16244 18544 16245 18584
rect 16203 18535 16245 18544
rect 16687 18584 16745 18585
rect 16687 18544 16696 18584
rect 16736 18544 16745 18584
rect 16687 18543 16745 18544
rect 16870 18584 16912 18593
rect 16870 18544 16871 18584
rect 16911 18544 16912 18584
rect 16870 18535 16912 18544
rect 17067 18584 17109 18593
rect 17067 18544 17068 18584
rect 17108 18544 17109 18584
rect 17067 18535 17109 18544
rect 17451 18584 17493 18593
rect 17835 18584 17877 18593
rect 17451 18544 17452 18584
rect 17492 18544 17493 18584
rect 17451 18535 17493 18544
rect 17547 18575 17589 18584
rect 17547 18535 17548 18575
rect 17588 18535 17589 18575
rect 17835 18544 17836 18584
rect 17876 18544 17877 18584
rect 17835 18535 17877 18544
rect 18349 18584 18407 18585
rect 18349 18544 18358 18584
rect 18398 18544 18407 18584
rect 18349 18543 18407 18544
rect 18916 18584 18974 18585
rect 18916 18544 18925 18584
rect 18965 18544 18974 18584
rect 18916 18543 18974 18544
rect 19179 18584 19221 18593
rect 19179 18544 19180 18584
rect 19220 18544 19221 18584
rect 19179 18535 19221 18544
rect 19467 18584 19509 18593
rect 19467 18544 19468 18584
rect 19508 18544 19509 18584
rect 19467 18535 19509 18544
rect 19659 18584 19701 18593
rect 19659 18544 19660 18584
rect 19700 18544 19701 18584
rect 19659 18535 19701 18544
rect 19834 18584 19892 18585
rect 20218 18584 20276 18585
rect 19834 18544 19843 18584
rect 19883 18544 19892 18584
rect 19834 18543 19892 18544
rect 19947 18575 19989 18584
rect 19947 18535 19948 18575
rect 19988 18535 19989 18575
rect 20218 18544 20227 18584
rect 20267 18544 20276 18584
rect 20218 18543 20276 18544
rect 20395 18584 20453 18585
rect 20395 18544 20404 18584
rect 20444 18544 20453 18584
rect 20395 18543 20453 18544
rect 20650 18584 20708 18585
rect 20650 18544 20659 18584
rect 20699 18544 20708 18584
rect 20650 18543 20708 18544
rect 20753 18584 20811 18585
rect 20753 18544 20762 18584
rect 20802 18544 20811 18584
rect 20753 18543 20811 18544
rect 21099 18584 21141 18593
rect 21099 18544 21100 18584
rect 21140 18544 21141 18584
rect 21099 18535 21141 18544
rect 21291 18584 21333 18593
rect 21291 18544 21292 18584
rect 21332 18544 21333 18584
rect 21291 18535 21333 18544
rect 21771 18584 21813 18593
rect 21771 18544 21772 18584
rect 21812 18544 21813 18584
rect 21771 18535 21813 18544
rect 21946 18584 22004 18585
rect 21946 18544 21955 18584
rect 21995 18544 22004 18584
rect 21946 18543 22004 18544
rect 22059 18584 22101 18593
rect 22059 18544 22060 18584
rect 22100 18544 22101 18584
rect 22059 18535 22101 18544
rect 22234 18584 22292 18585
rect 22234 18544 22243 18584
rect 22283 18544 22292 18584
rect 22234 18543 22292 18544
rect 22347 18584 22389 18593
rect 22347 18544 22348 18584
rect 22388 18544 22389 18584
rect 22347 18535 22389 18544
rect 22553 18584 22595 18593
rect 22553 18544 22554 18584
rect 22594 18544 22595 18584
rect 22553 18535 22595 18544
rect 22731 18584 22773 18593
rect 23062 18584 23120 18585
rect 24224 18584 24282 18585
rect 22731 18544 22732 18584
rect 22772 18544 22773 18584
rect 22731 18535 22773 18544
rect 22962 18575 23008 18584
rect 22962 18535 22963 18575
rect 23003 18535 23008 18575
rect 23062 18544 23071 18584
rect 23111 18544 23120 18584
rect 23062 18543 23120 18544
rect 23595 18575 23637 18584
rect 17547 18526 17589 18535
rect 19947 18526 19989 18535
rect 22962 18526 23008 18535
rect 23595 18535 23596 18575
rect 23636 18535 23637 18575
rect 23595 18526 23637 18535
rect 23706 18575 23748 18584
rect 23706 18535 23707 18575
rect 23747 18535 23748 18575
rect 23706 18526 23748 18535
rect 23826 18575 23872 18584
rect 23826 18535 23827 18575
rect 23867 18535 23872 18575
rect 24224 18544 24233 18584
rect 24273 18544 24282 18584
rect 24224 18543 24282 18544
rect 24555 18584 24597 18593
rect 24555 18544 24556 18584
rect 24596 18544 24597 18584
rect 24555 18535 24597 18544
rect 24747 18584 24789 18593
rect 24747 18544 24748 18584
rect 24788 18544 24789 18584
rect 24747 18535 24789 18544
rect 24862 18584 24904 18593
rect 24862 18544 24863 18584
rect 24903 18544 24904 18584
rect 24862 18535 24904 18544
rect 25035 18584 25077 18593
rect 25035 18544 25036 18584
rect 25076 18544 25077 18584
rect 25035 18535 25077 18544
rect 25227 18584 25269 18593
rect 25227 18544 25228 18584
rect 25268 18544 25269 18584
rect 25227 18535 25269 18544
rect 25402 18584 25460 18585
rect 25402 18544 25411 18584
rect 25451 18544 25460 18584
rect 25402 18543 25460 18544
rect 25594 18584 25652 18585
rect 25594 18544 25603 18584
rect 25643 18544 25652 18584
rect 25594 18543 25652 18544
rect 25910 18584 25952 18593
rect 25910 18544 25911 18584
rect 25951 18544 25952 18584
rect 25910 18535 25952 18544
rect 26187 18584 26229 18593
rect 26187 18544 26188 18584
rect 26228 18544 26229 18584
rect 26187 18535 26229 18544
rect 26379 18584 26421 18593
rect 26379 18544 26380 18584
rect 26420 18544 26421 18584
rect 26379 18535 26421 18544
rect 26859 18584 26901 18593
rect 26859 18544 26860 18584
rect 26900 18544 26901 18584
rect 26859 18535 26901 18544
rect 27034 18584 27092 18585
rect 27034 18544 27043 18584
rect 27083 18544 27092 18584
rect 27034 18543 27092 18544
rect 27147 18584 27189 18593
rect 27147 18544 27148 18584
rect 27188 18544 27189 18584
rect 27147 18535 27189 18544
rect 29242 18584 29300 18585
rect 29242 18544 29251 18584
rect 29291 18544 29300 18584
rect 29242 18543 29300 18544
rect 29626 18584 29684 18585
rect 29626 18544 29635 18584
rect 29675 18544 29684 18584
rect 29626 18543 29684 18544
rect 29821 18584 29863 18593
rect 29821 18544 29822 18584
rect 29862 18544 29863 18584
rect 29821 18535 29863 18544
rect 29931 18584 29973 18593
rect 29931 18544 29932 18584
rect 29972 18544 29973 18584
rect 29931 18535 29973 18544
rect 30123 18584 30165 18593
rect 30123 18544 30124 18584
rect 30164 18544 30165 18584
rect 30123 18535 30165 18544
rect 30315 18584 30357 18593
rect 30315 18544 30316 18584
rect 30356 18544 30357 18584
rect 30315 18535 30357 18544
rect 30603 18584 30645 18593
rect 30603 18544 30604 18584
rect 30644 18544 30645 18584
rect 30603 18535 30645 18544
rect 30786 18575 30832 18584
rect 30786 18535 30787 18575
rect 30827 18535 30832 18575
rect 23826 18526 23872 18535
rect 30786 18526 30832 18535
rect 10378 18501 10436 18502
rect 8619 18460 8620 18500
rect 8660 18460 8661 18500
rect 8619 18451 8661 18460
rect 8986 18500 9044 18501
rect 8986 18460 8995 18500
rect 9035 18460 9044 18500
rect 8986 18459 9044 18460
rect 10186 18500 10244 18501
rect 11626 18500 11684 18501
rect 10186 18460 10195 18500
rect 10235 18460 10244 18500
rect 10186 18459 10244 18460
rect 11250 18491 11296 18500
rect 11250 18451 11251 18491
rect 11291 18451 11296 18491
rect 11626 18460 11635 18500
rect 11675 18460 11684 18500
rect 11626 18459 11684 18460
rect 12795 18500 12837 18509
rect 12795 18460 12796 18500
rect 12836 18460 12837 18500
rect 12795 18451 12837 18460
rect 14938 18500 14996 18501
rect 14938 18460 14947 18500
rect 14987 18460 14996 18500
rect 14938 18459 14996 18460
rect 15147 18500 15189 18509
rect 15147 18460 15148 18500
rect 15188 18460 15189 18500
rect 15147 18451 15189 18460
rect 16522 18500 16580 18501
rect 16522 18460 16531 18500
rect 16571 18460 16580 18500
rect 16522 18459 16580 18460
rect 18154 18500 18212 18501
rect 18154 18460 18163 18500
rect 18203 18460 18212 18500
rect 18154 18459 18212 18460
rect 24326 18500 24384 18501
rect 24326 18460 24335 18500
rect 24375 18460 24384 18500
rect 24326 18459 24384 18460
rect 26074 18500 26132 18501
rect 26074 18460 26083 18500
rect 26123 18460 26132 18500
rect 26074 18459 26132 18460
rect 27706 18500 27764 18501
rect 27706 18460 27715 18500
rect 27755 18460 27764 18500
rect 27706 18459 27764 18460
rect 30939 18500 30981 18509
rect 30939 18460 30940 18500
rect 30980 18460 30981 18500
rect 30939 18451 30981 18460
rect 4338 18442 4384 18451
rect 11250 18442 11296 18451
rect 5914 18416 5972 18417
rect 5914 18376 5923 18416
rect 5963 18376 5972 18416
rect 5914 18375 5972 18376
rect 7179 18416 7221 18425
rect 7179 18376 7180 18416
rect 7220 18376 7221 18416
rect 7179 18367 7221 18376
rect 12459 18416 12501 18425
rect 12459 18376 12460 18416
rect 12500 18376 12501 18416
rect 12459 18367 12501 18376
rect 15723 18416 15765 18425
rect 15723 18376 15724 18416
rect 15764 18376 15765 18416
rect 15723 18367 15765 18376
rect 18507 18416 18549 18425
rect 18507 18376 18508 18416
rect 18548 18376 18549 18416
rect 18507 18367 18549 18376
rect 23979 18416 24021 18425
rect 23979 18376 23980 18416
rect 24020 18376 24021 18416
rect 23979 18367 24021 18376
rect 24747 18416 24789 18425
rect 24747 18376 24748 18416
rect 24788 18376 24789 18416
rect 24747 18367 24789 18376
rect 26955 18416 26997 18425
rect 26955 18376 26956 18416
rect 26996 18376 26997 18416
rect 26955 18367 26997 18376
rect 29835 18416 29877 18425
rect 29835 18376 29836 18416
rect 29876 18376 29877 18416
rect 29835 18367 29877 18376
rect 1131 18332 1173 18341
rect 1131 18292 1132 18332
rect 1172 18292 1173 18332
rect 1131 18283 1173 18292
rect 3243 18332 3285 18341
rect 3243 18292 3244 18332
rect 3284 18292 3285 18332
rect 3243 18283 3285 18292
rect 16971 18332 17013 18341
rect 16971 18292 16972 18332
rect 17012 18292 17013 18332
rect 16971 18283 17013 18292
rect 22827 18332 22869 18341
rect 22827 18292 22828 18332
rect 22868 18292 22869 18332
rect 22827 18283 22869 18292
rect 24459 18332 24501 18341
rect 24459 18292 24460 18332
rect 24500 18292 24501 18332
rect 24459 18283 24501 18292
rect 25402 18332 25460 18333
rect 25402 18292 25411 18332
rect 25451 18292 25460 18332
rect 25402 18291 25460 18292
rect 25899 18332 25941 18341
rect 25899 18292 25900 18332
rect 25940 18292 25941 18332
rect 25899 18283 25941 18292
rect 27339 18332 27381 18341
rect 27339 18292 27340 18332
rect 27380 18292 27381 18332
rect 27339 18283 27381 18292
rect 576 18164 31392 18188
rect 576 18124 3112 18164
rect 3480 18124 10886 18164
rect 11254 18124 18660 18164
rect 19028 18124 26434 18164
rect 26802 18124 31392 18164
rect 576 18100 31392 18124
rect 6315 17996 6357 18005
rect 6315 17956 6316 17996
rect 6356 17956 6357 17996
rect 6315 17947 6357 17956
rect 6970 17996 7028 17997
rect 6970 17956 6979 17996
rect 7019 17956 7028 17996
rect 6970 17955 7028 17956
rect 7546 17996 7604 17997
rect 7546 17956 7555 17996
rect 7595 17956 7604 17996
rect 7546 17955 7604 17956
rect 11979 17996 12021 18005
rect 11979 17956 11980 17996
rect 12020 17956 12021 17996
rect 11979 17947 12021 17956
rect 12747 17996 12789 18005
rect 12747 17956 12748 17996
rect 12788 17956 12789 17996
rect 12747 17947 12789 17956
rect 22635 17996 22677 18005
rect 22635 17956 22636 17996
rect 22676 17956 22677 17996
rect 22635 17947 22677 17956
rect 23499 17996 23541 18005
rect 23499 17956 23500 17996
rect 23540 17956 23541 17996
rect 23499 17947 23541 17956
rect 24555 17996 24597 18005
rect 24555 17956 24556 17996
rect 24596 17956 24597 17996
rect 24555 17947 24597 17956
rect 26170 17996 26228 17997
rect 26170 17956 26179 17996
rect 26219 17956 26228 17996
rect 26170 17955 26228 17956
rect 27723 17996 27765 18005
rect 27723 17956 27724 17996
rect 27764 17956 27765 17996
rect 27723 17947 27765 17956
rect 1995 17912 2037 17921
rect 1995 17872 1996 17912
rect 2036 17872 2037 17912
rect 1995 17863 2037 17872
rect 2379 17912 2421 17921
rect 2379 17872 2380 17912
rect 2420 17872 2421 17912
rect 2379 17863 2421 17872
rect 3723 17912 3765 17921
rect 3723 17872 3724 17912
rect 3764 17872 3765 17912
rect 3723 17863 3765 17872
rect 4203 17912 4245 17921
rect 4203 17872 4204 17912
rect 4244 17872 4245 17912
rect 4203 17863 4245 17872
rect 7179 17912 7221 17921
rect 7179 17872 7180 17912
rect 7220 17872 7221 17912
rect 7179 17863 7221 17872
rect 9099 17912 9141 17921
rect 9099 17872 9100 17912
rect 9140 17872 9141 17912
rect 9099 17863 9141 17872
rect 11499 17912 11541 17921
rect 11499 17872 11500 17912
rect 11540 17872 11541 17912
rect 11499 17863 11541 17872
rect 20043 17912 20085 17921
rect 20043 17872 20044 17912
rect 20084 17872 20085 17912
rect 20043 17863 20085 17872
rect 24778 17912 24836 17913
rect 24778 17872 24787 17912
rect 24827 17872 24836 17912
rect 24778 17871 24836 17872
rect 2763 17828 2805 17837
rect 2763 17788 2764 17828
rect 2804 17788 2805 17828
rect 2763 17779 2805 17788
rect 8571 17828 8613 17837
rect 8571 17788 8572 17828
rect 8612 17788 8613 17828
rect 8571 17779 8613 17788
rect 9003 17828 9045 17837
rect 9003 17788 9004 17828
rect 9044 17788 9045 17828
rect 9562 17828 9620 17829
rect 9003 17779 9045 17788
rect 9435 17786 9477 17795
rect 9562 17788 9571 17828
rect 9611 17788 9620 17828
rect 9562 17787 9620 17788
rect 9963 17828 10005 17837
rect 9963 17788 9964 17828
rect 10004 17788 10005 17828
rect 6198 17755 6256 17756
rect 2283 17744 2325 17753
rect 2283 17704 2284 17744
rect 2324 17704 2325 17744
rect 2283 17695 2325 17704
rect 2458 17744 2516 17745
rect 2458 17704 2467 17744
rect 2507 17704 2516 17744
rect 2458 17703 2516 17704
rect 2571 17744 2613 17753
rect 2571 17704 2572 17744
rect 2612 17704 2613 17744
rect 2571 17695 2613 17704
rect 2859 17744 2901 17753
rect 2859 17704 2860 17744
rect 2900 17704 2901 17744
rect 2859 17695 2901 17704
rect 2978 17744 3020 17753
rect 2978 17704 2979 17744
rect 3019 17704 3020 17744
rect 2978 17695 3020 17704
rect 3088 17744 3146 17745
rect 3088 17704 3097 17744
rect 3137 17704 3146 17744
rect 3088 17703 3146 17704
rect 3418 17744 3476 17745
rect 3418 17704 3427 17744
rect 3467 17704 3476 17744
rect 3418 17703 3476 17704
rect 3531 17744 3573 17753
rect 3531 17704 3532 17744
rect 3572 17704 3573 17744
rect 3531 17695 3573 17704
rect 4395 17744 4437 17753
rect 4395 17704 4396 17744
rect 4436 17704 4437 17744
rect 4395 17695 4437 17704
rect 4779 17744 4821 17753
rect 4779 17704 4780 17744
rect 4820 17704 4821 17744
rect 4779 17695 4821 17704
rect 4898 17744 4940 17753
rect 4898 17704 4899 17744
rect 4939 17704 4940 17744
rect 4898 17695 4940 17704
rect 5008 17744 5066 17745
rect 5008 17704 5017 17744
rect 5057 17704 5066 17744
rect 5008 17703 5066 17704
rect 5261 17744 5303 17753
rect 5261 17704 5262 17744
rect 5302 17704 5303 17744
rect 5261 17695 5303 17704
rect 5451 17744 5493 17753
rect 5451 17704 5452 17744
rect 5492 17704 5493 17744
rect 5451 17695 5493 17704
rect 5755 17744 5813 17745
rect 5755 17704 5764 17744
rect 5804 17704 5813 17744
rect 5755 17703 5813 17704
rect 5914 17744 5972 17745
rect 5914 17704 5923 17744
rect 5963 17704 5972 17744
rect 5914 17703 5972 17704
rect 6058 17744 6116 17745
rect 6058 17704 6067 17744
rect 6107 17704 6116 17744
rect 6198 17715 6207 17755
rect 6247 17715 6256 17755
rect 6198 17714 6256 17715
rect 6324 17755 6382 17756
rect 6324 17715 6333 17755
rect 6373 17715 6382 17755
rect 6324 17714 6382 17715
rect 6795 17744 6837 17753
rect 6058 17703 6116 17704
rect 6795 17704 6796 17744
rect 6836 17704 6837 17744
rect 6795 17695 6837 17704
rect 6964 17744 7006 17753
rect 6964 17704 6965 17744
rect 7005 17704 7006 17744
rect 6964 17695 7006 17704
rect 7179 17744 7221 17753
rect 7179 17704 7180 17744
rect 7220 17704 7221 17744
rect 7179 17695 7221 17704
rect 7371 17744 7413 17753
rect 7371 17704 7372 17744
rect 7412 17704 7413 17744
rect 7371 17695 7413 17704
rect 7546 17744 7604 17745
rect 7546 17704 7555 17744
rect 7595 17704 7604 17744
rect 7546 17703 7604 17704
rect 7664 17744 7722 17745
rect 7970 17744 8028 17745
rect 7664 17704 7673 17744
rect 7713 17704 7722 17744
rect 7664 17703 7722 17704
rect 7842 17735 7888 17744
rect 7842 17695 7843 17735
rect 7883 17695 7888 17735
rect 7970 17704 7979 17744
rect 8019 17704 8028 17744
rect 7970 17703 8028 17704
rect 8107 17744 8165 17745
rect 8107 17704 8116 17744
rect 8156 17704 8165 17744
rect 8107 17703 8165 17704
rect 8362 17744 8420 17745
rect 8362 17704 8371 17744
rect 8411 17704 8420 17744
rect 8362 17703 8420 17704
rect 8859 17744 8901 17753
rect 8859 17704 8860 17744
rect 8900 17704 8901 17744
rect 8859 17695 8901 17704
rect 9174 17744 9216 17753
rect 9174 17704 9175 17744
rect 9215 17704 9216 17744
rect 9174 17695 9216 17704
rect 9314 17744 9356 17753
rect 9314 17704 9315 17744
rect 9355 17704 9356 17744
rect 9435 17746 9436 17786
rect 9476 17746 9477 17786
rect 9963 17779 10005 17788
rect 11115 17828 11157 17837
rect 11115 17788 11116 17828
rect 11156 17788 11157 17828
rect 11115 17779 11157 17788
rect 13634 17828 13676 17837
rect 13634 17788 13635 17828
rect 13675 17788 13676 17828
rect 13634 17779 13676 17788
rect 14114 17828 14156 17837
rect 14114 17788 14115 17828
rect 14155 17788 14156 17828
rect 14114 17779 14156 17788
rect 14458 17828 14516 17829
rect 14458 17788 14467 17828
rect 14507 17788 14516 17828
rect 14458 17787 14516 17788
rect 15147 17828 15189 17837
rect 15147 17788 15148 17828
rect 15188 17788 15189 17828
rect 15147 17779 15189 17788
rect 16138 17828 16196 17829
rect 16138 17788 16147 17828
rect 16187 17788 16196 17828
rect 16138 17787 16196 17788
rect 18868 17828 18910 17837
rect 18868 17788 18869 17828
rect 18909 17788 18910 17828
rect 18868 17779 18910 17788
rect 19083 17828 19125 17837
rect 19083 17788 19084 17828
rect 19124 17788 19125 17828
rect 19083 17779 19125 17788
rect 20986 17828 21044 17829
rect 20986 17788 20995 17828
rect 21035 17788 21044 17828
rect 20986 17787 21044 17788
rect 25611 17828 25653 17837
rect 25611 17788 25612 17828
rect 25652 17788 25653 17828
rect 19594 17786 19652 17787
rect 9435 17737 9477 17746
rect 9656 17744 9698 17753
rect 9314 17695 9356 17704
rect 9656 17704 9657 17744
rect 9697 17704 9698 17744
rect 9656 17695 9698 17704
rect 10639 17744 10697 17745
rect 10639 17704 10648 17744
rect 10688 17704 10697 17744
rect 10639 17703 10697 17704
rect 10774 17744 10816 17753
rect 10774 17704 10775 17744
rect 10815 17704 10816 17744
rect 10774 17695 10816 17704
rect 10906 17744 10964 17745
rect 10906 17704 10915 17744
rect 10955 17704 10964 17744
rect 10906 17703 10964 17704
rect 11019 17744 11061 17753
rect 11019 17704 11020 17744
rect 11060 17704 11061 17744
rect 11019 17695 11061 17704
rect 11499 17744 11541 17753
rect 11499 17704 11500 17744
rect 11540 17704 11541 17744
rect 11499 17695 11541 17704
rect 11691 17744 11733 17753
rect 11691 17704 11692 17744
rect 11732 17704 11733 17744
rect 11691 17695 11733 17704
rect 11872 17744 11914 17753
rect 11872 17704 11873 17744
rect 11913 17704 11914 17744
rect 11872 17695 11914 17704
rect 12076 17744 12134 17745
rect 12076 17704 12085 17744
rect 12125 17704 12134 17744
rect 12076 17703 12134 17704
rect 12267 17744 12309 17753
rect 12267 17704 12268 17744
rect 12308 17704 12309 17744
rect 12267 17695 12309 17704
rect 12442 17744 12500 17745
rect 12442 17704 12451 17744
rect 12491 17704 12500 17744
rect 12442 17703 12500 17704
rect 12651 17744 12693 17753
rect 12651 17704 12652 17744
rect 12692 17704 12693 17744
rect 13035 17744 13077 17753
rect 12651 17695 12693 17704
rect 12830 17717 12888 17718
rect 7842 17686 7888 17695
rect 12830 17677 12839 17717
rect 12879 17677 12888 17717
rect 13035 17704 13036 17744
rect 13076 17704 13077 17744
rect 13035 17695 13077 17704
rect 13225 17744 13267 17753
rect 13225 17704 13226 17744
rect 13266 17704 13267 17744
rect 13225 17695 13267 17704
rect 13515 17744 13557 17753
rect 13515 17704 13516 17744
rect 13556 17704 13557 17744
rect 13515 17695 13557 17704
rect 13732 17744 13774 17753
rect 13732 17704 13733 17744
rect 13773 17704 13774 17744
rect 13732 17695 13774 17704
rect 13995 17744 14037 17753
rect 13995 17704 13996 17744
rect 14036 17704 14037 17744
rect 13995 17695 14037 17704
rect 14212 17744 14254 17753
rect 14212 17704 14213 17744
rect 14253 17704 14254 17744
rect 14212 17695 14254 17704
rect 14326 17744 14368 17753
rect 14326 17704 14327 17744
rect 14367 17704 14368 17744
rect 14326 17695 14368 17704
rect 14571 17744 14613 17753
rect 14571 17704 14572 17744
rect 14612 17704 14613 17744
rect 14571 17695 14613 17704
rect 14806 17744 14848 17753
rect 14806 17704 14807 17744
rect 14847 17704 14848 17744
rect 14806 17695 14848 17704
rect 14938 17744 14996 17745
rect 14938 17704 14947 17744
rect 14987 17704 14996 17744
rect 14938 17703 14996 17704
rect 15051 17744 15093 17753
rect 15051 17704 15052 17744
rect 15092 17704 15093 17744
rect 15051 17695 15093 17704
rect 15483 17744 15525 17753
rect 15483 17704 15484 17744
rect 15524 17704 15525 17744
rect 15483 17695 15525 17704
rect 15610 17744 15668 17745
rect 15610 17704 15619 17744
rect 15659 17704 15668 17744
rect 15610 17703 15668 17704
rect 15723 17744 15765 17753
rect 15723 17704 15724 17744
rect 15764 17704 15765 17744
rect 15723 17695 15765 17704
rect 16303 17744 16361 17745
rect 16303 17704 16312 17744
rect 16352 17704 16361 17744
rect 16303 17703 16361 17704
rect 16474 17744 16532 17745
rect 16474 17704 16483 17744
rect 16523 17704 16532 17744
rect 16474 17703 16532 17704
rect 16775 17744 16817 17753
rect 16775 17704 16776 17744
rect 16816 17704 16817 17744
rect 16775 17695 16817 17704
rect 16954 17744 17012 17745
rect 16954 17704 16963 17744
rect 17003 17704 17012 17744
rect 16954 17703 17012 17704
rect 17072 17744 17130 17745
rect 17072 17704 17081 17744
rect 17121 17704 17130 17744
rect 17072 17703 17130 17704
rect 17247 17744 17289 17753
rect 17247 17704 17248 17744
rect 17288 17704 17289 17744
rect 17247 17695 17289 17704
rect 17346 17744 17404 17745
rect 17346 17704 17355 17744
rect 17395 17704 17404 17744
rect 17346 17703 17404 17704
rect 17515 17744 17573 17745
rect 17515 17704 17524 17744
rect 17564 17704 17573 17744
rect 17515 17703 17573 17704
rect 17835 17744 17877 17753
rect 17835 17704 17836 17744
rect 17876 17704 17877 17744
rect 17835 17695 17877 17704
rect 18262 17744 18304 17753
rect 18262 17704 18263 17744
rect 18303 17704 18304 17744
rect 18262 17695 18304 17704
rect 18388 17744 18430 17753
rect 18388 17704 18389 17744
rect 18429 17704 18430 17744
rect 18388 17695 18430 17704
rect 18492 17744 18550 17745
rect 18492 17704 18501 17744
rect 18541 17704 18550 17744
rect 18492 17703 18550 17704
rect 18742 17744 18784 17753
rect 18742 17704 18743 17744
rect 18783 17704 18784 17744
rect 18742 17695 18784 17704
rect 18987 17744 19029 17753
rect 19594 17746 19603 17786
rect 19643 17746 19652 17786
rect 23742 17777 23784 17786
rect 25611 17779 25653 17788
rect 27706 17828 27764 17829
rect 27706 17788 27715 17828
rect 27755 17788 27764 17828
rect 27706 17787 27764 17788
rect 28090 17828 28148 17829
rect 28090 17788 28099 17828
rect 28139 17788 28148 17828
rect 28090 17787 28148 17788
rect 19594 17745 19652 17746
rect 18987 17704 18988 17744
rect 19028 17704 19029 17744
rect 18987 17695 19029 17704
rect 20043 17744 20085 17753
rect 20043 17704 20044 17744
rect 20084 17704 20085 17744
rect 20043 17695 20085 17704
rect 20160 17744 20218 17745
rect 20160 17704 20169 17744
rect 20209 17704 20218 17744
rect 20160 17703 20218 17704
rect 20331 17744 20373 17753
rect 20331 17704 20332 17744
rect 20372 17704 20373 17744
rect 20331 17695 20373 17704
rect 20506 17744 20564 17745
rect 20506 17704 20515 17744
rect 20555 17704 20564 17744
rect 20506 17703 20564 17704
rect 20811 17744 20853 17753
rect 20811 17704 20812 17744
rect 20852 17704 20853 17744
rect 20811 17695 20853 17704
rect 21675 17744 21717 17753
rect 21675 17704 21676 17744
rect 21716 17704 21717 17744
rect 21675 17695 21717 17704
rect 21963 17744 22005 17753
rect 21963 17704 21964 17744
rect 22004 17704 22005 17744
rect 21963 17695 22005 17704
rect 22155 17744 22197 17753
rect 22155 17704 22156 17744
rect 22196 17704 22197 17744
rect 22155 17695 22197 17704
rect 22810 17744 22868 17745
rect 22810 17704 22819 17744
rect 22859 17704 22868 17744
rect 22810 17703 22868 17704
rect 22915 17744 22973 17745
rect 22915 17704 22924 17744
rect 22964 17704 22973 17744
rect 22915 17703 22973 17704
rect 23050 17744 23108 17745
rect 23050 17704 23059 17744
rect 23099 17704 23108 17744
rect 23050 17703 23108 17704
rect 23211 17744 23253 17753
rect 23211 17704 23212 17744
rect 23252 17704 23253 17744
rect 23211 17695 23253 17704
rect 23403 17744 23445 17753
rect 23403 17704 23404 17744
rect 23444 17704 23445 17744
rect 23403 17695 23445 17704
rect 23517 17744 23575 17745
rect 23517 17704 23526 17744
rect 23566 17704 23575 17744
rect 23517 17703 23575 17704
rect 23643 17744 23685 17753
rect 23643 17704 23644 17744
rect 23684 17704 23685 17744
rect 23742 17737 23743 17777
rect 23783 17737 23784 17777
rect 23742 17728 23784 17737
rect 23979 17744 24021 17753
rect 23643 17695 23685 17704
rect 23979 17704 23980 17744
rect 24020 17704 24021 17744
rect 23979 17695 24021 17704
rect 24171 17744 24213 17753
rect 24171 17704 24172 17744
rect 24212 17704 24213 17744
rect 24171 17695 24213 17704
rect 24406 17744 24448 17753
rect 24651 17744 24693 17753
rect 24406 17704 24407 17744
rect 24447 17704 24448 17744
rect 24406 17695 24448 17704
rect 24546 17735 24592 17744
rect 24546 17695 24547 17735
rect 24587 17695 24592 17735
rect 24651 17704 24652 17744
rect 24692 17704 24693 17744
rect 24651 17695 24693 17704
rect 24987 17744 25029 17753
rect 24987 17704 24988 17744
rect 25028 17704 25029 17744
rect 24987 17695 25029 17704
rect 25131 17744 25173 17753
rect 25131 17704 25132 17744
rect 25172 17704 25173 17744
rect 25131 17695 25173 17704
rect 25707 17744 25749 17753
rect 25707 17704 25708 17744
rect 25748 17704 25749 17744
rect 25707 17695 25749 17704
rect 25826 17744 25868 17753
rect 25826 17704 25827 17744
rect 25867 17704 25868 17744
rect 25826 17695 25868 17704
rect 25938 17744 25980 17753
rect 25938 17704 25939 17744
rect 25979 17704 25980 17744
rect 25938 17695 25980 17704
rect 26571 17744 26613 17753
rect 26571 17704 26572 17744
rect 26612 17704 26613 17744
rect 26571 17695 26613 17704
rect 26842 17744 26900 17745
rect 26842 17704 26851 17744
rect 26891 17704 26900 17744
rect 26842 17703 26900 17704
rect 27531 17744 27573 17753
rect 27531 17704 27532 17744
rect 27572 17704 27573 17744
rect 27531 17695 27573 17704
rect 29626 17744 29684 17745
rect 29626 17704 29635 17744
rect 29675 17704 29684 17744
rect 29626 17703 29684 17704
rect 30199 17744 30257 17745
rect 30199 17704 30208 17744
rect 30248 17704 30257 17744
rect 30199 17703 30257 17704
rect 30679 17744 30737 17745
rect 30679 17704 30688 17744
rect 30728 17704 30737 17744
rect 30679 17703 30737 17704
rect 24546 17686 24592 17695
rect 12830 17676 12888 17677
rect 4683 17660 4725 17669
rect 4683 17620 4684 17660
rect 4724 17620 4725 17660
rect 4683 17611 4725 17620
rect 10474 17660 10532 17661
rect 10474 17620 10483 17660
rect 10523 17620 10532 17660
rect 10474 17619 10532 17620
rect 13899 17660 13941 17669
rect 13899 17620 13900 17660
rect 13940 17620 13941 17660
rect 13899 17611 13941 17620
rect 15802 17660 15860 17661
rect 15802 17620 15811 17660
rect 15851 17620 15860 17660
rect 15802 17619 15860 17620
rect 16683 17660 16725 17669
rect 16683 17620 16684 17660
rect 16724 17620 16725 17660
rect 16683 17611 16725 17620
rect 22042 17660 22100 17661
rect 22042 17620 22051 17660
rect 22091 17620 22100 17660
rect 22042 17619 22100 17620
rect 30010 17660 30068 17661
rect 30010 17620 30019 17660
rect 30059 17620 30068 17660
rect 30010 17619 30068 17620
rect 3435 17576 3477 17585
rect 3435 17536 3436 17576
rect 3476 17536 3477 17576
rect 3435 17527 3477 17536
rect 5451 17576 5493 17585
rect 5451 17536 5452 17576
rect 5492 17536 5493 17576
rect 5451 17527 5493 17536
rect 9754 17576 9812 17577
rect 9754 17536 9763 17576
rect 9803 17536 9812 17576
rect 9754 17535 9812 17536
rect 10203 17576 10245 17585
rect 10203 17536 10204 17576
rect 10244 17536 10245 17576
rect 10203 17527 10245 17536
rect 12363 17576 12405 17585
rect 12363 17536 12364 17576
rect 12404 17536 12405 17576
rect 12363 17527 12405 17536
rect 13131 17576 13173 17585
rect 13131 17536 13132 17576
rect 13172 17536 13173 17576
rect 13131 17527 13173 17536
rect 13419 17576 13461 17585
rect 13419 17536 13420 17576
rect 13460 17536 13461 17576
rect 13419 17527 13461 17536
rect 14650 17576 14708 17577
rect 14650 17536 14659 17576
rect 14699 17536 14708 17576
rect 14650 17535 14708 17536
rect 17434 17576 17492 17577
rect 17434 17536 17443 17576
rect 17483 17536 17492 17576
rect 17434 17535 17492 17536
rect 17722 17576 17780 17577
rect 17722 17536 17731 17576
rect 17771 17536 17780 17576
rect 17722 17535 17780 17536
rect 18010 17576 18068 17577
rect 18010 17536 18019 17576
rect 18059 17536 18068 17576
rect 18010 17535 18068 17536
rect 18586 17576 18644 17577
rect 18586 17536 18595 17576
rect 18635 17536 18644 17576
rect 18586 17535 18644 17536
rect 19402 17576 19460 17577
rect 19402 17536 19411 17576
rect 19451 17536 19460 17576
rect 19402 17535 19460 17536
rect 20715 17576 20757 17585
rect 20715 17536 20716 17576
rect 20756 17536 20757 17576
rect 20715 17527 20757 17536
rect 23979 17576 24021 17585
rect 23979 17536 23980 17576
rect 24020 17536 24021 17576
rect 23979 17527 24021 17536
rect 26379 17576 26421 17585
rect 26379 17536 26380 17576
rect 26420 17536 26421 17576
rect 26379 17527 26421 17536
rect 30363 17576 30405 17585
rect 30363 17536 30364 17576
rect 30404 17536 30405 17576
rect 30363 17527 30405 17536
rect 30843 17576 30885 17585
rect 30843 17536 30844 17576
rect 30884 17536 30885 17576
rect 30843 17527 30885 17536
rect 576 17408 31392 17432
rect 576 17368 4352 17408
rect 4720 17368 12126 17408
rect 12494 17368 19900 17408
rect 20268 17368 27674 17408
rect 28042 17368 31392 17408
rect 576 17344 31392 17368
rect 2170 17240 2228 17241
rect 2170 17200 2179 17240
rect 2219 17200 2228 17240
rect 2170 17199 2228 17200
rect 3322 17240 3380 17241
rect 3322 17200 3331 17240
rect 3371 17200 3380 17240
rect 3322 17199 3380 17200
rect 4282 17240 4340 17241
rect 4282 17200 4291 17240
rect 4331 17200 4340 17240
rect 4282 17199 4340 17200
rect 4474 17240 4532 17241
rect 4474 17200 4483 17240
rect 4523 17200 4532 17240
rect 4474 17199 4532 17200
rect 4954 17240 5012 17241
rect 4954 17200 4963 17240
rect 5003 17200 5012 17240
rect 4954 17199 5012 17200
rect 8314 17240 8372 17241
rect 8314 17200 8323 17240
rect 8363 17200 8372 17240
rect 8314 17199 8372 17200
rect 8794 17240 8852 17241
rect 8794 17200 8803 17240
rect 8843 17200 8852 17240
rect 8794 17199 8852 17200
rect 12730 17240 12788 17241
rect 12730 17200 12739 17240
rect 12779 17200 12788 17240
rect 12730 17199 12788 17200
rect 13882 17240 13940 17241
rect 13882 17200 13891 17240
rect 13931 17200 13940 17240
rect 13882 17199 13940 17200
rect 15898 17240 15956 17241
rect 15898 17200 15907 17240
rect 15947 17200 15956 17240
rect 15898 17199 15956 17200
rect 16299 17240 16341 17249
rect 16299 17200 16300 17240
rect 16340 17200 16341 17240
rect 16299 17191 16341 17200
rect 16762 17240 16820 17241
rect 16762 17200 16771 17240
rect 16811 17200 16820 17240
rect 16762 17199 16820 17200
rect 17716 17240 17774 17241
rect 17716 17200 17725 17240
rect 17765 17200 17774 17240
rect 17716 17199 17774 17200
rect 18891 17240 18933 17249
rect 18891 17200 18892 17240
rect 18932 17200 18933 17240
rect 18891 17191 18933 17200
rect 20602 17240 20660 17241
rect 20602 17200 20611 17240
rect 20651 17200 20660 17240
rect 20602 17199 20660 17200
rect 21195 17240 21237 17249
rect 21195 17200 21196 17240
rect 21236 17200 21237 17240
rect 21195 17191 21237 17200
rect 21946 17240 22004 17241
rect 21946 17200 21955 17240
rect 21995 17200 22004 17240
rect 21946 17199 22004 17200
rect 25131 17240 25173 17249
rect 25131 17200 25132 17240
rect 25172 17200 25173 17240
rect 25131 17191 25173 17200
rect 26164 17240 26222 17241
rect 26164 17200 26173 17240
rect 26213 17200 26222 17240
rect 26164 17199 26222 17200
rect 27147 17240 27189 17249
rect 27147 17200 27148 17240
rect 27188 17200 27189 17240
rect 27147 17191 27189 17200
rect 27531 17240 27573 17249
rect 27531 17200 27532 17240
rect 27572 17200 27573 17240
rect 27531 17191 27573 17200
rect 29547 17240 29589 17249
rect 29547 17200 29548 17240
rect 29588 17200 29589 17240
rect 29547 17191 29589 17200
rect 29722 17240 29780 17241
rect 29722 17200 29731 17240
rect 29771 17200 29780 17240
rect 29722 17199 29780 17200
rect 30027 17240 30069 17249
rect 30027 17200 30028 17240
rect 30068 17200 30069 17240
rect 30027 17191 30069 17200
rect 3034 17156 3092 17157
rect 3034 17116 3043 17156
rect 3083 17116 3092 17156
rect 3034 17115 3092 17116
rect 3802 17156 3860 17157
rect 6699 17156 6741 17165
rect 3802 17116 3811 17156
rect 3851 17116 3860 17156
rect 3802 17115 3860 17116
rect 5250 17147 5296 17156
rect 5250 17107 5251 17147
rect 5291 17107 5296 17147
rect 5250 17098 5296 17107
rect 6018 17147 6064 17156
rect 6018 17107 6019 17147
rect 6059 17107 6064 17147
rect 6699 17116 6700 17156
rect 6740 17116 6741 17156
rect 6699 17107 6741 17116
rect 10539 17156 10581 17165
rect 10539 17116 10540 17156
rect 10580 17116 10581 17156
rect 10539 17107 10581 17116
rect 13611 17156 13653 17165
rect 18490 17156 18548 17157
rect 13611 17116 13612 17156
rect 13652 17116 13653 17156
rect 13611 17107 13653 17116
rect 14178 17147 14224 17156
rect 14178 17107 14179 17147
rect 14219 17107 14224 17147
rect 6018 17098 6064 17107
rect 14178 17098 14224 17107
rect 15714 17147 15760 17156
rect 15714 17107 15715 17147
rect 15755 17107 15760 17147
rect 18490 17116 18499 17156
rect 18539 17116 18548 17156
rect 18490 17115 18548 17116
rect 19659 17156 19701 17165
rect 19659 17116 19660 17156
rect 19700 17116 19701 17156
rect 19659 17107 19701 17116
rect 21305 17156 21347 17165
rect 21305 17116 21306 17156
rect 21346 17116 21347 17156
rect 21305 17107 21347 17116
rect 22635 17156 22677 17165
rect 22635 17116 22636 17156
rect 22676 17116 22677 17156
rect 22635 17107 22677 17116
rect 26698 17156 26756 17157
rect 26698 17116 26707 17156
rect 26747 17116 26756 17156
rect 26698 17115 26756 17116
rect 15714 17098 15760 17107
rect 2283 17072 2325 17081
rect 2283 17032 2284 17072
rect 2324 17032 2325 17072
rect 2283 17023 2325 17032
rect 3243 17072 3285 17081
rect 3243 17032 3244 17072
rect 3284 17032 3285 17072
rect 3243 17023 3285 17032
rect 3478 17072 3520 17081
rect 3478 17032 3479 17072
rect 3519 17032 3520 17072
rect 3478 17023 3520 17032
rect 3723 17072 3765 17081
rect 3723 17032 3724 17072
rect 3764 17032 3765 17072
rect 3723 17023 3765 17032
rect 4203 17072 4245 17081
rect 4203 17032 4204 17072
rect 4244 17032 4245 17072
rect 4203 17023 4245 17032
rect 4587 17072 4629 17081
rect 4587 17032 4588 17072
rect 4628 17032 4629 17072
rect 4587 17023 4629 17032
rect 4954 17072 5012 17073
rect 5338 17072 5396 17073
rect 4954 17032 4963 17072
rect 5003 17032 5012 17072
rect 4954 17031 5012 17032
rect 5067 17063 5109 17072
rect 5067 17023 5068 17063
rect 5108 17023 5109 17063
rect 5338 17032 5347 17072
rect 5387 17032 5396 17072
rect 5338 17031 5396 17032
rect 5472 17072 5530 17073
rect 5472 17032 5481 17072
rect 5521 17032 5530 17072
rect 5472 17031 5530 17032
rect 5733 17072 5791 17073
rect 5733 17032 5742 17072
rect 5782 17032 5791 17072
rect 5733 17031 5791 17032
rect 5878 17072 5936 17073
rect 5878 17032 5887 17072
rect 5927 17032 5936 17072
rect 5878 17031 5936 17032
rect 6106 17072 6164 17073
rect 6106 17032 6115 17072
rect 6155 17032 6164 17072
rect 6106 17031 6164 17032
rect 6282 17072 6340 17073
rect 6795 17072 6837 17081
rect 6282 17032 6291 17072
rect 6331 17032 6340 17072
rect 6282 17031 6340 17032
rect 6490 17071 6548 17072
rect 6490 17031 6499 17071
rect 6539 17031 6548 17071
rect 6490 17030 6548 17031
rect 6795 17032 6796 17072
rect 6836 17032 6837 17072
rect 6795 17023 6837 17032
rect 7066 17072 7124 17073
rect 7453 17072 7495 17081
rect 7066 17032 7075 17072
rect 7115 17032 7124 17072
rect 7066 17031 7124 17032
rect 7179 17063 7221 17072
rect 7179 17023 7180 17063
rect 7220 17023 7221 17063
rect 5067 17014 5109 17023
rect 7179 17014 7221 17023
rect 7323 17063 7365 17072
rect 7323 17023 7324 17063
rect 7364 17023 7365 17063
rect 7453 17032 7454 17072
rect 7494 17032 7495 17072
rect 7453 17023 7495 17032
rect 7627 17072 7685 17073
rect 7627 17032 7636 17072
rect 7676 17032 7685 17072
rect 7627 17031 7685 17032
rect 7975 17072 8033 17073
rect 7975 17032 7984 17072
rect 8024 17032 8033 17072
rect 7975 17031 8033 17032
rect 8153 17072 8195 17081
rect 8153 17032 8154 17072
rect 8194 17032 8195 17072
rect 8153 17023 8195 17032
rect 8266 17072 8324 17073
rect 8266 17032 8275 17072
rect 8315 17032 8324 17072
rect 8731 17072 8789 17073
rect 8266 17031 8324 17032
rect 8395 17061 8437 17070
rect 7323 17014 7365 17023
rect 8395 17021 8396 17061
rect 8436 17021 8437 17061
rect 8395 17012 8437 17021
rect 8532 17061 8590 17062
rect 8532 17021 8541 17061
rect 8581 17021 8590 17061
rect 8731 17032 8740 17072
rect 8780 17032 8789 17072
rect 8731 17031 8789 17032
rect 8890 17072 8948 17073
rect 8890 17032 8899 17072
rect 8939 17032 8948 17072
rect 8890 17031 8948 17032
rect 9015 17072 9057 17081
rect 9015 17032 9016 17072
rect 9056 17032 9057 17072
rect 9015 17023 9057 17032
rect 9146 17072 9204 17073
rect 9146 17032 9155 17072
rect 9195 17032 9204 17072
rect 9146 17031 9204 17032
rect 9274 17072 9332 17073
rect 9274 17032 9283 17072
rect 9323 17032 9332 17072
rect 9274 17031 9332 17032
rect 9531 17072 9573 17081
rect 9531 17032 9532 17072
rect 9572 17032 9573 17072
rect 9994 17072 10052 17073
rect 9531 17023 9573 17032
rect 9675 17030 9717 17039
rect 9994 17032 10003 17072
rect 10043 17032 10052 17072
rect 9994 17031 10052 17032
rect 10618 17072 10676 17073
rect 10618 17032 10627 17072
rect 10667 17032 10676 17072
rect 10618 17031 10676 17032
rect 11019 17072 11061 17081
rect 11019 17032 11020 17072
rect 11060 17032 11061 17072
rect 8532 17020 8590 17021
rect 9675 16990 9676 17030
rect 9716 16990 9717 17030
rect 11019 17023 11061 17032
rect 11503 17072 11561 17073
rect 11503 17032 11512 17072
rect 11552 17032 11561 17072
rect 11503 17031 11561 17032
rect 11691 17072 11733 17081
rect 11691 17032 11692 17072
rect 11732 17032 11733 17072
rect 11691 17023 11733 17032
rect 12058 17072 12116 17073
rect 12058 17032 12067 17072
rect 12107 17032 12116 17072
rect 12058 17031 12116 17032
rect 12171 17072 12213 17081
rect 12171 17032 12172 17072
rect 12212 17032 12213 17072
rect 12171 17023 12213 17032
rect 12538 17072 12596 17073
rect 12538 17032 12547 17072
rect 12587 17032 12596 17072
rect 12538 17031 12596 17032
rect 12970 17072 13028 17073
rect 12970 17032 12979 17072
rect 13019 17032 13028 17072
rect 12970 17031 13028 17032
rect 13515 17072 13557 17081
rect 13515 17032 13516 17072
rect 13556 17032 13557 17072
rect 13515 17023 13557 17032
rect 13707 17072 13749 17081
rect 13707 17032 13708 17072
rect 13748 17032 13749 17072
rect 13707 17023 13749 17032
rect 13882 17072 13940 17073
rect 14266 17072 14324 17073
rect 13882 17032 13891 17072
rect 13931 17032 13940 17072
rect 13882 17031 13940 17032
rect 13995 17063 14037 17072
rect 13995 17023 13996 17063
rect 14036 17023 14037 17063
rect 14266 17032 14275 17072
rect 14315 17032 14324 17072
rect 14266 17031 14324 17032
rect 14400 17072 14458 17073
rect 14400 17032 14409 17072
rect 14449 17032 14458 17072
rect 14400 17031 14458 17032
rect 15247 17072 15305 17073
rect 15247 17032 15256 17072
rect 15296 17032 15305 17072
rect 15247 17031 15305 17032
rect 15429 17072 15487 17073
rect 15798 17072 15856 17073
rect 15429 17032 15438 17072
rect 15478 17032 15487 17072
rect 15429 17031 15487 17032
rect 15531 17063 15573 17072
rect 13995 17014 14037 17023
rect 15531 17023 15532 17063
rect 15572 17023 15573 17063
rect 15798 17032 15807 17072
rect 15847 17032 15856 17072
rect 15798 17031 15856 17032
rect 15979 17072 16037 17073
rect 15979 17032 15988 17072
rect 16028 17032 16037 17072
rect 15979 17031 16037 17032
rect 16210 17072 16268 17073
rect 16210 17032 16219 17072
rect 16259 17032 16268 17072
rect 16210 17031 16268 17032
rect 16395 17072 16437 17081
rect 16395 17032 16396 17072
rect 16436 17032 16437 17072
rect 16395 17023 16437 17032
rect 16603 17072 16661 17073
rect 16603 17032 16612 17072
rect 16652 17032 16661 17072
rect 16603 17031 16661 17032
rect 16762 17072 16820 17073
rect 16762 17032 16771 17072
rect 16811 17032 16820 17072
rect 16762 17031 16820 17032
rect 16887 17072 16929 17081
rect 17146 17072 17204 17073
rect 16887 17032 16888 17072
rect 16928 17032 16929 17072
rect 16887 17023 16929 17032
rect 17019 17063 17061 17072
rect 17019 17023 17020 17063
rect 17060 17023 17061 17063
rect 17146 17032 17155 17072
rect 17195 17032 17204 17072
rect 17146 17031 17204 17032
rect 17355 17072 17397 17081
rect 17355 17032 17356 17072
rect 17396 17032 17397 17072
rect 17355 17023 17397 17032
rect 17547 17072 17589 17081
rect 17547 17032 17548 17072
rect 17588 17032 17589 17072
rect 17547 17023 17589 17032
rect 17818 17072 17876 17073
rect 18397 17072 18439 17081
rect 17818 17032 17827 17072
rect 17867 17032 17876 17072
rect 17818 17031 17876 17032
rect 17931 17063 17973 17072
rect 17931 17023 17932 17063
rect 17972 17023 17973 17063
rect 18397 17032 18398 17072
rect 18438 17032 18439 17072
rect 18397 17023 18439 17032
rect 18603 17072 18645 17081
rect 18934 17072 18976 17081
rect 19179 17072 19221 17081
rect 18603 17032 18604 17072
rect 18644 17032 18645 17072
rect 18603 17023 18645 17032
rect 18699 17063 18741 17072
rect 18699 17023 18700 17063
rect 18740 17023 18741 17063
rect 18934 17032 18935 17072
rect 18975 17032 18976 17072
rect 18934 17023 18976 17032
rect 19074 17063 19120 17072
rect 19074 17023 19075 17063
rect 19115 17023 19120 17063
rect 19179 17032 19180 17072
rect 19220 17032 19221 17072
rect 19179 17023 19221 17032
rect 19467 17072 19509 17081
rect 19467 17032 19468 17072
rect 19508 17032 19509 17072
rect 19467 17023 19509 17032
rect 19786 17072 19844 17073
rect 19786 17032 19795 17072
rect 19835 17032 19844 17072
rect 19786 17031 19844 17032
rect 20251 17072 20309 17073
rect 20251 17032 20260 17072
rect 20300 17032 20309 17072
rect 20251 17031 20309 17032
rect 20410 17072 20468 17073
rect 20410 17032 20419 17072
rect 20459 17032 20468 17072
rect 20410 17031 20468 17032
rect 20535 17072 20577 17081
rect 20794 17072 20852 17073
rect 20535 17032 20536 17072
rect 20576 17032 20577 17072
rect 20535 17023 20577 17032
rect 20667 17063 20709 17072
rect 20667 17023 20668 17063
rect 20708 17023 20709 17063
rect 20794 17032 20803 17072
rect 20843 17032 20852 17072
rect 20794 17031 20852 17032
rect 20986 17072 21044 17073
rect 20986 17032 20995 17072
rect 21035 17032 21044 17072
rect 20986 17031 21044 17032
rect 21099 17072 21141 17081
rect 21099 17032 21100 17072
rect 21140 17032 21141 17072
rect 21099 17023 21141 17032
rect 21867 17072 21909 17081
rect 21867 17032 21868 17072
rect 21908 17032 21909 17072
rect 21867 17023 21909 17032
rect 22155 17072 22197 17081
rect 22155 17032 22156 17072
rect 22196 17032 22197 17072
rect 22155 17023 22197 17032
rect 22539 17072 22581 17081
rect 22539 17032 22540 17072
rect 22580 17032 22581 17072
rect 22539 17023 22581 17032
rect 22827 17072 22869 17081
rect 22827 17032 22828 17072
rect 22868 17032 22869 17072
rect 22827 17023 22869 17032
rect 23019 17072 23061 17081
rect 23019 17032 23020 17072
rect 23060 17032 23061 17072
rect 23019 17023 23061 17032
rect 23350 17072 23408 17073
rect 23350 17032 23359 17072
rect 23399 17032 23408 17072
rect 23350 17031 23408 17032
rect 23595 17072 23637 17081
rect 23595 17032 23596 17072
rect 23636 17032 23637 17072
rect 23595 17023 23637 17032
rect 23787 17072 23829 17081
rect 23787 17032 23788 17072
rect 23828 17032 23829 17072
rect 23787 17023 23829 17032
rect 24126 17072 24184 17073
rect 24359 17072 24417 17073
rect 24126 17032 24135 17072
rect 24175 17032 24184 17072
rect 24126 17031 24184 17032
rect 24258 17063 24304 17072
rect 24258 17023 24259 17063
rect 24299 17023 24304 17063
rect 24359 17032 24368 17072
rect 24408 17032 24417 17072
rect 24359 17031 24417 17032
rect 24651 17072 24693 17081
rect 24651 17032 24652 17072
rect 24692 17032 24693 17072
rect 24651 17023 24693 17032
rect 24768 17072 24826 17073
rect 24768 17032 24777 17072
rect 24817 17032 24826 17072
rect 24768 17031 24826 17032
rect 24939 17072 24981 17081
rect 24939 17032 24940 17072
rect 24980 17032 24981 17072
rect 24939 17023 24981 17032
rect 25227 17072 25269 17081
rect 25227 17032 25228 17072
rect 25268 17032 25269 17072
rect 25227 17023 25269 17032
rect 25456 17072 25514 17073
rect 25456 17032 25465 17072
rect 25505 17032 25514 17072
rect 25456 17031 25514 17032
rect 25707 17072 25749 17081
rect 25707 17032 25708 17072
rect 25748 17032 25749 17072
rect 25707 17023 25749 17032
rect 25821 17072 25879 17073
rect 25821 17032 25830 17072
rect 25870 17032 25879 17072
rect 25821 17031 25879 17032
rect 25948 17072 26006 17073
rect 25948 17032 25957 17072
rect 25997 17032 26006 17072
rect 25948 17031 26006 17032
rect 26266 17072 26324 17073
rect 27051 17072 27093 17081
rect 26266 17032 26275 17072
rect 26315 17032 26324 17072
rect 26266 17031 26324 17032
rect 26379 17063 26421 17072
rect 26379 17023 26380 17063
rect 26420 17023 26421 17063
rect 27051 17032 27052 17072
rect 27092 17032 27093 17072
rect 27051 17023 27093 17032
rect 27172 17072 27214 17081
rect 27172 17032 27173 17072
rect 27213 17032 27214 17072
rect 27172 17023 27214 17032
rect 27574 17072 27616 17081
rect 27574 17032 27575 17072
rect 27615 17032 27616 17072
rect 27574 17023 27616 17032
rect 27688 17072 27746 17073
rect 27688 17032 27697 17072
rect 27737 17032 27746 17072
rect 27688 17031 27746 17032
rect 27819 17072 27861 17081
rect 27819 17032 27820 17072
rect 27860 17032 27861 17072
rect 27819 17023 27861 17032
rect 28683 17072 28725 17081
rect 28683 17032 28684 17072
rect 28724 17032 28725 17072
rect 28683 17023 28725 17032
rect 28875 17072 28917 17081
rect 28875 17032 28876 17072
rect 28916 17032 28917 17072
rect 28875 17023 28917 17032
rect 29835 17072 29877 17081
rect 29835 17032 29836 17072
rect 29876 17032 29877 17072
rect 29835 17023 29877 17032
rect 30219 17072 30261 17081
rect 30219 17032 30220 17072
rect 30260 17032 30261 17072
rect 30219 17023 30261 17032
rect 15531 17014 15573 17023
rect 17019 17014 17061 17023
rect 17931 17014 17973 17023
rect 18699 17014 18741 17023
rect 19074 17014 19120 17023
rect 20667 17014 20709 17023
rect 24258 17014 24304 17023
rect 26379 17014 26421 17023
rect 3610 16988 3668 16989
rect 3610 16948 3619 16988
rect 3659 16948 3668 16988
rect 9675 16981 9717 16990
rect 9867 16988 9909 16997
rect 3610 16947 3668 16948
rect 9867 16948 9868 16988
rect 9908 16948 9909 16988
rect 9867 16939 9909 16948
rect 11338 16988 11396 16989
rect 11338 16948 11347 16988
rect 11387 16948 11396 16988
rect 11338 16947 11396 16948
rect 13179 16988 13221 16997
rect 13179 16948 13180 16988
rect 13220 16948 13221 16988
rect 13179 16939 13221 16948
rect 15082 16988 15140 16989
rect 15082 16948 15091 16988
rect 15131 16948 15140 16988
rect 15082 16947 15140 16948
rect 23241 16988 23283 16997
rect 23241 16948 23242 16988
rect 23282 16948 23283 16988
rect 23241 16939 23283 16948
rect 23691 16988 23733 16997
rect 23691 16948 23692 16988
rect 23732 16948 23733 16988
rect 23691 16939 23733 16948
rect 25362 16979 25408 16988
rect 25362 16939 25363 16979
rect 25403 16939 25408 16979
rect 25362 16930 25408 16939
rect 4011 16904 4053 16913
rect 4011 16864 4012 16904
rect 4052 16864 4053 16904
rect 4011 16855 4053 16864
rect 4779 16904 4821 16913
rect 4779 16864 4780 16904
rect 4820 16864 4821 16904
rect 4779 16855 4821 16864
rect 9771 16904 9813 16913
rect 9771 16864 9772 16904
rect 9812 16864 9813 16904
rect 9771 16855 9813 16864
rect 12518 16904 12560 16913
rect 12518 16864 12519 16904
rect 12559 16864 12560 16904
rect 12518 16855 12560 16864
rect 18219 16904 18261 16913
rect 18219 16864 18220 16904
rect 18260 16864 18261 16904
rect 18219 16855 18261 16864
rect 21483 16904 21525 16913
rect 21483 16864 21484 16904
rect 21524 16864 21525 16904
rect 21483 16855 21525 16864
rect 23115 16904 23157 16913
rect 23115 16864 23116 16904
rect 23156 16864 23157 16904
rect 23115 16855 23157 16864
rect 23403 16904 23445 16913
rect 23403 16864 23404 16904
rect 23444 16864 23445 16904
rect 23403 16855 23445 16864
rect 24747 16904 24789 16913
rect 24747 16864 24748 16904
rect 24788 16864 24789 16904
rect 24747 16855 24789 16864
rect 26842 16904 26900 16905
rect 26842 16864 26851 16904
rect 26891 16864 26900 16904
rect 26842 16863 26900 16864
rect 30603 16904 30645 16913
rect 30603 16864 30604 16904
rect 30644 16864 30645 16904
rect 30603 16855 30645 16864
rect 30987 16904 31029 16913
rect 30987 16864 30988 16904
rect 31028 16864 31029 16904
rect 30987 16855 31029 16864
rect 2475 16820 2517 16829
rect 2475 16780 2476 16820
rect 2516 16780 2517 16820
rect 2475 16771 2517 16780
rect 5722 16820 5780 16821
rect 5722 16780 5731 16820
rect 5771 16780 5780 16820
rect 5722 16779 5780 16780
rect 7066 16820 7124 16821
rect 7066 16780 7075 16820
rect 7115 16780 7124 16820
rect 7066 16779 7124 16780
rect 10539 16820 10581 16829
rect 10539 16780 10540 16820
rect 10580 16780 10581 16820
rect 10539 16771 10581 16780
rect 12171 16820 12213 16829
rect 12171 16780 12172 16820
rect 12212 16780 12213 16820
rect 12171 16771 12213 16780
rect 17451 16820 17493 16829
rect 17451 16780 17452 16820
rect 17492 16780 17493 16820
rect 17451 16771 17493 16780
rect 19659 16820 19701 16829
rect 19659 16780 19660 16820
rect 19700 16780 19701 16820
rect 19659 16771 19701 16780
rect 23979 16820 24021 16829
rect 23979 16780 23980 16820
rect 24020 16780 24021 16820
rect 23979 16771 24021 16780
rect 25995 16820 26037 16829
rect 25995 16780 25996 16820
rect 26036 16780 26037 16820
rect 25995 16771 26037 16780
rect 28011 16820 28053 16829
rect 28011 16780 28012 16820
rect 28052 16780 28053 16820
rect 28011 16771 28053 16780
rect 30315 16820 30357 16829
rect 30315 16780 30316 16820
rect 30356 16780 30357 16820
rect 30315 16771 30357 16780
rect 576 16652 31392 16676
rect 576 16612 3112 16652
rect 3480 16612 10886 16652
rect 11254 16612 18660 16652
rect 19028 16612 26434 16652
rect 26802 16612 31392 16652
rect 576 16588 31392 16612
rect 1515 16484 1557 16493
rect 1515 16444 1516 16484
rect 1556 16444 1557 16484
rect 1515 16435 1557 16444
rect 3627 16484 3669 16493
rect 3627 16444 3628 16484
rect 3668 16444 3669 16484
rect 3627 16435 3669 16444
rect 8523 16484 8565 16493
rect 8523 16444 8524 16484
rect 8564 16444 8565 16484
rect 8523 16435 8565 16444
rect 8890 16484 8948 16485
rect 8890 16444 8899 16484
rect 8939 16444 8948 16484
rect 8890 16443 8948 16444
rect 17259 16484 17301 16493
rect 17259 16444 17260 16484
rect 17300 16444 17301 16484
rect 17259 16435 17301 16444
rect 24075 16484 24117 16493
rect 24075 16444 24076 16484
rect 24116 16444 24117 16484
rect 24075 16435 24117 16444
rect 25402 16484 25460 16485
rect 25402 16444 25411 16484
rect 25451 16444 25460 16484
rect 25402 16443 25460 16444
rect 27435 16484 27477 16493
rect 27435 16444 27436 16484
rect 27476 16444 27477 16484
rect 27435 16435 27477 16444
rect 30795 16484 30837 16493
rect 30795 16444 30796 16484
rect 30836 16444 30837 16484
rect 30795 16435 30837 16444
rect 5547 16400 5589 16409
rect 5547 16360 5548 16400
rect 5588 16360 5589 16400
rect 5547 16351 5589 16360
rect 9291 16400 9333 16409
rect 9291 16360 9292 16400
rect 9332 16360 9333 16400
rect 9291 16351 9333 16360
rect 15147 16400 15189 16409
rect 15147 16360 15148 16400
rect 15188 16360 15189 16400
rect 15147 16351 15189 16360
rect 15723 16400 15765 16409
rect 15723 16360 15724 16400
rect 15764 16360 15765 16400
rect 15723 16351 15765 16360
rect 16395 16400 16437 16409
rect 16395 16360 16396 16400
rect 16436 16360 16437 16400
rect 16395 16351 16437 16360
rect 22251 16400 22293 16409
rect 22251 16360 22252 16400
rect 22292 16360 22293 16400
rect 22251 16351 22293 16360
rect 25035 16400 25077 16409
rect 25035 16360 25036 16400
rect 25076 16360 25077 16400
rect 25035 16351 25077 16360
rect 30315 16400 30357 16409
rect 30315 16360 30316 16400
rect 30356 16360 30357 16400
rect 30315 16351 30357 16360
rect 6699 16316 6741 16325
rect 4050 16307 4096 16316
rect 4050 16267 4051 16307
rect 4091 16267 4096 16307
rect 6699 16276 6700 16316
rect 6740 16276 6741 16316
rect 6699 16267 6741 16276
rect 9389 16316 9431 16325
rect 9389 16276 9390 16316
rect 9430 16276 9431 16316
rect 9389 16267 9431 16276
rect 10443 16316 10485 16325
rect 10443 16276 10444 16316
rect 10484 16276 10485 16316
rect 10443 16267 10485 16276
rect 10658 16316 10700 16325
rect 10658 16276 10659 16316
rect 10699 16276 10700 16316
rect 10658 16267 10700 16276
rect 11115 16316 11157 16325
rect 11115 16276 11116 16316
rect 11156 16276 11157 16316
rect 11115 16267 11157 16276
rect 12699 16316 12741 16325
rect 12699 16276 12700 16316
rect 12740 16276 12741 16316
rect 12699 16267 12741 16276
rect 15051 16316 15093 16325
rect 15051 16276 15052 16316
rect 15092 16276 15093 16316
rect 15051 16267 15093 16276
rect 15627 16316 15669 16325
rect 15627 16276 15628 16316
rect 15668 16276 15669 16316
rect 15627 16267 15669 16276
rect 16491 16316 16533 16325
rect 16491 16276 16492 16316
rect 16532 16276 16533 16316
rect 16491 16267 16533 16276
rect 16923 16316 16965 16325
rect 16923 16276 16924 16316
rect 16964 16276 16965 16316
rect 16923 16267 16965 16276
rect 19275 16316 19317 16325
rect 19275 16276 19276 16316
rect 19316 16276 19317 16316
rect 4050 16258 4096 16267
rect 17974 16265 18016 16274
rect 19275 16267 19317 16276
rect 19947 16316 19989 16325
rect 19947 16276 19948 16316
rect 19988 16276 19989 16316
rect 19947 16267 19989 16276
rect 21867 16316 21909 16325
rect 21867 16276 21868 16316
rect 21908 16276 21909 16316
rect 21867 16267 21909 16276
rect 25755 16316 25797 16325
rect 25755 16276 25756 16316
rect 25796 16276 25797 16316
rect 25402 16274 25460 16275
rect 9691 16243 9733 16252
rect 1419 16232 1461 16241
rect 1419 16192 1420 16232
rect 1460 16192 1461 16232
rect 1834 16232 1892 16233
rect 1419 16183 1461 16192
rect 1612 16205 1670 16206
rect 1612 16165 1621 16205
rect 1661 16165 1670 16205
rect 1834 16192 1843 16232
rect 1883 16192 1892 16232
rect 1834 16191 1892 16192
rect 2187 16232 2229 16241
rect 2187 16192 2188 16232
rect 2228 16192 2229 16232
rect 2187 16183 2229 16192
rect 2746 16232 2804 16233
rect 2746 16192 2755 16232
rect 2795 16192 2804 16232
rect 2746 16191 2804 16192
rect 2859 16232 2901 16241
rect 2859 16192 2860 16232
rect 2900 16192 2901 16232
rect 2859 16183 2901 16192
rect 3435 16232 3477 16241
rect 3435 16192 3436 16232
rect 3476 16192 3477 16232
rect 3435 16183 3477 16192
rect 3915 16232 3957 16241
rect 3915 16192 3916 16232
rect 3956 16192 3957 16232
rect 3915 16183 3957 16192
rect 4144 16232 4202 16233
rect 4144 16192 4153 16232
rect 4193 16192 4202 16232
rect 4144 16191 4202 16192
rect 4491 16232 4533 16241
rect 4491 16192 4492 16232
rect 4532 16192 4533 16232
rect 4491 16183 4533 16192
rect 5355 16232 5397 16241
rect 5355 16192 5356 16232
rect 5396 16192 5397 16232
rect 5355 16183 5397 16192
rect 5722 16232 5780 16233
rect 5722 16192 5731 16232
rect 5771 16192 5780 16232
rect 5722 16191 5780 16192
rect 5866 16232 5924 16233
rect 5866 16192 5875 16232
rect 5915 16192 5924 16232
rect 5866 16191 5924 16192
rect 5972 16232 6030 16233
rect 5972 16192 5981 16232
rect 6021 16192 6030 16232
rect 5972 16191 6030 16192
rect 6100 16232 6142 16241
rect 6100 16192 6101 16232
rect 6141 16192 6142 16232
rect 6100 16183 6142 16192
rect 6240 16232 6298 16233
rect 6240 16192 6249 16232
rect 6289 16192 6298 16232
rect 6240 16191 6298 16192
rect 6795 16232 6837 16241
rect 6795 16192 6796 16232
rect 6836 16192 6837 16232
rect 6795 16183 6837 16192
rect 6914 16232 6956 16241
rect 6914 16192 6915 16232
rect 6955 16192 6956 16232
rect 6914 16183 6956 16192
rect 7024 16232 7082 16233
rect 7024 16192 7033 16232
rect 7073 16192 7082 16232
rect 7024 16191 7082 16192
rect 7195 16232 7253 16233
rect 7195 16192 7204 16232
rect 7244 16192 7253 16232
rect 7195 16191 7253 16192
rect 7354 16232 7412 16233
rect 7354 16192 7363 16232
rect 7403 16192 7412 16232
rect 7354 16191 7412 16192
rect 7480 16232 7538 16233
rect 7480 16192 7489 16232
rect 7529 16192 7538 16232
rect 7480 16191 7538 16192
rect 7637 16232 7695 16233
rect 7637 16192 7646 16232
rect 7686 16192 7695 16232
rect 7637 16191 7695 16192
rect 7738 16232 7796 16233
rect 7738 16192 7747 16232
rect 7787 16192 7796 16232
rect 7738 16191 7796 16192
rect 7978 16232 8036 16233
rect 7978 16192 7987 16232
rect 8027 16192 8036 16232
rect 7978 16191 8036 16192
rect 8122 16232 8180 16233
rect 8122 16192 8131 16232
rect 8171 16192 8180 16232
rect 8122 16191 8180 16192
rect 8247 16232 8289 16241
rect 8247 16192 8248 16232
rect 8288 16192 8289 16232
rect 8247 16183 8289 16192
rect 8378 16232 8436 16233
rect 8378 16192 8387 16232
rect 8427 16192 8436 16232
rect 8378 16191 8436 16192
rect 8506 16232 8564 16233
rect 8506 16192 8515 16232
rect 8555 16192 8564 16232
rect 8506 16191 8564 16192
rect 8715 16232 8757 16241
rect 8715 16192 8716 16232
rect 8756 16192 8757 16232
rect 8715 16183 8757 16192
rect 8890 16232 8948 16233
rect 8890 16192 8899 16232
rect 8939 16192 8948 16232
rect 8890 16191 8948 16192
rect 9051 16232 9093 16241
rect 9051 16192 9052 16232
rect 9092 16192 9093 16232
rect 9051 16183 9093 16192
rect 9216 16232 9258 16241
rect 9216 16192 9217 16232
rect 9257 16192 9258 16232
rect 9216 16183 9258 16192
rect 9508 16232 9550 16241
rect 9508 16192 9509 16232
rect 9549 16192 9550 16232
rect 9691 16203 9692 16243
rect 9732 16203 9733 16243
rect 9691 16194 9733 16203
rect 9872 16232 9914 16241
rect 9508 16183 9550 16192
rect 9872 16192 9873 16232
rect 9913 16192 9914 16232
rect 9872 16183 9914 16192
rect 9994 16232 10052 16233
rect 9994 16192 10003 16232
rect 10043 16192 10052 16232
rect 9994 16191 10052 16192
rect 10099 16232 10157 16233
rect 10099 16192 10108 16232
rect 10148 16192 10157 16232
rect 10099 16191 10157 16192
rect 10234 16232 10292 16233
rect 10234 16192 10243 16232
rect 10283 16192 10292 16232
rect 10234 16191 10292 16192
rect 10539 16232 10581 16241
rect 10539 16192 10540 16232
rect 10580 16192 10581 16232
rect 10539 16183 10581 16192
rect 10768 16232 10826 16233
rect 10768 16192 10777 16232
rect 10817 16192 10826 16232
rect 10768 16191 10826 16192
rect 11211 16232 11253 16241
rect 11211 16192 11212 16232
rect 11252 16192 11253 16232
rect 11211 16183 11253 16192
rect 11330 16232 11372 16241
rect 11330 16192 11331 16232
rect 11371 16192 11372 16232
rect 11330 16183 11372 16192
rect 11440 16232 11498 16233
rect 11440 16192 11449 16232
rect 11489 16192 11498 16232
rect 11440 16191 11498 16192
rect 11595 16232 11637 16241
rect 11595 16192 11596 16232
rect 11636 16192 11637 16232
rect 11595 16183 11637 16192
rect 11787 16232 11829 16241
rect 11787 16192 11788 16232
rect 11828 16192 11829 16232
rect 11787 16183 11829 16192
rect 12535 16232 12593 16233
rect 12535 16192 12544 16232
rect 12584 16192 12593 16232
rect 12535 16191 12593 16192
rect 13453 16232 13511 16233
rect 13453 16192 13462 16232
rect 13502 16192 13511 16232
rect 13453 16191 13511 16192
rect 13611 16232 13653 16241
rect 13611 16192 13612 16232
rect 13652 16192 13653 16232
rect 13611 16183 13653 16192
rect 13899 16232 13941 16241
rect 13899 16192 13900 16232
rect 13940 16192 13941 16232
rect 13899 16183 13941 16192
rect 14266 16232 14324 16233
rect 14266 16192 14275 16232
rect 14315 16192 14324 16232
rect 14266 16191 14324 16192
rect 14571 16232 14613 16241
rect 14571 16192 14572 16232
rect 14612 16192 14613 16232
rect 14571 16183 14613 16192
rect 14907 16232 14949 16241
rect 14907 16192 14908 16232
rect 14948 16192 14949 16232
rect 14907 16183 14949 16192
rect 15222 16232 15264 16241
rect 15222 16192 15223 16232
rect 15263 16192 15264 16232
rect 15222 16183 15264 16192
rect 15362 16232 15404 16241
rect 15362 16192 15363 16232
rect 15403 16192 15404 16232
rect 15362 16183 15404 16192
rect 15483 16232 15525 16241
rect 15483 16192 15484 16232
rect 15524 16192 15525 16232
rect 15483 16183 15525 16192
rect 15784 16232 15826 16241
rect 15784 16192 15785 16232
rect 15825 16192 15826 16232
rect 15784 16183 15826 16192
rect 15946 16232 16004 16233
rect 15946 16192 15955 16232
rect 15995 16192 16004 16232
rect 15946 16191 16004 16192
rect 16155 16232 16197 16241
rect 16155 16192 16156 16232
rect 16196 16192 16197 16232
rect 16155 16183 16197 16192
rect 16320 16232 16362 16241
rect 16320 16192 16321 16232
rect 16361 16192 16362 16232
rect 16320 16183 16362 16192
rect 16612 16232 16654 16241
rect 16612 16192 16613 16232
rect 16653 16192 16654 16232
rect 16612 16183 16654 16192
rect 16759 16232 16817 16233
rect 16759 16192 16768 16232
rect 16808 16192 16817 16232
rect 16759 16191 16817 16192
rect 17451 16232 17493 16241
rect 17451 16192 17452 16232
rect 17492 16192 17493 16232
rect 17451 16183 17493 16192
rect 17835 16232 17877 16241
rect 17835 16192 17836 16232
rect 17876 16192 17877 16232
rect 17974 16225 17975 16265
rect 18015 16225 18016 16265
rect 25035 16265 25077 16274
rect 17974 16216 18016 16225
rect 18586 16232 18644 16233
rect 17835 16183 17877 16192
rect 18586 16192 18595 16232
rect 18635 16192 18644 16232
rect 18586 16191 18644 16192
rect 19371 16232 19413 16241
rect 19371 16192 19372 16232
rect 19412 16192 19413 16232
rect 19371 16183 19413 16192
rect 19490 16232 19532 16241
rect 19490 16192 19491 16232
rect 19531 16192 19532 16232
rect 19490 16183 19532 16192
rect 19605 16232 19647 16241
rect 19605 16192 19606 16232
rect 19646 16192 19647 16232
rect 19605 16183 19647 16192
rect 20314 16232 20372 16233
rect 20314 16192 20323 16232
rect 20363 16192 20372 16232
rect 20314 16191 20372 16192
rect 22378 16232 22436 16233
rect 22378 16192 22387 16232
rect 22427 16192 22436 16232
rect 22378 16191 22436 16192
rect 22923 16232 22965 16241
rect 22923 16192 22924 16232
rect 22964 16192 22965 16232
rect 22923 16183 22965 16192
rect 23115 16232 23157 16241
rect 23115 16192 23116 16232
rect 23156 16192 23157 16232
rect 23115 16183 23157 16192
rect 23595 16232 23637 16241
rect 23595 16192 23596 16232
rect 23636 16192 23637 16232
rect 23595 16183 23637 16192
rect 23787 16232 23829 16241
rect 23787 16192 23788 16232
rect 23828 16192 23829 16232
rect 23787 16183 23829 16192
rect 24075 16232 24117 16241
rect 24075 16192 24076 16232
rect 24116 16192 24117 16232
rect 24075 16183 24117 16192
rect 24267 16232 24309 16241
rect 24267 16192 24268 16232
rect 24308 16192 24309 16232
rect 24267 16183 24309 16192
rect 24737 16232 24779 16241
rect 24737 16192 24738 16232
rect 24778 16192 24779 16232
rect 24737 16183 24779 16192
rect 24922 16232 24980 16233
rect 24922 16192 24931 16232
rect 24971 16192 24980 16232
rect 25035 16225 25036 16265
rect 25076 16225 25077 16265
rect 25035 16216 25077 16225
rect 25227 16232 25269 16241
rect 25402 16234 25411 16274
rect 25451 16234 25460 16274
rect 25755 16267 25797 16276
rect 26170 16316 26228 16317
rect 26170 16276 26179 16316
rect 26219 16276 26228 16316
rect 26170 16275 26228 16276
rect 26379 16316 26421 16325
rect 26379 16276 26380 16316
rect 26420 16276 26421 16316
rect 26379 16267 26421 16276
rect 28186 16316 28244 16317
rect 28186 16276 28195 16316
rect 28235 16276 28244 16316
rect 28186 16275 28244 16276
rect 30106 16316 30164 16317
rect 30106 16276 30115 16316
rect 30155 16276 30164 16316
rect 30106 16275 30164 16276
rect 25402 16233 25460 16234
rect 24922 16191 24980 16192
rect 25227 16192 25228 16232
rect 25268 16192 25269 16232
rect 25227 16183 25269 16192
rect 25591 16232 25649 16233
rect 25591 16192 25600 16232
rect 25640 16192 25649 16232
rect 25591 16191 25649 16192
rect 26050 16232 26108 16233
rect 26050 16192 26059 16232
rect 26099 16192 26108 16232
rect 26050 16191 26108 16192
rect 26283 16232 26325 16241
rect 26955 16232 26997 16241
rect 26283 16192 26284 16232
rect 26324 16192 26325 16232
rect 26283 16183 26325 16192
rect 26658 16223 26704 16232
rect 26658 16183 26659 16223
rect 26699 16183 26704 16223
rect 26955 16192 26956 16232
rect 26996 16192 26997 16232
rect 26955 16183 26997 16192
rect 27435 16232 27477 16241
rect 27435 16192 27436 16232
rect 27476 16192 27477 16232
rect 27435 16183 27477 16192
rect 27627 16232 27669 16241
rect 27627 16192 27628 16232
rect 27668 16192 27669 16232
rect 27627 16183 27669 16192
rect 29722 16232 29780 16233
rect 29722 16192 29731 16232
rect 29771 16192 29780 16232
rect 29722 16191 29780 16192
rect 30699 16232 30741 16241
rect 30699 16192 30700 16232
rect 30740 16192 30741 16232
rect 30699 16183 30741 16192
rect 30891 16232 30933 16241
rect 30891 16192 30892 16232
rect 30932 16192 30933 16232
rect 30891 16183 30933 16192
rect 31072 16232 31114 16241
rect 31072 16192 31073 16232
rect 31113 16192 31114 16232
rect 31072 16183 31114 16192
rect 31275 16232 31317 16241
rect 31275 16192 31276 16232
rect 31316 16192 31317 16232
rect 31275 16183 31317 16192
rect 26658 16174 26704 16183
rect 1612 16164 1670 16165
rect 3819 16148 3861 16157
rect 3819 16108 3820 16148
rect 3860 16108 3861 16148
rect 3819 16099 3861 16108
rect 4282 16148 4340 16149
rect 4282 16108 4291 16148
rect 4331 16108 4340 16148
rect 4282 16107 4340 16108
rect 13707 16148 13749 16157
rect 13707 16108 13708 16148
rect 13748 16108 13749 16148
rect 13707 16099 13749 16108
rect 22587 16148 22629 16157
rect 22587 16108 22588 16148
rect 22628 16108 22629 16148
rect 22587 16099 22629 16108
rect 26763 16148 26805 16157
rect 26763 16108 26764 16148
rect 26804 16108 26805 16148
rect 26763 16099 26805 16108
rect 2283 16064 2325 16073
rect 2283 16024 2284 16064
rect 2324 16024 2325 16064
rect 2283 16015 2325 16024
rect 3147 16064 3189 16073
rect 3147 16024 3148 16064
rect 3188 16024 3189 16064
rect 3147 16015 3189 16024
rect 3322 16064 3380 16065
rect 3322 16024 3331 16064
rect 3371 16024 3380 16064
rect 3322 16023 3380 16024
rect 4570 16064 4628 16065
rect 4570 16024 4579 16064
rect 4619 16024 4628 16064
rect 4570 16023 4628 16024
rect 5242 16064 5300 16065
rect 5242 16024 5251 16064
rect 5291 16024 5300 16064
rect 5242 16023 5300 16024
rect 6202 16064 6260 16065
rect 6202 16024 6211 16064
rect 6251 16024 6260 16064
rect 6202 16023 6260 16024
rect 7354 16064 7412 16065
rect 7354 16024 7363 16064
rect 7403 16024 7412 16064
rect 7354 16023 7412 16024
rect 9754 16064 9812 16065
rect 9754 16024 9763 16064
rect 9803 16024 9812 16064
rect 9754 16023 9812 16024
rect 11691 16064 11733 16073
rect 11691 16024 11692 16064
rect 11732 16024 11733 16064
rect 11691 16015 11733 16024
rect 13258 16064 13316 16065
rect 13258 16024 13267 16064
rect 13307 16024 13316 16064
rect 13258 16023 13316 16024
rect 14475 16064 14517 16073
rect 14475 16024 14476 16064
rect 14516 16024 14517 16064
rect 14475 16015 14517 16024
rect 17530 16064 17588 16065
rect 17530 16024 17539 16064
rect 17579 16024 17588 16064
rect 17530 16023 17588 16024
rect 18123 16064 18165 16073
rect 18123 16024 18124 16064
rect 18164 16024 18165 16064
rect 18123 16015 18165 16024
rect 18795 16064 18837 16073
rect 18795 16024 18796 16064
rect 18836 16024 18837 16064
rect 18795 16015 18837 16024
rect 23019 16064 23061 16073
rect 23019 16024 23020 16064
rect 23060 16024 23061 16064
rect 23019 16015 23061 16024
rect 23595 16064 23637 16073
rect 23595 16024 23596 16064
rect 23636 16024 23637 16064
rect 23595 16015 23637 16024
rect 27819 16064 27861 16073
rect 27819 16024 27820 16064
rect 27860 16024 27861 16064
rect 27819 16015 27861 16024
rect 31083 16064 31125 16073
rect 31083 16024 31084 16064
rect 31124 16024 31125 16064
rect 31083 16015 31125 16024
rect 576 15896 31392 15920
rect 576 15856 4352 15896
rect 4720 15856 12126 15896
rect 12494 15856 19900 15896
rect 20268 15856 27674 15896
rect 28042 15856 31392 15896
rect 576 15832 31392 15856
rect 7738 15770 7796 15771
rect 1995 15728 2037 15737
rect 1995 15688 1996 15728
rect 2036 15688 2037 15728
rect 1995 15679 2037 15688
rect 2356 15728 2414 15729
rect 2356 15688 2365 15728
rect 2405 15688 2414 15728
rect 2356 15687 2414 15688
rect 3418 15728 3476 15729
rect 3418 15688 3427 15728
rect 3467 15688 3476 15728
rect 3418 15687 3476 15688
rect 3898 15728 3956 15729
rect 3898 15688 3907 15728
rect 3947 15688 3956 15728
rect 3898 15687 3956 15688
rect 4107 15728 4149 15737
rect 7738 15730 7747 15770
rect 7787 15730 7796 15770
rect 7738 15729 7796 15730
rect 4107 15688 4108 15728
rect 4148 15688 4149 15728
rect 4107 15679 4149 15688
rect 5242 15728 5300 15729
rect 5242 15688 5251 15728
rect 5291 15688 5300 15728
rect 5242 15687 5300 15688
rect 5434 15728 5492 15729
rect 5434 15688 5443 15728
rect 5483 15688 5492 15728
rect 5434 15687 5492 15688
rect 7354 15728 7412 15729
rect 7354 15688 7363 15728
rect 7403 15688 7412 15728
rect 11770 15728 11828 15729
rect 7354 15687 7412 15688
rect 10935 15686 10977 15695
rect 11770 15688 11779 15728
rect 11819 15688 11828 15728
rect 11770 15687 11828 15688
rect 13498 15728 13556 15729
rect 13498 15688 13507 15728
rect 13547 15688 13556 15728
rect 13498 15687 13556 15688
rect 14283 15728 14325 15737
rect 14283 15688 14284 15728
rect 14324 15688 14325 15728
rect 3610 15644 3668 15645
rect 3610 15604 3619 15644
rect 3659 15604 3668 15644
rect 9675 15644 9717 15653
rect 10935 15646 10936 15686
rect 10976 15646 10977 15686
rect 14283 15679 14325 15688
rect 15915 15728 15957 15737
rect 15915 15688 15916 15728
rect 15956 15688 15957 15728
rect 15915 15679 15957 15688
rect 16762 15728 16820 15729
rect 16762 15688 16771 15728
rect 16811 15688 16820 15728
rect 16762 15687 16820 15688
rect 18987 15728 19029 15737
rect 18987 15688 18988 15728
rect 19028 15688 19029 15728
rect 18987 15679 19029 15688
rect 20523 15728 20565 15737
rect 20523 15688 20524 15728
rect 20564 15688 20565 15728
rect 20523 15679 20565 15688
rect 20890 15728 20948 15729
rect 20890 15688 20899 15728
rect 20939 15688 20948 15728
rect 20890 15687 20948 15688
rect 25227 15728 25269 15737
rect 25227 15688 25228 15728
rect 25268 15688 25269 15728
rect 25227 15679 25269 15688
rect 27051 15728 27093 15737
rect 27051 15688 27052 15728
rect 27092 15688 27093 15728
rect 27051 15679 27093 15688
rect 27418 15728 27476 15729
rect 27418 15688 27427 15728
rect 27467 15688 27476 15728
rect 27418 15687 27476 15688
rect 29818 15728 29876 15729
rect 29818 15688 29827 15728
rect 29867 15688 29876 15728
rect 29818 15687 29876 15688
rect 3610 15603 3668 15604
rect 7783 15602 7825 15611
rect 1594 15560 1652 15561
rect 1594 15520 1603 15560
rect 1643 15520 1652 15560
rect 1594 15519 1652 15520
rect 1707 15560 1749 15569
rect 1707 15520 1708 15560
rect 1748 15520 1749 15560
rect 1707 15511 1749 15520
rect 2458 15560 2516 15561
rect 3094 15560 3136 15569
rect 2458 15520 2467 15560
rect 2507 15520 2516 15560
rect 2458 15519 2516 15520
rect 2571 15551 2613 15560
rect 2571 15511 2572 15551
rect 2612 15511 2613 15551
rect 3094 15520 3095 15560
rect 3135 15520 3136 15560
rect 3094 15511 3136 15520
rect 3339 15560 3381 15569
rect 3339 15520 3340 15560
rect 3380 15520 3381 15560
rect 3339 15511 3381 15520
rect 3819 15560 3861 15569
rect 3819 15520 3820 15560
rect 3860 15520 3861 15560
rect 4322 15560 4364 15569
rect 3819 15511 3861 15520
rect 4203 15518 4245 15527
rect 2571 15502 2613 15511
rect 4203 15478 4204 15518
rect 4244 15478 4245 15518
rect 4322 15520 4323 15560
rect 4363 15520 4364 15560
rect 4322 15511 4364 15520
rect 4432 15560 4490 15561
rect 4432 15520 4441 15560
rect 4481 15520 4490 15560
rect 4432 15519 4490 15520
rect 4587 15560 4629 15569
rect 4587 15520 4588 15560
rect 4628 15520 4629 15560
rect 4587 15511 4629 15520
rect 4779 15560 4821 15569
rect 4779 15520 4780 15560
rect 4820 15520 4821 15560
rect 4779 15511 4821 15520
rect 5163 15560 5205 15569
rect 5163 15520 5164 15560
rect 5204 15520 5205 15560
rect 5163 15511 5205 15520
rect 5547 15560 5589 15569
rect 5547 15520 5548 15560
rect 5588 15520 5589 15560
rect 5547 15511 5589 15520
rect 6315 15560 6357 15569
rect 6315 15520 6316 15560
rect 6356 15520 6357 15560
rect 6315 15511 6357 15520
rect 7035 15560 7077 15569
rect 7035 15520 7036 15560
rect 7076 15520 7077 15560
rect 6922 15518 6980 15519
rect 3226 15476 3284 15477
rect 3226 15436 3235 15476
rect 3275 15436 3284 15476
rect 4203 15469 4245 15478
rect 4683 15476 4725 15485
rect 6922 15478 6931 15518
rect 6971 15478 6980 15518
rect 7035 15511 7077 15520
rect 7162 15560 7220 15561
rect 7162 15520 7171 15560
rect 7211 15520 7220 15560
rect 7162 15519 7220 15520
rect 7275 15560 7317 15569
rect 7275 15520 7276 15560
rect 7316 15520 7317 15560
rect 7783 15562 7784 15602
rect 7824 15562 7825 15602
rect 9675 15604 9676 15644
rect 9716 15604 9717 15644
rect 9675 15595 9717 15604
rect 10282 15644 10340 15645
rect 10282 15604 10291 15644
rect 10331 15604 10340 15644
rect 10935 15637 10977 15646
rect 15387 15644 15429 15653
rect 10282 15603 10340 15604
rect 11586 15635 11632 15644
rect 11586 15595 11587 15635
rect 11627 15595 11632 15635
rect 13794 15635 13840 15644
rect 11586 15586 11632 15595
rect 13199 15602 13241 15611
rect 7783 15553 7825 15562
rect 8074 15560 8132 15561
rect 7275 15511 7317 15520
rect 8074 15520 8083 15560
rect 8123 15520 8132 15560
rect 8074 15519 8132 15520
rect 8331 15560 8373 15569
rect 8331 15520 8332 15560
rect 8372 15520 8373 15560
rect 8331 15511 8373 15520
rect 8523 15560 8565 15569
rect 8523 15520 8524 15560
rect 8564 15520 8565 15560
rect 8523 15511 8565 15520
rect 9099 15560 9141 15569
rect 9099 15520 9100 15560
rect 9140 15520 9141 15560
rect 9099 15511 9141 15520
rect 9291 15560 9333 15569
rect 9291 15520 9292 15560
rect 9332 15520 9333 15560
rect 9291 15511 9333 15520
rect 9771 15560 9813 15569
rect 9771 15520 9772 15560
rect 9812 15520 9813 15560
rect 9771 15511 9813 15520
rect 10000 15560 10058 15561
rect 10000 15520 10009 15560
rect 10049 15520 10058 15560
rect 10000 15519 10058 15520
rect 10447 15560 10505 15561
rect 10447 15520 10456 15560
rect 10496 15520 10505 15560
rect 10447 15519 10505 15520
rect 10692 15560 10750 15561
rect 10692 15520 10701 15560
rect 10741 15520 10750 15560
rect 11140 15560 11182 15569
rect 10692 15519 10750 15520
rect 10855 15518 10897 15527
rect 6922 15477 6980 15478
rect 3226 15435 3284 15436
rect 4683 15436 4684 15476
rect 4724 15436 4725 15476
rect 4683 15427 4725 15436
rect 6730 15476 6788 15477
rect 6730 15436 6739 15476
rect 6779 15436 6788 15476
rect 6730 15435 6788 15436
rect 7947 15476 7989 15485
rect 10855 15478 10856 15518
rect 10896 15478 10897 15518
rect 11140 15520 11141 15560
rect 11181 15520 11182 15560
rect 11140 15511 11182 15520
rect 11290 15560 11348 15561
rect 11674 15560 11732 15561
rect 11290 15520 11299 15560
rect 11339 15520 11348 15560
rect 11290 15519 11348 15520
rect 11403 15551 11445 15560
rect 11403 15511 11404 15551
rect 11444 15511 11445 15551
rect 11674 15520 11683 15560
rect 11723 15520 11732 15560
rect 11674 15519 11732 15520
rect 11851 15560 11909 15561
rect 11851 15520 11860 15560
rect 11900 15520 11909 15560
rect 11851 15519 11909 15520
rect 12363 15560 12405 15569
rect 12363 15520 12364 15560
rect 12404 15520 12405 15560
rect 12363 15511 12405 15520
rect 12592 15560 12650 15561
rect 12592 15520 12601 15560
rect 12641 15520 12650 15560
rect 12592 15519 12650 15520
rect 12891 15560 12933 15569
rect 12891 15520 12892 15560
rect 12932 15520 12933 15560
rect 13199 15562 13200 15602
rect 13240 15562 13241 15602
rect 13794 15595 13795 15635
rect 13835 15595 13840 15635
rect 13794 15586 13840 15595
rect 14946 15635 14992 15644
rect 14946 15595 14947 15635
rect 14987 15595 14992 15635
rect 15387 15604 15388 15644
rect 15428 15604 15429 15644
rect 15387 15595 15429 15604
rect 21483 15644 21525 15653
rect 21483 15604 21484 15644
rect 21524 15604 21525 15644
rect 21483 15595 21525 15604
rect 22522 15644 22580 15645
rect 22522 15604 22531 15644
rect 22571 15604 22580 15644
rect 22522 15603 22580 15604
rect 14946 15586 14992 15595
rect 13199 15553 13241 15562
rect 13354 15560 13412 15561
rect 12891 15511 12933 15520
rect 13354 15520 13363 15560
rect 13403 15520 13412 15560
rect 13354 15519 13412 15520
rect 13498 15560 13556 15561
rect 13882 15560 13940 15561
rect 13498 15520 13507 15560
rect 13547 15520 13556 15560
rect 13498 15519 13556 15520
rect 13611 15551 13653 15560
rect 13611 15511 13612 15551
rect 13652 15511 13653 15551
rect 13882 15520 13891 15560
rect 13931 15520 13940 15560
rect 13882 15519 13940 15520
rect 14028 15560 14086 15561
rect 14028 15520 14037 15560
rect 14077 15520 14086 15560
rect 14028 15519 14086 15520
rect 14272 15560 14314 15569
rect 14272 15520 14273 15560
rect 14313 15520 14314 15560
rect 14272 15511 14314 15520
rect 14475 15560 14517 15569
rect 14475 15520 14476 15560
rect 14516 15520 14517 15560
rect 14475 15511 14517 15520
rect 14650 15560 14708 15561
rect 15034 15560 15092 15561
rect 14650 15520 14659 15560
rect 14699 15520 14708 15560
rect 14650 15519 14708 15520
rect 14763 15551 14805 15560
rect 14763 15511 14764 15551
rect 14804 15511 14805 15551
rect 15034 15520 15043 15560
rect 15083 15520 15092 15560
rect 15034 15519 15092 15520
rect 15211 15560 15269 15561
rect 15211 15520 15220 15560
rect 15260 15520 15269 15560
rect 15211 15519 15269 15520
rect 15915 15560 15957 15569
rect 15915 15520 15916 15560
rect 15956 15520 15957 15560
rect 15915 15511 15957 15520
rect 16105 15560 16147 15569
rect 16105 15520 16106 15560
rect 16146 15520 16147 15560
rect 16105 15511 16147 15520
rect 16411 15560 16469 15561
rect 16411 15520 16420 15560
rect 16460 15520 16469 15560
rect 16411 15519 16469 15520
rect 16570 15560 16628 15561
rect 16570 15520 16579 15560
rect 16619 15520 16628 15560
rect 16570 15519 16628 15520
rect 16695 15560 16737 15569
rect 16695 15520 16696 15560
rect 16736 15520 16737 15560
rect 16695 15511 16737 15520
rect 16858 15560 16916 15561
rect 16858 15520 16867 15560
rect 16907 15520 16916 15560
rect 17242 15560 17300 15561
rect 16858 15519 16916 15520
rect 16971 15549 17013 15558
rect 11403 15502 11445 15511
rect 13611 15502 13653 15511
rect 14763 15502 14805 15511
rect 16971 15509 16972 15549
rect 17012 15509 17013 15549
rect 17242 15520 17251 15560
rect 17291 15520 17300 15560
rect 17242 15519 17300 15520
rect 17355 15560 17397 15569
rect 17355 15520 17356 15560
rect 17396 15520 17397 15560
rect 17355 15511 17397 15520
rect 17739 15560 17781 15569
rect 19563 15560 19605 15569
rect 17739 15520 17740 15560
rect 17780 15520 17781 15560
rect 17739 15511 17781 15520
rect 18315 15551 18357 15560
rect 18315 15511 18316 15551
rect 18356 15511 18357 15551
rect 16971 15500 17013 15509
rect 18315 15502 18357 15511
rect 18795 15551 18837 15560
rect 18795 15511 18796 15551
rect 18836 15511 18837 15551
rect 19563 15520 19564 15560
rect 19604 15520 19605 15560
rect 19563 15511 19605 15520
rect 19664 15560 19722 15561
rect 19664 15520 19673 15560
rect 19713 15520 19722 15560
rect 19664 15519 19722 15520
rect 19947 15560 19989 15569
rect 19947 15520 19948 15560
rect 19988 15520 19989 15560
rect 19947 15511 19989 15520
rect 20235 15560 20277 15569
rect 20235 15520 20236 15560
rect 20276 15520 20277 15560
rect 20235 15511 20277 15520
rect 20369 15560 20427 15561
rect 20369 15520 20378 15560
rect 20418 15520 20427 15560
rect 20369 15519 20427 15520
rect 21003 15560 21045 15569
rect 21003 15520 21004 15560
rect 21044 15520 21045 15560
rect 21003 15511 21045 15520
rect 21387 15560 21429 15569
rect 21387 15520 21388 15560
rect 21428 15520 21429 15560
rect 21387 15511 21429 15520
rect 21562 15560 21620 15561
rect 21562 15520 21571 15560
rect 21611 15520 21620 15560
rect 21562 15519 21620 15520
rect 21946 15560 22004 15561
rect 21946 15520 21955 15560
rect 21995 15520 22004 15560
rect 21946 15519 22004 15520
rect 22059 15560 22101 15569
rect 22059 15520 22060 15560
rect 22100 15520 22101 15560
rect 22059 15511 22101 15520
rect 22906 15560 22964 15561
rect 22906 15520 22915 15560
rect 22955 15520 22964 15560
rect 22906 15519 22964 15520
rect 25483 15560 25541 15561
rect 25483 15520 25492 15560
rect 25532 15520 25541 15560
rect 25483 15519 25541 15520
rect 25594 15560 25652 15561
rect 25594 15520 25603 15560
rect 25643 15520 25652 15560
rect 25594 15519 25652 15520
rect 26043 15560 26085 15569
rect 26043 15520 26044 15560
rect 26084 15520 26085 15560
rect 25380 15518 25438 15519
rect 18795 15502 18837 15511
rect 7947 15436 7948 15476
rect 7988 15436 7989 15476
rect 7947 15427 7989 15436
rect 9906 15467 9952 15476
rect 10855 15469 10897 15478
rect 11019 15476 11061 15485
rect 9906 15427 9907 15467
rect 9947 15427 9952 15467
rect 11019 15436 11020 15476
rect 11060 15436 11061 15476
rect 11019 15427 11061 15436
rect 12267 15476 12309 15485
rect 13035 15476 13077 15485
rect 12267 15436 12268 15476
rect 12308 15436 12309 15476
rect 12267 15427 12309 15436
rect 12498 15467 12544 15476
rect 12498 15427 12499 15467
rect 12539 15427 12544 15467
rect 13035 15436 13036 15476
rect 13076 15436 13077 15476
rect 13035 15427 13077 15436
rect 15627 15476 15669 15485
rect 15627 15436 15628 15476
rect 15668 15436 15669 15476
rect 15627 15427 15669 15436
rect 17835 15476 17877 15485
rect 25380 15478 25389 15518
rect 25429 15478 25438 15518
rect 26043 15511 26085 15520
rect 26187 15560 26229 15569
rect 26187 15520 26188 15560
rect 26228 15520 26229 15560
rect 26187 15511 26229 15520
rect 26763 15560 26805 15569
rect 26763 15520 26764 15560
rect 26804 15520 26805 15560
rect 26763 15511 26805 15520
rect 26890 15560 26948 15561
rect 26890 15520 26899 15560
rect 26939 15520 26948 15560
rect 26890 15519 26948 15520
rect 27004 15560 27062 15561
rect 27004 15520 27013 15560
rect 27053 15520 27062 15560
rect 27004 15519 27062 15520
rect 27531 15560 27573 15569
rect 27531 15520 27532 15560
rect 27572 15520 27573 15560
rect 27531 15511 27573 15520
rect 27915 15560 27957 15569
rect 27915 15520 27916 15560
rect 27956 15520 27957 15560
rect 27915 15511 27957 15520
rect 28779 15560 28821 15569
rect 28779 15520 28780 15560
rect 28820 15520 28821 15560
rect 28779 15511 28821 15520
rect 28971 15560 29013 15569
rect 28971 15520 28972 15560
rect 29012 15520 29013 15560
rect 28971 15511 29013 15520
rect 30123 15560 30165 15569
rect 30123 15520 30124 15560
rect 30164 15520 30165 15560
rect 30123 15511 30165 15520
rect 30594 15551 30640 15560
rect 30594 15511 30595 15551
rect 30635 15511 30640 15551
rect 30594 15502 30640 15511
rect 25380 15477 25438 15478
rect 17835 15436 17836 15476
rect 17876 15436 17877 15476
rect 17835 15427 17877 15436
rect 30033 15476 30075 15485
rect 30033 15436 30034 15476
rect 30074 15436 30075 15476
rect 30033 15427 30075 15436
rect 30747 15476 30789 15485
rect 30747 15436 30748 15476
rect 30788 15436 30789 15476
rect 30747 15427 30789 15436
rect 9906 15418 9952 15427
rect 12498 15418 12544 15427
rect 6459 15392 6501 15401
rect 6459 15352 6460 15392
rect 6500 15352 6501 15392
rect 6459 15343 6501 15352
rect 7851 15392 7893 15401
rect 7851 15352 7852 15392
rect 7892 15352 7893 15392
rect 7851 15343 7893 15352
rect 13131 15392 13173 15401
rect 13131 15352 13132 15392
rect 13172 15352 13173 15392
rect 13131 15343 13173 15352
rect 25834 15392 25892 15393
rect 25834 15352 25843 15392
rect 25883 15352 25892 15392
rect 25834 15351 25892 15352
rect 26379 15392 26421 15401
rect 26379 15352 26380 15392
rect 26420 15352 26421 15392
rect 26379 15343 26421 15352
rect 31083 15392 31125 15401
rect 31083 15352 31084 15392
rect 31124 15352 31125 15392
rect 31083 15343 31125 15352
rect 2859 15308 2901 15317
rect 2859 15268 2860 15308
rect 2900 15268 2901 15308
rect 2859 15259 2901 15268
rect 4971 15308 5013 15317
rect 4971 15268 4972 15308
rect 5012 15268 5013 15308
rect 4971 15259 5013 15268
rect 5739 15308 5781 15317
rect 5739 15268 5740 15308
rect 5780 15268 5781 15308
rect 5739 15259 5781 15268
rect 8331 15308 8373 15317
rect 8331 15268 8332 15308
rect 8372 15268 8373 15308
rect 8331 15259 8373 15268
rect 9099 15308 9141 15317
rect 9099 15268 9100 15308
rect 9140 15268 9141 15308
rect 9099 15259 9141 15268
rect 14650 15308 14708 15309
rect 14650 15268 14659 15308
rect 14699 15268 14708 15308
rect 14650 15267 14708 15268
rect 19275 15308 19317 15317
rect 19275 15268 19276 15308
rect 19316 15268 19317 15308
rect 19275 15259 19317 15268
rect 21195 15308 21237 15317
rect 21195 15268 21196 15308
rect 21236 15268 21237 15308
rect 21195 15259 21237 15268
rect 22234 15308 22292 15309
rect 22234 15268 22243 15308
rect 22283 15268 22292 15308
rect 22234 15267 22292 15268
rect 24459 15308 24501 15317
rect 24459 15268 24460 15308
rect 24500 15268 24501 15308
rect 24459 15259 24501 15268
rect 24843 15308 24885 15317
rect 24843 15268 24844 15308
rect 24884 15268 24885 15308
rect 24843 15259 24885 15268
rect 28107 15308 28149 15317
rect 28107 15268 28108 15308
rect 28148 15268 28149 15308
rect 28107 15259 28149 15268
rect 29643 15308 29685 15317
rect 29643 15268 29644 15308
rect 29684 15268 29685 15308
rect 29643 15259 29685 15268
rect 576 15140 31392 15164
rect 576 15100 3112 15140
rect 3480 15100 10886 15140
rect 11254 15100 18660 15140
rect 19028 15100 26434 15140
rect 26802 15100 31392 15140
rect 576 15076 31392 15100
rect 1947 14972 1989 14981
rect 1947 14932 1948 14972
rect 1988 14932 1989 14972
rect 1947 14923 1989 14932
rect 4186 14972 4244 14973
rect 4186 14932 4195 14972
rect 4235 14932 4244 14972
rect 4186 14931 4244 14932
rect 10330 14972 10388 14973
rect 10330 14932 10339 14972
rect 10379 14932 10388 14972
rect 10330 14931 10388 14932
rect 12538 14972 12596 14973
rect 12538 14932 12547 14972
rect 12587 14932 12596 14972
rect 12538 14931 12596 14932
rect 13515 14972 13557 14981
rect 13515 14932 13516 14972
rect 13556 14932 13557 14972
rect 13515 14923 13557 14932
rect 16683 14972 16725 14981
rect 16683 14932 16684 14972
rect 16724 14932 16725 14972
rect 16683 14923 16725 14932
rect 19659 14972 19701 14981
rect 19659 14932 19660 14972
rect 19700 14932 19701 14972
rect 19659 14923 19701 14932
rect 23115 14972 23157 14981
rect 23115 14932 23116 14972
rect 23156 14932 23157 14972
rect 23115 14923 23157 14932
rect 24939 14972 24981 14981
rect 24939 14932 24940 14972
rect 24980 14932 24981 14972
rect 24939 14923 24981 14932
rect 25227 14972 25269 14981
rect 25227 14932 25228 14972
rect 25268 14932 25269 14972
rect 25227 14923 25269 14932
rect 27627 14972 27669 14981
rect 27627 14932 27628 14972
rect 27668 14932 27669 14972
rect 27627 14923 27669 14932
rect 30699 14972 30741 14981
rect 30699 14932 30700 14972
rect 30740 14932 30741 14972
rect 30699 14923 30741 14932
rect 8102 14888 8144 14897
rect 3979 14879 4021 14888
rect 3979 14839 3980 14879
rect 4020 14839 4021 14879
rect 8102 14848 8103 14888
rect 8143 14848 8144 14888
rect 8102 14839 8144 14848
rect 8715 14888 8757 14897
rect 15034 14888 15092 14889
rect 8715 14848 8716 14888
rect 8756 14848 8757 14888
rect 8715 14839 8757 14848
rect 11659 14879 11701 14888
rect 11659 14839 11660 14879
rect 11700 14839 11701 14879
rect 15034 14848 15043 14888
rect 15083 14848 15092 14888
rect 15034 14847 15092 14848
rect 16011 14888 16053 14897
rect 16011 14848 16012 14888
rect 16052 14848 16053 14888
rect 16011 14839 16053 14848
rect 18315 14888 18357 14897
rect 18315 14848 18316 14888
rect 18356 14848 18357 14888
rect 18315 14839 18357 14848
rect 20619 14888 20661 14897
rect 20619 14848 20620 14888
rect 20660 14848 20661 14888
rect 20619 14839 20661 14848
rect 21178 14888 21236 14889
rect 21178 14848 21187 14888
rect 21227 14848 21236 14888
rect 21178 14847 21236 14848
rect 21867 14888 21909 14897
rect 21867 14848 21868 14888
rect 21908 14848 21909 14888
rect 21867 14839 21909 14848
rect 24058 14888 24116 14889
rect 24058 14848 24067 14888
rect 24107 14848 24116 14888
rect 24058 14847 24116 14848
rect 25899 14888 25941 14897
rect 25899 14848 25900 14888
rect 25940 14848 25941 14888
rect 25899 14839 25941 14848
rect 30987 14888 31029 14897
rect 30987 14848 30988 14888
rect 31028 14848 31029 14888
rect 30987 14839 31029 14848
rect 3979 14830 4021 14839
rect 11659 14830 11701 14839
rect 14794 14832 14852 14833
rect 7083 14804 7125 14813
rect 8811 14804 8853 14813
rect 7083 14764 7084 14804
rect 7124 14764 7125 14804
rect 7083 14755 7125 14764
rect 7314 14795 7360 14804
rect 7314 14755 7315 14795
rect 7355 14755 7360 14795
rect 7314 14746 7360 14755
rect 8647 14762 8689 14771
rect 5067 14731 5109 14740
rect 1323 14720 1365 14729
rect 1323 14680 1324 14720
rect 1364 14680 1365 14720
rect 1323 14671 1365 14680
rect 1611 14720 1653 14729
rect 1611 14680 1612 14720
rect 1652 14680 1653 14720
rect 1611 14671 1653 14680
rect 2091 14720 2133 14729
rect 2091 14680 2092 14720
rect 2132 14680 2133 14720
rect 2091 14671 2133 14680
rect 2283 14720 2325 14729
rect 2283 14680 2284 14720
rect 2324 14680 2325 14720
rect 2283 14671 2325 14680
rect 3243 14720 3285 14729
rect 3243 14680 3244 14720
rect 3284 14680 3285 14720
rect 3243 14671 3285 14680
rect 3331 14720 3389 14721
rect 3331 14680 3340 14720
rect 3380 14680 3389 14720
rect 3331 14679 3389 14680
rect 3994 14720 4052 14721
rect 3994 14680 4003 14720
rect 4043 14680 4052 14720
rect 3994 14679 4052 14680
rect 4587 14720 4629 14729
rect 4587 14680 4588 14720
rect 4628 14680 4629 14720
rect 4587 14671 4629 14680
rect 4954 14720 5012 14721
rect 4954 14680 4963 14720
rect 5003 14680 5012 14720
rect 5067 14691 5068 14731
rect 5108 14691 5109 14731
rect 5931 14731 5973 14740
rect 5377 14720 5435 14721
rect 5067 14682 5109 14691
rect 5250 14711 5296 14720
rect 4954 14679 5012 14680
rect 5250 14671 5251 14711
rect 5291 14671 5296 14711
rect 5377 14680 5386 14720
rect 5426 14680 5435 14720
rect 5377 14679 5435 14680
rect 5515 14720 5573 14721
rect 5515 14680 5524 14720
rect 5564 14680 5573 14720
rect 5931 14691 5932 14731
rect 5972 14691 5973 14731
rect 6475 14731 6533 14732
rect 5931 14682 5973 14691
rect 6070 14720 6128 14721
rect 5515 14679 5573 14680
rect 6070 14680 6079 14720
rect 6119 14680 6128 14720
rect 6070 14679 6128 14680
rect 6198 14720 6256 14721
rect 6198 14680 6207 14720
rect 6247 14680 6256 14720
rect 6198 14679 6256 14680
rect 6298 14720 6356 14721
rect 6298 14680 6307 14720
rect 6347 14680 6356 14720
rect 6475 14691 6484 14731
rect 6524 14691 6533 14731
rect 6475 14690 6533 14691
rect 7179 14720 7221 14729
rect 8647 14722 8648 14762
rect 8688 14722 8689 14762
rect 8811 14764 8812 14804
rect 8852 14764 8853 14804
rect 8811 14755 8853 14764
rect 9602 14804 9644 14813
rect 9602 14764 9603 14804
rect 9643 14764 9644 14804
rect 9602 14755 9644 14764
rect 12075 14804 12117 14813
rect 12075 14764 12076 14804
rect 12116 14764 12117 14804
rect 12075 14755 12117 14764
rect 12290 14804 12332 14813
rect 12290 14764 12291 14804
rect 12331 14764 12332 14804
rect 14794 14792 14803 14832
rect 14843 14792 14852 14832
rect 14794 14791 14852 14792
rect 21082 14804 21140 14805
rect 12290 14755 12332 14764
rect 21082 14764 21091 14804
rect 21131 14764 21140 14804
rect 21082 14763 21140 14764
rect 21658 14804 21716 14805
rect 21658 14764 21667 14804
rect 21707 14764 21716 14804
rect 21658 14763 21716 14764
rect 25056 14804 25098 14813
rect 25056 14764 25057 14804
rect 25097 14764 25098 14804
rect 25056 14755 25098 14764
rect 25419 14804 25461 14813
rect 25419 14764 25420 14804
rect 25460 14764 25461 14804
rect 25174 14753 25216 14762
rect 25419 14755 25461 14764
rect 25634 14804 25676 14813
rect 25634 14764 25635 14804
rect 25675 14764 25676 14804
rect 25634 14755 25676 14764
rect 26746 14804 26804 14805
rect 26746 14764 26755 14804
rect 26795 14764 26804 14804
rect 26746 14763 26804 14764
rect 28474 14804 28532 14805
rect 28474 14764 28483 14804
rect 28523 14764 28532 14804
rect 28474 14763 28532 14764
rect 6298 14679 6356 14680
rect 7179 14680 7180 14720
rect 7220 14680 7221 14720
rect 7179 14671 7221 14680
rect 7408 14720 7466 14721
rect 7408 14680 7417 14720
rect 7457 14680 7466 14720
rect 7408 14679 7466 14680
rect 7543 14720 7601 14721
rect 7543 14680 7552 14720
rect 7592 14680 7601 14720
rect 7543 14679 7601 14680
rect 8136 14720 8194 14721
rect 8136 14680 8145 14720
rect 8185 14680 8194 14720
rect 8136 14679 8194 14680
rect 8484 14720 8542 14721
rect 8484 14680 8493 14720
rect 8533 14680 8542 14720
rect 8647 14713 8689 14722
rect 8938 14720 8996 14721
rect 8484 14679 8542 14680
rect 8938 14680 8947 14720
rect 8987 14680 8996 14720
rect 8938 14679 8996 14680
rect 9483 14720 9525 14729
rect 9483 14680 9484 14720
rect 9524 14680 9525 14720
rect 9483 14671 9525 14680
rect 9700 14720 9742 14729
rect 9700 14680 9701 14720
rect 9741 14680 9742 14720
rect 9700 14671 9742 14680
rect 9850 14720 9908 14721
rect 9850 14680 9859 14720
rect 9899 14680 9908 14720
rect 9850 14679 9908 14680
rect 10155 14720 10197 14729
rect 10155 14680 10156 14720
rect 10196 14680 10197 14720
rect 10155 14671 10197 14680
rect 10330 14720 10388 14721
rect 10330 14680 10339 14720
rect 10379 14680 10388 14720
rect 10330 14679 10388 14680
rect 10474 14720 10532 14721
rect 10474 14680 10483 14720
rect 10523 14680 10532 14720
rect 10474 14679 10532 14680
rect 10616 14720 10658 14729
rect 10616 14680 10617 14720
rect 10657 14680 10658 14720
rect 10616 14671 10658 14680
rect 10717 14720 10759 14729
rect 10717 14680 10718 14720
rect 10758 14680 10759 14720
rect 10717 14671 10759 14680
rect 10891 14720 10949 14721
rect 10891 14680 10900 14720
rect 10940 14680 10949 14720
rect 10891 14679 10949 14680
rect 11674 14720 11732 14721
rect 11674 14680 11683 14720
rect 11723 14680 11732 14720
rect 11674 14679 11732 14680
rect 11883 14720 11925 14729
rect 11883 14680 11884 14720
rect 11924 14680 11925 14720
rect 11883 14671 11925 14680
rect 12171 14720 12213 14729
rect 12831 14727 12873 14736
rect 13995 14731 14037 14740
rect 12171 14680 12172 14720
rect 12212 14680 12213 14720
rect 12171 14671 12213 14680
rect 12400 14720 12458 14721
rect 12400 14680 12409 14720
rect 12449 14680 12458 14720
rect 12400 14679 12458 14680
rect 12831 14687 12832 14727
rect 12872 14687 12873 14727
rect 12831 14678 12873 14687
rect 12923 14720 12981 14721
rect 12923 14680 12932 14720
rect 12972 14680 12981 14720
rect 12923 14679 12981 14680
rect 13323 14720 13365 14729
rect 13323 14680 13324 14720
rect 13364 14680 13365 14720
rect 13323 14671 13365 14680
rect 13882 14720 13940 14721
rect 13882 14680 13891 14720
rect 13931 14680 13940 14720
rect 13995 14691 13996 14731
rect 14036 14691 14037 14731
rect 13995 14682 14037 14691
rect 14132 14720 14190 14721
rect 13882 14679 13940 14680
rect 14132 14680 14141 14720
rect 14181 14680 14190 14720
rect 14132 14679 14190 14680
rect 14269 14720 14311 14729
rect 14269 14680 14270 14720
rect 14310 14680 14311 14720
rect 14269 14671 14311 14680
rect 14443 14720 14501 14721
rect 14443 14680 14452 14720
rect 14492 14680 14501 14720
rect 14443 14679 14501 14680
rect 14842 14720 14900 14721
rect 14842 14680 14851 14720
rect 14891 14680 14900 14720
rect 14842 14679 14900 14680
rect 15243 14720 15285 14729
rect 15243 14680 15244 14720
rect 15284 14680 15285 14720
rect 15243 14671 15285 14680
rect 15435 14720 15477 14729
rect 15435 14680 15436 14720
rect 15476 14680 15477 14720
rect 15435 14671 15477 14680
rect 16011 14720 16053 14729
rect 16011 14680 16012 14720
rect 16052 14680 16053 14720
rect 16011 14671 16053 14680
rect 16203 14720 16245 14729
rect 16203 14680 16204 14720
rect 16244 14680 16245 14720
rect 16203 14671 16245 14680
rect 16491 14720 16533 14729
rect 16491 14680 16492 14720
rect 16532 14680 16533 14720
rect 16491 14671 16533 14680
rect 16875 14720 16917 14729
rect 16875 14680 16876 14720
rect 16916 14680 16917 14720
rect 16875 14671 16917 14680
rect 17067 14720 17109 14729
rect 17067 14680 17068 14720
rect 17108 14680 17109 14720
rect 17067 14671 17109 14680
rect 18507 14720 18549 14729
rect 18507 14680 18508 14720
rect 18548 14680 18549 14720
rect 18507 14671 18549 14680
rect 18699 14720 18741 14729
rect 18699 14680 18700 14720
rect 18740 14680 18741 14720
rect 18699 14671 18741 14680
rect 18987 14720 19029 14729
rect 18987 14680 18988 14720
rect 19028 14680 19029 14720
rect 19947 14720 19989 14729
rect 18987 14671 19029 14680
rect 19258 14702 19316 14703
rect 5250 14662 5296 14671
rect 19258 14662 19267 14702
rect 19307 14662 19316 14702
rect 19947 14680 19948 14720
rect 19988 14680 19989 14720
rect 19947 14671 19989 14680
rect 20218 14720 20276 14721
rect 20218 14680 20227 14720
rect 20267 14680 20276 14720
rect 20218 14679 20276 14680
rect 21466 14720 21524 14721
rect 21466 14680 21475 14720
rect 21515 14680 21524 14720
rect 21466 14679 21524 14680
rect 21867 14720 21909 14729
rect 21867 14680 21868 14720
rect 21908 14680 21909 14720
rect 21867 14671 21909 14680
rect 22155 14720 22197 14729
rect 22155 14680 22156 14720
rect 22196 14680 22197 14720
rect 22155 14671 22197 14680
rect 22443 14720 22485 14729
rect 22443 14680 22444 14720
rect 22484 14680 22485 14720
rect 22443 14671 22485 14680
rect 23482 14720 23540 14721
rect 23482 14680 23491 14720
rect 23531 14680 23540 14720
rect 23482 14679 23540 14680
rect 23595 14720 23637 14729
rect 23595 14680 23596 14720
rect 23636 14680 23637 14720
rect 23595 14671 23637 14680
rect 24459 14720 24501 14729
rect 24459 14680 24460 14720
rect 24500 14680 24501 14720
rect 24459 14671 24501 14680
rect 24843 14720 24885 14729
rect 24843 14680 24844 14720
rect 24884 14680 24885 14720
rect 25174 14713 25175 14753
rect 25215 14713 25216 14753
rect 25174 14704 25216 14713
rect 25515 14720 25557 14729
rect 24843 14671 24885 14680
rect 25515 14680 25516 14720
rect 25556 14680 25557 14720
rect 25515 14671 25557 14680
rect 25749 14720 25791 14729
rect 25749 14680 25750 14720
rect 25790 14680 25791 14720
rect 25749 14671 25791 14680
rect 25920 14720 25962 14729
rect 25920 14680 25921 14720
rect 25961 14680 25962 14720
rect 25920 14671 25962 14680
rect 26187 14720 26229 14729
rect 26187 14680 26188 14720
rect 26228 14680 26229 14720
rect 26187 14671 26229 14680
rect 26379 14720 26421 14729
rect 26379 14680 26380 14720
rect 26420 14680 26421 14720
rect 26379 14671 26421 14680
rect 26614 14720 26656 14729
rect 26614 14680 26615 14720
rect 26655 14680 26656 14720
rect 26614 14671 26656 14680
rect 26859 14720 26901 14729
rect 26859 14680 26860 14720
rect 26900 14680 26901 14720
rect 26859 14671 26901 14680
rect 27339 14720 27381 14729
rect 27339 14680 27340 14720
rect 27380 14680 27381 14720
rect 27339 14671 27381 14680
rect 27427 14720 27485 14721
rect 27427 14680 27436 14720
rect 27476 14680 27485 14720
rect 27427 14679 27485 14680
rect 27627 14720 27669 14729
rect 27627 14680 27628 14720
rect 27668 14680 27669 14720
rect 27627 14671 27669 14680
rect 27808 14720 27866 14721
rect 27808 14680 27817 14720
rect 27857 14680 27866 14720
rect 27808 14679 27866 14680
rect 30010 14720 30068 14721
rect 30010 14680 30019 14720
rect 30059 14680 30068 14720
rect 30010 14679 30068 14680
rect 30603 14720 30645 14729
rect 30603 14680 30604 14720
rect 30644 14680 30645 14720
rect 30603 14671 30645 14680
rect 30795 14720 30837 14729
rect 30795 14680 30796 14720
rect 30836 14680 30837 14720
rect 30795 14671 30837 14680
rect 19258 14661 19316 14662
rect 3037 14636 3079 14645
rect 3037 14596 3038 14636
rect 3078 14596 3079 14636
rect 3037 14587 3079 14596
rect 9387 14636 9429 14645
rect 9387 14596 9388 14636
rect 9428 14596 9429 14636
rect 9387 14587 9429 14596
rect 10059 14636 10101 14645
rect 10059 14596 10060 14636
rect 10100 14596 10101 14636
rect 10059 14587 10101 14596
rect 19371 14636 19413 14645
rect 19371 14596 19372 14636
rect 19412 14596 19413 14636
rect 19371 14587 19413 14596
rect 20331 14636 20373 14645
rect 20331 14596 20332 14636
rect 20372 14596 20373 14636
rect 20331 14587 20373 14596
rect 23770 14636 23828 14637
rect 23770 14596 23779 14636
rect 23819 14596 23828 14636
rect 23770 14595 23828 14596
rect 26938 14636 26996 14637
rect 26938 14596 26947 14636
rect 26987 14596 26996 14636
rect 26938 14595 26996 14596
rect 27133 14636 27175 14645
rect 27133 14596 27134 14636
rect 27174 14596 27175 14636
rect 27133 14587 27175 14596
rect 28090 14636 28148 14637
rect 28090 14596 28099 14636
rect 28139 14596 28148 14636
rect 28090 14595 28148 14596
rect 30394 14636 30452 14637
rect 30394 14596 30403 14636
rect 30443 14596 30452 14636
rect 30394 14595 30452 14596
rect 2091 14552 2133 14561
rect 2091 14512 2092 14552
rect 2132 14512 2133 14552
rect 2091 14503 2133 14512
rect 3130 14552 3188 14553
rect 3130 14512 3139 14552
rect 3179 14512 3188 14552
rect 3130 14511 3188 14512
rect 4474 14552 4532 14553
rect 4474 14512 4483 14552
rect 4523 14512 4532 14552
rect 4474 14511 4532 14512
rect 4779 14552 4821 14561
rect 4779 14512 4780 14552
rect 4820 14512 4821 14552
rect 4779 14503 4821 14512
rect 5163 14552 5205 14561
rect 5163 14512 5164 14552
rect 5204 14512 5205 14552
rect 5163 14503 5205 14512
rect 6394 14552 6452 14553
rect 6394 14512 6403 14552
rect 6443 14512 6452 14552
rect 6394 14511 6452 14512
rect 7707 14552 7749 14561
rect 7707 14512 7708 14552
rect 7748 14512 7749 14552
rect 7707 14503 7749 14512
rect 8314 14552 8372 14553
rect 8314 14512 8323 14552
rect 8363 14512 8372 14552
rect 8314 14511 8372 14512
rect 13210 14552 13268 14553
rect 13210 14512 13219 14552
rect 13259 14512 13268 14552
rect 13210 14511 13268 14512
rect 14362 14552 14420 14553
rect 14362 14512 14371 14552
rect 14411 14512 14420 14552
rect 14362 14511 14420 14512
rect 15339 14552 15381 14561
rect 15339 14512 15340 14552
rect 15380 14512 15381 14552
rect 13066 14510 13124 14511
rect 13066 14470 13075 14510
rect 13115 14470 13124 14510
rect 15339 14503 15381 14512
rect 16378 14552 16436 14553
rect 16378 14512 16387 14552
rect 16427 14512 16436 14552
rect 16378 14511 16436 14512
rect 16971 14552 17013 14561
rect 16971 14512 16972 14552
rect 17012 14512 17013 14552
rect 16971 14503 17013 14512
rect 18682 14552 18740 14553
rect 18682 14512 18691 14552
rect 18731 14512 18740 14552
rect 18682 14511 18740 14512
rect 23499 14552 23541 14561
rect 23499 14512 23500 14552
rect 23540 14512 23541 14552
rect 23499 14503 23541 14512
rect 27226 14552 27284 14553
rect 27226 14512 27235 14552
rect 27275 14512 27284 14552
rect 27226 14511 27284 14512
rect 13066 14469 13124 14470
rect 576 14384 31392 14408
rect 576 14344 4352 14384
rect 4720 14344 12126 14384
rect 12494 14344 19900 14384
rect 20268 14344 27674 14384
rect 28042 14344 31392 14384
rect 576 14320 31392 14344
rect 1546 14216 1604 14217
rect 1546 14176 1555 14216
rect 1595 14176 1604 14216
rect 1546 14175 1604 14176
rect 2091 14216 2133 14225
rect 2091 14176 2092 14216
rect 2132 14176 2133 14216
rect 2091 14167 2133 14176
rect 3627 14216 3669 14225
rect 3627 14176 3628 14216
rect 3668 14176 3669 14216
rect 3627 14167 3669 14176
rect 3994 14216 4052 14217
rect 3994 14176 4003 14216
rect 4043 14176 4052 14216
rect 3994 14175 4052 14176
rect 5434 14216 5492 14217
rect 5434 14176 5443 14216
rect 5483 14176 5492 14216
rect 5434 14175 5492 14176
rect 5818 14216 5876 14217
rect 5818 14176 5827 14216
rect 5867 14176 5876 14216
rect 5818 14175 5876 14176
rect 6171 14216 6213 14225
rect 6171 14176 6172 14216
rect 6212 14176 6213 14216
rect 6171 14167 6213 14176
rect 7738 14216 7796 14217
rect 7738 14176 7747 14216
rect 7787 14176 7796 14216
rect 7738 14175 7796 14176
rect 9771 14216 9813 14225
rect 9771 14176 9772 14216
rect 9812 14176 9813 14216
rect 9771 14167 9813 14176
rect 10042 14216 10100 14217
rect 10042 14176 10051 14216
rect 10091 14176 10100 14216
rect 10042 14175 10100 14176
rect 13210 14216 13268 14217
rect 13210 14176 13219 14216
rect 13259 14176 13268 14216
rect 13210 14175 13268 14176
rect 13515 14216 13557 14225
rect 13515 14176 13516 14216
rect 13556 14176 13557 14216
rect 13515 14167 13557 14176
rect 15898 14216 15956 14217
rect 15898 14176 15907 14216
rect 15947 14176 15956 14216
rect 15898 14175 15956 14176
rect 16587 14216 16629 14225
rect 16587 14176 16588 14216
rect 16628 14176 16629 14216
rect 16587 14167 16629 14176
rect 21195 14216 21237 14225
rect 21195 14176 21196 14216
rect 21236 14176 21237 14216
rect 21195 14167 21237 14176
rect 23883 14216 23925 14225
rect 23883 14176 23884 14216
rect 23924 14176 23925 14216
rect 23883 14167 23925 14176
rect 29643 14216 29685 14225
rect 29643 14176 29644 14216
rect 29684 14176 29685 14216
rect 29643 14167 29685 14176
rect 30843 14216 30885 14225
rect 30843 14176 30844 14216
rect 30884 14176 30885 14216
rect 30843 14167 30885 14176
rect 10810 14132 10868 14133
rect 5250 14123 5296 14132
rect 5250 14083 5251 14123
rect 5291 14083 5296 14123
rect 10810 14092 10819 14132
rect 10859 14092 10868 14132
rect 10810 14091 10868 14092
rect 11115 14132 11157 14141
rect 11115 14092 11116 14132
rect 11156 14092 11157 14132
rect 11115 14083 11157 14092
rect 13899 14132 13941 14141
rect 13899 14092 13900 14132
rect 13940 14092 13941 14132
rect 11578 14090 11636 14091
rect 5250 14074 5296 14083
rect 1035 14048 1077 14057
rect 1035 14008 1036 14048
rect 1076 14008 1077 14048
rect 1035 13999 1077 14008
rect 1210 14048 1268 14049
rect 1210 14008 1219 14048
rect 1259 14008 1268 14048
rect 1210 14007 1268 14008
rect 1711 14048 1769 14049
rect 1711 14008 1720 14048
rect 1760 14008 1769 14048
rect 1711 14007 1769 14008
rect 1882 14048 1940 14049
rect 1882 14008 1891 14048
rect 1931 14008 1940 14048
rect 1882 14007 1940 14008
rect 2187 14048 2229 14057
rect 2187 14008 2188 14048
rect 2228 14008 2229 14048
rect 2187 13999 2229 14008
rect 2554 14048 2612 14049
rect 2554 14008 2563 14048
rect 2603 14008 2612 14048
rect 2554 14007 2612 14008
rect 2667 14048 2709 14057
rect 2667 14008 2668 14048
rect 2708 14008 2709 14048
rect 2667 13999 2709 14008
rect 3147 14048 3189 14057
rect 3147 14008 3148 14048
rect 3188 14008 3189 14048
rect 3147 13999 3189 14008
rect 3435 14048 3477 14057
rect 3435 14008 3436 14048
rect 3476 14008 3477 14048
rect 3435 13999 3477 14008
rect 4299 14048 4341 14057
rect 4299 14008 4300 14048
rect 4340 14008 4341 14048
rect 4299 13999 4341 14008
rect 4954 14048 5012 14049
rect 5334 14048 5392 14049
rect 4954 14008 4963 14048
rect 5003 14008 5012 14048
rect 4954 14007 5012 14008
rect 5067 14039 5109 14048
rect 5067 13999 5068 14039
rect 5108 13999 5109 14039
rect 5334 14008 5343 14048
rect 5383 14008 5392 14048
rect 5334 14007 5392 14008
rect 5515 14048 5573 14049
rect 5515 14008 5524 14048
rect 5564 14008 5573 14048
rect 5515 14007 5573 14008
rect 5728 14048 5770 14057
rect 5728 14008 5729 14048
rect 5769 14008 5770 14048
rect 5728 13999 5770 14008
rect 5931 14048 5973 14057
rect 7066 14048 7124 14049
rect 5931 14008 5932 14048
rect 5972 14008 5973 14048
rect 5931 13999 5973 14008
rect 6027 14039 6069 14048
rect 6027 13999 6028 14039
rect 6068 13999 6069 14039
rect 7066 14008 7075 14048
rect 7115 14008 7124 14048
rect 7066 14007 7124 14008
rect 7179 14048 7221 14057
rect 7179 14008 7180 14048
rect 7220 14008 7221 14048
rect 7179 13999 7221 14008
rect 7675 14048 7733 14049
rect 7675 14008 7684 14048
rect 7724 14008 7733 14048
rect 7675 14007 7733 14008
rect 7812 14048 7870 14049
rect 7812 14008 7821 14048
rect 7861 14008 7870 14048
rect 7812 14007 7870 14008
rect 7978 14048 8036 14049
rect 7978 14008 7987 14048
rect 8027 14008 8036 14048
rect 7978 14007 8036 14008
rect 8122 14048 8180 14049
rect 8122 14008 8131 14048
rect 8171 14008 8180 14048
rect 8122 14007 8180 14008
rect 8244 14048 8302 14049
rect 8244 14008 8253 14048
rect 8293 14008 8302 14048
rect 8244 14007 8302 14008
rect 8811 14048 8853 14057
rect 8811 14008 8812 14048
rect 8852 14008 8853 14048
rect 8811 13999 8853 14008
rect 8986 14048 9044 14049
rect 8986 14008 8995 14048
rect 9035 14008 9044 14048
rect 8986 14007 9044 14008
rect 9099 14048 9141 14057
rect 9099 14008 9100 14048
rect 9140 14008 9141 14048
rect 9099 13999 9141 14008
rect 9291 14048 9333 14057
rect 9291 14008 9292 14048
rect 9332 14008 9333 14048
rect 9291 13999 9333 14008
rect 9408 14048 9466 14049
rect 9408 14008 9417 14048
rect 9457 14008 9466 14048
rect 9408 14007 9466 14008
rect 9579 14048 9621 14057
rect 9579 14008 9580 14048
rect 9620 14008 9621 14048
rect 9579 13999 9621 14008
rect 9963 14048 10005 14057
rect 9963 14008 9964 14048
rect 10004 14008 10005 14048
rect 9963 13999 10005 14008
rect 10486 14048 10528 14057
rect 10486 14008 10487 14048
rect 10527 14008 10528 14048
rect 10486 13999 10528 14008
rect 10712 14048 10754 14057
rect 10712 14008 10713 14048
rect 10753 14008 10754 14048
rect 10712 13999 10754 14008
rect 11019 14048 11061 14057
rect 11019 14008 11020 14048
rect 11060 14008 11061 14048
rect 11019 13999 11061 14008
rect 11211 14048 11253 14057
rect 11578 14050 11587 14090
rect 11627 14050 11636 14090
rect 13899 14083 13941 14092
rect 14009 14132 14051 14141
rect 14009 14092 14010 14132
rect 14050 14092 14051 14132
rect 14009 14083 14051 14092
rect 15808 14132 15850 14141
rect 15808 14092 15809 14132
rect 15849 14092 15850 14132
rect 15808 14083 15850 14092
rect 21370 14132 21428 14133
rect 21370 14092 21379 14132
rect 21419 14092 21428 14132
rect 21370 14091 21428 14092
rect 29211 14132 29253 14141
rect 29211 14092 29212 14132
rect 29252 14092 29253 14132
rect 29211 14083 29253 14092
rect 12742 14067 12784 14076
rect 11578 14049 11636 14050
rect 11211 14008 11212 14048
rect 11252 14008 11253 14048
rect 11211 13999 11253 14008
rect 11712 14048 11754 14057
rect 11712 14008 11713 14048
rect 11753 14008 11754 14048
rect 11712 13999 11754 14008
rect 12004 14048 12046 14057
rect 12004 14008 12005 14048
rect 12045 14008 12046 14048
rect 12004 13999 12046 14008
rect 12363 14048 12405 14057
rect 12363 14008 12364 14048
rect 12404 14008 12405 14048
rect 12363 13999 12405 14008
rect 12555 14048 12597 14057
rect 12555 14008 12556 14048
rect 12596 14008 12597 14048
rect 12742 14027 12743 14067
rect 12783 14027 12784 14067
rect 12742 14018 12784 14027
rect 12939 14048 12981 14057
rect 12555 13999 12597 14008
rect 12939 14008 12940 14048
rect 12980 14008 12981 14048
rect 12939 13999 12981 14008
rect 13323 14048 13365 14057
rect 13323 14008 13324 14048
rect 13364 14008 13365 14048
rect 13323 13999 13365 14008
rect 13690 14048 13748 14049
rect 13690 14008 13699 14048
rect 13739 14008 13748 14048
rect 13690 14007 13748 14008
rect 13803 14048 13845 14057
rect 13803 14008 13804 14048
rect 13844 14008 13845 14048
rect 13803 13999 13845 14008
rect 14283 14048 14325 14057
rect 14283 14008 14284 14048
rect 14324 14008 14325 14048
rect 14283 13999 14325 14008
rect 14464 14048 14522 14049
rect 14464 14008 14473 14048
rect 14513 14008 14522 14048
rect 14464 14007 14522 14008
rect 14619 14048 14661 14057
rect 14619 14008 14620 14048
rect 14660 14008 14661 14048
rect 15076 14048 15118 14057
rect 14619 13999 14661 14008
rect 14763 14006 14805 14015
rect 5067 13990 5109 13999
rect 6027 13990 6069 13999
rect 4209 13964 4251 13973
rect 4209 13924 4210 13964
rect 4250 13924 4251 13964
rect 4209 13915 4251 13924
rect 6411 13964 6453 13973
rect 6411 13924 6412 13964
rect 6452 13924 6453 13964
rect 6411 13915 6453 13924
rect 10612 13964 10654 13973
rect 10612 13924 10613 13964
rect 10653 13924 10654 13964
rect 10612 13915 10654 13924
rect 11883 13964 11925 13973
rect 11883 13924 11884 13964
rect 11924 13924 11925 13964
rect 11883 13915 11925 13924
rect 12843 13964 12885 13973
rect 12843 13924 12844 13964
rect 12884 13924 12885 13964
rect 14763 13966 14764 14006
rect 14804 13966 14805 14006
rect 15076 14008 15077 14048
rect 15117 14008 15118 14048
rect 15076 13999 15118 14008
rect 15435 14048 15477 14057
rect 15435 14008 15436 14048
rect 15476 14008 15477 14048
rect 15435 13999 15477 14008
rect 15616 14048 15674 14049
rect 15616 14008 15625 14048
rect 15665 14008 15674 14048
rect 15616 14007 15674 14008
rect 16011 14048 16053 14057
rect 16011 14008 16012 14048
rect 16052 14008 16053 14048
rect 16762 14048 16820 14049
rect 17739 14048 17781 14057
rect 16011 13999 16053 14008
rect 16105 14045 16163 14046
rect 16105 14005 16114 14045
rect 16154 14005 16163 14045
rect 16762 14008 16771 14048
rect 16811 14008 16820 14048
rect 16762 14007 16820 14008
rect 17259 14039 17301 14048
rect 16105 14004 16163 14005
rect 17259 13999 17260 14039
rect 17300 13999 17301 14039
rect 17739 14008 17740 14048
rect 17780 14008 17781 14048
rect 17739 13999 17781 14008
rect 18219 14048 18261 14057
rect 18219 14008 18220 14048
rect 18260 14008 18261 14048
rect 18219 13999 18261 14008
rect 18329 14048 18387 14049
rect 18329 14008 18338 14048
rect 18378 14008 18387 14048
rect 18329 14007 18387 14008
rect 18682 14048 18740 14049
rect 18682 14008 18691 14048
rect 18731 14008 18740 14048
rect 18682 14007 18740 14008
rect 19851 14048 19893 14057
rect 19851 14008 19852 14048
rect 19892 14008 19893 14048
rect 19851 13999 19893 14008
rect 19952 14048 20010 14049
rect 19952 14008 19961 14048
rect 20001 14008 20010 14048
rect 19952 14007 20010 14008
rect 20235 14048 20277 14057
rect 20235 14008 20236 14048
rect 20276 14008 20277 14048
rect 20235 13999 20277 14008
rect 20523 14048 20565 14057
rect 20523 14008 20524 14048
rect 20564 14008 20565 14048
rect 20523 13999 20565 14008
rect 21562 14048 21620 14049
rect 22539 14048 22581 14057
rect 21562 14008 21571 14048
rect 21611 14008 21620 14048
rect 21562 14007 21620 14008
rect 22059 14039 22101 14048
rect 22059 13999 22060 14039
rect 22100 13999 22101 14039
rect 22539 14008 22540 14048
rect 22580 14008 22581 14048
rect 22539 13999 22581 14008
rect 23019 14048 23061 14057
rect 23019 14008 23020 14048
rect 23060 14008 23061 14048
rect 23403 14048 23445 14057
rect 23019 13999 23061 14008
rect 23132 14029 23174 14038
rect 17259 13990 17301 13999
rect 22059 13990 22101 13999
rect 23132 13989 23133 14029
rect 23173 13989 23174 14029
rect 23403 14008 23404 14048
rect 23444 14008 23445 14048
rect 23403 13999 23445 14008
rect 23787 14048 23829 14057
rect 23787 14008 23788 14048
rect 23828 14008 23829 14048
rect 23787 13999 23829 14008
rect 26170 14048 26228 14049
rect 26170 14008 26179 14048
rect 26219 14008 26228 14048
rect 26170 14007 26228 14008
rect 27034 14048 27092 14049
rect 27034 14008 27043 14048
rect 27083 14008 27092 14048
rect 27034 14007 27092 14008
rect 27147 14048 27189 14057
rect 27147 14008 27148 14048
rect 27188 14008 27189 14048
rect 27147 13999 27189 14008
rect 27610 14048 27668 14049
rect 27610 14008 27619 14048
rect 27659 14008 27668 14048
rect 27610 14007 27668 14008
rect 27915 14048 27957 14057
rect 27915 14008 27916 14048
rect 27956 14008 27957 14048
rect 27915 13999 27957 14008
rect 28186 14048 28244 14049
rect 28186 14008 28195 14048
rect 28235 14008 28244 14048
rect 28186 14007 28244 14008
rect 28875 14048 28917 14057
rect 28875 14008 28876 14048
rect 28916 14008 28917 14048
rect 28875 13999 28917 14008
rect 29023 14048 29081 14049
rect 29023 14008 29032 14048
rect 29072 14008 29081 14048
rect 29023 14007 29081 14008
rect 29547 14048 29589 14057
rect 29547 14008 29548 14048
rect 29588 14008 29589 14048
rect 29547 13999 29589 14008
rect 29738 14048 29780 14057
rect 29738 14008 29739 14048
rect 29779 14008 29780 14048
rect 30112 14048 30170 14049
rect 29738 13999 29780 14008
rect 29931 14006 29973 14015
rect 30112 14008 30121 14048
rect 30161 14008 30170 14048
rect 30112 14007 30170 14008
rect 23132 13980 23174 13989
rect 14763 13957 14805 13966
rect 14955 13964 14997 13973
rect 12843 13915 12885 13924
rect 14955 13924 14956 13964
rect 14996 13924 14997 13964
rect 14955 13915 14997 13924
rect 17835 13964 17877 13973
rect 17835 13924 17836 13964
rect 17876 13924 17877 13964
rect 17835 13915 17877 13924
rect 22635 13964 22677 13973
rect 29931 13966 29932 14006
rect 29972 13966 29973 14006
rect 22635 13924 22636 13964
rect 22676 13924 22677 13964
rect 22635 13915 22677 13924
rect 24634 13964 24692 13965
rect 24634 13924 24643 13964
rect 24683 13924 24692 13964
rect 24634 13923 24692 13924
rect 26554 13964 26612 13965
rect 26554 13924 26563 13964
rect 26603 13924 26612 13964
rect 29931 13957 29973 13966
rect 31083 13964 31125 13973
rect 26554 13923 26612 13924
rect 31083 13924 31084 13964
rect 31124 13924 31125 13964
rect 31083 13915 31125 13924
rect 2842 13880 2900 13881
rect 2842 13840 2851 13880
rect 2891 13840 2900 13880
rect 2842 13839 2900 13840
rect 8907 13880 8949 13889
rect 8907 13840 8908 13880
rect 8948 13840 8949 13880
rect 8907 13831 8949 13840
rect 9291 13880 9333 13889
rect 9291 13840 9292 13880
rect 9332 13840 9333 13880
rect 9291 13831 9333 13840
rect 11787 13880 11829 13889
rect 11787 13840 11788 13880
rect 11828 13840 11829 13880
rect 11787 13831 11829 13840
rect 12363 13880 12405 13889
rect 12363 13840 12364 13880
rect 12404 13840 12405 13880
rect 12363 13831 12405 13840
rect 14859 13880 14901 13889
rect 14859 13840 14860 13880
rect 14900 13840 14901 13880
rect 14859 13831 14901 13840
rect 27915 13880 27957 13889
rect 27915 13840 27916 13880
rect 27956 13840 27957 13880
rect 27915 13831 27957 13840
rect 30315 13880 30357 13889
rect 30315 13840 30316 13880
rect 30356 13840 30357 13880
rect 30315 13831 30357 13840
rect 1210 13796 1268 13797
rect 1210 13756 1219 13796
rect 1259 13756 1268 13796
rect 1210 13755 1268 13756
rect 7354 13796 7412 13797
rect 7354 13756 7363 13796
rect 7403 13756 7412 13796
rect 7354 13755 7412 13756
rect 14283 13796 14325 13805
rect 14283 13756 14284 13796
rect 14324 13756 14325 13796
rect 14283 13747 14325 13756
rect 15435 13796 15477 13805
rect 15435 13756 15436 13796
rect 15476 13756 15477 13796
rect 15435 13747 15477 13756
rect 19083 13796 19125 13805
rect 19083 13756 19084 13796
rect 19124 13756 19125 13796
rect 19083 13747 19125 13756
rect 19563 13796 19605 13805
rect 19563 13756 19564 13796
rect 19604 13756 19605 13796
rect 19563 13747 19605 13756
rect 24267 13796 24309 13805
rect 24267 13756 24268 13796
rect 24308 13756 24309 13796
rect 24267 13747 24309 13756
rect 27322 13796 27380 13797
rect 27322 13756 27331 13796
rect 27371 13756 27380 13796
rect 27322 13755 27380 13756
rect 29931 13796 29973 13805
rect 29931 13756 29932 13796
rect 29972 13756 29973 13796
rect 29931 13747 29973 13756
rect 576 13628 31392 13652
rect 576 13588 3112 13628
rect 3480 13588 10886 13628
rect 11254 13588 18660 13628
rect 19028 13588 26434 13628
rect 26802 13588 31392 13628
rect 576 13564 31392 13588
rect 8122 13460 8180 13461
rect 8122 13420 8131 13460
rect 8171 13420 8180 13460
rect 8122 13419 8180 13420
rect 9562 13460 9620 13461
rect 9562 13420 9571 13460
rect 9611 13420 9620 13460
rect 9562 13419 9620 13420
rect 10330 13460 10388 13461
rect 10330 13420 10339 13460
rect 10379 13420 10388 13460
rect 10330 13419 10388 13420
rect 12747 13460 12789 13469
rect 12747 13420 12748 13460
rect 12788 13420 12789 13460
rect 12747 13411 12789 13420
rect 14266 13460 14324 13461
rect 14266 13420 14275 13460
rect 14315 13420 14324 13460
rect 14266 13419 14324 13420
rect 15243 13460 15285 13469
rect 15243 13420 15244 13460
rect 15284 13420 15285 13460
rect 15243 13411 15285 13420
rect 19851 13460 19893 13469
rect 19851 13420 19852 13460
rect 19892 13420 19893 13460
rect 19851 13411 19893 13420
rect 21099 13460 21141 13469
rect 21099 13420 21100 13460
rect 21140 13420 21141 13460
rect 21099 13411 21141 13420
rect 23482 13460 23540 13461
rect 23482 13420 23491 13460
rect 23531 13420 23540 13460
rect 23482 13419 23540 13420
rect 24459 13460 24501 13469
rect 24459 13420 24460 13460
rect 24500 13420 24501 13460
rect 24459 13411 24501 13420
rect 25803 13460 25845 13469
rect 25803 13420 25804 13460
rect 25844 13420 25845 13460
rect 25803 13411 25845 13420
rect 27819 13460 27861 13469
rect 27819 13420 27820 13460
rect 27860 13420 27861 13460
rect 27819 13411 27861 13420
rect 11866 13376 11924 13377
rect 11866 13336 11875 13376
rect 11915 13336 11924 13376
rect 11866 13335 11924 13336
rect 21483 13376 21525 13385
rect 21483 13336 21484 13376
rect 21524 13336 21525 13376
rect 21483 13327 21525 13336
rect 24075 13376 24117 13385
rect 24075 13336 24076 13376
rect 24116 13336 24117 13376
rect 24075 13327 24117 13336
rect 30795 13376 30837 13385
rect 30795 13336 30796 13376
rect 30836 13336 30837 13376
rect 30795 13327 30837 13336
rect 2074 13292 2132 13293
rect 2074 13252 2083 13292
rect 2123 13252 2132 13292
rect 2074 13251 2132 13252
rect 2283 13292 2325 13301
rect 2283 13252 2284 13292
rect 2324 13252 2325 13292
rect 2283 13243 2325 13252
rect 5739 13292 5781 13301
rect 6778 13292 6836 13293
rect 5739 13252 5740 13292
rect 5780 13252 5781 13292
rect 5739 13243 5781 13252
rect 5970 13283 6016 13292
rect 5970 13243 5971 13283
rect 6011 13243 6016 13283
rect 6778 13252 6787 13292
rect 6827 13252 6836 13292
rect 6778 13251 6836 13252
rect 6987 13292 7029 13301
rect 6987 13252 6988 13292
rect 7028 13252 7029 13292
rect 6987 13243 7029 13252
rect 8890 13292 8948 13293
rect 8890 13252 8899 13292
rect 8939 13252 8948 13292
rect 8890 13251 8948 13252
rect 9099 13292 9141 13301
rect 13707 13292 13749 13301
rect 9099 13252 9100 13292
rect 9140 13252 9141 13292
rect 5970 13234 6016 13243
rect 8415 13241 8457 13250
rect 9099 13243 9141 13252
rect 11538 13283 11584 13292
rect 5242 13219 5300 13220
rect 1549 13208 1607 13209
rect 1549 13168 1558 13208
rect 1598 13168 1607 13208
rect 1549 13167 1607 13168
rect 1942 13208 1984 13217
rect 1942 13168 1943 13208
rect 1983 13168 1984 13208
rect 1942 13159 1984 13168
rect 2187 13208 2229 13217
rect 2187 13168 2188 13208
rect 2228 13168 2229 13208
rect 2187 13159 2229 13168
rect 3034 13208 3092 13209
rect 3034 13168 3043 13208
rect 3083 13168 3092 13208
rect 3034 13167 3092 13168
rect 3147 13208 3189 13217
rect 3147 13168 3148 13208
rect 3188 13168 3189 13208
rect 3147 13159 3189 13168
rect 4299 13208 4341 13217
rect 4299 13168 4300 13208
rect 4340 13168 4341 13208
rect 4299 13159 4341 13168
rect 4426 13208 4484 13209
rect 4426 13168 4435 13208
rect 4475 13168 4484 13208
rect 4426 13167 4484 13168
rect 4795 13208 4853 13209
rect 4795 13168 4804 13208
rect 4844 13168 4853 13208
rect 4795 13167 4853 13168
rect 4976 13208 5018 13217
rect 4976 13168 4977 13208
rect 5017 13168 5018 13208
rect 4976 13159 5018 13168
rect 5080 13208 5138 13209
rect 5080 13168 5089 13208
rect 5129 13168 5138 13208
rect 5242 13179 5251 13219
rect 5291 13179 5300 13219
rect 5242 13178 5300 13179
rect 5364 13208 5422 13209
rect 5080 13167 5138 13168
rect 5364 13168 5373 13208
rect 5413 13168 5422 13208
rect 5364 13167 5422 13168
rect 5835 13208 5877 13217
rect 5835 13168 5836 13208
rect 5876 13168 5877 13208
rect 5835 13159 5877 13168
rect 6075 13208 6117 13217
rect 6075 13168 6076 13208
rect 6116 13168 6117 13208
rect 6075 13159 6117 13168
rect 6214 13208 6256 13217
rect 6214 13168 6215 13208
rect 6255 13168 6256 13208
rect 6214 13159 6256 13168
rect 6394 13208 6452 13209
rect 6394 13168 6403 13208
rect 6443 13168 6452 13208
rect 6394 13167 6452 13168
rect 6646 13208 6688 13217
rect 6646 13168 6647 13208
rect 6687 13168 6688 13208
rect 6646 13159 6688 13168
rect 6891 13208 6933 13217
rect 6891 13168 6892 13208
rect 6932 13168 6933 13208
rect 6891 13159 6933 13168
rect 7459 13208 7517 13209
rect 7459 13168 7468 13208
rect 7508 13168 7517 13208
rect 7459 13167 7517 13168
rect 7642 13208 7700 13209
rect 7642 13168 7651 13208
rect 7691 13168 7700 13208
rect 7642 13167 7700 13168
rect 7755 13208 7797 13217
rect 7755 13168 7756 13208
rect 7796 13168 7797 13208
rect 8415 13201 8416 13241
rect 8456 13201 8457 13241
rect 10623 13241 10665 13250
rect 8415 13192 8457 13201
rect 8506 13208 8564 13209
rect 7755 13159 7797 13168
rect 8506 13168 8515 13208
rect 8555 13168 8564 13208
rect 8506 13167 8564 13168
rect 8758 13208 8800 13217
rect 8758 13168 8759 13208
rect 8799 13168 8800 13208
rect 8758 13159 8800 13168
rect 9003 13208 9045 13217
rect 9003 13168 9004 13208
rect 9044 13168 9045 13208
rect 9003 13159 9045 13168
rect 9859 13208 9917 13209
rect 9859 13168 9868 13208
rect 9908 13168 9917 13208
rect 10623 13201 10624 13241
rect 10664 13201 10665 13241
rect 11538 13243 11539 13283
rect 11579 13243 11584 13283
rect 13707 13252 13708 13292
rect 13748 13252 13749 13292
rect 13707 13243 13749 13252
rect 14763 13292 14805 13301
rect 14763 13252 14764 13292
rect 14804 13252 14805 13292
rect 14763 13243 14805 13252
rect 16034 13292 16076 13301
rect 16034 13252 16035 13292
rect 16075 13252 16076 13292
rect 16378 13292 16436 13293
rect 16034 13243 16076 13252
rect 16155 13250 16197 13259
rect 16378 13252 16387 13292
rect 16427 13252 16436 13292
rect 16378 13251 16436 13252
rect 17931 13292 17973 13301
rect 17931 13252 17932 13292
rect 17972 13252 17973 13292
rect 11538 13234 11584 13243
rect 10623 13192 10665 13201
rect 10714 13208 10772 13209
rect 9859 13167 9917 13168
rect 10714 13168 10723 13208
rect 10763 13168 10772 13208
rect 10714 13167 10772 13168
rect 11403 13208 11445 13217
rect 11403 13168 11404 13208
rect 11444 13168 11445 13208
rect 11403 13159 11445 13168
rect 11632 13208 11690 13209
rect 11632 13168 11641 13208
rect 11681 13168 11690 13208
rect 11632 13167 11690 13168
rect 12267 13208 12309 13217
rect 12267 13168 12268 13208
rect 12308 13168 12309 13208
rect 12267 13159 12309 13168
rect 12922 13208 12980 13209
rect 12922 13168 12931 13208
rect 12971 13168 12980 13208
rect 12922 13167 12980 13168
rect 13227 13208 13269 13217
rect 13227 13168 13228 13208
rect 13268 13168 13269 13208
rect 13227 13159 13269 13168
rect 13786 13208 13844 13209
rect 13786 13168 13795 13208
rect 13835 13168 13844 13208
rect 13786 13167 13844 13168
rect 14269 13208 14311 13217
rect 14269 13168 14270 13208
rect 14310 13168 14311 13208
rect 14269 13159 14311 13168
rect 14563 13208 14621 13209
rect 14563 13168 14572 13208
rect 14612 13168 14621 13208
rect 14563 13167 14621 13168
rect 14859 13208 14901 13217
rect 14859 13168 14860 13208
rect 14900 13168 14901 13208
rect 14859 13159 14901 13168
rect 14978 13208 15020 13217
rect 14978 13168 14979 13208
rect 15019 13168 15020 13208
rect 14978 13159 15020 13168
rect 15088 13208 15146 13209
rect 15088 13168 15097 13208
rect 15137 13168 15146 13208
rect 15088 13167 15146 13168
rect 15243 13208 15285 13217
rect 15243 13168 15244 13208
rect 15284 13168 15285 13208
rect 15243 13159 15285 13168
rect 15360 13208 15418 13209
rect 15360 13168 15369 13208
rect 15409 13168 15418 13208
rect 15360 13167 15418 13168
rect 15531 13208 15573 13217
rect 15531 13168 15532 13208
rect 15572 13168 15573 13208
rect 15531 13159 15573 13168
rect 15915 13208 15957 13217
rect 15915 13168 15916 13208
rect 15956 13168 15957 13208
rect 16155 13210 16156 13250
rect 16196 13210 16197 13250
rect 17931 13243 17973 13252
rect 26410 13292 26468 13293
rect 26410 13252 26419 13292
rect 26459 13252 26468 13292
rect 26410 13251 26468 13252
rect 26907 13292 26949 13301
rect 26907 13252 26908 13292
rect 26948 13252 26949 13292
rect 26907 13243 26949 13252
rect 29722 13292 29780 13293
rect 29722 13252 29731 13292
rect 29771 13252 29780 13292
rect 29722 13251 29780 13252
rect 16155 13201 16197 13210
rect 16258 13208 16316 13209
rect 15915 13159 15957 13168
rect 16258 13168 16267 13208
rect 16307 13168 16316 13208
rect 16258 13167 16316 13168
rect 16491 13208 16533 13217
rect 16491 13168 16492 13208
rect 16532 13168 16533 13208
rect 16491 13159 16533 13168
rect 16954 13208 17012 13209
rect 16954 13168 16963 13208
rect 17003 13168 17012 13208
rect 16954 13167 17012 13168
rect 17443 13208 17501 13209
rect 17443 13168 17452 13208
rect 17492 13168 17501 13208
rect 17443 13167 17501 13168
rect 18027 13208 18069 13217
rect 18027 13168 18028 13208
rect 18068 13168 18069 13208
rect 18027 13159 18069 13168
rect 18411 13208 18453 13217
rect 18411 13168 18412 13208
rect 18452 13168 18453 13208
rect 18411 13159 18453 13168
rect 18512 13208 18554 13217
rect 18512 13168 18513 13208
rect 18553 13168 18554 13208
rect 18512 13159 18554 13168
rect 19179 13208 19221 13217
rect 19179 13168 19180 13208
rect 19220 13168 19221 13208
rect 19179 13159 19221 13168
rect 19450 13208 19508 13209
rect 19450 13168 19459 13208
rect 19499 13168 19508 13208
rect 19450 13167 19508 13168
rect 20427 13208 20469 13217
rect 20811 13208 20853 13217
rect 20427 13168 20428 13208
rect 20468 13168 20469 13208
rect 20427 13159 20469 13168
rect 20523 13199 20565 13208
rect 20523 13159 20524 13199
rect 20564 13159 20565 13199
rect 20811 13168 20812 13208
rect 20852 13168 20853 13208
rect 20811 13159 20853 13168
rect 21099 13208 21141 13217
rect 21099 13168 21100 13208
rect 21140 13168 21141 13208
rect 21099 13159 21141 13168
rect 21291 13208 21333 13217
rect 21291 13168 21292 13208
rect 21332 13168 21333 13208
rect 21291 13159 21333 13168
rect 21771 13208 21813 13217
rect 22155 13208 22197 13217
rect 21771 13168 21772 13208
rect 21812 13168 21813 13208
rect 21771 13159 21813 13168
rect 21867 13199 21909 13208
rect 21867 13159 21868 13199
rect 21908 13159 21909 13199
rect 22155 13168 22156 13208
rect 22196 13168 22197 13208
rect 22155 13159 22197 13168
rect 22443 13208 22485 13217
rect 22443 13168 22444 13208
rect 22484 13168 22485 13208
rect 22443 13159 22485 13168
rect 23451 13208 23493 13217
rect 23451 13168 23452 13208
rect 23492 13168 23493 13208
rect 23451 13159 23493 13168
rect 23595 13208 23637 13217
rect 23595 13168 23596 13208
rect 23636 13168 23637 13208
rect 23595 13159 23637 13168
rect 25131 13208 25173 13217
rect 25131 13168 25132 13208
rect 25172 13168 25173 13208
rect 25131 13159 25173 13168
rect 25306 13208 25364 13209
rect 25306 13168 25315 13208
rect 25355 13168 25364 13208
rect 25306 13167 25364 13168
rect 25803 13208 25845 13217
rect 25803 13168 25804 13208
rect 25844 13168 25845 13208
rect 25803 13159 25845 13168
rect 25920 13208 25978 13209
rect 25920 13168 25929 13208
rect 25969 13168 25978 13208
rect 25920 13167 25978 13168
rect 26091 13208 26133 13217
rect 26091 13168 26092 13208
rect 26132 13168 26133 13208
rect 26091 13159 26133 13168
rect 26575 13208 26633 13209
rect 26575 13168 26584 13208
rect 26624 13168 26633 13208
rect 26575 13167 26633 13168
rect 26743 13208 26801 13209
rect 26743 13168 26752 13208
rect 26792 13168 26801 13208
rect 26743 13167 26801 13168
rect 29338 13208 29396 13209
rect 29338 13168 29347 13208
rect 29387 13168 29396 13208
rect 29338 13167 29396 13168
rect 29866 13208 29924 13209
rect 29866 13168 29875 13208
rect 29915 13168 29924 13208
rect 29866 13167 29924 13168
rect 30411 13208 30453 13217
rect 30411 13168 30412 13208
rect 30452 13168 30453 13208
rect 30411 13159 30453 13168
rect 30603 13208 30645 13217
rect 30603 13168 30604 13208
rect 30644 13168 30645 13208
rect 30603 13159 30645 13168
rect 31179 13208 31221 13217
rect 31179 13168 31180 13208
rect 31220 13168 31221 13208
rect 31179 13159 31221 13168
rect 20523 13150 20565 13159
rect 21867 13150 21909 13159
rect 7165 13124 7207 13133
rect 7165 13084 7166 13124
rect 7206 13084 7207 13124
rect 7165 13075 7207 13084
rect 7258 13124 7316 13125
rect 7258 13084 7267 13124
rect 7307 13084 7316 13124
rect 7258 13083 7316 13084
rect 7961 13124 8003 13133
rect 7961 13084 7962 13124
rect 8002 13084 8003 13124
rect 7961 13075 8003 13084
rect 9565 13124 9607 13133
rect 9565 13084 9566 13124
rect 9606 13084 9607 13124
rect 9565 13075 9607 13084
rect 11307 13124 11349 13133
rect 11307 13084 11308 13124
rect 11348 13084 11349 13124
rect 11307 13075 11349 13084
rect 11962 13124 12020 13125
rect 11962 13084 11971 13124
rect 12011 13084 12020 13124
rect 11962 13083 12020 13084
rect 12747 13124 12789 13133
rect 12747 13084 12748 13124
rect 12788 13084 12789 13124
rect 12747 13075 12789 13084
rect 14475 13124 14517 13133
rect 14475 13084 14476 13124
rect 14516 13084 14517 13124
rect 14475 13075 14517 13084
rect 15819 13124 15861 13133
rect 15819 13084 15820 13124
rect 15860 13084 15861 13124
rect 15819 13075 15861 13084
rect 16570 13124 16628 13125
rect 16570 13084 16579 13124
rect 16619 13084 16628 13124
rect 16570 13083 16628 13084
rect 19563 13124 19605 13133
rect 19563 13084 19564 13124
rect 19604 13084 19605 13124
rect 19563 13075 19605 13084
rect 25622 13124 25664 13133
rect 25622 13084 25623 13124
rect 25663 13084 25664 13124
rect 25622 13075 25664 13084
rect 27418 13124 27476 13125
rect 27418 13084 27427 13124
rect 27467 13084 27476 13124
rect 27418 13083 27476 13084
rect 1354 13040 1412 13041
rect 1354 13000 1363 13040
rect 1403 13000 1412 13040
rect 1354 12999 1412 13000
rect 3435 13040 3477 13049
rect 3435 13000 3436 13040
rect 3476 13000 3477 13040
rect 3435 12991 3477 13000
rect 4587 13040 4629 13049
rect 4587 13000 4588 13040
rect 4628 13000 4629 13040
rect 4587 12991 4629 13000
rect 4858 13040 4916 13041
rect 4858 13000 4867 13040
rect 4907 13000 4916 13040
rect 4858 12999 4916 13000
rect 6315 13040 6357 13049
rect 6315 13000 6316 13040
rect 6356 13000 6357 13040
rect 6315 12991 6357 13000
rect 7371 13040 7413 13049
rect 7371 13000 7372 13040
rect 7412 13000 7413 13040
rect 7371 12991 7413 13000
rect 7851 13040 7893 13049
rect 7851 13000 7852 13040
rect 7892 13000 7893 13040
rect 7851 12991 7893 13000
rect 8649 13040 8707 13041
rect 8649 13000 8658 13040
rect 8698 13000 8707 13040
rect 8649 12999 8707 13000
rect 9771 13040 9813 13049
rect 9771 13000 9772 13040
rect 9812 13000 9813 13040
rect 9771 12991 9813 13000
rect 10834 13040 10892 13041
rect 10834 13000 10843 13040
rect 10883 13000 10892 13040
rect 10834 12999 10892 13000
rect 13402 13040 13460 13041
rect 13402 13000 13411 13040
rect 13451 13000 13460 13040
rect 13402 12999 13460 13000
rect 13611 13040 13653 13049
rect 13611 13000 13612 13040
rect 13652 13000 13653 13040
rect 13611 12991 13653 13000
rect 16779 13040 16821 13049
rect 16779 13000 16780 13040
rect 16820 13000 16821 13040
rect 16779 12991 16821 13000
rect 20091 13040 20133 13049
rect 20091 13000 20092 13040
rect 20132 13000 20133 13040
rect 20091 12991 20133 13000
rect 23115 13040 23157 13049
rect 23115 13000 23116 13040
rect 23156 13000 23157 13040
rect 23115 12991 23157 13000
rect 25402 13040 25460 13041
rect 25402 13000 25411 13040
rect 25451 13000 25460 13040
rect 25402 12999 25460 13000
rect 25515 13040 25557 13049
rect 25515 13000 25516 13040
rect 25556 13000 25557 13040
rect 25515 12991 25557 13000
rect 30075 13040 30117 13049
rect 30075 13000 30076 13040
rect 30116 13000 30117 13040
rect 30075 12991 30117 13000
rect 30586 13040 30644 13041
rect 30586 13000 30595 13040
rect 30635 13000 30644 13040
rect 30586 12999 30644 13000
rect 576 12872 31392 12896
rect 576 12832 4352 12872
rect 4720 12832 12126 12872
rect 12494 12832 19900 12872
rect 20268 12832 27674 12872
rect 28042 12832 31392 12872
rect 576 12808 31392 12832
rect 1227 12704 1269 12713
rect 1227 12664 1228 12704
rect 1268 12664 1269 12704
rect 1227 12655 1269 12664
rect 1995 12704 2037 12713
rect 1995 12664 1996 12704
rect 2036 12664 2037 12704
rect 1995 12655 2037 12664
rect 2379 12704 2421 12713
rect 2379 12664 2380 12704
rect 2420 12664 2421 12704
rect 2379 12655 2421 12664
rect 4282 12704 4340 12705
rect 4282 12664 4291 12704
rect 4331 12664 4340 12704
rect 4282 12663 4340 12664
rect 4570 12704 4628 12705
rect 4570 12664 4579 12704
rect 4619 12664 4628 12704
rect 4570 12663 4628 12664
rect 5931 12704 5973 12713
rect 5931 12664 5932 12704
rect 5972 12664 5973 12704
rect 5931 12655 5973 12664
rect 6315 12704 6357 12713
rect 6315 12664 6316 12704
rect 6356 12664 6357 12704
rect 6315 12655 6357 12664
rect 7563 12704 7605 12713
rect 7563 12664 7564 12704
rect 7604 12664 7605 12704
rect 7563 12655 7605 12664
rect 9562 12704 9620 12705
rect 9562 12664 9571 12704
rect 9611 12664 9620 12704
rect 9562 12663 9620 12664
rect 11002 12704 11060 12705
rect 11002 12664 11011 12704
rect 11051 12664 11060 12704
rect 11002 12663 11060 12664
rect 11499 12704 11541 12713
rect 11499 12664 11500 12704
rect 11540 12664 11541 12704
rect 11499 12655 11541 12664
rect 12795 12704 12837 12713
rect 12795 12664 12796 12704
rect 12836 12664 12837 12704
rect 12795 12655 12837 12664
rect 13707 12704 13749 12713
rect 13707 12664 13708 12704
rect 13748 12664 13749 12704
rect 13707 12655 13749 12664
rect 15051 12704 15093 12713
rect 15051 12664 15052 12704
rect 15092 12664 15093 12704
rect 15051 12655 15093 12664
rect 15730 12704 15788 12705
rect 15730 12664 15739 12704
rect 15779 12664 15788 12704
rect 15730 12663 15788 12664
rect 16011 12704 16053 12713
rect 16011 12664 16012 12704
rect 16052 12664 16053 12704
rect 16011 12655 16053 12664
rect 17019 12704 17061 12713
rect 17019 12664 17020 12704
rect 17060 12664 17061 12704
rect 17019 12655 17061 12664
rect 18682 12704 18740 12705
rect 18682 12664 18691 12704
rect 18731 12664 18740 12704
rect 18682 12663 18740 12664
rect 20235 12704 20277 12713
rect 20235 12664 20236 12704
rect 20276 12664 20277 12704
rect 20235 12655 20277 12664
rect 29739 12704 29781 12713
rect 29739 12664 29740 12704
rect 29780 12664 29781 12704
rect 29739 12655 29781 12664
rect 2489 12620 2531 12629
rect 2489 12580 2490 12620
rect 2530 12580 2531 12620
rect 2489 12571 2531 12580
rect 2938 12620 2996 12621
rect 16714 12620 16772 12621
rect 2938 12580 2947 12620
rect 2987 12580 2996 12620
rect 2938 12579 2996 12580
rect 9858 12611 9904 12620
rect 9858 12571 9859 12611
rect 9899 12571 9904 12611
rect 16714 12580 16723 12620
rect 16763 12580 16772 12620
rect 16714 12579 16772 12580
rect 18795 12620 18837 12629
rect 18795 12580 18796 12620
rect 18836 12580 18837 12620
rect 18795 12571 18837 12580
rect 30123 12620 30165 12629
rect 30123 12580 30124 12620
rect 30164 12580 30165 12620
rect 30123 12571 30165 12580
rect 9858 12562 9904 12571
rect 939 12536 981 12545
rect 939 12496 940 12536
rect 980 12496 981 12536
rect 939 12487 981 12496
rect 1066 12536 1124 12537
rect 1066 12496 1075 12536
rect 1115 12496 1124 12536
rect 1066 12495 1124 12496
rect 1594 12536 1652 12537
rect 1594 12496 1603 12536
rect 1643 12496 1652 12536
rect 1594 12495 1652 12496
rect 1707 12536 1749 12545
rect 1707 12496 1708 12536
rect 1748 12496 1749 12536
rect 1707 12487 1749 12496
rect 2170 12536 2228 12537
rect 2170 12496 2179 12536
rect 2219 12496 2228 12536
rect 2170 12495 2228 12496
rect 2283 12536 2325 12545
rect 2283 12496 2284 12536
rect 2324 12496 2325 12536
rect 2283 12487 2325 12496
rect 2614 12536 2656 12545
rect 2614 12496 2615 12536
rect 2655 12496 2656 12536
rect 2614 12487 2656 12496
rect 2859 12536 2901 12545
rect 2859 12496 2860 12536
rect 2900 12496 2901 12536
rect 2859 12487 2901 12496
rect 3958 12536 4000 12545
rect 3958 12496 3959 12536
rect 3999 12496 4000 12536
rect 3958 12487 4000 12496
rect 4090 12536 4148 12537
rect 4090 12496 4099 12536
rect 4139 12496 4148 12536
rect 4090 12495 4148 12496
rect 4203 12536 4245 12545
rect 4203 12496 4204 12536
rect 4244 12496 4245 12536
rect 4203 12487 4245 12496
rect 4779 12536 4821 12545
rect 4779 12496 4780 12536
rect 4820 12496 4821 12536
rect 4779 12487 4821 12496
rect 5067 12536 5109 12545
rect 5067 12496 5068 12536
rect 5108 12496 5109 12536
rect 5067 12487 5109 12496
rect 5259 12536 5301 12545
rect 5259 12496 5260 12536
rect 5300 12496 5301 12536
rect 5259 12487 5301 12496
rect 5451 12536 5493 12545
rect 5451 12496 5452 12536
rect 5492 12496 5493 12536
rect 5451 12487 5493 12496
rect 5835 12536 5877 12545
rect 5835 12496 5836 12536
rect 5876 12496 5877 12536
rect 5835 12487 5877 12496
rect 6010 12536 6068 12537
rect 6010 12496 6019 12536
rect 6059 12496 6068 12536
rect 6010 12495 6068 12496
rect 6222 12536 6280 12537
rect 6222 12496 6231 12536
rect 6271 12496 6280 12536
rect 6222 12495 6280 12496
rect 6394 12536 6452 12537
rect 6394 12496 6403 12536
rect 6443 12496 6452 12536
rect 6394 12495 6452 12496
rect 7083 12536 7125 12545
rect 7083 12496 7084 12536
rect 7124 12496 7125 12536
rect 7083 12487 7125 12496
rect 7467 12536 7509 12545
rect 7467 12496 7468 12536
rect 7508 12496 7509 12536
rect 7467 12487 7509 12496
rect 8314 12536 8372 12537
rect 8314 12496 8323 12536
rect 8363 12496 8372 12536
rect 8314 12495 8372 12496
rect 8667 12536 8709 12545
rect 8667 12496 8668 12536
rect 8708 12496 8709 12536
rect 8667 12487 8709 12496
rect 8968 12536 9010 12545
rect 8968 12496 8969 12536
rect 9009 12496 9010 12536
rect 8968 12487 9010 12496
rect 9130 12536 9188 12537
rect 9130 12496 9139 12536
rect 9179 12496 9188 12536
rect 9130 12495 9188 12496
rect 9562 12536 9620 12537
rect 9942 12536 10000 12537
rect 9562 12496 9571 12536
rect 9611 12496 9620 12536
rect 9562 12495 9620 12496
rect 9675 12527 9717 12536
rect 9675 12487 9676 12527
rect 9716 12487 9717 12527
rect 9942 12496 9951 12536
rect 9991 12496 10000 12536
rect 10347 12536 10389 12545
rect 9942 12495 10000 12496
rect 10123 12525 10181 12526
rect 9675 12478 9717 12487
rect 10123 12485 10132 12525
rect 10172 12485 10181 12525
rect 10347 12496 10348 12536
rect 10388 12496 10389 12536
rect 10347 12487 10389 12496
rect 10462 12536 10504 12545
rect 10462 12496 10463 12536
rect 10503 12496 10504 12536
rect 10462 12487 10504 12496
rect 10635 12536 10677 12545
rect 10635 12496 10636 12536
rect 10676 12496 10677 12536
rect 10635 12487 10677 12496
rect 11163 12536 11205 12545
rect 11163 12496 11164 12536
rect 11204 12496 11205 12536
rect 11163 12487 11205 12496
rect 11307 12536 11349 12545
rect 11307 12496 11308 12536
rect 11348 12496 11349 12536
rect 11307 12487 11349 12496
rect 11595 12536 11637 12545
rect 11595 12496 11596 12536
rect 11636 12496 11637 12536
rect 11595 12487 11637 12496
rect 11824 12536 11882 12537
rect 11824 12496 11833 12536
rect 11873 12496 11882 12536
rect 11824 12495 11882 12496
rect 11979 12536 12021 12545
rect 11979 12496 11980 12536
rect 12020 12496 12021 12536
rect 11979 12487 12021 12496
rect 12171 12536 12213 12545
rect 12171 12496 12172 12536
rect 12212 12496 12213 12536
rect 12171 12487 12213 12496
rect 12607 12536 12665 12537
rect 12607 12496 12616 12536
rect 12656 12496 12665 12536
rect 12607 12495 12665 12496
rect 13083 12536 13125 12545
rect 13083 12496 13084 12536
rect 13124 12496 13125 12536
rect 13083 12487 13125 12496
rect 13419 12536 13461 12545
rect 13419 12496 13420 12536
rect 13460 12496 13461 12536
rect 13419 12487 13461 12496
rect 13803 12536 13845 12545
rect 13803 12496 13804 12536
rect 13844 12496 13845 12536
rect 13803 12487 13845 12496
rect 14032 12536 14090 12537
rect 14032 12496 14041 12536
rect 14081 12496 14090 12536
rect 14032 12495 14090 12496
rect 14650 12536 14708 12537
rect 14650 12496 14659 12536
rect 14699 12496 14708 12536
rect 14650 12495 14708 12496
rect 14763 12536 14805 12545
rect 15915 12536 15957 12545
rect 14763 12496 14764 12536
rect 14804 12496 14805 12536
rect 14763 12487 14805 12496
rect 15519 12527 15561 12536
rect 15519 12487 15520 12527
rect 15560 12487 15561 12527
rect 15915 12496 15916 12536
rect 15956 12496 15957 12536
rect 10123 12484 10181 12485
rect 15519 12478 15561 12487
rect 15610 12494 15668 12495
rect 2746 12452 2804 12453
rect 2746 12412 2755 12452
rect 2795 12412 2804 12452
rect 2746 12411 2804 12412
rect 7930 12452 7988 12453
rect 7930 12412 7939 12452
rect 7979 12412 7988 12452
rect 7930 12411 7988 12412
rect 8506 12452 8564 12453
rect 8506 12412 8515 12452
rect 8555 12412 8564 12452
rect 8506 12411 8564 12412
rect 8811 12452 8853 12461
rect 13922 12452 13964 12461
rect 15610 12454 15619 12494
rect 15659 12454 15668 12494
rect 15915 12487 15957 12496
rect 16107 12536 16149 12545
rect 16107 12496 16108 12536
rect 16148 12496 16149 12536
rect 16107 12487 16149 12496
rect 16909 12536 16967 12537
rect 16909 12496 16918 12536
rect 16958 12496 16967 12536
rect 16909 12495 16967 12496
rect 17163 12536 17205 12545
rect 17163 12496 17164 12536
rect 17204 12496 17205 12536
rect 17163 12487 17205 12496
rect 17878 12536 17920 12545
rect 17878 12496 17879 12536
rect 17919 12496 17920 12536
rect 17878 12487 17920 12496
rect 18123 12536 18165 12545
rect 18123 12496 18124 12536
rect 18164 12496 18165 12536
rect 18123 12487 18165 12496
rect 18589 12536 18631 12545
rect 19659 12536 19701 12545
rect 18589 12496 18590 12536
rect 18630 12496 18631 12536
rect 18589 12487 18631 12496
rect 18891 12527 18933 12536
rect 18891 12487 18892 12527
rect 18932 12487 18933 12527
rect 19659 12496 19660 12536
rect 19700 12496 19701 12536
rect 19659 12487 19701 12496
rect 22138 12536 22196 12537
rect 22138 12496 22147 12536
rect 22187 12496 22196 12536
rect 22138 12495 22196 12496
rect 23053 12536 23111 12537
rect 23053 12496 23062 12536
rect 23102 12496 23111 12536
rect 23053 12495 23111 12496
rect 25402 12536 25460 12537
rect 25402 12496 25411 12536
rect 25451 12496 25460 12536
rect 25402 12495 25460 12496
rect 25995 12536 26037 12545
rect 25995 12496 25996 12536
rect 26036 12496 26037 12536
rect 25995 12487 26037 12496
rect 26187 12536 26229 12545
rect 26187 12496 26188 12536
rect 26228 12496 26229 12536
rect 26187 12487 26229 12496
rect 26746 12536 26804 12537
rect 26746 12496 26755 12536
rect 26795 12496 26804 12536
rect 26746 12495 26804 12496
rect 29643 12536 29685 12545
rect 29643 12496 29644 12536
rect 29684 12496 29685 12536
rect 29643 12487 29685 12496
rect 29816 12536 29858 12545
rect 29816 12496 29817 12536
rect 29857 12496 29858 12536
rect 29816 12487 29858 12496
rect 30027 12536 30069 12545
rect 30027 12496 30028 12536
rect 30068 12496 30069 12536
rect 30027 12487 30069 12496
rect 30219 12536 30261 12545
rect 30219 12496 30220 12536
rect 30260 12496 30261 12536
rect 30219 12487 30261 12496
rect 18891 12478 18933 12487
rect 15610 12453 15668 12454
rect 8811 12412 8812 12452
rect 8852 12412 8853 12452
rect 8811 12403 8853 12412
rect 11730 12443 11776 12452
rect 11730 12403 11731 12443
rect 11771 12403 11776 12443
rect 13922 12412 13923 12452
rect 13963 12412 13964 12452
rect 13922 12403 13964 12412
rect 18010 12452 18068 12453
rect 18010 12412 18019 12452
rect 18059 12412 18068 12452
rect 18010 12411 18068 12412
rect 18219 12452 18261 12461
rect 18219 12412 18220 12452
rect 18260 12412 18261 12452
rect 18219 12403 18261 12412
rect 19569 12452 19611 12461
rect 19569 12412 19570 12452
rect 19610 12412 19611 12452
rect 19569 12403 19611 12412
rect 20602 12452 20660 12453
rect 20602 12412 20611 12452
rect 20651 12412 20660 12452
rect 20602 12411 20660 12412
rect 22522 12452 22580 12453
rect 22522 12412 22531 12452
rect 22571 12412 22580 12452
rect 22522 12411 22580 12412
rect 22858 12452 22916 12453
rect 22858 12412 22867 12452
rect 22907 12412 22916 12452
rect 22858 12411 22916 12412
rect 23866 12452 23924 12453
rect 23866 12412 23875 12452
rect 23915 12412 23924 12452
rect 23866 12411 23924 12412
rect 25786 12452 25844 12453
rect 25786 12412 25795 12452
rect 25835 12412 25844 12452
rect 25786 12411 25844 12412
rect 26379 12452 26421 12461
rect 26379 12412 26380 12452
rect 26420 12412 26421 12452
rect 26379 12403 26421 12412
rect 28299 12452 28341 12461
rect 28299 12412 28300 12452
rect 28340 12412 28341 12452
rect 28299 12403 28341 12412
rect 11730 12394 11776 12403
rect 8026 12368 8084 12369
rect 8026 12328 8035 12368
rect 8075 12328 8084 12368
rect 8026 12327 8084 12328
rect 8907 12368 8949 12377
rect 8907 12328 8908 12368
rect 8948 12328 8949 12368
rect 8907 12319 8949 12328
rect 10347 12368 10389 12377
rect 10347 12328 10348 12368
rect 10388 12328 10389 12368
rect 10347 12319 10389 12328
rect 11979 12368 12021 12377
rect 11979 12328 11980 12368
rect 12020 12328 12021 12368
rect 11979 12319 12021 12328
rect 15226 12368 15284 12369
rect 15226 12328 15235 12368
rect 15275 12328 15284 12368
rect 15226 12327 15284 12328
rect 20235 12368 20277 12377
rect 20235 12328 20236 12368
rect 20276 12328 20277 12368
rect 20235 12319 20277 12328
rect 25995 12368 26037 12377
rect 25995 12328 25996 12368
rect 26036 12328 26037 12368
rect 25995 12319 26037 12328
rect 28875 12368 28917 12377
rect 28875 12328 28876 12368
rect 28916 12328 28917 12368
rect 28875 12319 28917 12328
rect 29259 12368 29301 12377
rect 29259 12328 29260 12368
rect 29300 12328 29301 12368
rect 29259 12319 29301 12328
rect 30507 12368 30549 12377
rect 30507 12328 30508 12368
rect 30548 12328 30549 12368
rect 30507 12319 30549 12328
rect 30891 12368 30933 12377
rect 30891 12328 30892 12368
rect 30932 12328 30933 12368
rect 30891 12319 30933 12328
rect 5259 12284 5301 12293
rect 5259 12244 5260 12284
rect 5300 12244 5301 12284
rect 5259 12235 5301 12244
rect 13210 12284 13268 12285
rect 13210 12244 13219 12284
rect 13259 12244 13268 12284
rect 13210 12243 13268 12244
rect 19467 12284 19509 12293
rect 19467 12244 19468 12284
rect 19508 12244 19509 12284
rect 19467 12235 19509 12244
rect 23499 12284 23541 12293
rect 23499 12244 23500 12284
rect 23540 12244 23541 12284
rect 23499 12235 23541 12244
rect 28683 12284 28725 12293
rect 28683 12244 28684 12284
rect 28724 12244 28725 12284
rect 28683 12235 28725 12244
rect 576 12116 31392 12140
rect 576 12076 3112 12116
rect 3480 12076 10886 12116
rect 11254 12076 18660 12116
rect 19028 12076 26434 12116
rect 26802 12076 31392 12116
rect 576 12052 31392 12076
rect 1419 11948 1461 11957
rect 1419 11908 1420 11948
rect 1460 11908 1461 11948
rect 1419 11899 1461 11908
rect 2283 11948 2325 11957
rect 2283 11908 2284 11948
rect 2324 11908 2325 11948
rect 2283 11899 2325 11908
rect 4779 11948 4821 11957
rect 4779 11908 4780 11948
rect 4820 11908 4821 11948
rect 4779 11899 4821 11908
rect 5643 11948 5685 11957
rect 5643 11908 5644 11948
rect 5684 11908 5685 11948
rect 5643 11899 5685 11908
rect 6603 11948 6645 11957
rect 6603 11908 6604 11948
rect 6644 11908 6645 11948
rect 6603 11899 6645 11908
rect 9466 11948 9524 11949
rect 9466 11908 9475 11948
rect 9515 11908 9524 11948
rect 9466 11907 9524 11908
rect 10059 11948 10101 11957
rect 10059 11908 10060 11948
rect 10100 11908 10101 11948
rect 10059 11899 10101 11908
rect 11770 11948 11828 11949
rect 11770 11908 11779 11948
rect 11819 11908 11828 11948
rect 11770 11907 11828 11908
rect 12922 11948 12980 11949
rect 12922 11908 12931 11948
rect 12971 11908 12980 11948
rect 12922 11907 12980 11908
rect 15339 11948 15381 11957
rect 15339 11908 15340 11948
rect 15380 11908 15381 11948
rect 15339 11899 15381 11908
rect 16090 11948 16148 11949
rect 16090 11908 16099 11948
rect 16139 11908 16148 11948
rect 16090 11907 16148 11908
rect 17355 11948 17397 11957
rect 17355 11908 17356 11948
rect 17396 11908 17397 11948
rect 17355 11899 17397 11908
rect 18106 11948 18164 11949
rect 18106 11908 18115 11948
rect 18155 11908 18164 11948
rect 18106 11907 18164 11908
rect 18586 11948 18644 11949
rect 18586 11908 18595 11948
rect 18635 11908 18644 11948
rect 18586 11907 18644 11908
rect 20427 11948 20469 11957
rect 20427 11908 20428 11948
rect 20468 11908 20469 11948
rect 20427 11899 20469 11908
rect 21675 11948 21717 11957
rect 21675 11908 21676 11948
rect 21716 11908 21717 11948
rect 21675 11899 21717 11908
rect 23482 11948 23540 11949
rect 23482 11908 23491 11948
rect 23531 11908 23540 11948
rect 23482 11907 23540 11908
rect 24075 11948 24117 11957
rect 24075 11908 24076 11948
rect 24116 11908 24117 11948
rect 24075 11899 24117 11908
rect 27147 11948 27189 11957
rect 27147 11908 27148 11948
rect 27188 11908 27189 11948
rect 27147 11899 27189 11908
rect 28587 11948 28629 11957
rect 28587 11908 28588 11948
rect 28628 11908 28629 11948
rect 28587 11899 28629 11908
rect 29146 11948 29204 11949
rect 29146 11908 29155 11948
rect 29195 11908 29204 11948
rect 29146 11907 29204 11908
rect 30315 11948 30357 11957
rect 30315 11908 30316 11948
rect 30356 11908 30357 11948
rect 30315 11899 30357 11908
rect 30699 11948 30741 11957
rect 30699 11908 30700 11948
rect 30740 11908 30741 11948
rect 30699 11899 30741 11908
rect 3339 11864 3381 11873
rect 3339 11824 3340 11864
rect 3380 11824 3381 11864
rect 3339 11815 3381 11824
rect 6123 11864 6165 11873
rect 6123 11824 6124 11864
rect 6164 11824 6165 11864
rect 6123 11815 6165 11824
rect 7258 11864 7316 11865
rect 7258 11824 7267 11864
rect 7307 11824 7316 11864
rect 7258 11823 7316 11824
rect 21963 11864 22005 11873
rect 29355 11864 29397 11873
rect 21963 11824 21964 11864
rect 22004 11824 22005 11864
rect 21963 11815 22005 11824
rect 24315 11855 24357 11864
rect 24315 11815 24316 11855
rect 24356 11815 24357 11855
rect 29355 11824 29356 11864
rect 29396 11824 29397 11864
rect 29355 11815 29397 11824
rect 30987 11864 31029 11873
rect 30987 11824 30988 11864
rect 31028 11824 31029 11864
rect 30987 11815 31029 11824
rect 24315 11806 24357 11815
rect 1995 11780 2037 11789
rect 1995 11740 1996 11780
rect 2036 11740 2037 11780
rect 1995 11731 2037 11740
rect 7761 11780 7803 11789
rect 7761 11740 7762 11780
rect 7802 11740 7803 11780
rect 4495 11729 4537 11738
rect 7761 11731 7803 11740
rect 10587 11780 10629 11789
rect 12945 11780 12987 11789
rect 10587 11740 10588 11780
rect 10628 11740 10629 11780
rect 8650 11738 8708 11739
rect 939 11696 981 11705
rect 939 11656 940 11696
rect 980 11656 981 11696
rect 939 11647 981 11656
rect 1114 11696 1172 11697
rect 1114 11656 1123 11696
rect 1163 11656 1172 11696
rect 1114 11655 1172 11656
rect 1314 11696 1372 11697
rect 1314 11656 1323 11696
rect 1363 11656 1372 11696
rect 1314 11655 1372 11656
rect 1514 11696 1556 11705
rect 1514 11656 1515 11696
rect 1555 11656 1556 11696
rect 1514 11647 1556 11656
rect 1659 11696 1701 11705
rect 1659 11656 1660 11696
rect 1700 11656 1701 11696
rect 1659 11647 1701 11656
rect 1786 11696 1844 11697
rect 1786 11656 1795 11696
rect 1835 11656 1844 11696
rect 1786 11655 1844 11656
rect 1899 11696 1941 11705
rect 1899 11656 1900 11696
rect 1940 11656 1941 11696
rect 1899 11647 1941 11656
rect 2187 11696 2229 11705
rect 2187 11656 2188 11696
rect 2228 11656 2229 11696
rect 2187 11647 2229 11656
rect 2379 11696 2421 11705
rect 2379 11656 2380 11696
rect 2420 11656 2421 11696
rect 2379 11647 2421 11656
rect 2667 11696 2709 11705
rect 2667 11656 2668 11696
rect 2708 11656 2709 11696
rect 2667 11647 2709 11656
rect 3147 11696 3189 11705
rect 3147 11656 3148 11696
rect 3188 11656 3189 11696
rect 3147 11647 3189 11656
rect 3531 11696 3573 11705
rect 3531 11656 3532 11696
rect 3572 11656 3573 11696
rect 3531 11647 3573 11656
rect 3915 11696 3957 11705
rect 3915 11656 3916 11696
rect 3956 11656 3957 11696
rect 3915 11647 3957 11656
rect 4378 11696 4436 11697
rect 4378 11656 4387 11696
rect 4427 11656 4436 11696
rect 4495 11689 4496 11729
rect 4536 11689 4537 11729
rect 4495 11680 4537 11689
rect 4971 11696 5013 11705
rect 4378 11655 4436 11656
rect 4971 11656 4972 11696
rect 5012 11656 5013 11696
rect 4971 11647 5013 11656
rect 5163 11696 5205 11705
rect 5163 11656 5164 11696
rect 5204 11656 5205 11696
rect 5163 11647 5205 11656
rect 5338 11696 5396 11697
rect 5338 11656 5347 11696
rect 5387 11656 5396 11696
rect 5338 11655 5396 11656
rect 5931 11696 5973 11705
rect 5931 11656 5932 11696
rect 5972 11656 5973 11696
rect 5931 11647 5973 11656
rect 6298 11696 6356 11697
rect 6298 11656 6307 11696
rect 6347 11656 6356 11696
rect 6298 11655 6356 11656
rect 6970 11696 7028 11697
rect 6970 11656 6979 11696
rect 7019 11656 7028 11696
rect 6970 11655 7028 11656
rect 7083 11696 7125 11705
rect 7083 11656 7084 11696
rect 7124 11656 7125 11696
rect 7083 11647 7125 11656
rect 7851 11696 7893 11705
rect 8650 11698 8659 11738
rect 8699 11698 8708 11738
rect 10587 11731 10629 11740
rect 12498 11771 12544 11780
rect 12498 11731 12499 11771
rect 12539 11731 12544 11771
rect 12945 11740 12946 11780
rect 12986 11740 12987 11780
rect 12945 11731 12987 11740
rect 13594 11780 13652 11781
rect 13594 11740 13603 11780
rect 13643 11740 13652 11780
rect 13594 11739 13652 11740
rect 15915 11780 15957 11789
rect 15915 11740 15916 11780
rect 15956 11740 15957 11780
rect 15915 11731 15957 11740
rect 19210 11780 19268 11781
rect 19210 11740 19219 11780
rect 19259 11740 19268 11780
rect 19210 11739 19268 11740
rect 19978 11780 20036 11781
rect 19978 11740 19987 11780
rect 20027 11740 20036 11780
rect 19978 11739 20036 11740
rect 20529 11780 20571 11789
rect 20529 11740 20530 11780
rect 20570 11740 20571 11780
rect 20170 11738 20228 11739
rect 12498 11722 12544 11731
rect 17067 11717 17109 11726
rect 8650 11697 8708 11698
rect 7851 11656 7852 11696
rect 7892 11656 7893 11696
rect 7851 11647 7893 11656
rect 8791 11696 8849 11697
rect 8791 11656 8800 11696
rect 8840 11656 8849 11696
rect 8791 11655 8849 11656
rect 9291 11696 9333 11705
rect 9291 11656 9292 11696
rect 9332 11656 9333 11696
rect 9291 11647 9333 11656
rect 9466 11696 9524 11697
rect 9466 11656 9475 11696
rect 9515 11656 9524 11696
rect 9466 11655 9524 11656
rect 9850 11696 9908 11697
rect 9850 11656 9859 11696
rect 9899 11656 9908 11696
rect 9850 11655 9908 11656
rect 9963 11696 10005 11705
rect 9963 11656 9964 11696
rect 10004 11656 10005 11696
rect 9963 11647 10005 11656
rect 10423 11696 10481 11697
rect 10423 11656 10432 11696
rect 10472 11656 10481 11696
rect 10423 11655 10481 11656
rect 11019 11696 11061 11705
rect 11019 11656 11020 11696
rect 11060 11656 11061 11696
rect 11019 11647 11061 11656
rect 11307 11696 11349 11705
rect 11307 11656 11308 11696
rect 11348 11656 11349 11696
rect 11307 11647 11349 11656
rect 12067 11696 12125 11697
rect 12067 11656 12076 11696
rect 12116 11656 12125 11696
rect 12067 11655 12125 11656
rect 12363 11696 12405 11705
rect 12363 11656 12364 11696
rect 12404 11656 12405 11696
rect 12363 11647 12405 11656
rect 12592 11696 12650 11697
rect 12592 11656 12601 11696
rect 12641 11656 12650 11696
rect 12592 11655 12650 11656
rect 13035 11696 13077 11705
rect 13035 11656 13036 11696
rect 13076 11656 13077 11696
rect 13035 11647 13077 11656
rect 13474 11696 13532 11697
rect 13474 11656 13483 11696
rect 13523 11656 13532 11696
rect 13474 11655 13532 11656
rect 13707 11696 13749 11705
rect 13707 11656 13708 11696
rect 13748 11656 13749 11696
rect 13707 11647 13749 11656
rect 14475 11696 14517 11705
rect 14475 11656 14476 11696
rect 14516 11656 14517 11696
rect 14475 11647 14517 11656
rect 14563 11696 14621 11697
rect 14563 11656 14572 11696
rect 14612 11656 14621 11696
rect 14563 11655 14621 11656
rect 14822 11696 14880 11697
rect 14822 11656 14831 11696
rect 14871 11656 14880 11696
rect 14822 11655 14880 11656
rect 14960 11696 15002 11705
rect 14960 11656 14961 11696
rect 15001 11656 15002 11696
rect 14960 11647 15002 11656
rect 15082 11696 15140 11697
rect 15082 11656 15091 11696
rect 15131 11656 15140 11696
rect 15082 11655 15140 11656
rect 15226 11696 15284 11697
rect 15226 11656 15235 11696
rect 15275 11656 15284 11696
rect 15226 11655 15284 11656
rect 15348 11696 15406 11697
rect 15348 11656 15357 11696
rect 15397 11656 15406 11696
rect 15348 11655 15406 11656
rect 15574 11696 15616 11705
rect 15574 11656 15575 11696
rect 15615 11656 15616 11696
rect 15574 11647 15616 11656
rect 15706 11696 15764 11697
rect 15706 11656 15715 11696
rect 15755 11656 15764 11696
rect 15706 11655 15764 11656
rect 15819 11696 15861 11705
rect 15819 11656 15820 11696
rect 15860 11656 15861 11696
rect 15819 11647 15861 11656
rect 16101 11696 16159 11697
rect 16101 11656 16110 11696
rect 16150 11656 16159 11696
rect 16101 11655 16159 11656
rect 16208 11696 16266 11697
rect 16208 11656 16217 11696
rect 16257 11656 16266 11696
rect 16208 11655 16266 11656
rect 16348 11696 16406 11697
rect 16348 11656 16357 11696
rect 16397 11656 16406 11696
rect 16348 11655 16406 11656
rect 16474 11696 16532 11697
rect 16474 11656 16483 11696
rect 16523 11656 16532 11696
rect 16474 11655 16532 11656
rect 16651 11696 16709 11697
rect 16651 11656 16660 11696
rect 16700 11656 16709 11696
rect 16651 11655 16709 11656
rect 16954 11696 17012 11697
rect 16954 11656 16963 11696
rect 17003 11656 17012 11696
rect 17067 11677 17068 11717
rect 17108 11677 17109 11717
rect 17067 11668 17109 11677
rect 17547 11696 17589 11705
rect 16954 11655 17012 11656
rect 17547 11656 17548 11696
rect 17588 11656 17589 11696
rect 17547 11647 17589 11656
rect 17722 11696 17780 11697
rect 17722 11656 17731 11696
rect 17771 11656 17780 11696
rect 17722 11655 17780 11656
rect 18405 11696 18463 11697
rect 18405 11656 18414 11696
rect 18454 11656 18463 11696
rect 18405 11655 18463 11656
rect 18795 11696 18837 11705
rect 20170 11698 20179 11738
rect 20219 11698 20228 11738
rect 20529 11731 20571 11740
rect 21243 11780 21285 11789
rect 21243 11740 21244 11780
rect 21284 11740 21285 11780
rect 21243 11731 21285 11740
rect 25594 11780 25652 11781
rect 25594 11740 25603 11780
rect 25643 11740 25652 11780
rect 25594 11739 25652 11740
rect 27249 11780 27291 11789
rect 27249 11740 27250 11780
rect 27290 11740 27291 11780
rect 27249 11731 27291 11740
rect 20170 11697 20228 11698
rect 18795 11656 18796 11696
rect 18836 11656 18837 11696
rect 18795 11647 18837 11656
rect 18883 11696 18941 11697
rect 18883 11656 18892 11696
rect 18932 11656 18941 11696
rect 18883 11655 18941 11656
rect 19375 11696 19433 11697
rect 19375 11656 19384 11696
rect 19424 11656 19433 11696
rect 19375 11655 19433 11656
rect 20619 11696 20661 11705
rect 20619 11656 20620 11696
rect 20660 11656 20661 11696
rect 20619 11647 20661 11656
rect 21034 11696 21092 11697
rect 21034 11656 21043 11696
rect 21083 11656 21092 11696
rect 21034 11655 21092 11656
rect 21771 11696 21813 11705
rect 21771 11656 21772 11696
rect 21812 11656 21813 11696
rect 21771 11647 21813 11656
rect 22827 11696 22869 11705
rect 22827 11656 22828 11696
rect 22868 11656 22869 11696
rect 22827 11647 22869 11656
rect 23115 11696 23157 11705
rect 23115 11656 23116 11696
rect 23156 11656 23157 11696
rect 23115 11647 23157 11656
rect 23307 11696 23349 11705
rect 23307 11656 23308 11696
rect 23348 11656 23349 11696
rect 23307 11647 23349 11656
rect 23482 11696 23540 11697
rect 23482 11656 23491 11696
rect 23531 11656 23540 11696
rect 23482 11655 23540 11656
rect 24250 11696 24308 11697
rect 24250 11656 24259 11696
rect 24299 11656 24308 11696
rect 24250 11655 24308 11656
rect 25131 11696 25173 11705
rect 25131 11656 25132 11696
rect 25172 11656 25173 11696
rect 25131 11647 25173 11656
rect 25995 11696 26037 11705
rect 25995 11656 25996 11696
rect 26036 11656 26037 11696
rect 25995 11647 26037 11656
rect 26475 11696 26517 11705
rect 26475 11656 26476 11696
rect 26516 11656 26517 11696
rect 26475 11647 26517 11656
rect 26859 11696 26901 11705
rect 26859 11656 26860 11696
rect 26900 11656 26901 11696
rect 26859 11647 26901 11656
rect 27339 11696 27381 11705
rect 27339 11656 27340 11696
rect 27380 11656 27381 11696
rect 27339 11647 27381 11656
rect 27963 11696 28005 11705
rect 27963 11656 27964 11696
rect 28004 11656 28005 11696
rect 27963 11647 28005 11656
rect 28107 11696 28149 11705
rect 28107 11656 28108 11696
rect 28148 11656 28149 11696
rect 28107 11647 28149 11656
rect 28587 11696 28629 11705
rect 28587 11656 28588 11696
rect 28628 11656 28629 11696
rect 28587 11647 28629 11656
rect 28779 11696 28821 11705
rect 28779 11656 28780 11696
rect 28820 11656 28821 11696
rect 28779 11647 28821 11656
rect 28971 11696 29013 11705
rect 28971 11656 28972 11696
rect 29012 11656 29013 11696
rect 28971 11647 29013 11656
rect 29140 11696 29182 11705
rect 29140 11656 29141 11696
rect 29181 11656 29182 11696
rect 29140 11647 29182 11656
rect 29355 11696 29397 11705
rect 29355 11656 29356 11696
rect 29396 11656 29397 11696
rect 29355 11647 29397 11656
rect 29547 11696 29589 11705
rect 29547 11656 29548 11696
rect 29588 11656 29589 11696
rect 29547 11647 29589 11656
rect 29739 11696 29781 11705
rect 29739 11656 29740 11696
rect 29780 11656 29781 11696
rect 29739 11647 29781 11656
rect 29931 11696 29973 11705
rect 29931 11656 29932 11696
rect 29972 11656 29973 11696
rect 29931 11647 29973 11656
rect 30219 11696 30261 11705
rect 30219 11656 30220 11696
rect 30260 11656 30261 11696
rect 30219 11647 30261 11656
rect 30411 11696 30453 11705
rect 30411 11656 30412 11696
rect 30452 11656 30453 11696
rect 30411 11647 30453 11656
rect 30603 11696 30645 11705
rect 30603 11656 30604 11696
rect 30644 11656 30645 11696
rect 30603 11647 30645 11656
rect 30795 11696 30837 11705
rect 30795 11656 30796 11696
rect 30836 11656 30837 11696
rect 30795 11647 30837 11656
rect 2283 11612 2325 11621
rect 2283 11572 2284 11612
rect 2324 11572 2325 11612
rect 2283 11563 2325 11572
rect 5067 11612 5109 11621
rect 5067 11572 5068 11612
rect 5108 11572 5109 11612
rect 5067 11563 5109 11572
rect 5451 11612 5493 11621
rect 5451 11572 5452 11612
rect 5492 11572 5493 11612
rect 5451 11563 5493 11572
rect 5657 11612 5699 11621
rect 5657 11572 5658 11612
rect 5698 11572 5699 11612
rect 5657 11563 5699 11572
rect 6411 11612 6453 11621
rect 6411 11572 6412 11612
rect 6452 11572 6453 11612
rect 6411 11563 6453 11572
rect 6617 11612 6659 11621
rect 6617 11572 6618 11612
rect 6658 11572 6659 11612
rect 6617 11563 6659 11572
rect 11776 11612 11818 11621
rect 11776 11572 11777 11612
rect 11817 11572 11818 11612
rect 11776 11563 11818 11572
rect 13786 11612 13844 11613
rect 13786 11572 13795 11612
rect 13835 11572 13844 11612
rect 13786 11571 13844 11572
rect 14270 11612 14312 11621
rect 14270 11572 14271 11612
rect 14311 11572 14312 11612
rect 14270 11563 14312 11572
rect 14362 11612 14420 11613
rect 14362 11572 14371 11612
rect 14411 11572 14420 11612
rect 14362 11571 14420 11572
rect 17643 11612 17685 11621
rect 17643 11572 17644 11612
rect 17684 11572 17685 11612
rect 17643 11563 17685 11572
rect 18109 11612 18151 11621
rect 18109 11572 18110 11612
rect 18150 11572 18151 11612
rect 18109 11563 18151 11572
rect 18589 11612 18631 11621
rect 18589 11572 18590 11612
rect 18630 11572 18631 11612
rect 18589 11563 18631 11572
rect 22491 11612 22533 11621
rect 22491 11572 22492 11612
rect 22532 11572 22533 11612
rect 22491 11563 22533 11572
rect 29835 11612 29877 11621
rect 29835 11572 29836 11612
rect 29876 11572 29877 11612
rect 29835 11563 29877 11572
rect 1035 11528 1077 11537
rect 1035 11488 1036 11528
rect 1076 11488 1077 11528
rect 1035 11479 1077 11488
rect 2554 11528 2612 11529
rect 2554 11488 2563 11528
rect 2603 11488 2612 11528
rect 2554 11487 2612 11488
rect 2859 11528 2901 11537
rect 2859 11488 2860 11528
rect 2900 11488 2901 11528
rect 2859 11479 2901 11488
rect 3034 11528 3092 11529
rect 3034 11488 3043 11528
rect 3083 11488 3092 11528
rect 3034 11487 3092 11488
rect 4011 11528 4053 11537
rect 5818 11528 5876 11529
rect 4011 11488 4012 11528
rect 4052 11488 4053 11528
rect 4011 11479 4053 11488
rect 4290 11519 4336 11528
rect 4290 11479 4291 11519
rect 4331 11479 4336 11519
rect 5818 11488 5827 11528
rect 5867 11488 5876 11528
rect 5818 11487 5876 11488
rect 7546 11528 7604 11529
rect 7546 11488 7555 11528
rect 7595 11488 7604 11528
rect 7546 11487 7604 11488
rect 8458 11528 8516 11529
rect 8458 11488 8467 11528
rect 8507 11488 8516 11528
rect 8458 11487 8516 11488
rect 8955 11528 8997 11537
rect 8955 11488 8956 11528
rect 8996 11488 8997 11528
rect 8955 11479 8997 11488
rect 11499 11528 11541 11537
rect 11499 11488 11500 11528
rect 11540 11488 11541 11528
rect 11499 11479 11541 11488
rect 11979 11528 12021 11537
rect 11979 11488 11980 11528
rect 12020 11488 12021 11528
rect 11979 11479 12021 11488
rect 12267 11528 12309 11537
rect 18315 11528 18357 11537
rect 12267 11488 12268 11528
rect 12308 11488 12309 11528
rect 12267 11479 12309 11488
rect 16866 11519 16912 11528
rect 16866 11479 16867 11519
rect 16907 11479 16912 11519
rect 18315 11488 18316 11528
rect 18356 11488 18357 11528
rect 18315 11479 18357 11488
rect 24939 11528 24981 11537
rect 24939 11488 24940 11528
rect 24980 11488 24981 11528
rect 24939 11479 24981 11488
rect 26362 11528 26420 11529
rect 26362 11488 26371 11528
rect 26411 11488 26420 11528
rect 26362 11487 26420 11488
rect 27802 11528 27860 11529
rect 27802 11488 27811 11528
rect 27851 11488 27860 11528
rect 27802 11487 27860 11488
rect 4290 11470 4336 11479
rect 16866 11470 16912 11479
rect 576 11360 31392 11384
rect 576 11320 4352 11360
rect 4720 11320 12126 11360
rect 12494 11320 19900 11360
rect 20268 11320 27674 11360
rect 28042 11320 31392 11360
rect 576 11296 31392 11320
rect 3802 11234 3860 11235
rect 1803 11192 1845 11201
rect 1803 11152 1804 11192
rect 1844 11152 1845 11192
rect 1803 11143 1845 11152
rect 2763 11192 2805 11201
rect 3802 11194 3811 11234
rect 3851 11194 3860 11234
rect 3802 11193 3860 11194
rect 2763 11152 2764 11192
rect 2804 11152 2805 11192
rect 2763 11143 2805 11152
rect 5146 11192 5204 11193
rect 5146 11152 5155 11192
rect 5195 11152 5204 11192
rect 5146 11151 5204 11152
rect 5914 11192 5972 11193
rect 5914 11152 5923 11192
rect 5963 11152 5972 11192
rect 5914 11151 5972 11152
rect 7659 11192 7701 11201
rect 7659 11152 7660 11192
rect 7700 11152 7701 11192
rect 7659 11143 7701 11152
rect 8427 11192 8469 11201
rect 8427 11152 8428 11192
rect 8468 11152 8469 11192
rect 8427 11143 8469 11152
rect 9466 11192 9524 11193
rect 9466 11152 9475 11192
rect 9515 11152 9524 11192
rect 9466 11151 9524 11152
rect 10042 11192 10100 11193
rect 10042 11152 10051 11192
rect 10091 11152 10100 11192
rect 10042 11151 10100 11152
rect 10731 11192 10773 11201
rect 10731 11152 10732 11192
rect 10772 11152 10773 11192
rect 10731 11143 10773 11152
rect 11307 11192 11349 11201
rect 11307 11152 11308 11192
rect 11348 11152 11349 11192
rect 11307 11143 11349 11152
rect 11883 11192 11925 11201
rect 11883 11152 11884 11192
rect 11924 11152 11925 11192
rect 11883 11143 11925 11152
rect 13323 11192 13365 11201
rect 13323 11152 13324 11192
rect 13364 11152 13365 11192
rect 13323 11143 13365 11152
rect 13594 11192 13652 11193
rect 13594 11152 13603 11192
rect 13643 11152 13652 11192
rect 13594 11151 13652 11152
rect 14475 11192 14517 11201
rect 14475 11152 14476 11192
rect 14516 11152 14517 11192
rect 14475 11143 14517 11152
rect 15819 11192 15861 11201
rect 15819 11152 15820 11192
rect 15860 11152 15861 11192
rect 15819 11143 15861 11152
rect 18394 11192 18452 11193
rect 18394 11152 18403 11192
rect 18443 11152 18452 11192
rect 18394 11151 18452 11152
rect 18795 11192 18837 11201
rect 18795 11152 18796 11192
rect 18836 11152 18837 11192
rect 18795 11143 18837 11152
rect 21082 11192 21140 11193
rect 21082 11152 21091 11192
rect 21131 11152 21140 11192
rect 21082 11151 21140 11152
rect 22570 11192 22628 11193
rect 22570 11152 22579 11192
rect 22619 11152 22628 11192
rect 22570 11151 22628 11152
rect 24363 11192 24405 11201
rect 24363 11152 24364 11192
rect 24404 11152 24405 11192
rect 24363 11143 24405 11152
rect 25402 11192 25460 11193
rect 25402 11152 25411 11192
rect 25451 11152 25460 11192
rect 25402 11151 25460 11152
rect 26667 11192 26709 11201
rect 26667 11152 26668 11192
rect 26708 11152 26709 11192
rect 26667 11143 26709 11152
rect 27130 11192 27188 11193
rect 27130 11152 27139 11192
rect 27179 11152 27188 11192
rect 27130 11151 27188 11152
rect 29355 11192 29397 11201
rect 29355 11152 29356 11192
rect 29396 11152 29397 11192
rect 29355 11143 29397 11152
rect 29643 11192 29685 11201
rect 29643 11152 29644 11192
rect 29684 11152 29685 11192
rect 29643 11143 29685 11152
rect 30123 11192 30165 11201
rect 30123 11152 30124 11192
rect 30164 11152 30165 11192
rect 30123 11143 30165 11152
rect 939 11108 981 11117
rect 939 11068 940 11108
rect 980 11068 981 11108
rect 939 11059 981 11068
rect 14266 11108 14324 11109
rect 14266 11068 14275 11108
rect 14315 11068 14324 11108
rect 14266 11067 14324 11068
rect 15339 11108 15381 11117
rect 15339 11068 15340 11108
rect 15380 11068 15381 11108
rect 15339 11059 15381 11068
rect 17835 11108 17877 11117
rect 17835 11068 17836 11108
rect 17876 11068 17877 11108
rect 17835 11059 17877 11068
rect 18507 11108 18549 11117
rect 18507 11068 18508 11108
rect 18548 11068 18549 11108
rect 18507 11059 18549 11068
rect 23355 11108 23397 11117
rect 23355 11068 23356 11108
rect 23396 11068 23397 11108
rect 23355 11059 23397 11068
rect 24250 11108 24308 11109
rect 24250 11068 24259 11108
rect 24299 11068 24308 11108
rect 24250 11067 24308 11068
rect 29828 11043 29870 11052
rect 843 11024 885 11033
rect 843 10984 844 11024
rect 884 10984 885 11024
rect 843 10975 885 10984
rect 1035 11024 1077 11033
rect 1035 10984 1036 11024
rect 1076 10984 1077 11024
rect 1035 10975 1077 10984
rect 1402 11024 1460 11025
rect 1402 10984 1411 11024
rect 1451 10984 1460 11024
rect 1402 10983 1460 10984
rect 1515 11024 1557 11033
rect 1515 10984 1516 11024
rect 1556 10984 1557 11024
rect 1515 10975 1557 10984
rect 2475 11024 2517 11033
rect 2475 10984 2476 11024
rect 2516 10984 2517 11024
rect 2475 10975 2517 10984
rect 2602 11024 2660 11025
rect 2602 10984 2611 11024
rect 2651 10984 2660 11024
rect 2602 10983 2660 10984
rect 3130 11024 3188 11025
rect 3130 10984 3139 11024
rect 3179 10984 3188 11024
rect 3130 10983 3188 10984
rect 3243 11024 3285 11033
rect 3243 10984 3244 11024
rect 3284 10984 3285 11024
rect 3243 10975 3285 10984
rect 3840 11024 3882 11033
rect 3840 10984 3841 11024
rect 3881 10984 3882 11024
rect 3840 10975 3882 10984
rect 4138 11024 4196 11025
rect 4138 10984 4147 11024
rect 4187 10984 4196 11024
rect 4138 10983 4196 10984
rect 4834 11024 4892 11025
rect 4834 10984 4843 11024
rect 4883 10984 4892 11024
rect 4834 10983 4892 10984
rect 5067 11024 5109 11033
rect 5067 10984 5068 11024
rect 5108 10984 5109 11024
rect 5067 10975 5109 10984
rect 5590 11024 5632 11033
rect 5590 10984 5591 11024
rect 5631 10984 5632 11024
rect 5590 10975 5632 10984
rect 5835 11024 5877 11033
rect 5835 10984 5836 11024
rect 5876 10984 5877 11024
rect 5835 10975 5877 10984
rect 6699 11024 6741 11033
rect 6699 10984 6700 11024
rect 6740 10984 6741 11024
rect 6699 10975 6741 10984
rect 6874 11024 6932 11025
rect 6874 10984 6883 11024
rect 6923 10984 6932 11024
rect 6874 10983 6932 10984
rect 7035 11024 7077 11033
rect 7035 10984 7036 11024
rect 7076 10984 7077 11024
rect 7035 10975 7077 10984
rect 7200 11024 7242 11033
rect 7200 10984 7201 11024
rect 7241 10984 7242 11024
rect 7200 10975 7242 10984
rect 7492 11024 7534 11033
rect 7492 10984 7493 11024
rect 7533 10984 7534 11024
rect 7492 10975 7534 10984
rect 7755 11024 7797 11033
rect 7755 10984 7756 11024
rect 7796 10984 7797 11024
rect 7755 10975 7797 10984
rect 7972 11024 8014 11033
rect 7972 10984 7973 11024
rect 8013 10984 8014 11024
rect 7972 10975 8014 10984
rect 8523 11024 8565 11033
rect 8523 10984 8524 11024
rect 8564 10984 8565 11024
rect 8523 10975 8565 10984
rect 8752 11024 8810 11025
rect 8752 10984 8761 11024
rect 8801 10984 8810 11024
rect 8752 10983 8810 10984
rect 9579 11024 9621 11033
rect 9579 10984 9580 11024
rect 9620 10984 9621 11024
rect 9579 10975 9621 10984
rect 9946 11024 10004 11025
rect 9946 10984 9955 11024
rect 9995 10984 10004 11024
rect 9946 10983 10004 10984
rect 10265 11024 10307 11033
rect 10265 10984 10266 11024
rect 10306 10984 10307 11024
rect 10265 10975 10307 10984
rect 10443 11024 10485 11033
rect 10443 10984 10444 11024
rect 10484 10984 10485 11024
rect 10443 10975 10485 10984
rect 10582 11024 10624 11033
rect 10582 10984 10583 11024
rect 10623 10984 10624 11024
rect 10582 10975 10624 10984
rect 11403 11024 11445 11033
rect 11632 11024 11690 11025
rect 11403 10984 11404 11024
rect 11444 10984 11445 11024
rect 11403 10975 11445 10984
rect 11538 11015 11584 11024
rect 11538 10975 11539 11015
rect 11579 10975 11584 11015
rect 11632 10984 11641 11024
rect 11681 10984 11690 11024
rect 11632 10983 11690 10984
rect 11787 11024 11829 11033
rect 11787 10984 11788 11024
rect 11828 10984 11829 11024
rect 11787 10975 11829 10984
rect 11979 11024 12021 11033
rect 11979 10984 11980 11024
rect 12020 10984 12021 11024
rect 11979 10975 12021 10984
rect 12202 11024 12260 11025
rect 12202 10984 12211 11024
rect 12251 10984 12260 11024
rect 12202 10983 12260 10984
rect 12922 11024 12980 11025
rect 12922 10984 12931 11024
rect 12971 10984 12980 11024
rect 12922 10983 12980 10984
rect 13035 11024 13077 11033
rect 13035 10984 13036 11024
rect 13076 10984 13077 11024
rect 13035 10975 13077 10984
rect 13504 11024 13546 11033
rect 13504 10984 13505 11024
rect 13545 10984 13546 11024
rect 13504 10975 13546 10984
rect 13707 11024 13749 11033
rect 13942 11024 13984 11033
rect 13707 10984 13708 11024
rect 13748 10984 13749 11024
rect 13707 10975 13749 10984
rect 13803 11015 13845 11024
rect 13803 10975 13804 11015
rect 13844 10975 13845 11015
rect 13942 10984 13943 11024
rect 13983 10984 13984 11024
rect 13942 10975 13984 10984
rect 14187 11024 14229 11033
rect 14187 10984 14188 11024
rect 14228 10984 14229 11024
rect 14187 10975 14229 10984
rect 14475 11024 14517 11033
rect 14475 10984 14476 11024
rect 14516 10984 14517 11024
rect 14475 10975 14517 10984
rect 14667 11024 14709 11033
rect 14667 10984 14668 11024
rect 14708 10984 14709 11024
rect 14667 10975 14709 10984
rect 14859 11024 14901 11033
rect 14859 10984 14860 11024
rect 14900 10984 14901 11024
rect 14859 10975 14901 10984
rect 15034 11024 15092 11025
rect 15034 10984 15043 11024
rect 15083 10984 15092 11024
rect 15034 10983 15092 10984
rect 15226 11024 15284 11025
rect 15226 10984 15235 11024
rect 15275 10984 15284 11024
rect 15226 10983 15284 10984
rect 15542 11024 15584 11033
rect 15542 10984 15543 11024
rect 15583 10984 15584 11024
rect 15542 10975 15584 10984
rect 15723 11024 15765 11033
rect 15723 10984 15724 11024
rect 15764 10984 15765 11024
rect 15723 10975 15765 10984
rect 15915 11024 15957 11033
rect 15915 10984 15916 11024
rect 15956 10984 15957 11024
rect 15915 10975 15957 10984
rect 16762 11024 16820 11025
rect 16762 10984 16771 11024
rect 16811 10984 16820 11024
rect 16762 10983 16820 10984
rect 16875 11024 16917 11033
rect 16875 10984 16876 11024
rect 16916 10984 16917 11024
rect 16875 10975 16917 10984
rect 17451 11024 17493 11033
rect 17451 10984 17452 11024
rect 17492 10984 17493 11024
rect 17451 10975 17493 10984
rect 17722 11024 17780 11025
rect 17722 10984 17731 11024
rect 17771 10984 17780 11024
rect 17722 10983 17780 10984
rect 18301 11024 18343 11033
rect 18970 11024 19028 11025
rect 18301 10984 18302 11024
rect 18342 10984 18343 11024
rect 18301 10975 18343 10984
rect 18603 11015 18645 11024
rect 18603 10975 18604 11015
rect 18644 10975 18645 11015
rect 18970 10984 18979 11024
rect 19019 10984 19028 11024
rect 18970 10983 19028 10984
rect 19947 11024 19989 11033
rect 19947 10984 19948 11024
rect 19988 10984 19989 11024
rect 19947 10975 19989 10984
rect 20715 11024 20757 11033
rect 20715 10984 20716 11024
rect 20756 10984 20757 11024
rect 20715 10975 20757 10984
rect 21195 11024 21237 11033
rect 21195 10984 21196 11024
rect 21236 10984 21237 11024
rect 21195 10975 21237 10984
rect 21579 11024 21621 11033
rect 22435 11024 22493 11025
rect 21579 10984 21580 11024
rect 21620 10984 21621 11024
rect 21579 10975 21621 10984
rect 22338 11015 22384 11024
rect 22338 10975 22339 11015
rect 22379 10975 22384 11015
rect 22435 10984 22444 11024
rect 22484 10984 22493 11024
rect 22435 10983 22493 10984
rect 22827 11024 22869 11033
rect 22827 10984 22828 11024
rect 22868 10984 22869 11024
rect 22827 10975 22869 10984
rect 22946 11024 22988 11033
rect 22946 10984 22947 11024
rect 22987 10984 22988 11024
rect 22946 10975 22988 10984
rect 23067 11024 23109 11033
rect 23638 11024 23680 11033
rect 23067 10984 23068 11024
rect 23108 10984 23109 11024
rect 23067 10975 23109 10984
rect 23202 11015 23248 11024
rect 23202 10975 23203 11015
rect 23243 10975 23248 11015
rect 23638 10984 23639 11024
rect 23679 10984 23680 11024
rect 23638 10975 23680 10984
rect 23883 11024 23925 11033
rect 23883 10984 23884 11024
rect 23924 10984 23925 11024
rect 23883 10975 23925 10984
rect 24160 11024 24202 11033
rect 24637 11024 24679 11033
rect 24160 10984 24161 11024
rect 24201 10984 24202 11024
rect 24160 10975 24202 10984
rect 24459 11015 24501 11024
rect 24459 10975 24460 11015
rect 24500 10975 24501 11015
rect 24637 10984 24638 11024
rect 24678 10984 24679 11024
rect 24637 10975 24679 10984
rect 24747 11024 24789 11033
rect 24747 10984 24748 11024
rect 24788 10984 24789 11024
rect 24747 10975 24789 10984
rect 25090 11024 25148 11025
rect 25090 10984 25099 11024
rect 25139 10984 25148 11024
rect 25090 10983 25148 10984
rect 25323 11024 25365 11033
rect 25323 10984 25324 11024
rect 25364 10984 25365 11024
rect 24936 10982 24994 10983
rect 11538 10966 11584 10975
rect 13803 10966 13845 10975
rect 18603 10966 18645 10975
rect 22338 10966 22384 10975
rect 23202 10966 23248 10975
rect 24459 10966 24501 10975
rect 4011 10940 4053 10949
rect 4011 10900 4012 10940
rect 4052 10900 4053 10940
rect 4011 10891 4053 10900
rect 4954 10940 5012 10941
rect 4954 10900 4963 10940
rect 5003 10900 5012 10940
rect 4954 10899 5012 10900
rect 5722 10940 5780 10941
rect 5722 10900 5731 10940
rect 5771 10900 5780 10940
rect 5722 10899 5780 10900
rect 7371 10940 7413 10949
rect 7371 10900 7372 10940
rect 7412 10900 7413 10940
rect 7371 10891 7413 10900
rect 7874 10940 7916 10949
rect 7874 10900 7875 10940
rect 7915 10900 7916 10940
rect 7874 10891 7916 10900
rect 8642 10940 8684 10949
rect 8642 10900 8643 10940
rect 8683 10900 8684 10940
rect 8642 10891 8684 10900
rect 14074 10940 14132 10941
rect 14074 10900 14083 10940
rect 14123 10900 14132 10940
rect 14074 10899 14132 10900
rect 22731 10940 22773 10949
rect 22731 10900 22732 10940
rect 22772 10900 22773 10940
rect 22731 10891 22773 10900
rect 23770 10940 23828 10941
rect 23770 10900 23779 10940
rect 23819 10900 23828 10940
rect 23770 10899 23828 10900
rect 23979 10940 24021 10949
rect 24936 10942 24945 10982
rect 24985 10942 24994 10982
rect 25323 10975 25365 10984
rect 25611 11024 25653 11033
rect 25611 10984 25612 11024
rect 25652 10984 25653 11024
rect 25611 10975 25653 10984
rect 25899 11024 25941 11033
rect 25899 10984 25900 11024
rect 25940 10984 25941 11024
rect 25899 10975 25941 10984
rect 26266 11024 26324 11025
rect 26266 10984 26275 11024
rect 26315 10984 26324 11024
rect 26266 10983 26324 10984
rect 26379 11024 26421 11033
rect 26379 10984 26380 11024
rect 26420 10984 26421 11024
rect 26379 10975 26421 10984
rect 27435 11024 27477 11033
rect 27435 10984 27436 11024
rect 27476 10984 27477 11024
rect 27435 10975 27477 10984
rect 28587 11024 28629 11033
rect 28587 10984 28588 11024
rect 28628 10984 28629 11024
rect 28587 10975 28629 10984
rect 29259 11024 29301 11033
rect 29259 10984 29260 11024
rect 29300 10984 29301 11024
rect 29259 10975 29301 10984
rect 29434 11024 29492 11025
rect 29434 10984 29443 11024
rect 29483 10984 29492 11024
rect 29434 10983 29492 10984
rect 29643 11024 29685 11033
rect 29643 10984 29644 11024
rect 29684 10984 29685 11024
rect 29828 11003 29829 11043
rect 29869 11003 29870 11043
rect 29828 10994 29870 11003
rect 30219 11024 30261 11033
rect 29643 10975 29685 10984
rect 30027 10982 30069 10991
rect 24936 10941 24994 10942
rect 23979 10900 23980 10940
rect 24020 10900 24021 10940
rect 23979 10891 24021 10900
rect 25210 10940 25268 10941
rect 25210 10900 25219 10940
rect 25259 10900 25268 10940
rect 25210 10899 25268 10900
rect 27345 10940 27387 10949
rect 27345 10900 27346 10940
rect 27386 10900 27387 10940
rect 30027 10942 30028 10982
rect 30068 10942 30069 10982
rect 30219 10984 30220 11024
rect 30260 10984 30261 11024
rect 30219 10975 30261 10984
rect 30027 10933 30069 10942
rect 27345 10891 27387 10900
rect 3915 10856 3957 10865
rect 3915 10816 3916 10856
rect 3956 10816 3957 10856
rect 3915 10807 3957 10816
rect 7275 10856 7317 10865
rect 7275 10816 7276 10856
rect 7316 10816 7317 10856
rect 7275 10807 7317 10816
rect 9771 10856 9813 10865
rect 9771 10816 9772 10856
rect 9812 10816 9813 10856
rect 9771 10807 9813 10816
rect 15034 10856 15092 10857
rect 15034 10816 15043 10856
rect 15083 10816 15092 10856
rect 15034 10815 15092 10816
rect 18123 10856 18165 10865
rect 18123 10816 18124 10856
rect 18164 10816 18165 10856
rect 18123 10807 18165 10816
rect 19023 10856 19065 10865
rect 19023 10816 19024 10856
rect 19064 10816 19065 10856
rect 19023 10807 19065 10816
rect 22042 10856 22100 10857
rect 22042 10816 22051 10856
rect 22091 10816 22100 10856
rect 22042 10815 22100 10816
rect 24843 10856 24885 10865
rect 24843 10816 24844 10856
rect 24884 10816 24885 10856
rect 24843 10807 24885 10816
rect 28875 10856 28917 10865
rect 28875 10816 28876 10856
rect 28916 10816 28917 10856
rect 28875 10807 28917 10816
rect 30411 10856 30453 10865
rect 30411 10816 30412 10856
rect 30452 10816 30453 10856
rect 30411 10807 30453 10816
rect 30795 10856 30837 10865
rect 30795 10816 30796 10856
rect 30836 10816 30837 10856
rect 30795 10807 30837 10816
rect 3418 10772 3476 10773
rect 3418 10732 3427 10772
rect 3467 10732 3476 10772
rect 3418 10731 3476 10732
rect 6874 10772 6932 10773
rect 6874 10732 6883 10772
rect 6923 10732 6932 10772
rect 6874 10731 6932 10732
rect 10251 10772 10293 10781
rect 10251 10732 10252 10772
rect 10292 10732 10293 10772
rect 10251 10723 10293 10732
rect 12315 10772 12357 10781
rect 12315 10732 12316 10772
rect 12356 10732 12357 10772
rect 12315 10723 12357 10732
rect 15531 10772 15573 10781
rect 15531 10732 15532 10772
rect 15572 10732 15573 10772
rect 15531 10723 15573 10732
rect 16971 10772 17013 10781
rect 16971 10732 16972 10772
rect 17012 10732 17013 10772
rect 16971 10723 17013 10732
rect 19546 10772 19604 10773
rect 19546 10732 19555 10772
rect 19595 10732 19604 10772
rect 19546 10731 19604 10732
rect 20314 10772 20372 10773
rect 20314 10732 20323 10772
rect 20363 10732 20372 10772
rect 20314 10731 20372 10732
rect 25611 10772 25653 10781
rect 25611 10732 25612 10772
rect 25652 10732 25653 10772
rect 25611 10723 25653 10732
rect 28186 10772 28244 10773
rect 28186 10732 28195 10772
rect 28235 10732 28244 10772
rect 28186 10731 28244 10732
rect 576 10604 31392 10628
rect 576 10564 3112 10604
rect 3480 10564 10886 10604
rect 11254 10564 18660 10604
rect 19028 10564 26434 10604
rect 26802 10564 31392 10604
rect 576 10540 31392 10564
rect 1659 10436 1701 10445
rect 1659 10396 1660 10436
rect 1700 10396 1701 10436
rect 1659 10387 1701 10396
rect 3339 10436 3381 10445
rect 3339 10396 3340 10436
rect 3380 10396 3381 10436
rect 3339 10387 3381 10396
rect 5242 10436 5300 10437
rect 5242 10396 5251 10436
rect 5291 10396 5300 10436
rect 5242 10395 5300 10396
rect 6411 10436 6453 10445
rect 6411 10396 6412 10436
rect 6452 10396 6453 10436
rect 6411 10387 6453 10396
rect 9051 10436 9093 10445
rect 9051 10396 9052 10436
rect 9092 10396 9093 10436
rect 9051 10387 9093 10396
rect 9483 10436 9525 10445
rect 9483 10396 9484 10436
rect 9524 10396 9525 10436
rect 9483 10387 9525 10396
rect 10138 10436 10196 10437
rect 10138 10396 10147 10436
rect 10187 10396 10196 10436
rect 10138 10395 10196 10396
rect 11403 10436 11445 10445
rect 11403 10396 11404 10436
rect 11444 10396 11445 10436
rect 11403 10387 11445 10396
rect 13306 10436 13364 10437
rect 13306 10396 13315 10436
rect 13355 10396 13364 10436
rect 13306 10395 13364 10396
rect 14907 10436 14949 10445
rect 14907 10396 14908 10436
rect 14948 10396 14949 10436
rect 14907 10387 14949 10396
rect 16635 10436 16677 10445
rect 16635 10396 16636 10436
rect 16676 10396 16677 10436
rect 16635 10387 16677 10396
rect 17242 10436 17300 10437
rect 17242 10396 17251 10436
rect 17291 10396 17300 10436
rect 17242 10395 17300 10396
rect 20667 10436 20709 10445
rect 20667 10396 20668 10436
rect 20708 10396 20709 10436
rect 20667 10387 20709 10396
rect 22042 10436 22100 10437
rect 22042 10396 22051 10436
rect 22091 10396 22100 10436
rect 22042 10395 22100 10396
rect 23979 10436 24021 10445
rect 23979 10396 23980 10436
rect 24020 10396 24021 10436
rect 23979 10387 24021 10396
rect 25035 10436 25077 10445
rect 25035 10396 25036 10436
rect 25076 10396 25077 10436
rect 25035 10387 25077 10396
rect 27802 10436 27860 10437
rect 27802 10396 27811 10436
rect 27851 10396 27860 10436
rect 27802 10395 27860 10396
rect 2266 10352 2324 10353
rect 2266 10312 2275 10352
rect 2315 10312 2324 10352
rect 19354 10352 19412 10353
rect 2266 10311 2324 10312
rect 9915 10326 9957 10335
rect 9915 10286 9916 10326
rect 9956 10286 9957 10326
rect 19354 10312 19363 10352
rect 19403 10312 19412 10352
rect 19354 10311 19412 10312
rect 23146 10352 23204 10353
rect 23146 10312 23155 10352
rect 23195 10312 23204 10352
rect 23146 10311 23204 10312
rect 28491 10352 28533 10361
rect 28491 10312 28492 10352
rect 28532 10312 28533 10352
rect 28491 10303 28533 10312
rect 30411 10352 30453 10361
rect 30411 10312 30412 10352
rect 30452 10312 30453 10352
rect 30411 10303 30453 10312
rect 30795 10352 30837 10361
rect 30795 10312 30796 10352
rect 30836 10312 30837 10352
rect 30795 10303 30837 10312
rect 9915 10277 9957 10286
rect 2650 10268 2708 10269
rect 2650 10228 2659 10268
rect 2699 10228 2708 10268
rect 2650 10227 2708 10228
rect 3610 10268 3668 10269
rect 3610 10228 3619 10268
rect 3659 10228 3668 10268
rect 3610 10227 3668 10228
rect 3819 10268 3861 10277
rect 3819 10228 3820 10268
rect 3860 10228 3861 10268
rect 3819 10219 3861 10228
rect 7162 10268 7220 10269
rect 7162 10228 7171 10268
rect 7211 10228 7220 10268
rect 7162 10227 7220 10228
rect 11505 10268 11547 10277
rect 11505 10228 11506 10268
rect 11546 10228 11547 10268
rect 11505 10219 11547 10228
rect 12010 10268 12068 10269
rect 12010 10228 12019 10268
rect 12059 10228 12068 10268
rect 12010 10227 12068 10228
rect 17547 10268 17589 10277
rect 17547 10228 17548 10268
rect 17588 10228 17589 10268
rect 17547 10219 17589 10228
rect 17762 10268 17804 10277
rect 17762 10228 17763 10268
rect 17803 10228 17804 10268
rect 17762 10219 17804 10228
rect 18027 10268 18069 10277
rect 18027 10228 18028 10268
rect 18068 10228 18069 10268
rect 22731 10268 22773 10277
rect 23643 10268 23685 10277
rect 18027 10219 18069 10228
rect 19995 10226 20037 10235
rect 651 10184 693 10193
rect 651 10144 652 10184
rect 692 10144 693 10184
rect 651 10135 693 10144
rect 843 10184 885 10193
rect 843 10144 844 10184
rect 884 10144 885 10184
rect 843 10135 885 10144
rect 1035 10184 1077 10193
rect 1035 10144 1036 10184
rect 1076 10144 1077 10184
rect 1035 10135 1077 10144
rect 1419 10184 1461 10193
rect 1419 10144 1420 10184
rect 1460 10144 1461 10184
rect 1419 10135 1461 10144
rect 1978 10184 2036 10185
rect 1978 10144 1987 10184
rect 2027 10144 2036 10184
rect 1978 10143 2036 10144
rect 2091 10184 2133 10193
rect 2091 10144 2092 10184
rect 2132 10144 2133 10184
rect 2091 10135 2133 10144
rect 2523 10184 2565 10193
rect 2523 10144 2524 10184
rect 2564 10144 2565 10184
rect 2523 10135 2565 10144
rect 2763 10184 2805 10193
rect 2763 10144 2764 10184
rect 2804 10144 2805 10184
rect 2763 10135 2805 10144
rect 3034 10184 3092 10185
rect 3034 10144 3043 10184
rect 3083 10144 3092 10184
rect 3034 10143 3092 10144
rect 3147 10184 3189 10193
rect 3147 10144 3148 10184
rect 3188 10144 3189 10184
rect 3147 10135 3189 10144
rect 3490 10184 3548 10185
rect 3490 10144 3499 10184
rect 3539 10144 3548 10184
rect 3490 10143 3548 10144
rect 3723 10184 3765 10193
rect 3723 10144 3724 10184
rect 3764 10144 3765 10184
rect 3723 10135 3765 10144
rect 4011 10184 4053 10193
rect 4011 10144 4012 10184
rect 4052 10144 4053 10184
rect 4011 10135 4053 10144
rect 4395 10184 4437 10193
rect 4395 10144 4396 10184
rect 4436 10144 4437 10184
rect 4395 10135 4437 10144
rect 4954 10184 5012 10185
rect 4954 10144 4963 10184
rect 5003 10144 5012 10184
rect 4954 10143 5012 10144
rect 5067 10184 5109 10193
rect 5067 10144 5068 10184
rect 5108 10144 5109 10184
rect 5067 10135 5109 10144
rect 5547 10184 5589 10193
rect 5547 10144 5548 10184
rect 5588 10144 5589 10184
rect 5547 10135 5589 10144
rect 5835 10184 5877 10193
rect 5835 10144 5836 10184
rect 5876 10144 5877 10184
rect 5835 10135 5877 10144
rect 6459 10184 6501 10193
rect 6459 10144 6460 10184
rect 6500 10144 6501 10184
rect 6459 10135 6501 10144
rect 6603 10184 6645 10193
rect 6603 10144 6604 10184
rect 6644 10144 6645 10184
rect 6603 10135 6645 10144
rect 7030 10184 7072 10193
rect 7030 10144 7031 10184
rect 7071 10144 7072 10184
rect 7030 10135 7072 10144
rect 7275 10184 7317 10193
rect 7275 10144 7276 10184
rect 7316 10144 7317 10184
rect 7275 10135 7317 10144
rect 7947 10184 7989 10193
rect 7947 10144 7948 10184
rect 7988 10144 7989 10184
rect 7947 10135 7989 10144
rect 8427 10184 8469 10193
rect 8427 10144 8428 10184
rect 8468 10144 8469 10184
rect 8427 10135 8469 10144
rect 8811 10184 8853 10193
rect 8811 10144 8812 10184
rect 8852 10144 8853 10184
rect 8811 10135 8853 10144
rect 9178 10184 9236 10185
rect 9178 10144 9187 10184
rect 9227 10144 9236 10184
rect 9178 10143 9236 10144
rect 9291 10184 9333 10193
rect 9291 10144 9292 10184
rect 9332 10144 9333 10184
rect 9291 10135 9333 10144
rect 9494 10184 9536 10193
rect 9494 10144 9495 10184
rect 9535 10144 9536 10184
rect 9494 10135 9536 10144
rect 9946 10184 10004 10185
rect 9946 10144 9955 10184
rect 9995 10144 10004 10184
rect 9946 10143 10004 10144
rect 10615 10184 10673 10185
rect 10615 10144 10624 10184
rect 10664 10144 10673 10184
rect 10615 10143 10673 10144
rect 11595 10184 11637 10193
rect 11595 10144 11596 10184
rect 11636 10144 11637 10184
rect 11595 10135 11637 10144
rect 12363 10184 12405 10193
rect 12363 10144 12364 10184
rect 12404 10144 12405 10184
rect 12363 10135 12405 10144
rect 12651 10184 12693 10193
rect 12651 10144 12652 10184
rect 12692 10144 12693 10184
rect 12651 10135 12693 10144
rect 13018 10184 13076 10185
rect 13018 10144 13027 10184
rect 13067 10144 13076 10184
rect 13018 10143 13076 10144
rect 13131 10184 13173 10193
rect 13131 10144 13132 10184
rect 13172 10144 13173 10184
rect 13131 10135 13173 10144
rect 13687 10184 13745 10185
rect 13687 10144 13696 10184
rect 13736 10144 13745 10184
rect 13687 10143 13745 10144
rect 14475 10184 14517 10193
rect 14475 10144 14476 10184
rect 14516 10144 14517 10184
rect 14475 10135 14517 10144
rect 14763 10184 14805 10193
rect 14763 10144 14764 10184
rect 14804 10144 14805 10184
rect 14763 10135 14805 10144
rect 15147 10184 15189 10193
rect 15147 10144 15148 10184
rect 15188 10144 15189 10184
rect 15147 10135 15189 10144
rect 15531 10184 15573 10193
rect 15531 10144 15532 10184
rect 15572 10144 15573 10184
rect 15531 10135 15573 10144
rect 16011 10184 16053 10193
rect 16011 10144 16012 10184
rect 16052 10144 16053 10184
rect 16011 10135 16053 10144
rect 16395 10184 16437 10193
rect 16395 10144 16396 10184
rect 16436 10144 16437 10184
rect 16395 10135 16437 10144
rect 16954 10184 17012 10185
rect 16954 10144 16963 10184
rect 17003 10144 17012 10184
rect 16954 10143 17012 10144
rect 17067 10184 17109 10193
rect 17067 10144 17068 10184
rect 17108 10144 17109 10184
rect 17067 10135 17109 10144
rect 17643 10184 17685 10193
rect 17643 10144 17644 10184
rect 17684 10144 17685 10184
rect 17643 10135 17685 10144
rect 17860 10184 17902 10193
rect 17860 10144 17861 10184
rect 17901 10144 17902 10184
rect 17860 10135 17902 10144
rect 18123 10184 18165 10193
rect 18123 10144 18124 10184
rect 18164 10144 18165 10184
rect 18123 10135 18165 10144
rect 18242 10184 18284 10193
rect 18242 10144 18243 10184
rect 18283 10144 18284 10184
rect 18242 10135 18284 10144
rect 18352 10184 18410 10185
rect 18352 10144 18361 10184
rect 18401 10144 18410 10184
rect 18352 10143 18410 10144
rect 19179 10184 19221 10193
rect 19179 10144 19180 10184
rect 19220 10144 19221 10184
rect 19179 10135 19221 10144
rect 19354 10184 19412 10185
rect 19354 10144 19363 10184
rect 19403 10144 19412 10184
rect 19354 10143 19412 10144
rect 19755 10184 19797 10193
rect 19755 10144 19756 10184
rect 19796 10144 19797 10184
rect 19755 10135 19797 10144
rect 19874 10184 19916 10193
rect 19874 10144 19875 10184
rect 19915 10144 19916 10184
rect 19995 10186 19996 10226
rect 20036 10186 20037 10226
rect 22731 10228 22732 10268
rect 22772 10228 22773 10268
rect 22731 10219 22773 10228
rect 22962 10259 23008 10268
rect 22962 10219 22963 10259
rect 23003 10219 23008 10259
rect 23643 10228 23644 10268
rect 23684 10228 23685 10268
rect 23643 10219 23685 10228
rect 25137 10268 25179 10277
rect 25137 10228 25138 10268
rect 25178 10228 25179 10268
rect 25137 10219 25179 10228
rect 26001 10268 26043 10277
rect 26001 10228 26002 10268
rect 26042 10228 26043 10268
rect 26001 10219 26043 10228
rect 22962 10210 23008 10219
rect 19995 10177 20037 10186
rect 21003 10184 21045 10193
rect 19874 10135 19916 10144
rect 21003 10144 21004 10184
rect 21044 10144 21045 10184
rect 21003 10135 21045 10144
rect 21291 10184 21333 10193
rect 21291 10144 21292 10184
rect 21332 10144 21333 10184
rect 21291 10135 21333 10144
rect 21579 10184 21621 10193
rect 21579 10144 21580 10184
rect 21620 10144 21621 10184
rect 21579 10135 21621 10144
rect 22443 10184 22485 10193
rect 22443 10144 22444 10184
rect 22484 10144 22485 10184
rect 22443 10135 22485 10144
rect 22827 10184 22869 10193
rect 22827 10144 22828 10184
rect 22868 10144 22869 10184
rect 22827 10135 22869 10144
rect 23056 10184 23114 10185
rect 23056 10144 23065 10184
rect 23105 10144 23114 10184
rect 23056 10143 23114 10144
rect 23355 10184 23397 10193
rect 23355 10144 23356 10184
rect 23396 10144 23397 10184
rect 23355 10135 23397 10144
rect 23499 10184 23541 10193
rect 23499 10144 23500 10184
rect 23540 10144 23541 10184
rect 23499 10135 23541 10144
rect 23787 10184 23829 10193
rect 23787 10144 23788 10184
rect 23828 10144 23829 10184
rect 23787 10135 23829 10144
rect 24132 10184 24190 10185
rect 24132 10144 24141 10184
rect 24181 10144 24190 10184
rect 24132 10143 24190 10144
rect 24235 10184 24293 10185
rect 24235 10144 24244 10184
rect 24284 10144 24293 10184
rect 24235 10143 24293 10144
rect 24359 10184 24417 10185
rect 24359 10144 24368 10184
rect 24408 10144 24417 10184
rect 24359 10143 24417 10144
rect 25227 10184 25269 10193
rect 25227 10144 25228 10184
rect 25268 10144 25269 10184
rect 25227 10135 25269 10144
rect 26091 10184 26133 10193
rect 26091 10144 26092 10184
rect 26132 10144 26133 10184
rect 26091 10135 26133 10144
rect 26859 10184 26901 10193
rect 26859 10144 26860 10184
rect 26900 10144 26901 10184
rect 26859 10135 26901 10144
rect 27147 10184 27189 10193
rect 27147 10144 27148 10184
rect 27188 10144 27189 10184
rect 27147 10135 27189 10144
rect 27322 10184 27380 10185
rect 27322 10144 27331 10184
rect 27371 10144 27380 10184
rect 27322 10143 27380 10144
rect 27627 10184 27669 10193
rect 27627 10144 27628 10184
rect 27668 10144 27669 10184
rect 27627 10135 27669 10144
rect 28011 10184 28053 10193
rect 28011 10144 28012 10184
rect 28052 10144 28053 10184
rect 28011 10135 28053 10144
rect 28099 10184 28157 10185
rect 28099 10144 28108 10184
rect 28148 10144 28157 10184
rect 28099 10143 28157 10144
rect 29355 10184 29397 10193
rect 29355 10144 29356 10184
rect 29396 10144 29397 10184
rect 29355 10135 29397 10144
rect 2842 10100 2900 10101
rect 2842 10060 2851 10100
rect 2891 10060 2900 10100
rect 2842 10059 2900 10060
rect 3353 10100 3395 10109
rect 3353 10060 3354 10100
rect 3394 10060 3395 10100
rect 3353 10051 3395 10060
rect 6171 10100 6213 10109
rect 6171 10060 6172 10100
rect 6212 10060 6213 10100
rect 6171 10051 6213 10060
rect 19659 10100 19701 10109
rect 19659 10060 19660 10100
rect 19700 10060 19701 10100
rect 19659 10051 19701 10060
rect 22234 10100 22292 10101
rect 22234 10060 22243 10100
rect 22283 10060 22292 10100
rect 22234 10059 22292 10060
rect 27531 10100 27573 10109
rect 27531 10060 27532 10100
rect 27572 10060 27573 10100
rect 27531 10051 27573 10060
rect 27805 10100 27847 10109
rect 27805 10060 27806 10100
rect 27846 10060 27847 10100
rect 27805 10051 27847 10060
rect 826 10016 884 10017
rect 826 9976 835 10016
rect 875 9976 884 10016
rect 826 9975 884 9976
rect 4491 10016 4533 10025
rect 4491 9976 4492 10016
rect 4532 9976 4533 10016
rect 4491 9967 4533 9976
rect 7354 10016 7412 10017
rect 7354 9976 7363 10016
rect 7403 9976 7412 10016
rect 7354 9975 7412 9976
rect 7834 10016 7892 10017
rect 7834 9976 7843 10016
rect 7883 9976 7892 10016
rect 7834 9975 7892 9976
rect 8139 10016 8181 10025
rect 8139 9976 8140 10016
rect 8180 9976 8181 10016
rect 8139 9967 8181 9976
rect 10779 10016 10821 10025
rect 10779 9976 10780 10016
rect 10820 9976 10821 10016
rect 10779 9967 10821 9976
rect 13851 10016 13893 10025
rect 13851 9976 13852 10016
rect 13892 9976 13893 10016
rect 13851 9967 13893 9976
rect 14266 10016 14324 10017
rect 14266 9976 14275 10016
rect 14315 9976 14324 10016
rect 14266 9975 14324 9976
rect 21675 10016 21717 10025
rect 21675 9976 21676 10016
rect 21716 9976 21717 10016
rect 21675 9967 21717 9976
rect 25786 10016 25844 10017
rect 25786 9976 25795 10016
rect 25835 9976 25844 10016
rect 25786 9975 25844 9976
rect 26650 10016 26708 10017
rect 26650 9976 26659 10016
rect 26699 9976 26708 10016
rect 26650 9975 26708 9976
rect 28011 10016 28053 10025
rect 28011 9976 28012 10016
rect 28052 9976 28053 10016
rect 28011 9967 28053 9976
rect 28683 10016 28725 10025
rect 28683 9976 28684 10016
rect 28724 9976 28725 10016
rect 28683 9967 28725 9976
rect 576 9848 31392 9872
rect 576 9808 4352 9848
rect 4720 9808 12126 9848
rect 12494 9808 19900 9848
rect 20268 9808 27674 9848
rect 28042 9808 31392 9848
rect 576 9784 31392 9808
rect 939 9680 981 9689
rect 939 9640 940 9680
rect 980 9640 981 9680
rect 939 9631 981 9640
rect 1803 9680 1845 9689
rect 1803 9640 1804 9680
rect 1844 9640 1845 9680
rect 1803 9631 1845 9640
rect 4203 9680 4245 9689
rect 4203 9640 4204 9680
rect 4244 9640 4245 9680
rect 4203 9631 4245 9640
rect 4762 9680 4820 9681
rect 4762 9640 4771 9680
rect 4811 9640 4820 9680
rect 4762 9639 4820 9640
rect 6970 9680 7028 9681
rect 6970 9640 6979 9680
rect 7019 9640 7028 9680
rect 6970 9639 7028 9640
rect 7659 9680 7701 9689
rect 7659 9640 7660 9680
rect 7700 9640 7701 9680
rect 7659 9631 7701 9640
rect 8523 9680 8565 9689
rect 8523 9640 8524 9680
rect 8564 9640 8565 9680
rect 8523 9631 8565 9640
rect 9195 9680 9237 9689
rect 9195 9640 9196 9680
rect 9236 9640 9237 9680
rect 9195 9631 9237 9640
rect 9754 9680 9812 9681
rect 9754 9640 9763 9680
rect 9803 9640 9812 9680
rect 9754 9639 9812 9640
rect 10443 9680 10485 9689
rect 10443 9640 10444 9680
rect 10484 9640 10485 9680
rect 10443 9631 10485 9640
rect 10906 9680 10964 9681
rect 10906 9640 10915 9680
rect 10955 9640 10964 9680
rect 10906 9639 10964 9640
rect 12267 9680 12309 9689
rect 12267 9640 12268 9680
rect 12308 9640 12309 9680
rect 12267 9631 12309 9640
rect 13690 9680 13748 9681
rect 13690 9640 13699 9680
rect 13739 9640 13748 9680
rect 13690 9639 13748 9640
rect 13995 9680 14037 9689
rect 13995 9640 13996 9680
rect 14036 9640 14037 9680
rect 13995 9631 14037 9640
rect 14667 9680 14709 9689
rect 14667 9640 14668 9680
rect 14708 9640 14709 9680
rect 14667 9631 14709 9640
rect 15147 9680 15189 9689
rect 15147 9640 15148 9680
rect 15188 9640 15189 9680
rect 15147 9631 15189 9640
rect 15802 9680 15860 9681
rect 15802 9640 15811 9680
rect 15851 9640 15860 9680
rect 15802 9639 15860 9640
rect 17643 9680 17685 9689
rect 17643 9640 17644 9680
rect 17684 9640 17685 9680
rect 17643 9631 17685 9640
rect 17818 9680 17876 9681
rect 17818 9640 17827 9680
rect 17867 9640 17876 9680
rect 17818 9639 17876 9640
rect 18682 9680 18740 9681
rect 18682 9640 18691 9680
rect 18731 9640 18740 9680
rect 18682 9639 18740 9640
rect 20218 9680 20276 9681
rect 20218 9640 20227 9680
rect 20267 9640 20276 9680
rect 20218 9639 20276 9640
rect 20890 9680 20948 9681
rect 20890 9640 20899 9680
rect 20939 9640 20948 9680
rect 20890 9639 20948 9640
rect 21658 9680 21716 9681
rect 21658 9640 21667 9680
rect 21707 9640 21716 9680
rect 21658 9639 21716 9640
rect 23019 9680 23061 9689
rect 23019 9640 23020 9680
rect 23060 9640 23061 9680
rect 23019 9631 23061 9640
rect 23403 9680 23445 9689
rect 23403 9640 23404 9680
rect 23444 9640 23445 9680
rect 23403 9631 23445 9640
rect 24267 9680 24309 9689
rect 24267 9640 24268 9680
rect 24308 9640 24309 9680
rect 24267 9631 24309 9640
rect 24442 9680 24500 9681
rect 24442 9640 24451 9680
rect 24491 9640 24500 9680
rect 24442 9639 24500 9640
rect 25834 9680 25892 9681
rect 25834 9640 25843 9680
rect 25883 9640 25892 9680
rect 25834 9639 25892 9640
rect 27435 9680 27477 9689
rect 27435 9640 27436 9680
rect 27476 9640 27477 9680
rect 27435 9631 27477 9640
rect 2379 9596 2421 9605
rect 2379 9556 2380 9596
rect 2420 9556 2421 9596
rect 2379 9547 2421 9556
rect 6315 9596 6357 9605
rect 6315 9556 6316 9596
rect 6356 9556 6357 9596
rect 6315 9547 6357 9556
rect 13323 9596 13365 9605
rect 13323 9556 13324 9596
rect 13364 9556 13365 9596
rect 13323 9547 13365 9556
rect 15254 9596 15296 9605
rect 15254 9556 15255 9596
rect 15295 9556 15296 9596
rect 15254 9547 15296 9556
rect 15531 9596 15573 9605
rect 15531 9556 15532 9596
rect 15572 9556 15573 9596
rect 15531 9547 15573 9556
rect 25213 9596 25255 9605
rect 25213 9556 25214 9596
rect 25254 9556 25255 9596
rect 25213 9547 25255 9556
rect 25306 9596 25364 9597
rect 25306 9556 25315 9596
rect 25355 9556 25364 9596
rect 25306 9555 25364 9556
rect 26283 9596 26325 9605
rect 26283 9556 26284 9596
rect 26324 9556 26325 9596
rect 26283 9547 26325 9556
rect 26955 9596 26997 9605
rect 26955 9556 26956 9596
rect 26996 9556 26997 9596
rect 26955 9547 26997 9556
rect 939 9512 981 9521
rect 939 9472 940 9512
rect 980 9472 981 9512
rect 939 9463 981 9472
rect 1131 9512 1173 9521
rect 1131 9472 1132 9512
rect 1172 9472 1173 9512
rect 1131 9463 1173 9472
rect 1323 9512 1365 9521
rect 1323 9472 1324 9512
rect 1364 9472 1365 9512
rect 1323 9463 1365 9472
rect 1707 9512 1749 9521
rect 1707 9472 1708 9512
rect 1748 9472 1749 9512
rect 1707 9463 1749 9472
rect 2283 9512 2325 9521
rect 2283 9472 2284 9512
rect 2324 9472 2325 9512
rect 2283 9463 2325 9472
rect 2479 9512 2521 9521
rect 2479 9472 2480 9512
rect 2520 9472 2521 9512
rect 2479 9463 2521 9472
rect 2667 9512 2709 9521
rect 2667 9472 2668 9512
rect 2708 9472 2709 9512
rect 2667 9463 2709 9472
rect 2955 9512 2997 9521
rect 2955 9472 2956 9512
rect 2996 9472 2997 9512
rect 2955 9463 2997 9472
rect 3094 9512 3136 9521
rect 3094 9472 3095 9512
rect 3135 9472 3136 9512
rect 3094 9463 3136 9472
rect 3339 9512 3381 9521
rect 3339 9472 3340 9512
rect 3380 9472 3381 9512
rect 3339 9463 3381 9472
rect 3627 9512 3669 9521
rect 3627 9472 3628 9512
rect 3668 9472 3669 9512
rect 3627 9463 3669 9472
rect 3744 9512 3802 9513
rect 3744 9472 3753 9512
rect 3793 9472 3802 9512
rect 3744 9471 3802 9472
rect 3915 9512 3957 9521
rect 3915 9472 3916 9512
rect 3956 9472 3957 9512
rect 3915 9463 3957 9472
rect 4107 9512 4149 9521
rect 4107 9472 4108 9512
rect 4148 9472 4149 9512
rect 4107 9463 4149 9472
rect 4299 9512 4341 9521
rect 4299 9472 4300 9512
rect 4340 9472 4341 9512
rect 4683 9512 4725 9521
rect 4299 9463 4341 9472
rect 4443 9470 4485 9479
rect 3220 9428 3262 9437
rect 3220 9388 3221 9428
rect 3261 9388 3262 9428
rect 3220 9379 3262 9388
rect 3435 9428 3477 9437
rect 3435 9388 3436 9428
rect 3476 9388 3477 9428
rect 4443 9430 4444 9470
rect 4484 9430 4485 9470
rect 4683 9472 4684 9512
rect 4724 9472 4725 9512
rect 4683 9463 4725 9472
rect 5110 9512 5152 9521
rect 5110 9472 5111 9512
rect 5151 9472 5152 9512
rect 5110 9463 5152 9472
rect 5355 9512 5397 9521
rect 5355 9472 5356 9512
rect 5396 9472 5397 9512
rect 5355 9463 5397 9472
rect 5643 9512 5685 9521
rect 5643 9472 5644 9512
rect 5684 9472 5685 9512
rect 5643 9463 5685 9472
rect 5818 9512 5876 9513
rect 5818 9472 5827 9512
rect 5867 9472 5876 9512
rect 5818 9471 5876 9472
rect 6219 9512 6261 9521
rect 6219 9472 6220 9512
rect 6260 9472 6261 9512
rect 6219 9463 6261 9472
rect 6411 9512 6453 9521
rect 6411 9472 6412 9512
rect 6452 9472 6453 9512
rect 6411 9463 6453 9472
rect 6795 9512 6837 9521
rect 6795 9472 6796 9512
rect 6836 9472 6837 9512
rect 6795 9463 6837 9472
rect 6987 9512 7029 9521
rect 6987 9472 6988 9512
rect 7028 9472 7029 9512
rect 6987 9463 7029 9472
rect 7210 9512 7268 9513
rect 7210 9472 7219 9512
rect 7259 9472 7268 9512
rect 7210 9471 7268 9472
rect 7467 9512 7509 9521
rect 7467 9472 7468 9512
rect 7508 9472 7509 9512
rect 7467 9463 7509 9472
rect 8122 9512 8180 9513
rect 8122 9472 8131 9512
rect 8171 9472 8180 9512
rect 8122 9471 8180 9472
rect 8235 9512 8277 9521
rect 8235 9472 8236 9512
rect 8276 9472 8277 9512
rect 8235 9463 8277 9472
rect 8715 9512 8757 9521
rect 8715 9472 8716 9512
rect 8756 9472 8757 9512
rect 8715 9463 8757 9472
rect 9099 9512 9141 9521
rect 9099 9472 9100 9512
rect 9140 9472 9141 9512
rect 9099 9463 9141 9472
rect 9430 9512 9472 9521
rect 9430 9472 9431 9512
rect 9471 9472 9472 9512
rect 9430 9463 9472 9472
rect 9562 9512 9620 9513
rect 9562 9472 9571 9512
rect 9611 9472 9620 9512
rect 9562 9471 9620 9472
rect 9675 9512 9717 9521
rect 9675 9472 9676 9512
rect 9716 9472 9717 9512
rect 9675 9463 9717 9472
rect 10285 9512 10343 9513
rect 10285 9472 10294 9512
rect 10334 9472 10343 9512
rect 10285 9471 10343 9472
rect 10539 9512 10581 9521
rect 10539 9472 10540 9512
rect 10580 9472 10581 9512
rect 10539 9463 10581 9472
rect 10658 9512 10700 9521
rect 10658 9472 10659 9512
rect 10699 9472 10700 9512
rect 10658 9463 10700 9472
rect 10768 9512 10826 9513
rect 10768 9472 10777 9512
rect 10817 9472 10826 9512
rect 10768 9471 10826 9472
rect 11211 9512 11253 9521
rect 11211 9472 11212 9512
rect 11252 9472 11253 9512
rect 11211 9463 11253 9472
rect 11979 9512 12021 9521
rect 11979 9472 11980 9512
rect 12020 9472 12021 9512
rect 11979 9463 12021 9472
rect 12118 9512 12160 9521
rect 12118 9472 12119 9512
rect 12159 9472 12160 9512
rect 12118 9463 12160 9472
rect 12406 9512 12448 9521
rect 12406 9472 12407 9512
rect 12447 9472 12448 9512
rect 12406 9463 12448 9472
rect 12651 9512 12693 9521
rect 12651 9472 12652 9512
rect 12692 9472 12693 9512
rect 12651 9463 12693 9472
rect 13227 9512 13269 9521
rect 13227 9472 13228 9512
rect 13268 9472 13269 9512
rect 13227 9463 13269 9472
rect 13419 9512 13461 9521
rect 13419 9472 13420 9512
rect 13460 9472 13461 9512
rect 13419 9463 13461 9472
rect 13803 9512 13845 9521
rect 13803 9472 13804 9512
rect 13844 9472 13845 9512
rect 13803 9463 13845 9472
rect 14187 9512 14229 9521
rect 14187 9472 14188 9512
rect 14228 9472 14229 9512
rect 14187 9463 14229 9472
rect 14571 9512 14613 9521
rect 14571 9472 14572 9512
rect 14612 9472 14613 9512
rect 14571 9463 14613 9472
rect 14938 9512 14996 9513
rect 14938 9472 14947 9512
rect 14987 9472 14996 9512
rect 14938 9471 14996 9472
rect 15051 9512 15093 9521
rect 15051 9472 15052 9512
rect 15092 9472 15093 9512
rect 15051 9463 15093 9472
rect 15435 9512 15477 9521
rect 15435 9472 15436 9512
rect 15476 9472 15477 9512
rect 15435 9463 15477 9472
rect 15627 9512 15669 9521
rect 15627 9472 15628 9512
rect 15668 9472 15669 9512
rect 15627 9463 15669 9472
rect 16107 9512 16149 9521
rect 16107 9472 16108 9512
rect 16148 9472 16149 9512
rect 16107 9463 16149 9472
rect 17242 9512 17300 9513
rect 17242 9472 17251 9512
rect 17291 9472 17300 9512
rect 17242 9471 17300 9472
rect 17355 9512 17397 9521
rect 17355 9472 17356 9512
rect 17396 9472 17397 9512
rect 17355 9463 17397 9472
rect 18012 9512 18054 9521
rect 18012 9472 18013 9512
rect 18053 9472 18054 9512
rect 18012 9463 18054 9472
rect 18123 9512 18165 9521
rect 18123 9472 18124 9512
rect 18164 9472 18165 9512
rect 18123 9463 18165 9472
rect 18795 9512 18837 9521
rect 18795 9472 18796 9512
rect 18836 9472 18837 9512
rect 18795 9463 18837 9472
rect 19179 9512 19221 9521
rect 19179 9472 19180 9512
rect 19220 9472 19221 9512
rect 19179 9463 19221 9472
rect 19371 9512 19413 9521
rect 19371 9472 19372 9512
rect 19412 9472 19413 9512
rect 19371 9463 19413 9472
rect 19659 9512 19701 9521
rect 19659 9472 19660 9512
rect 19700 9472 19701 9512
rect 19659 9463 19701 9472
rect 20506 9512 20564 9513
rect 20506 9472 20515 9512
rect 20555 9472 20564 9512
rect 20506 9471 20564 9472
rect 21084 9512 21126 9521
rect 21084 9472 21085 9512
rect 21125 9472 21126 9512
rect 21084 9463 21126 9472
rect 21195 9512 21237 9521
rect 21195 9472 21196 9512
rect 21236 9472 21237 9512
rect 21195 9463 21237 9472
rect 21963 9512 22005 9521
rect 21963 9472 21964 9512
rect 22004 9472 22005 9512
rect 21963 9463 22005 9472
rect 22618 9512 22676 9513
rect 22618 9472 22627 9512
rect 22667 9472 22676 9512
rect 22618 9471 22676 9472
rect 22731 9512 22773 9521
rect 22731 9472 22732 9512
rect 22772 9472 22773 9512
rect 22731 9463 22773 9472
rect 23194 9512 23252 9513
rect 23194 9472 23203 9512
rect 23243 9472 23252 9512
rect 23194 9471 23252 9472
rect 23499 9512 23541 9521
rect 23499 9472 23500 9512
rect 23540 9472 23541 9512
rect 23499 9463 23541 9472
rect 23866 9512 23924 9513
rect 23866 9472 23875 9512
rect 23915 9472 23924 9512
rect 23866 9471 23924 9472
rect 23979 9512 24021 9521
rect 23979 9472 23980 9512
rect 24020 9472 24021 9512
rect 23979 9463 24021 9472
rect 24603 9512 24645 9521
rect 24603 9472 24604 9512
rect 24644 9472 24645 9512
rect 24603 9463 24645 9472
rect 24747 9512 24789 9521
rect 24747 9472 24748 9512
rect 24788 9472 24789 9512
rect 24747 9463 24789 9472
rect 25419 9512 25461 9521
rect 25999 9512 26057 9513
rect 25419 9472 25420 9512
rect 25460 9472 25461 9512
rect 25419 9463 25461 9472
rect 25515 9503 25557 9512
rect 25515 9463 25516 9503
rect 25556 9463 25557 9503
rect 25999 9472 26008 9512
rect 26048 9472 26057 9512
rect 25999 9471 26057 9472
rect 26170 9512 26212 9521
rect 26170 9472 26171 9512
rect 26211 9472 26212 9512
rect 26170 9463 26212 9472
rect 26374 9512 26432 9513
rect 26374 9472 26383 9512
rect 26423 9472 26432 9512
rect 26374 9471 26432 9472
rect 26571 9512 26613 9521
rect 26571 9472 26572 9512
rect 26612 9472 26613 9512
rect 26571 9463 26613 9472
rect 26746 9512 26804 9513
rect 26746 9472 26755 9512
rect 26795 9472 26804 9512
rect 26746 9471 26804 9472
rect 27051 9512 27093 9521
rect 27051 9472 27052 9512
rect 27092 9472 27093 9512
rect 27051 9463 27093 9472
rect 27280 9512 27338 9513
rect 27280 9472 27289 9512
rect 27329 9472 27338 9512
rect 27280 9471 27338 9472
rect 29338 9512 29396 9513
rect 29338 9472 29347 9512
rect 29387 9472 29396 9512
rect 29338 9471 29396 9472
rect 25515 9454 25557 9463
rect 4443 9421 4485 9430
rect 4570 9428 4628 9429
rect 3435 9379 3477 9388
rect 4570 9388 4579 9428
rect 4619 9388 4628 9428
rect 4570 9387 4628 9388
rect 5242 9428 5300 9429
rect 5242 9388 5251 9428
rect 5291 9388 5300 9428
rect 5242 9387 5300 9388
rect 5451 9428 5493 9437
rect 5451 9388 5452 9428
rect 5492 9388 5493 9428
rect 5451 9379 5493 9388
rect 10090 9428 10148 9429
rect 10090 9388 10099 9428
rect 10139 9388 10148 9428
rect 10090 9387 10148 9388
rect 11121 9428 11163 9437
rect 11121 9388 11122 9428
rect 11162 9388 11163 9428
rect 11121 9379 11163 9388
rect 12532 9428 12574 9437
rect 12532 9388 12533 9428
rect 12573 9388 12574 9428
rect 12532 9379 12574 9388
rect 12747 9428 12789 9437
rect 12747 9388 12748 9428
rect 12788 9388 12789 9428
rect 12747 9379 12789 9388
rect 16017 9428 16059 9437
rect 16017 9388 16018 9428
rect 16058 9388 16059 9428
rect 16017 9379 16059 9388
rect 20122 9428 20180 9429
rect 20122 9388 20131 9428
rect 20171 9388 20180 9428
rect 20122 9387 20180 9388
rect 20698 9428 20756 9429
rect 20698 9388 20707 9428
rect 20747 9388 20756 9428
rect 20698 9387 20756 9388
rect 21873 9428 21915 9437
rect 29722 9428 29780 9429
rect 21873 9388 21874 9428
rect 21914 9388 21915 9428
rect 21873 9379 21915 9388
rect 27186 9419 27232 9428
rect 27186 9379 27187 9419
rect 27227 9379 27232 9419
rect 29722 9388 29731 9428
rect 29771 9388 29780 9428
rect 29722 9387 29780 9388
rect 27186 9370 27232 9379
rect 5871 9344 5913 9353
rect 5871 9304 5872 9344
rect 5912 9304 5913 9344
rect 5871 9295 5913 9304
rect 26746 9344 26804 9345
rect 26746 9304 26755 9344
rect 26795 9304 26804 9344
rect 26746 9303 26804 9304
rect 2667 9260 2709 9269
rect 2667 9220 2668 9260
rect 2708 9220 2709 9260
rect 2667 9211 2709 9220
rect 3627 9260 3669 9269
rect 3627 9220 3628 9260
rect 3668 9220 3669 9260
rect 3627 9211 3669 9220
rect 11019 9260 11061 9269
rect 11019 9220 11020 9260
rect 11060 9220 11061 9260
rect 11019 9211 11061 9220
rect 19995 9260 20037 9269
rect 19995 9220 19996 9260
rect 20036 9220 20037 9260
rect 19995 9211 20037 9220
rect 576 9092 31392 9116
rect 576 9052 3112 9092
rect 3480 9052 10886 9092
rect 11254 9052 18660 9092
rect 19028 9052 26434 9092
rect 26802 9052 31392 9092
rect 576 9028 31392 9052
rect 1035 8924 1077 8933
rect 1035 8884 1036 8924
rect 1076 8884 1077 8924
rect 1035 8875 1077 8884
rect 3322 8924 3380 8925
rect 3322 8884 3331 8924
rect 3371 8884 3380 8924
rect 3322 8883 3380 8884
rect 6363 8924 6405 8933
rect 6363 8884 6364 8924
rect 6404 8884 6405 8924
rect 6363 8875 6405 8884
rect 7659 8924 7701 8933
rect 7659 8884 7660 8924
rect 7700 8884 7701 8924
rect 7659 8875 7701 8884
rect 8427 8924 8469 8933
rect 8427 8884 8428 8924
rect 8468 8884 8469 8924
rect 8427 8875 8469 8884
rect 11115 8924 11157 8933
rect 11115 8884 11116 8924
rect 11156 8884 11157 8924
rect 11115 8875 11157 8884
rect 13515 8924 13557 8933
rect 13515 8884 13516 8924
rect 13556 8884 13557 8924
rect 13515 8875 13557 8884
rect 16491 8924 16533 8933
rect 16491 8884 16492 8924
rect 16532 8884 16533 8924
rect 16491 8875 16533 8884
rect 17242 8924 17300 8925
rect 17242 8884 17251 8924
rect 17291 8884 17300 8924
rect 17242 8883 17300 8884
rect 20026 8924 20084 8925
rect 20026 8884 20035 8924
rect 20075 8884 20084 8924
rect 20026 8883 20084 8884
rect 20907 8924 20949 8933
rect 20907 8884 20908 8924
rect 20948 8884 20949 8924
rect 20907 8875 20949 8884
rect 23019 8924 23061 8933
rect 23019 8884 23020 8924
rect 23060 8884 23061 8924
rect 23019 8875 23061 8884
rect 28203 8924 28245 8933
rect 28203 8884 28204 8924
rect 28244 8884 28245 8924
rect 28203 8875 28245 8884
rect 651 8840 693 8849
rect 12442 8840 12500 8841
rect 651 8800 652 8840
rect 692 8800 693 8840
rect 651 8791 693 8800
rect 9243 8831 9285 8840
rect 9243 8791 9244 8831
rect 9284 8791 9285 8831
rect 9243 8782 9285 8791
rect 12219 8831 12261 8840
rect 12219 8791 12220 8831
rect 12260 8791 12261 8831
rect 12442 8800 12451 8840
rect 12491 8800 12500 8840
rect 12442 8799 12500 8800
rect 14187 8840 14229 8849
rect 14187 8800 14188 8840
rect 14228 8800 14229 8840
rect 14187 8791 14229 8800
rect 16858 8840 16916 8841
rect 16858 8800 16867 8840
rect 16907 8800 16916 8840
rect 16858 8799 16916 8800
rect 19738 8840 19796 8841
rect 19738 8800 19747 8840
rect 19787 8800 19796 8840
rect 19738 8799 19796 8800
rect 23403 8840 23445 8849
rect 23403 8800 23404 8840
rect 23444 8800 23445 8840
rect 23403 8791 23445 8800
rect 28395 8840 28437 8849
rect 28395 8800 28396 8840
rect 28436 8800 28437 8840
rect 28395 8791 28437 8800
rect 12219 8782 12261 8791
rect 2938 8756 2996 8757
rect 2938 8716 2947 8756
rect 2987 8716 2996 8756
rect 2938 8715 2996 8716
rect 4785 8756 4827 8765
rect 4785 8716 4786 8756
rect 4826 8716 4827 8756
rect 4785 8707 4827 8716
rect 9963 8756 10005 8765
rect 9963 8716 9964 8756
rect 10004 8716 10005 8756
rect 9963 8707 10005 8716
rect 12651 8756 12693 8765
rect 12651 8716 12652 8756
rect 12692 8716 12693 8756
rect 12651 8707 12693 8716
rect 13227 8756 13269 8765
rect 13227 8716 13228 8756
rect 13268 8716 13269 8756
rect 13227 8707 13269 8716
rect 15531 8756 15573 8765
rect 15531 8716 15532 8756
rect 15572 8716 15573 8756
rect 15531 8707 15573 8716
rect 25137 8756 25179 8765
rect 25137 8716 25138 8756
rect 25178 8716 25179 8756
rect 25137 8707 25179 8716
rect 25947 8756 25989 8765
rect 25947 8716 25948 8756
rect 25988 8716 25989 8756
rect 25947 8707 25989 8716
rect 2554 8672 2612 8673
rect 2554 8632 2563 8672
rect 2603 8632 2612 8672
rect 2554 8631 2612 8632
rect 3328 8672 3370 8681
rect 3328 8632 3329 8672
rect 3369 8632 3370 8672
rect 3328 8623 3370 8632
rect 3619 8672 3677 8673
rect 3619 8632 3628 8672
rect 3668 8632 3677 8672
rect 3619 8631 3677 8632
rect 3819 8672 3861 8681
rect 3819 8632 3820 8672
rect 3860 8632 3861 8672
rect 3819 8623 3861 8632
rect 4203 8672 4245 8681
rect 4203 8632 4204 8672
rect 4244 8632 4245 8672
rect 4203 8623 4245 8632
rect 4875 8672 4917 8681
rect 4875 8632 4876 8672
rect 4916 8632 4917 8672
rect 4875 8623 4917 8632
rect 5451 8672 5493 8681
rect 5451 8632 5452 8672
rect 5492 8632 5493 8672
rect 5451 8623 5493 8632
rect 5674 8672 5732 8673
rect 5674 8632 5683 8672
rect 5723 8632 5732 8672
rect 5674 8631 5732 8632
rect 6027 8672 6069 8681
rect 6027 8632 6028 8672
rect 6068 8632 6069 8672
rect 6027 8623 6069 8632
rect 6603 8672 6645 8681
rect 6603 8632 6604 8672
rect 6644 8632 6645 8672
rect 6603 8623 6645 8632
rect 6987 8672 7029 8681
rect 7375 8679 7417 8688
rect 6987 8632 6988 8672
rect 7028 8632 7029 8672
rect 6987 8623 7029 8632
rect 7258 8672 7316 8673
rect 7258 8632 7267 8672
rect 7307 8632 7316 8672
rect 7258 8631 7316 8632
rect 7375 8639 7376 8679
rect 7416 8639 7417 8679
rect 7375 8630 7417 8639
rect 8122 8672 8180 8673
rect 8122 8632 8131 8672
rect 8171 8632 8180 8672
rect 8122 8631 8180 8632
rect 8235 8672 8277 8681
rect 8235 8632 8236 8672
rect 8276 8632 8277 8672
rect 8235 8623 8277 8632
rect 9274 8672 9332 8673
rect 9274 8632 9283 8672
rect 9323 8632 9332 8672
rect 9274 8631 9332 8632
rect 9634 8672 9692 8673
rect 9634 8632 9643 8672
rect 9683 8632 9692 8672
rect 9634 8631 9692 8632
rect 9754 8672 9812 8673
rect 9754 8632 9763 8672
rect 9803 8632 9812 8672
rect 9754 8631 9812 8632
rect 9867 8672 9909 8681
rect 9867 8632 9868 8672
rect 9908 8632 9909 8672
rect 9867 8623 9909 8632
rect 10327 8672 10385 8673
rect 10327 8632 10336 8672
rect 10376 8632 10385 8672
rect 10327 8631 10385 8632
rect 10810 8672 10868 8673
rect 10810 8632 10819 8672
rect 10859 8632 10868 8672
rect 10810 8631 10868 8632
rect 11787 8672 11829 8681
rect 11787 8632 11788 8672
rect 11828 8632 11829 8672
rect 11787 8623 11829 8632
rect 12250 8672 12308 8673
rect 12250 8632 12259 8672
rect 12299 8632 12308 8672
rect 12250 8631 12308 8632
rect 12826 8672 12884 8673
rect 12826 8632 12835 8672
rect 12875 8632 12884 8672
rect 12826 8631 12884 8632
rect 13563 8672 13605 8681
rect 13563 8632 13564 8672
rect 13604 8632 13605 8672
rect 13563 8623 13605 8632
rect 13707 8672 13749 8681
rect 13707 8632 13708 8672
rect 13748 8632 13749 8672
rect 13707 8623 13749 8632
rect 14187 8672 14229 8681
rect 14187 8632 14188 8672
rect 14228 8632 14229 8672
rect 14187 8623 14229 8632
rect 14379 8672 14421 8681
rect 14379 8632 14380 8672
rect 14420 8632 14421 8672
rect 14379 8623 14421 8632
rect 15034 8672 15092 8673
rect 15034 8632 15043 8672
rect 15083 8632 15092 8672
rect 15034 8631 15092 8632
rect 15147 8672 15189 8681
rect 15147 8632 15148 8672
rect 15188 8632 15189 8672
rect 15147 8623 15189 8632
rect 15627 8672 15669 8681
rect 15627 8632 15628 8672
rect 15668 8632 15669 8672
rect 15627 8623 15669 8632
rect 15746 8672 15788 8681
rect 15746 8632 15747 8672
rect 15787 8632 15788 8672
rect 15746 8623 15788 8632
rect 15856 8672 15914 8673
rect 15856 8632 15865 8672
rect 15905 8632 15914 8672
rect 15856 8631 15914 8632
rect 16186 8672 16244 8673
rect 16186 8632 16195 8672
rect 16235 8632 16244 8672
rect 16186 8631 16244 8632
rect 16491 8672 16533 8681
rect 16491 8632 16492 8672
rect 16532 8632 16533 8672
rect 16491 8623 16533 8632
rect 16683 8672 16725 8681
rect 16683 8632 16684 8672
rect 16724 8632 16725 8672
rect 16683 8623 16725 8632
rect 16858 8672 16916 8673
rect 16858 8632 16867 8672
rect 16907 8632 16916 8672
rect 16858 8631 16916 8632
rect 17067 8672 17109 8681
rect 17067 8632 17068 8672
rect 17108 8632 17109 8672
rect 17067 8623 17109 8632
rect 17242 8672 17300 8673
rect 17242 8632 17251 8672
rect 17291 8632 17300 8672
rect 17242 8631 17300 8632
rect 17869 8672 17927 8673
rect 17869 8632 17878 8672
rect 17918 8632 17927 8672
rect 17869 8631 17927 8632
rect 18507 8672 18549 8681
rect 18507 8632 18508 8672
rect 18548 8632 18549 8672
rect 18507 8623 18549 8632
rect 18641 8672 18699 8673
rect 18641 8632 18650 8672
rect 18690 8632 18699 8672
rect 18641 8631 18699 8632
rect 19450 8672 19508 8673
rect 19450 8632 19459 8672
rect 19499 8632 19508 8672
rect 19450 8631 19508 8632
rect 19563 8672 19605 8681
rect 19563 8632 19564 8672
rect 19604 8632 19605 8672
rect 19563 8623 19605 8632
rect 20235 8672 20277 8681
rect 20235 8632 20236 8672
rect 20276 8632 20277 8672
rect 20235 8623 20277 8632
rect 20323 8672 20381 8673
rect 20323 8632 20332 8672
rect 20372 8632 20381 8672
rect 20323 8631 20381 8632
rect 20602 8672 20660 8673
rect 20602 8632 20611 8672
rect 20651 8632 20660 8672
rect 20602 8631 20660 8632
rect 21466 8672 21524 8673
rect 21466 8632 21475 8672
rect 21515 8632 21524 8672
rect 21466 8631 21524 8632
rect 24171 8672 24213 8681
rect 24171 8632 24172 8672
rect 24212 8632 24213 8672
rect 24171 8623 24213 8632
rect 24555 8672 24597 8681
rect 24555 8632 24556 8672
rect 24596 8632 24597 8672
rect 24555 8623 24597 8632
rect 25227 8672 25269 8681
rect 25227 8632 25228 8672
rect 25268 8632 25269 8672
rect 25227 8623 25269 8632
rect 25803 8672 25845 8681
rect 25803 8632 25804 8672
rect 25844 8632 25845 8672
rect 25803 8623 25845 8632
rect 26763 8672 26805 8681
rect 26763 8632 26764 8672
rect 26804 8632 26805 8672
rect 26763 8623 26805 8632
rect 27147 8672 27189 8681
rect 27147 8632 27148 8672
rect 27188 8632 27189 8672
rect 27147 8623 27189 8632
rect 27235 8672 27293 8673
rect 27235 8632 27244 8672
rect 27284 8632 27293 8672
rect 27235 8631 27293 8632
rect 27531 8672 27573 8681
rect 27531 8632 27532 8672
rect 27572 8632 27573 8672
rect 27531 8623 27573 8632
rect 29067 8672 29109 8681
rect 29067 8632 29068 8672
rect 29108 8632 29109 8672
rect 29067 8623 29109 8632
rect 8438 8588 8480 8597
rect 8438 8548 8439 8588
rect 8479 8548 8480 8588
rect 8438 8539 8480 8548
rect 9483 8588 9525 8597
rect 9483 8548 9484 8588
rect 9524 8548 9525 8588
rect 9483 8539 9525 8548
rect 10491 8588 10533 8597
rect 10491 8548 10492 8588
rect 10532 8548 10533 8588
rect 10491 8539 10533 8548
rect 11129 8588 11171 8597
rect 11129 8548 11130 8588
rect 11170 8548 11171 8588
rect 11129 8539 11171 8548
rect 13131 8588 13173 8597
rect 13131 8548 13132 8588
rect 13172 8548 13173 8588
rect 13131 8539 13173 8548
rect 15243 8588 15285 8597
rect 15243 8548 15244 8588
rect 15284 8548 15285 8588
rect 15243 8539 15285 8548
rect 15350 8588 15392 8597
rect 15350 8548 15351 8588
rect 15391 8548 15392 8588
rect 15350 8539 15392 8548
rect 17674 8588 17732 8589
rect 17674 8548 17683 8588
rect 17723 8548 17732 8588
rect 17674 8547 17732 8548
rect 20029 8588 20071 8597
rect 20029 8548 20030 8588
rect 20070 8548 20071 8588
rect 20029 8539 20071 8548
rect 20918 8588 20960 8597
rect 20918 8548 20919 8588
rect 20959 8548 20960 8588
rect 20918 8539 20960 8548
rect 21082 8588 21140 8589
rect 21082 8548 21091 8588
rect 21131 8548 21140 8588
rect 21082 8547 21140 8548
rect 26941 8588 26983 8597
rect 26941 8548 26942 8588
rect 26982 8548 26983 8588
rect 26941 8539 26983 8548
rect 27034 8588 27092 8589
rect 27034 8548 27043 8588
rect 27083 8548 27092 8588
rect 27034 8547 27092 8548
rect 3531 8504 3573 8513
rect 3531 8464 3532 8504
rect 3572 8464 3573 8504
rect 3531 8455 3573 8464
rect 4299 8504 4341 8513
rect 4299 8464 4300 8504
rect 4340 8464 4341 8504
rect 4299 8455 4341 8464
rect 4570 8504 4628 8505
rect 4570 8464 4579 8504
rect 4619 8464 4628 8504
rect 4570 8463 4628 8464
rect 5307 8504 5349 8513
rect 5307 8464 5308 8504
rect 5348 8464 5349 8504
rect 5307 8455 5349 8464
rect 6123 8504 6165 8513
rect 10906 8504 10964 8505
rect 6123 8464 6124 8504
rect 6164 8464 6165 8504
rect 6123 8455 6165 8464
rect 7170 8495 7216 8504
rect 7170 8455 7171 8495
rect 7211 8455 7216 8495
rect 10906 8464 10915 8504
rect 10955 8464 10964 8504
rect 10906 8463 10964 8464
rect 11674 8504 11732 8505
rect 11674 8464 11683 8504
rect 11723 8464 11732 8504
rect 11674 8463 11732 8464
rect 11979 8504 12021 8513
rect 11979 8464 11980 8504
rect 12020 8464 12021 8504
rect 11979 8455 12021 8464
rect 18795 8504 18837 8513
rect 18795 8464 18796 8504
rect 18836 8464 18837 8504
rect 18795 8455 18837 8464
rect 20698 8504 20756 8505
rect 20698 8464 20707 8504
rect 20747 8464 20756 8504
rect 20698 8463 20756 8464
rect 24651 8504 24693 8513
rect 24651 8464 24652 8504
rect 24692 8464 24693 8504
rect 24651 8455 24693 8464
rect 24922 8504 24980 8505
rect 24922 8464 24931 8504
rect 24971 8464 24980 8504
rect 24922 8463 24980 8464
rect 26091 8504 26133 8513
rect 26091 8464 26092 8504
rect 26132 8464 26133 8504
rect 26091 8455 26133 8464
rect 7170 8446 7216 8455
rect 576 8336 31392 8360
rect 576 8296 4352 8336
rect 4720 8296 12126 8336
rect 12494 8296 19900 8336
rect 20268 8296 27674 8336
rect 28042 8296 31392 8336
rect 576 8272 31392 8296
rect 1467 8168 1509 8177
rect 1467 8128 1468 8168
rect 1508 8128 1509 8168
rect 1467 8119 1509 8128
rect 3034 8168 3092 8169
rect 3034 8128 3043 8168
rect 3083 8128 3092 8168
rect 3034 8127 3092 8128
rect 3339 8168 3381 8177
rect 3339 8128 3340 8168
rect 3380 8128 3381 8168
rect 3339 8119 3381 8128
rect 3802 8168 3860 8169
rect 3802 8128 3811 8168
rect 3851 8128 3860 8168
rect 3802 8127 3860 8128
rect 5818 8168 5876 8169
rect 5818 8128 5827 8168
rect 5867 8128 5876 8168
rect 5818 8127 5876 8128
rect 6298 8168 6356 8169
rect 6298 8128 6307 8168
rect 6347 8128 6356 8168
rect 6298 8127 6356 8128
rect 6603 8168 6645 8177
rect 6603 8128 6604 8168
rect 6644 8128 6645 8168
rect 6603 8119 6645 8128
rect 7659 8168 7701 8177
rect 7659 8128 7660 8168
rect 7700 8128 7701 8168
rect 7659 8119 7701 8128
rect 9082 8168 9140 8169
rect 9082 8128 9091 8168
rect 9131 8128 9140 8168
rect 9082 8127 9140 8128
rect 9850 8168 9908 8169
rect 9850 8128 9859 8168
rect 9899 8128 9908 8168
rect 9850 8127 9908 8128
rect 9963 8168 10005 8177
rect 9963 8128 9964 8168
rect 10004 8128 10005 8168
rect 9963 8119 10005 8128
rect 10731 8168 10773 8177
rect 10731 8128 10732 8168
rect 10772 8128 10773 8168
rect 10731 8119 10773 8128
rect 11403 8168 11445 8177
rect 11403 8128 11404 8168
rect 11444 8128 11445 8168
rect 11403 8119 11445 8128
rect 15819 8168 15861 8177
rect 15819 8128 15820 8168
rect 15860 8128 15861 8168
rect 15819 8119 15861 8128
rect 16186 8168 16244 8169
rect 16186 8128 16195 8168
rect 16235 8128 16244 8168
rect 16186 8127 16244 8128
rect 17530 8168 17588 8169
rect 17530 8128 17539 8168
rect 17579 8128 17588 8168
rect 17530 8127 17588 8128
rect 18202 8168 18260 8169
rect 18202 8128 18211 8168
rect 18251 8128 18260 8168
rect 18202 8127 18260 8128
rect 20122 8168 20180 8169
rect 20122 8128 20131 8168
rect 20171 8128 20180 8168
rect 20122 8127 20180 8128
rect 20331 8168 20373 8177
rect 20331 8128 20332 8168
rect 20372 8128 20373 8168
rect 20331 8119 20373 8128
rect 21099 8168 21141 8177
rect 21099 8128 21100 8168
rect 21140 8128 21141 8168
rect 21099 8119 21141 8128
rect 28107 8168 28149 8177
rect 28107 8128 28108 8168
rect 28148 8128 28149 8168
rect 28107 8119 28149 8128
rect 2763 8084 2805 8093
rect 2763 8044 2764 8084
rect 2804 8044 2805 8084
rect 2763 8035 2805 8044
rect 11979 8084 12021 8093
rect 11979 8044 11980 8084
rect 12020 8044 12021 8084
rect 11979 8035 12021 8044
rect 12183 8084 12225 8093
rect 12183 8044 12184 8084
rect 12224 8044 12225 8084
rect 12183 8035 12225 8044
rect 13018 8084 13076 8085
rect 13018 8044 13027 8084
rect 13067 8044 13076 8084
rect 13018 8043 13076 8044
rect 22138 8084 22196 8085
rect 25131 8084 25173 8093
rect 22138 8044 22147 8084
rect 22187 8044 22196 8084
rect 22138 8043 22196 8044
rect 24066 8075 24112 8084
rect 24066 8035 24067 8075
rect 24107 8035 24112 8075
rect 25131 8044 25132 8084
rect 25172 8044 25173 8084
rect 25131 8035 25173 8044
rect 25786 8084 25844 8085
rect 25786 8044 25795 8084
rect 25835 8044 25844 8084
rect 25786 8043 25844 8044
rect 24066 8026 24112 8035
rect 2667 8000 2709 8009
rect 1314 7991 1360 8000
rect 1314 7951 1315 7991
rect 1355 7951 1360 7991
rect 2667 7960 2668 8000
rect 2708 7960 2709 8000
rect 2667 7951 2709 7960
rect 2842 8000 2900 8001
rect 2842 7960 2851 8000
rect 2891 7960 2900 8000
rect 2842 7959 2900 7960
rect 3147 8000 3189 8009
rect 3147 7960 3148 8000
rect 3188 7960 3189 8000
rect 3147 7951 3189 7960
rect 4107 8000 4149 8009
rect 4107 7960 4108 8000
rect 4148 7960 4149 8000
rect 4107 7951 4149 7960
rect 4836 8000 4894 8001
rect 4836 7960 4845 8000
rect 4885 7960 4894 8000
rect 4836 7959 4894 7960
rect 4992 8000 5034 8009
rect 4992 7960 4993 8000
rect 5033 7960 5034 8000
rect 4992 7951 5034 7960
rect 5284 8000 5326 8009
rect 5284 7960 5285 8000
rect 5325 7960 5326 8000
rect 5284 7951 5326 7960
rect 5931 8000 5973 8009
rect 5931 7960 5932 8000
rect 5972 7960 5973 8000
rect 5931 7951 5973 7960
rect 6411 8000 6453 8009
rect 6411 7960 6412 8000
rect 6452 7960 6453 8000
rect 6411 7951 6453 7960
rect 7258 8000 7316 8001
rect 7258 7960 7267 8000
rect 7307 7960 7316 8000
rect 7258 7959 7316 7960
rect 7371 8000 7413 8009
rect 7371 7960 7372 8000
rect 7412 7960 7413 8000
rect 7371 7951 7413 7960
rect 8026 8000 8084 8001
rect 8026 7960 8035 8000
rect 8075 7960 8084 8000
rect 8026 7959 8084 7960
rect 8139 8000 8181 8009
rect 8139 7960 8140 8000
rect 8180 7960 8181 8000
rect 8139 7951 8181 7960
rect 8619 8000 8661 8009
rect 8619 7960 8620 8000
rect 8660 7960 8661 8000
rect 8619 7951 8661 7960
rect 8811 8000 8853 8009
rect 8811 7960 8812 8000
rect 8852 7960 8853 8000
rect 8811 7951 8853 7960
rect 9291 8000 9333 8009
rect 9291 7960 9292 8000
rect 9332 7960 9333 8000
rect 9291 7951 9333 7960
rect 9579 8000 9621 8009
rect 9579 7960 9580 8000
rect 9620 7960 9621 8000
rect 9579 7951 9621 7960
rect 9754 8000 9812 8001
rect 9754 7960 9763 8000
rect 9803 7960 9812 8000
rect 9754 7959 9812 7960
rect 10073 8000 10115 8009
rect 10073 7960 10074 8000
rect 10114 7960 10115 8000
rect 10073 7951 10115 7960
rect 10251 8000 10293 8009
rect 10251 7960 10252 8000
rect 10292 7960 10293 8000
rect 10251 7951 10293 7960
rect 10635 8000 10677 8009
rect 10635 7960 10636 8000
rect 10676 7960 10677 8000
rect 10635 7951 10677 7960
rect 11499 8000 11541 8009
rect 11499 7960 11500 8000
rect 11540 7960 11541 8000
rect 11499 7951 11541 7960
rect 11716 8000 11758 8009
rect 11716 7960 11717 8000
rect 11757 7960 11758 8000
rect 11716 7951 11758 7960
rect 11866 8000 11924 8001
rect 11866 7960 11875 8000
rect 11915 7960 11924 8000
rect 11866 7959 11924 7960
rect 12694 8000 12736 8009
rect 12694 7960 12695 8000
rect 12735 7960 12736 8000
rect 12694 7951 12736 7960
rect 12930 8000 12972 8009
rect 12930 7960 12931 8000
rect 12971 7960 12972 8000
rect 12930 7951 12972 7960
rect 13275 8000 13317 8009
rect 13275 7960 13276 8000
rect 13316 7960 13317 8000
rect 13275 7951 13317 7960
rect 13576 8000 13618 8009
rect 13576 7960 13577 8000
rect 13617 7960 13618 8000
rect 13576 7951 13618 7960
rect 13730 8000 13772 8009
rect 13730 7960 13731 8000
rect 13771 7960 13772 8000
rect 13730 7951 13772 7960
rect 14475 8000 14517 8009
rect 14475 7960 14476 8000
rect 14516 7960 14517 8000
rect 14475 7951 14517 7960
rect 14602 8000 14660 8001
rect 14602 7960 14611 8000
rect 14651 7960 14660 8000
rect 14602 7959 14660 7960
rect 14955 8000 14997 8009
rect 14955 7960 14956 8000
rect 14996 7960 14997 8000
rect 14955 7951 14997 7960
rect 15147 8000 15189 8009
rect 15147 7960 15148 8000
rect 15188 7960 15189 8000
rect 15147 7951 15189 7960
rect 15370 8000 15428 8001
rect 15370 7960 15379 8000
rect 15419 7960 15428 8000
rect 15370 7959 15428 7960
rect 15723 8000 15765 8009
rect 15723 7960 15724 8000
rect 15764 7960 15765 8000
rect 15723 7951 15765 7960
rect 16395 8000 16437 8009
rect 16395 7960 16396 8000
rect 16436 7960 16437 8000
rect 16395 7951 16437 7960
rect 16683 8000 16725 8009
rect 16683 7960 16684 8000
rect 16724 7960 16725 8000
rect 16683 7951 16725 7960
rect 17206 8000 17248 8009
rect 17206 7960 17207 8000
rect 17247 7960 17248 8000
rect 17206 7951 17248 7960
rect 17451 8000 17493 8009
rect 17451 7960 17452 8000
rect 17492 7960 17493 8000
rect 17451 7951 17493 7960
rect 17739 8000 17781 8009
rect 17739 7960 17740 8000
rect 17780 7960 17781 8000
rect 17739 7951 17781 7960
rect 18027 8000 18069 8009
rect 18027 7960 18028 8000
rect 18068 7960 18069 8000
rect 18027 7951 18069 7960
rect 18363 8000 18405 8009
rect 18363 7960 18364 8000
rect 18404 7960 18405 8000
rect 18363 7951 18405 7960
rect 18507 8000 18549 8009
rect 18507 7960 18508 8000
rect 18548 7960 18549 8000
rect 18507 7951 18549 7960
rect 19258 8000 19316 8001
rect 19258 7960 19267 8000
rect 19307 7960 19316 8000
rect 19258 7959 19316 7960
rect 19371 8000 19413 8009
rect 19371 7960 19372 8000
rect 19412 7960 19413 8000
rect 19371 7951 19413 7960
rect 19798 8000 19840 8009
rect 19798 7960 19799 8000
rect 19839 7960 19840 8000
rect 19798 7951 19840 7960
rect 20043 8000 20085 8009
rect 20043 7960 20044 8000
rect 20084 7960 20085 8000
rect 20043 7951 20085 7960
rect 20427 8000 20469 8009
rect 20427 7960 20428 8000
rect 20468 7960 20469 8000
rect 20427 7951 20469 7960
rect 20658 8000 20700 8009
rect 20658 7960 20659 8000
rect 20699 7960 20700 8000
rect 20658 7951 20700 7960
rect 21771 8000 21813 8009
rect 21771 7960 21772 8000
rect 21812 7960 21813 8000
rect 21771 7951 21813 7960
rect 22827 8000 22869 8009
rect 22827 7960 22828 8000
rect 22868 7960 22869 8000
rect 22827 7951 22869 7960
rect 23307 8000 23349 8009
rect 23307 7960 23308 8000
rect 23348 7960 23349 8000
rect 23307 7951 23349 7960
rect 23770 8000 23828 8001
rect 24162 8000 24220 8001
rect 23770 7960 23779 8000
rect 23819 7960 23828 8000
rect 23770 7959 23828 7960
rect 23883 7991 23925 8000
rect 23883 7951 23884 7991
rect 23924 7951 23925 7991
rect 24162 7960 24171 8000
rect 24211 7960 24220 8000
rect 24541 8000 24583 8009
rect 24162 7959 24220 7960
rect 24331 7989 24389 7990
rect 1314 7942 1360 7951
rect 23883 7942 23925 7951
rect 24331 7949 24340 7989
rect 24380 7949 24389 7989
rect 24541 7960 24542 8000
rect 24582 7960 24583 8000
rect 24541 7951 24583 7960
rect 24651 8000 24693 8009
rect 24651 7960 24652 8000
rect 24692 7960 24693 8000
rect 24651 7951 24693 7960
rect 24843 8000 24885 8009
rect 24843 7960 24844 8000
rect 24884 7960 24885 8000
rect 24843 7951 24885 7960
rect 25030 8000 25072 8009
rect 25030 7960 25031 8000
rect 25071 7960 25072 8000
rect 25030 7951 25072 7960
rect 25215 8000 25257 8009
rect 25215 7960 25216 8000
rect 25256 7960 25257 8000
rect 25215 7951 25257 7960
rect 25419 8000 25461 8009
rect 25419 7960 25420 8000
rect 25460 7960 25461 8000
rect 25419 7951 25461 7960
rect 25611 8000 25653 8009
rect 25611 7960 25612 8000
rect 25652 7960 25653 8000
rect 25611 7951 25653 7960
rect 26170 8000 26228 8001
rect 26170 7960 26179 8000
rect 26219 7960 26228 8000
rect 26170 7959 26228 7960
rect 24331 7948 24389 7949
rect 4017 7916 4059 7925
rect 4017 7876 4018 7916
rect 4058 7876 4059 7916
rect 4017 7867 4059 7876
rect 5163 7916 5205 7925
rect 5163 7876 5164 7916
rect 5204 7876 5205 7916
rect 5163 7867 5205 7876
rect 11618 7916 11660 7925
rect 11618 7876 11619 7916
rect 11659 7876 11660 7916
rect 11618 7867 11660 7876
rect 12826 7916 12884 7917
rect 12826 7876 12835 7916
rect 12875 7876 12884 7916
rect 12826 7875 12884 7876
rect 13419 7916 13461 7925
rect 13419 7876 13420 7916
rect 13460 7876 13461 7916
rect 13419 7867 13461 7876
rect 17338 7916 17396 7917
rect 17338 7876 17347 7916
rect 17387 7876 17396 7916
rect 17338 7875 17396 7876
rect 19930 7916 19988 7917
rect 23217 7916 23259 7925
rect 19930 7876 19939 7916
rect 19979 7876 19988 7916
rect 19930 7875 19988 7876
rect 20562 7907 20608 7916
rect 20562 7867 20563 7907
rect 20603 7867 20608 7907
rect 23217 7876 23218 7916
rect 23258 7876 23259 7916
rect 23217 7867 23259 7876
rect 20562 7858 20608 7867
rect 1995 7832 2037 7841
rect 1995 7792 1996 7832
rect 2036 7792 2037 7832
rect 1995 7783 2037 7792
rect 5067 7832 5109 7841
rect 5067 7792 5068 7832
rect 5108 7792 5109 7832
rect 5067 7783 5109 7792
rect 13515 7832 13557 7841
rect 13515 7792 13516 7832
rect 13556 7792 13557 7832
rect 13515 7783 13557 7792
rect 17739 7832 17781 7841
rect 17739 7792 17740 7832
rect 17780 7792 17781 7832
rect 17739 7783 17781 7792
rect 19546 7832 19604 7833
rect 19546 7792 19555 7832
rect 19595 7792 19604 7832
rect 19546 7791 19604 7792
rect 24555 7832 24597 7841
rect 24555 7792 24556 7832
rect 24596 7792 24597 7832
rect 24555 7783 24597 7792
rect 25210 7832 25268 7833
rect 25210 7792 25219 7832
rect 25259 7792 25268 7832
rect 25210 7791 25268 7792
rect 28299 7832 28341 7841
rect 28299 7792 28300 7832
rect 28340 7792 28341 7832
rect 28299 7783 28341 7792
rect 6123 7748 6165 7757
rect 6123 7708 6124 7748
rect 6164 7708 6165 7748
rect 6123 7699 6165 7708
rect 8314 7748 8372 7749
rect 8314 7708 8323 7748
rect 8363 7708 8372 7748
rect 8314 7707 8372 7708
rect 8619 7748 8661 7757
rect 8619 7708 8620 7748
rect 8660 7708 8661 7748
rect 8619 7699 8661 7708
rect 12171 7748 12213 7757
rect 12171 7708 12172 7748
rect 12212 7708 12213 7748
rect 12171 7699 12213 7708
rect 14650 7748 14708 7749
rect 14650 7708 14659 7748
rect 14699 7708 14708 7748
rect 14650 7707 14708 7708
rect 14955 7748 14997 7757
rect 14955 7708 14956 7748
rect 14996 7708 14997 7748
rect 14955 7699 14997 7708
rect 23115 7748 23157 7757
rect 23115 7708 23116 7748
rect 23156 7708 23157 7748
rect 23115 7699 23157 7708
rect 23770 7748 23828 7749
rect 23770 7708 23779 7748
rect 23819 7708 23828 7748
rect 23770 7707 23828 7708
rect 25419 7748 25461 7757
rect 25419 7708 25420 7748
rect 25460 7708 25461 7748
rect 25419 7699 25461 7708
rect 27723 7748 27765 7757
rect 27723 7708 27724 7748
rect 27764 7708 27765 7748
rect 27723 7699 27765 7708
rect 576 7580 31392 7604
rect 576 7540 3112 7580
rect 3480 7540 10886 7580
rect 11254 7540 18660 7580
rect 19028 7540 26434 7580
rect 26802 7540 31392 7580
rect 576 7516 31392 7540
rect 6027 7412 6069 7421
rect 6027 7372 6028 7412
rect 6068 7372 6069 7412
rect 6027 7363 6069 7372
rect 8026 7412 8084 7413
rect 8026 7372 8035 7412
rect 8075 7372 8084 7412
rect 8026 7371 8084 7372
rect 9387 7412 9429 7421
rect 9387 7372 9388 7412
rect 9428 7372 9429 7412
rect 9387 7363 9429 7372
rect 10251 7412 10293 7421
rect 10251 7372 10252 7412
rect 10292 7372 10293 7412
rect 10251 7363 10293 7372
rect 14475 7412 14517 7421
rect 14475 7372 14476 7412
rect 14516 7372 14517 7412
rect 14475 7363 14517 7372
rect 18970 7412 19028 7413
rect 18970 7372 18979 7412
rect 19019 7372 19028 7412
rect 18970 7371 19028 7372
rect 19659 7412 19701 7421
rect 19659 7372 19660 7412
rect 19700 7372 19701 7412
rect 19659 7363 19701 7372
rect 20811 7412 20853 7421
rect 20811 7372 20812 7412
rect 20852 7372 20853 7412
rect 20811 7363 20853 7372
rect 21178 7412 21236 7413
rect 21178 7372 21187 7412
rect 21227 7372 21236 7412
rect 21178 7371 21236 7372
rect 23355 7412 23397 7421
rect 23355 7372 23356 7412
rect 23396 7372 23397 7412
rect 23355 7363 23397 7372
rect 4203 7328 4245 7337
rect 7179 7328 7221 7337
rect 4203 7288 4204 7328
rect 4244 7288 4245 7328
rect 4203 7279 4245 7288
rect 4651 7319 4693 7328
rect 4651 7279 4652 7319
rect 4692 7279 4693 7319
rect 7179 7288 7180 7328
rect 7220 7288 7221 7328
rect 7179 7279 7221 7288
rect 12891 7328 12933 7337
rect 12891 7288 12892 7328
rect 12932 7288 12933 7328
rect 12891 7279 12933 7288
rect 18490 7328 18548 7329
rect 23499 7328 23541 7337
rect 18490 7288 18499 7328
rect 18539 7288 18548 7328
rect 18490 7287 18548 7288
rect 22379 7319 22421 7328
rect 22379 7279 22380 7319
rect 22420 7279 22421 7319
rect 23499 7288 23500 7328
rect 23540 7288 23541 7328
rect 23499 7279 23541 7288
rect 4651 7270 4693 7279
rect 22379 7270 22421 7279
rect 2122 7244 2180 7245
rect 2122 7204 2131 7244
rect 2171 7204 2180 7244
rect 2122 7203 2180 7204
rect 10353 7244 10395 7253
rect 10353 7204 10354 7244
rect 10394 7204 10395 7244
rect 6891 7193 6933 7202
rect 10353 7195 10395 7204
rect 16203 7244 16245 7253
rect 16203 7204 16204 7244
rect 16244 7204 16245 7244
rect 16203 7195 16245 7204
rect 21675 7244 21717 7253
rect 21675 7204 21676 7244
rect 21716 7204 21717 7244
rect 21675 7195 21717 7204
rect 26475 7244 26517 7253
rect 26475 7204 26476 7244
rect 26516 7204 26517 7244
rect 25066 7202 25124 7203
rect 2317 7160 2375 7161
rect 2317 7120 2326 7160
rect 2366 7120 2375 7160
rect 2317 7119 2375 7120
rect 2571 7160 2613 7169
rect 2571 7120 2572 7160
rect 2612 7120 2613 7160
rect 2571 7111 2613 7120
rect 3235 7160 3293 7161
rect 3235 7120 3244 7160
rect 3284 7120 3293 7160
rect 3235 7119 3293 7120
rect 3435 7160 3477 7169
rect 3435 7120 3436 7160
rect 3476 7120 3477 7160
rect 3435 7111 3477 7120
rect 3819 7160 3861 7169
rect 3819 7120 3820 7160
rect 3860 7120 3861 7160
rect 3819 7111 3861 7120
rect 4666 7160 4724 7161
rect 4666 7120 4675 7160
rect 4715 7120 4724 7160
rect 4666 7119 4724 7120
rect 5067 7160 5109 7169
rect 5067 7120 5068 7160
rect 5108 7120 5109 7160
rect 5067 7111 5109 7120
rect 6108 7160 6150 7169
rect 6108 7120 6109 7160
rect 6149 7120 6150 7160
rect 6108 7111 6150 7120
rect 6214 7160 6272 7161
rect 6214 7120 6223 7160
rect 6263 7120 6272 7160
rect 6214 7119 6272 7120
rect 6778 7160 6836 7161
rect 6778 7120 6787 7160
rect 6827 7120 6836 7160
rect 6891 7153 6892 7193
rect 6932 7153 6933 7193
rect 6891 7144 6933 7153
rect 7738 7160 7796 7161
rect 6778 7119 6836 7120
rect 7738 7120 7747 7160
rect 7787 7120 7796 7160
rect 7738 7119 7796 7120
rect 7851 7160 7893 7169
rect 7851 7120 7852 7160
rect 7892 7120 7893 7160
rect 7851 7111 7893 7120
rect 8314 7160 8372 7161
rect 8314 7120 8323 7160
rect 8363 7120 8372 7160
rect 8314 7119 8372 7120
rect 8630 7160 8672 7169
rect 8630 7120 8631 7160
rect 8671 7120 8672 7160
rect 8630 7111 8672 7120
rect 9178 7160 9236 7161
rect 9178 7120 9187 7160
rect 9227 7120 9236 7160
rect 9178 7119 9236 7120
rect 9297 7160 9339 7169
rect 9297 7120 9298 7160
rect 9338 7120 9339 7160
rect 9297 7111 9339 7120
rect 9771 7160 9813 7169
rect 9771 7120 9772 7160
rect 9812 7120 9813 7160
rect 9771 7111 9813 7120
rect 9963 7160 10005 7169
rect 9963 7120 9964 7160
rect 10004 7120 10005 7160
rect 9963 7111 10005 7120
rect 10443 7160 10485 7169
rect 10443 7120 10444 7160
rect 10484 7120 10485 7160
rect 10443 7111 10485 7120
rect 11115 7160 11157 7169
rect 11115 7120 11116 7160
rect 11156 7120 11157 7160
rect 11115 7111 11157 7120
rect 11499 7160 11541 7169
rect 11499 7120 11500 7160
rect 11540 7120 11541 7160
rect 11499 7111 11541 7120
rect 12267 7160 12309 7169
rect 12267 7120 12268 7160
rect 12308 7120 12309 7160
rect 12267 7111 12309 7120
rect 12651 7160 12693 7169
rect 12651 7120 12652 7160
rect 12692 7120 12693 7160
rect 12651 7111 12693 7120
rect 13210 7160 13268 7161
rect 13210 7120 13219 7160
rect 13259 7120 13268 7160
rect 13210 7119 13268 7120
rect 13323 7160 13365 7169
rect 13323 7120 13324 7160
rect 13364 7120 13365 7160
rect 13323 7111 13365 7120
rect 14170 7160 14228 7161
rect 14170 7120 14179 7160
rect 14219 7120 14228 7160
rect 14170 7119 14228 7120
rect 14842 7160 14900 7161
rect 14842 7120 14851 7160
rect 14891 7120 14900 7160
rect 14842 7119 14900 7120
rect 14955 7160 14997 7169
rect 14955 7120 14956 7160
rect 14996 7120 14997 7160
rect 14955 7111 14997 7120
rect 15627 7160 15669 7169
rect 15627 7120 15628 7160
rect 15668 7120 15669 7160
rect 15627 7111 15669 7120
rect 15715 7160 15773 7161
rect 15715 7120 15724 7160
rect 15764 7120 15773 7160
rect 15715 7119 15773 7120
rect 15862 7160 15904 7169
rect 15862 7120 15863 7160
rect 15903 7120 15904 7160
rect 15862 7111 15904 7120
rect 15994 7160 16052 7161
rect 15994 7120 16003 7160
rect 16043 7120 16052 7160
rect 15994 7119 16052 7120
rect 16107 7160 16149 7169
rect 16107 7120 16108 7160
rect 16148 7120 16149 7160
rect 16107 7111 16149 7120
rect 16395 7160 16437 7169
rect 16395 7120 16396 7160
rect 16436 7120 16437 7160
rect 16395 7111 16437 7120
rect 16587 7160 16629 7169
rect 16587 7120 16588 7160
rect 16628 7120 16629 7160
rect 16587 7111 16629 7120
rect 17434 7160 17492 7161
rect 17434 7120 17443 7160
rect 17483 7120 17492 7160
rect 17434 7119 17492 7120
rect 17547 7160 17589 7169
rect 17547 7120 17548 7160
rect 17588 7120 17589 7160
rect 17547 7111 17589 7120
rect 18202 7160 18260 7161
rect 18202 7120 18211 7160
rect 18251 7120 18260 7160
rect 18202 7119 18260 7120
rect 18315 7160 18357 7169
rect 18315 7120 18316 7160
rect 18356 7120 18357 7160
rect 18315 7111 18357 7120
rect 18939 7160 18981 7169
rect 18939 7120 18940 7160
rect 18980 7120 18981 7160
rect 18939 7111 18981 7120
rect 19083 7160 19125 7169
rect 19083 7120 19084 7160
rect 19124 7120 19125 7160
rect 19083 7111 19125 7120
rect 19707 7160 19749 7169
rect 19707 7120 19708 7160
rect 19748 7120 19749 7160
rect 19707 7111 19749 7120
rect 19851 7160 19893 7169
rect 19851 7120 19852 7160
rect 19892 7120 19893 7160
rect 19851 7111 19893 7120
rect 20602 7160 20660 7161
rect 20602 7120 20611 7160
rect 20651 7120 20660 7160
rect 20602 7119 20660 7120
rect 20715 7160 20757 7169
rect 20715 7120 20716 7160
rect 20756 7120 20757 7160
rect 20715 7111 20757 7120
rect 21181 7160 21223 7169
rect 21181 7120 21182 7160
rect 21222 7120 21223 7160
rect 21181 7111 21223 7120
rect 21475 7160 21533 7161
rect 21475 7120 21484 7160
rect 21524 7120 21533 7160
rect 21475 7119 21533 7120
rect 21771 7160 21813 7169
rect 21771 7120 21772 7160
rect 21812 7120 21813 7160
rect 21771 7111 21813 7120
rect 21890 7160 21932 7169
rect 21890 7120 21891 7160
rect 21931 7120 21932 7160
rect 21890 7111 21932 7120
rect 22000 7160 22058 7161
rect 22000 7120 22009 7160
rect 22049 7120 22058 7160
rect 22000 7119 22058 7120
rect 22330 7160 22388 7161
rect 22330 7120 22339 7160
rect 22379 7120 22388 7160
rect 22330 7119 22388 7120
rect 22731 7160 22773 7169
rect 22731 7120 22732 7160
rect 22772 7120 22773 7160
rect 22731 7111 22773 7120
rect 23019 7160 23061 7169
rect 25066 7162 25075 7202
rect 25115 7162 25124 7202
rect 26475 7195 26517 7204
rect 25066 7161 25124 7162
rect 23019 7120 23020 7160
rect 23060 7120 23061 7160
rect 23019 7111 23061 7120
rect 24055 7160 24113 7161
rect 24055 7120 24064 7160
rect 24104 7120 24113 7160
rect 24055 7119 24113 7120
rect 25227 7160 25269 7169
rect 25227 7120 25228 7160
rect 25268 7120 25269 7160
rect 25227 7111 25269 7120
rect 25419 7160 25461 7169
rect 25419 7120 25420 7160
rect 25460 7120 25461 7160
rect 25419 7111 25461 7120
rect 26134 7160 26176 7169
rect 26134 7120 26135 7160
rect 26175 7120 26176 7160
rect 26134 7111 26176 7120
rect 26266 7160 26324 7161
rect 26266 7120 26275 7160
rect 26315 7120 26324 7160
rect 26266 7119 26324 7120
rect 26379 7160 26421 7169
rect 26379 7120 26380 7160
rect 26420 7120 26421 7160
rect 26379 7111 26421 7120
rect 27226 7160 27284 7161
rect 27226 7120 27235 7160
rect 27275 7120 27284 7160
rect 27226 7119 27284 7120
rect 27542 7160 27584 7169
rect 27542 7120 27543 7160
rect 27583 7120 27584 7160
rect 27542 7111 27584 7120
rect 2941 7076 2983 7085
rect 2941 7036 2942 7076
rect 2982 7036 2983 7076
rect 2941 7027 2983 7036
rect 4875 7076 4917 7085
rect 4875 7036 4876 7076
rect 4916 7036 4917 7076
rect 4875 7027 4917 7036
rect 8523 7076 8565 7085
rect 8523 7036 8524 7076
rect 8564 7036 8565 7076
rect 8523 7027 8565 7036
rect 14283 7076 14325 7085
rect 14283 7036 14284 7076
rect 14324 7036 14325 7076
rect 14283 7027 14325 7036
rect 14489 7076 14531 7085
rect 14489 7036 14490 7076
rect 14530 7036 14531 7076
rect 14489 7027 14531 7036
rect 15424 7076 15466 7085
rect 15424 7036 15425 7076
rect 15465 7036 15466 7076
rect 15424 7027 15466 7036
rect 21387 7076 21429 7085
rect 21387 7036 21388 7076
rect 21428 7036 21429 7076
rect 21387 7027 21429 7036
rect 24219 7076 24261 7085
rect 24219 7036 24220 7076
rect 24260 7036 24261 7076
rect 24219 7027 24261 7036
rect 25323 7076 25365 7085
rect 25323 7036 25324 7076
rect 25364 7036 25365 7076
rect 25323 7027 25365 7036
rect 27435 7076 27477 7085
rect 27435 7036 27436 7076
rect 27476 7036 27477 7076
rect 27435 7027 27477 7036
rect 2458 6992 2516 6993
rect 2458 6952 2467 6992
rect 2507 6952 2516 6992
rect 2458 6951 2516 6952
rect 2763 6992 2805 7001
rect 2763 6952 2764 6992
rect 2804 6952 2805 6992
rect 2763 6943 2805 6952
rect 3034 6992 3092 6993
rect 3034 6952 3043 6992
rect 3083 6952 3092 6992
rect 3034 6951 3092 6952
rect 3147 6992 3189 7001
rect 3147 6952 3148 6992
rect 3188 6952 3189 6992
rect 3147 6943 3189 6952
rect 3915 6992 3957 7001
rect 3915 6952 3916 6992
rect 3956 6952 3957 6992
rect 3915 6943 3957 6952
rect 5739 6992 5781 7001
rect 8410 6992 8468 6993
rect 5739 6952 5740 6992
rect 5780 6952 5781 6992
rect 5739 6943 5781 6952
rect 6690 6983 6736 6992
rect 6690 6943 6691 6983
rect 6731 6943 6736 6983
rect 8410 6952 8419 6992
rect 8459 6952 8468 6992
rect 8410 6951 8468 6952
rect 9946 6992 10004 6993
rect 9946 6952 9955 6992
rect 9995 6952 10004 6992
rect 9946 6951 10004 6952
rect 10138 6992 10196 6993
rect 10138 6952 10147 6992
rect 10187 6952 10196 6992
rect 10138 6951 10196 6952
rect 11595 6992 11637 7001
rect 11595 6952 11596 6992
rect 11636 6952 11637 6992
rect 11595 6943 11637 6952
rect 13611 6992 13653 7001
rect 13611 6952 13612 6992
rect 13652 6952 13653 6992
rect 13611 6943 13653 6952
rect 15243 6992 15285 7001
rect 15243 6952 15244 6992
rect 15284 6952 15285 6992
rect 15243 6943 15285 6952
rect 15514 6992 15572 6993
rect 15514 6952 15523 6992
rect 15563 6952 15572 6992
rect 15514 6951 15572 6952
rect 15627 6992 15669 7001
rect 15627 6952 15628 6992
rect 15668 6952 15669 6992
rect 15627 6943 15669 6952
rect 16395 6992 16437 7001
rect 16395 6952 16396 6992
rect 16436 6952 16437 6992
rect 16395 6943 16437 6952
rect 17835 6992 17877 7001
rect 17835 6952 17836 6992
rect 17876 6952 17877 6992
rect 17835 6943 17877 6952
rect 21003 6992 21045 7001
rect 21003 6952 21004 6992
rect 21044 6952 21045 6992
rect 21003 6943 21045 6952
rect 22155 6992 22197 7001
rect 22155 6952 22156 6992
rect 22196 6952 22197 6992
rect 22155 6943 22197 6952
rect 24874 6992 24932 6993
rect 24874 6952 24883 6992
rect 24923 6952 24932 6992
rect 24874 6951 24932 6952
rect 27322 6992 27380 6993
rect 27322 6952 27331 6992
rect 27371 6952 27380 6992
rect 27322 6951 27380 6952
rect 6690 6934 6736 6943
rect 576 6824 31392 6848
rect 576 6784 4352 6824
rect 4720 6784 12126 6824
rect 12494 6784 19900 6824
rect 20268 6784 27674 6824
rect 28042 6784 31392 6824
rect 576 6760 31392 6784
rect 5067 6656 5109 6665
rect 5067 6616 5068 6656
rect 5108 6616 5109 6656
rect 5067 6607 5109 6616
rect 6219 6656 6261 6665
rect 6219 6616 6220 6656
rect 6260 6616 6261 6656
rect 6219 6607 6261 6616
rect 7659 6656 7701 6665
rect 7659 6616 7660 6656
rect 7700 6616 7701 6656
rect 7659 6607 7701 6616
rect 8811 6656 8853 6665
rect 8811 6616 8812 6656
rect 8852 6616 8853 6656
rect 8811 6607 8853 6616
rect 9675 6656 9717 6665
rect 9675 6616 9676 6656
rect 9716 6616 9717 6656
rect 9675 6607 9717 6616
rect 9850 6656 9908 6657
rect 9850 6616 9859 6656
rect 9899 6616 9908 6656
rect 9850 6615 9908 6616
rect 11787 6656 11829 6665
rect 11787 6616 11788 6656
rect 11828 6616 11829 6656
rect 11787 6607 11829 6616
rect 12250 6656 12308 6657
rect 12250 6616 12259 6656
rect 12299 6616 12308 6656
rect 12250 6615 12308 6616
rect 13323 6656 13365 6665
rect 13323 6616 13324 6656
rect 13364 6616 13365 6656
rect 13323 6607 13365 6616
rect 13690 6656 13748 6657
rect 13690 6616 13699 6656
rect 13739 6616 13748 6656
rect 13690 6615 13748 6616
rect 16107 6656 16149 6665
rect 16107 6616 16108 6656
rect 16148 6616 16149 6656
rect 16107 6607 16149 6616
rect 16779 6656 16821 6665
rect 16779 6616 16780 6656
rect 16820 6616 16821 6656
rect 16779 6607 16821 6616
rect 19162 6656 19220 6657
rect 19162 6616 19171 6656
rect 19211 6616 19220 6656
rect 19162 6615 19220 6616
rect 19930 6656 19988 6657
rect 19930 6616 19939 6656
rect 19979 6616 19988 6656
rect 19930 6615 19988 6616
rect 20986 6656 21044 6657
rect 20986 6616 20995 6656
rect 21035 6616 21044 6656
rect 20986 6615 21044 6616
rect 21754 6656 21812 6657
rect 21754 6616 21763 6656
rect 21803 6616 21812 6656
rect 21754 6615 21812 6616
rect 22234 6656 22292 6657
rect 22234 6616 22243 6656
rect 22283 6616 22292 6656
rect 22234 6615 22292 6616
rect 23866 6656 23924 6657
rect 23866 6616 23875 6656
rect 23915 6616 23924 6656
rect 23866 6615 23924 6616
rect 23979 6656 24021 6665
rect 23979 6616 23980 6656
rect 24020 6616 24021 6656
rect 23979 6607 24021 6616
rect 24363 6656 24405 6665
rect 24363 6616 24364 6656
rect 24404 6616 24405 6656
rect 24363 6607 24405 6616
rect 2746 6572 2804 6573
rect 2746 6532 2755 6572
rect 2795 6532 2804 6572
rect 2746 6531 2804 6532
rect 8122 6572 8180 6573
rect 8122 6532 8131 6572
rect 8171 6532 8180 6572
rect 8122 6531 8180 6532
rect 13913 6572 13955 6581
rect 13913 6532 13914 6572
rect 13954 6532 13955 6572
rect 13913 6523 13955 6532
rect 15243 6572 15285 6581
rect 15243 6532 15244 6572
rect 15284 6532 15285 6572
rect 15243 6523 15285 6532
rect 2379 6488 2421 6497
rect 2379 6448 2380 6488
rect 2420 6448 2421 6488
rect 2379 6439 2421 6448
rect 2596 6488 2638 6497
rect 2596 6448 2597 6488
rect 2637 6448 2638 6488
rect 2596 6439 2638 6448
rect 3130 6488 3188 6489
rect 3130 6448 3139 6488
rect 3179 6448 3188 6488
rect 3130 6447 3188 6448
rect 5581 6488 5639 6489
rect 5581 6448 5590 6488
rect 5630 6448 5639 6488
rect 5581 6447 5639 6448
rect 5931 6488 5973 6497
rect 5931 6448 5932 6488
rect 5972 6448 5973 6488
rect 5931 6439 5973 6448
rect 6070 6488 6112 6497
rect 6070 6448 6071 6488
rect 6111 6448 6112 6488
rect 6070 6439 6112 6448
rect 6411 6488 6453 6497
rect 6411 6448 6412 6488
rect 6452 6448 6453 6488
rect 6411 6439 6453 6448
rect 6526 6488 6568 6497
rect 6526 6448 6527 6488
rect 6567 6448 6568 6488
rect 6526 6439 6568 6448
rect 6699 6488 6741 6497
rect 7377 6490 7419 6499
rect 6699 6448 6700 6488
rect 6740 6448 6741 6488
rect 6699 6439 6741 6448
rect 7258 6488 7316 6489
rect 7258 6448 7267 6488
rect 7307 6448 7316 6488
rect 7258 6447 7316 6448
rect 7377 6450 7378 6490
rect 7418 6450 7419 6490
rect 7377 6441 7419 6450
rect 7810 6488 7868 6489
rect 7810 6448 7819 6488
rect 7859 6448 7868 6488
rect 7810 6447 7868 6448
rect 8043 6488 8085 6497
rect 8043 6448 8044 6488
rect 8084 6448 8085 6488
rect 8043 6439 8085 6448
rect 8331 6488 8373 6497
rect 8331 6448 8332 6488
rect 8372 6448 8373 6488
rect 8331 6439 8373 6448
rect 8715 6488 8757 6497
rect 8715 6448 8716 6488
rect 8756 6448 8757 6488
rect 8715 6439 8757 6448
rect 9387 6488 9429 6497
rect 9387 6448 9388 6488
rect 9428 6448 9429 6488
rect 9387 6439 9429 6448
rect 9514 6488 9572 6489
rect 9514 6448 9523 6488
rect 9563 6448 9572 6488
rect 9514 6447 9572 6448
rect 10011 6488 10053 6497
rect 10011 6448 10012 6488
rect 10052 6448 10053 6488
rect 10011 6439 10053 6448
rect 10155 6488 10197 6497
rect 10155 6448 10156 6488
rect 10196 6448 10197 6488
rect 10155 6439 10197 6448
rect 10582 6488 10624 6497
rect 10582 6448 10583 6488
rect 10623 6448 10624 6488
rect 10582 6439 10624 6448
rect 10827 6488 10869 6497
rect 10827 6448 10828 6488
rect 10868 6448 10869 6488
rect 10827 6439 10869 6448
rect 11386 6488 11444 6489
rect 11386 6448 11395 6488
rect 11435 6448 11444 6488
rect 11386 6447 11444 6448
rect 11499 6488 11541 6497
rect 11499 6448 11500 6488
rect 11540 6448 11541 6488
rect 11499 6439 11541 6448
rect 11926 6488 11968 6497
rect 11926 6448 11927 6488
rect 11967 6448 11968 6488
rect 11926 6439 11968 6448
rect 12171 6488 12213 6497
rect 12171 6448 12172 6488
rect 12212 6448 12213 6488
rect 12171 6439 12213 6448
rect 12843 6488 12885 6497
rect 12843 6448 12844 6488
rect 12884 6448 12885 6488
rect 12843 6439 12885 6448
rect 13131 6488 13173 6497
rect 13131 6448 13132 6488
rect 13172 6448 13173 6488
rect 13131 6439 13173 6448
rect 13594 6488 13652 6489
rect 13594 6448 13603 6488
rect 13643 6448 13652 6488
rect 13594 6447 13652 6448
rect 13707 6488 13749 6497
rect 13707 6448 13708 6488
rect 13748 6448 13749 6488
rect 13707 6439 13749 6448
rect 14038 6488 14080 6497
rect 14038 6448 14039 6488
rect 14079 6448 14080 6488
rect 14038 6439 14080 6448
rect 14283 6488 14325 6497
rect 14283 6448 14284 6488
rect 14324 6448 14325 6488
rect 14283 6439 14325 6448
rect 15037 6488 15079 6497
rect 15706 6488 15764 6489
rect 15037 6448 15038 6488
rect 15078 6448 15079 6488
rect 15037 6439 15079 6448
rect 15339 6479 15381 6488
rect 15339 6439 15340 6479
rect 15380 6439 15381 6479
rect 15706 6448 15715 6488
rect 15755 6448 15764 6488
rect 15706 6447 15764 6448
rect 15819 6488 15861 6497
rect 15819 6448 15820 6488
rect 15860 6448 15861 6488
rect 15819 6439 15861 6448
rect 16299 6488 16341 6497
rect 16299 6448 16300 6488
rect 16340 6448 16341 6488
rect 16299 6439 16341 6448
rect 16683 6488 16725 6497
rect 16683 6448 16684 6488
rect 16724 6448 16725 6488
rect 16683 6439 16725 6448
rect 17163 6488 17205 6497
rect 17163 6448 17164 6488
rect 17204 6448 17205 6488
rect 17163 6439 17205 6448
rect 17392 6488 17450 6489
rect 17392 6448 17401 6488
rect 17441 6448 17450 6488
rect 17392 6447 17450 6448
rect 17931 6488 17973 6497
rect 17931 6448 17932 6488
rect 17972 6448 17973 6488
rect 17931 6439 17973 6448
rect 18315 6488 18357 6497
rect 18315 6448 18316 6488
rect 18356 6448 18357 6488
rect 18315 6439 18357 6448
rect 19467 6488 19509 6497
rect 19467 6448 19468 6488
rect 19508 6448 19509 6488
rect 19467 6439 19509 6448
rect 20124 6488 20166 6497
rect 20124 6448 20125 6488
rect 20165 6448 20166 6488
rect 20124 6439 20166 6448
rect 20235 6488 20277 6497
rect 20235 6448 20236 6488
rect 20276 6448 20277 6488
rect 20235 6439 20277 6448
rect 20662 6488 20704 6497
rect 20662 6448 20663 6488
rect 20703 6448 20704 6488
rect 20662 6439 20704 6448
rect 20907 6488 20949 6497
rect 20907 6448 20908 6488
rect 20948 6448 20949 6488
rect 20907 6439 20949 6448
rect 21195 6488 21237 6497
rect 21195 6448 21196 6488
rect 21236 6448 21237 6488
rect 21195 6439 21237 6448
rect 21370 6488 21428 6489
rect 21370 6448 21379 6488
rect 21419 6448 21428 6488
rect 21370 6447 21428 6448
rect 21483 6488 21525 6497
rect 21483 6448 21484 6488
rect 21524 6448 21525 6488
rect 21483 6439 21525 6448
rect 21915 6488 21973 6489
rect 21915 6448 21924 6488
rect 21964 6448 21973 6488
rect 21915 6447 21973 6448
rect 22059 6488 22101 6497
rect 22059 6448 22060 6488
rect 22100 6448 22101 6488
rect 22059 6439 22101 6448
rect 22347 6488 22389 6497
rect 22347 6448 22348 6488
rect 22388 6448 22389 6488
rect 22347 6439 22389 6448
rect 23595 6488 23637 6497
rect 23595 6448 23596 6488
rect 23636 6448 23637 6488
rect 23595 6439 23637 6448
rect 23776 6488 23818 6497
rect 24262 6488 24304 6497
rect 23776 6448 23777 6488
rect 23817 6448 23818 6488
rect 23776 6439 23818 6448
rect 24075 6479 24117 6488
rect 24075 6439 24076 6479
rect 24116 6439 24117 6479
rect 24262 6448 24263 6488
rect 24303 6448 24304 6488
rect 24262 6439 24304 6448
rect 24442 6488 24500 6489
rect 24442 6448 24451 6488
rect 24491 6448 24500 6488
rect 24442 6447 24500 6448
rect 15339 6430 15381 6439
rect 24075 6430 24117 6439
rect 2283 6404 2325 6413
rect 5386 6404 5444 6405
rect 2283 6364 2284 6404
rect 2324 6364 2325 6404
rect 2283 6355 2325 6364
rect 2514 6395 2560 6404
rect 2514 6355 2515 6395
rect 2555 6355 2560 6395
rect 5386 6364 5395 6404
rect 5435 6364 5444 6404
rect 5386 6363 5444 6364
rect 7930 6404 7988 6405
rect 7930 6364 7939 6404
rect 7979 6364 7988 6404
rect 7930 6363 7988 6364
rect 10714 6404 10772 6405
rect 10714 6364 10723 6404
rect 10763 6364 10772 6404
rect 10714 6363 10772 6364
rect 10923 6404 10965 6413
rect 10923 6364 10924 6404
rect 10964 6364 10965 6404
rect 10923 6355 10965 6364
rect 12058 6404 12116 6405
rect 12058 6364 12067 6404
rect 12107 6364 12116 6404
rect 12058 6363 12116 6364
rect 14170 6404 14228 6405
rect 14170 6364 14179 6404
rect 14219 6364 14228 6404
rect 14170 6363 14228 6364
rect 14379 6404 14421 6413
rect 14379 6364 14380 6404
rect 14420 6364 14421 6404
rect 14379 6355 14421 6364
rect 17067 6404 17109 6413
rect 17067 6364 17068 6404
rect 17108 6364 17109 6404
rect 17067 6355 17109 6364
rect 17282 6404 17324 6413
rect 17282 6364 17283 6404
rect 17323 6364 17324 6404
rect 17282 6355 17324 6364
rect 19377 6404 19419 6413
rect 19377 6364 19378 6404
rect 19418 6364 19419 6404
rect 19377 6355 19419 6364
rect 20794 6404 20852 6405
rect 20794 6364 20803 6404
rect 20843 6364 20852 6404
rect 20794 6363 20852 6364
rect 2514 6346 2560 6355
rect 15994 6320 16052 6321
rect 15994 6280 16003 6320
rect 16043 6280 16052 6320
rect 15994 6279 16052 6280
rect 21291 6320 21333 6329
rect 21291 6280 21292 6320
rect 21332 6280 21333 6320
rect 21291 6271 21333 6280
rect 22539 6320 22581 6329
rect 22539 6280 22540 6320
rect 22580 6280 22581 6320
rect 22539 6271 22581 6280
rect 4683 6236 4725 6245
rect 4683 6196 4684 6236
rect 4724 6196 4725 6236
rect 4683 6187 4725 6196
rect 6411 6236 6453 6245
rect 6411 6196 6412 6236
rect 6452 6196 6453 6236
rect 6411 6187 6453 6196
rect 13899 6236 13941 6245
rect 13899 6196 13900 6236
rect 13940 6196 13941 6236
rect 13899 6187 13941 6196
rect 15034 6236 15092 6237
rect 15034 6196 15043 6236
rect 15083 6196 15092 6236
rect 15034 6195 15092 6196
rect 18555 6236 18597 6245
rect 18555 6196 18556 6236
rect 18596 6196 18597 6236
rect 18555 6187 18597 6196
rect 22923 6236 22965 6245
rect 22923 6196 22924 6236
rect 22964 6196 22965 6236
rect 22923 6187 22965 6196
rect 24442 6236 24500 6237
rect 24442 6196 24451 6236
rect 24491 6196 24500 6236
rect 24442 6195 24500 6196
rect 576 6068 31392 6092
rect 576 6028 3112 6068
rect 3480 6028 10886 6068
rect 11254 6028 18660 6068
rect 19028 6028 26434 6068
rect 26802 6028 31392 6068
rect 576 6004 31392 6028
rect 5739 5900 5781 5909
rect 5739 5860 5740 5900
rect 5780 5860 5781 5900
rect 5739 5851 5781 5860
rect 9675 5900 9717 5909
rect 9675 5860 9676 5900
rect 9716 5860 9717 5900
rect 9675 5851 9717 5860
rect 14379 5900 14421 5909
rect 14379 5860 14380 5900
rect 14420 5860 14421 5900
rect 14379 5851 14421 5860
rect 15034 5900 15092 5901
rect 15034 5860 15043 5900
rect 15083 5860 15092 5900
rect 15034 5859 15092 5860
rect 20602 5900 20660 5901
rect 20602 5860 20611 5900
rect 20651 5860 20660 5900
rect 20602 5859 20660 5860
rect 20907 5900 20949 5909
rect 20907 5860 20908 5900
rect 20948 5860 20949 5900
rect 20907 5851 20949 5860
rect 23211 5900 23253 5909
rect 23211 5860 23212 5900
rect 23252 5860 23253 5900
rect 23211 5851 23253 5860
rect 23595 5900 23637 5909
rect 23595 5860 23596 5900
rect 23636 5860 23637 5900
rect 23595 5851 23637 5860
rect 4875 5816 4917 5825
rect 4875 5776 4876 5816
rect 4916 5776 4917 5816
rect 4875 5767 4917 5776
rect 9003 5816 9045 5825
rect 9003 5776 9004 5816
rect 9044 5776 9045 5816
rect 9003 5767 9045 5776
rect 13419 5816 13461 5825
rect 13419 5776 13420 5816
rect 13460 5776 13461 5816
rect 13419 5767 13461 5776
rect 23787 5816 23829 5825
rect 23787 5776 23788 5816
rect 23828 5776 23829 5816
rect 23787 5767 23829 5776
rect 6699 5732 6741 5741
rect 6699 5692 6700 5732
rect 6740 5692 6741 5732
rect 6699 5683 6741 5692
rect 10658 5732 10700 5741
rect 10658 5692 10659 5732
rect 10699 5692 10700 5732
rect 10658 5683 10700 5692
rect 21291 5732 21333 5741
rect 21291 5692 21292 5732
rect 21332 5692 21333 5732
rect 21291 5683 21333 5692
rect 2461 5648 2503 5657
rect 2461 5608 2462 5648
rect 2502 5608 2503 5648
rect 2461 5599 2503 5608
rect 2755 5648 2813 5649
rect 2755 5608 2764 5648
rect 2804 5608 2813 5648
rect 2755 5607 2813 5608
rect 2938 5648 2996 5649
rect 2938 5608 2947 5648
rect 2987 5608 2996 5648
rect 2938 5607 2996 5608
rect 3627 5648 3669 5657
rect 3627 5608 3628 5648
rect 3668 5608 3669 5648
rect 3627 5599 3669 5608
rect 3898 5648 3956 5649
rect 3898 5608 3907 5648
rect 3947 5608 3956 5648
rect 3898 5607 3956 5608
rect 4562 5648 4604 5657
rect 4562 5608 4563 5648
rect 4603 5608 4604 5648
rect 4562 5599 4604 5608
rect 4674 5648 4732 5649
rect 4674 5608 4683 5648
rect 4723 5608 4732 5648
rect 4674 5607 4732 5608
rect 5067 5648 5109 5657
rect 5067 5608 5068 5648
rect 5108 5608 5109 5648
rect 5067 5599 5109 5608
rect 6106 5648 6164 5649
rect 6106 5608 6115 5648
rect 6155 5608 6164 5648
rect 6106 5607 6164 5608
rect 6219 5648 6261 5657
rect 6219 5608 6220 5648
rect 6260 5608 6261 5648
rect 6219 5599 6261 5608
rect 6603 5648 6645 5657
rect 6603 5608 6604 5648
rect 6644 5608 6645 5648
rect 6603 5599 6645 5608
rect 6795 5648 6837 5657
rect 6795 5608 6796 5648
rect 6836 5608 6837 5648
rect 6795 5599 6837 5608
rect 7114 5648 7172 5649
rect 7114 5608 7123 5648
rect 7163 5608 7172 5648
rect 7114 5607 7172 5608
rect 7309 5648 7367 5649
rect 7309 5608 7318 5648
rect 7358 5608 7367 5648
rect 7309 5607 7367 5608
rect 7450 5648 7508 5649
rect 7450 5608 7459 5648
rect 7499 5608 7508 5648
rect 7450 5607 7508 5608
rect 8139 5648 8181 5657
rect 8139 5608 8140 5648
rect 8180 5608 8181 5648
rect 8139 5599 8181 5608
rect 8619 5648 8661 5657
rect 8619 5608 8620 5648
rect 8660 5608 8661 5648
rect 8619 5599 8661 5608
rect 9370 5648 9428 5649
rect 9370 5608 9379 5648
rect 9419 5608 9428 5648
rect 9370 5607 9428 5608
rect 10059 5648 10101 5657
rect 10059 5608 10060 5648
rect 10100 5608 10101 5648
rect 10059 5599 10101 5608
rect 10539 5648 10581 5657
rect 10539 5608 10540 5648
rect 10580 5608 10581 5648
rect 10539 5599 10581 5608
rect 10768 5648 10826 5649
rect 10768 5608 10777 5648
rect 10817 5608 10826 5648
rect 10768 5607 10826 5608
rect 11098 5648 11156 5649
rect 11098 5608 11107 5648
rect 11147 5608 11156 5648
rect 11098 5607 11156 5608
rect 11211 5648 11253 5657
rect 11211 5608 11212 5648
rect 11252 5608 11253 5648
rect 11211 5599 11253 5608
rect 11643 5648 11685 5657
rect 11643 5608 11644 5648
rect 11684 5608 11685 5648
rect 11643 5599 11685 5608
rect 11825 5648 11883 5649
rect 11825 5608 11834 5648
rect 11874 5608 11883 5648
rect 11825 5607 11883 5608
rect 12171 5648 12213 5657
rect 12171 5608 12172 5648
rect 12212 5608 12213 5648
rect 12171 5599 12213 5608
rect 12555 5648 12597 5657
rect 13143 5655 13185 5664
rect 12555 5608 12556 5648
rect 12596 5608 12597 5648
rect 12555 5599 12597 5608
rect 13018 5648 13076 5649
rect 13018 5608 13027 5648
rect 13067 5608 13076 5648
rect 13018 5607 13076 5608
rect 13143 5615 13144 5655
rect 13184 5615 13185 5655
rect 13143 5606 13185 5615
rect 13803 5648 13845 5657
rect 13803 5608 13804 5648
rect 13844 5608 13845 5648
rect 13803 5599 13845 5608
rect 14074 5648 14132 5649
rect 14074 5608 14083 5648
rect 14123 5608 14132 5648
rect 14074 5607 14132 5608
rect 14379 5648 14421 5657
rect 14379 5608 14380 5648
rect 14420 5608 14421 5648
rect 14379 5599 14421 5608
rect 14746 5648 14804 5649
rect 14746 5608 14755 5648
rect 14795 5608 14804 5648
rect 14746 5607 14804 5608
rect 14859 5648 14901 5657
rect 14859 5608 14860 5648
rect 14900 5608 14901 5648
rect 14859 5599 14901 5608
rect 15483 5648 15525 5657
rect 15483 5608 15484 5648
rect 15524 5608 15525 5648
rect 15483 5599 15525 5608
rect 15627 5648 15669 5657
rect 15627 5608 15628 5648
rect 15668 5608 15669 5648
rect 15627 5599 15669 5608
rect 16203 5648 16245 5657
rect 16203 5608 16204 5648
rect 16244 5608 16245 5648
rect 16203 5599 16245 5608
rect 16322 5648 16364 5657
rect 16322 5608 16323 5648
rect 16363 5608 16364 5648
rect 16322 5599 16364 5608
rect 16432 5648 16490 5649
rect 16432 5608 16441 5648
rect 16481 5608 16490 5648
rect 16432 5607 16490 5608
rect 16683 5648 16725 5657
rect 16683 5608 16684 5648
rect 16724 5608 16725 5648
rect 16683 5599 16725 5608
rect 17067 5648 17109 5657
rect 17067 5608 17068 5648
rect 17108 5608 17109 5648
rect 17067 5599 17109 5608
rect 17626 5648 17684 5649
rect 17626 5608 17635 5648
rect 17675 5608 17684 5648
rect 17626 5607 17684 5608
rect 17739 5648 17781 5657
rect 17739 5608 17740 5648
rect 17780 5608 17781 5648
rect 17739 5599 17781 5608
rect 18411 5648 18453 5657
rect 18411 5608 18412 5648
rect 18452 5608 18453 5648
rect 18411 5599 18453 5608
rect 18795 5648 18837 5657
rect 18795 5608 18796 5648
rect 18836 5608 18837 5648
rect 18795 5599 18837 5608
rect 19179 5648 19221 5657
rect 19179 5608 19180 5648
rect 19220 5608 19221 5648
rect 19179 5599 19221 5608
rect 19563 5648 19605 5657
rect 19563 5608 19564 5648
rect 19604 5608 19605 5648
rect 19563 5599 19605 5608
rect 20427 5648 20469 5657
rect 20427 5608 20428 5648
rect 20468 5608 20469 5648
rect 20427 5599 20469 5608
rect 20602 5648 20660 5649
rect 20602 5608 20611 5648
rect 20651 5608 20660 5648
rect 20602 5607 20660 5608
rect 20811 5648 20853 5657
rect 20811 5608 20812 5648
rect 20852 5608 20853 5648
rect 20811 5599 20853 5608
rect 21003 5648 21045 5657
rect 21003 5608 21004 5648
rect 21044 5608 21045 5648
rect 21003 5599 21045 5608
rect 21658 5648 21716 5649
rect 21658 5608 21667 5648
rect 21707 5608 21716 5648
rect 21658 5607 21716 5608
rect 2554 5564 2612 5565
rect 2554 5524 2563 5564
rect 2603 5524 2612 5564
rect 2554 5523 2612 5524
rect 4107 5564 4149 5573
rect 4107 5524 4108 5564
rect 4148 5524 4149 5564
rect 4107 5515 4149 5524
rect 4217 5564 4259 5573
rect 4217 5524 4218 5564
rect 4258 5524 4259 5564
rect 4217 5515 4259 5524
rect 6394 5564 6452 5565
rect 6394 5524 6403 5564
rect 6443 5524 6452 5564
rect 6394 5523 6452 5524
rect 9483 5564 9525 5573
rect 9483 5524 9484 5564
rect 9524 5524 9525 5564
rect 9483 5515 9525 5524
rect 9689 5564 9731 5573
rect 9689 5524 9690 5564
rect 9730 5524 9731 5564
rect 9689 5515 9731 5524
rect 9850 5564 9908 5565
rect 9850 5524 9859 5564
rect 9899 5524 9908 5564
rect 9850 5523 9908 5524
rect 10443 5564 10485 5573
rect 10443 5524 10444 5564
rect 10484 5524 10485 5564
rect 10443 5515 10485 5524
rect 2667 5480 2709 5489
rect 2667 5440 2668 5480
rect 2708 5440 2709 5480
rect 2667 5431 2709 5440
rect 3994 5480 4052 5481
rect 3994 5440 4003 5480
rect 4043 5440 4052 5480
rect 3994 5439 4052 5440
rect 4587 5480 4629 5489
rect 4587 5440 4588 5480
rect 4628 5440 4629 5480
rect 4587 5431 4629 5440
rect 6123 5480 6165 5489
rect 6123 5440 6124 5480
rect 6164 5440 6165 5480
rect 6123 5431 6165 5440
rect 8506 5480 8564 5481
rect 8506 5440 8515 5480
rect 8555 5440 8564 5480
rect 8506 5439 8564 5440
rect 8811 5480 8853 5489
rect 8811 5440 8812 5480
rect 8852 5440 8853 5480
rect 8811 5431 8853 5440
rect 10138 5480 10196 5481
rect 10138 5440 10147 5480
rect 10187 5440 10196 5480
rect 10138 5439 10196 5440
rect 11499 5480 11541 5489
rect 11499 5440 11500 5480
rect 11540 5440 11541 5480
rect 11499 5431 11541 5440
rect 11979 5480 12021 5489
rect 11979 5440 11980 5480
rect 12020 5440 12021 5480
rect 11979 5431 12021 5440
rect 12651 5480 12693 5489
rect 13611 5480 13653 5489
rect 12651 5440 12652 5480
rect 12692 5440 12693 5480
rect 12651 5431 12693 5440
rect 12930 5471 12976 5480
rect 12930 5431 12931 5471
rect 12971 5431 12976 5471
rect 13611 5440 13612 5480
rect 13652 5440 13653 5480
rect 13611 5431 13653 5440
rect 13882 5480 13940 5481
rect 13882 5440 13891 5480
rect 13931 5440 13940 5480
rect 13882 5439 13940 5440
rect 15322 5480 15380 5481
rect 15322 5440 15331 5480
rect 15371 5440 15380 5480
rect 15322 5439 15380 5440
rect 16107 5480 16149 5489
rect 16107 5440 16108 5480
rect 16148 5440 16149 5480
rect 16107 5431 16149 5440
rect 17163 5480 17205 5489
rect 17163 5440 17164 5480
rect 17204 5440 17205 5480
rect 17163 5431 17205 5440
rect 18027 5480 18069 5489
rect 18027 5440 18028 5480
rect 18068 5440 18069 5480
rect 18027 5431 18069 5440
rect 18298 5480 18356 5481
rect 18298 5440 18307 5480
rect 18347 5440 18356 5480
rect 18298 5439 18356 5440
rect 18987 5480 19029 5489
rect 18987 5440 18988 5480
rect 19028 5440 19029 5480
rect 18987 5431 19029 5440
rect 19258 5480 19316 5481
rect 19258 5440 19267 5480
rect 19307 5440 19316 5480
rect 19258 5439 19316 5440
rect 20235 5480 20277 5489
rect 20235 5440 20236 5480
rect 20276 5440 20277 5480
rect 20235 5431 20277 5440
rect 12930 5422 12976 5431
rect 576 5312 31392 5336
rect 576 5272 4352 5312
rect 4720 5272 12126 5312
rect 12494 5272 19900 5312
rect 20268 5272 27674 5312
rect 28042 5272 31392 5312
rect 576 5248 31392 5272
rect 7371 5144 7413 5153
rect 7371 5104 7372 5144
rect 7412 5104 7413 5144
rect 7371 5095 7413 5104
rect 10347 5144 10389 5153
rect 10347 5104 10348 5144
rect 10388 5104 10389 5144
rect 10347 5095 10389 5104
rect 11386 5144 11444 5145
rect 11386 5104 11395 5144
rect 11435 5104 11444 5144
rect 11386 5103 11444 5104
rect 12250 5144 12308 5145
rect 12250 5104 12259 5144
rect 12299 5104 12308 5144
rect 12250 5103 12308 5104
rect 12555 5144 12597 5153
rect 12555 5104 12556 5144
rect 12596 5104 12597 5144
rect 12555 5095 12597 5104
rect 15531 5144 15573 5153
rect 15531 5104 15532 5144
rect 15572 5104 15573 5144
rect 15531 5095 15573 5104
rect 18411 5144 18453 5153
rect 18411 5104 18412 5144
rect 18452 5104 18453 5144
rect 18411 5095 18453 5104
rect 18682 5144 18740 5145
rect 18682 5104 18691 5144
rect 18731 5104 18740 5144
rect 18682 5103 18740 5104
rect 21435 5144 21477 5153
rect 21435 5104 21436 5144
rect 21476 5104 21477 5144
rect 21435 5095 21477 5104
rect 21867 5144 21909 5153
rect 21867 5104 21868 5144
rect 21908 5104 21909 5144
rect 21867 5095 21909 5104
rect 22251 5144 22293 5153
rect 22251 5104 22252 5144
rect 22292 5104 22293 5144
rect 22251 5095 22293 5104
rect 5050 5060 5108 5061
rect 5050 5020 5059 5060
rect 5099 5020 5108 5060
rect 5050 5019 5108 5020
rect 12826 5060 12884 5061
rect 12826 5020 12835 5060
rect 12875 5020 12884 5060
rect 12826 5019 12884 5020
rect 13210 5060 13268 5061
rect 13210 5020 13219 5060
rect 13259 5020 13268 5060
rect 13210 5019 13268 5020
rect 18905 5060 18947 5069
rect 18905 5020 18906 5060
rect 18946 5020 18947 5060
rect 18905 5011 18947 5020
rect 21977 5060 22019 5069
rect 21977 5020 21978 5060
rect 22018 5020 22019 5060
rect 21977 5011 22019 5020
rect 5434 4976 5492 4977
rect 8410 4976 8468 4977
rect 5434 4936 5443 4976
rect 5483 4936 5492 4976
rect 5434 4935 5492 4936
rect 7554 4967 7600 4976
rect 7554 4927 7555 4967
rect 7595 4927 7600 4967
rect 8410 4936 8419 4976
rect 8459 4936 8468 4976
rect 8410 4935 8468 4936
rect 11211 4976 11253 4985
rect 11211 4936 11212 4976
rect 11252 4936 11253 4976
rect 11211 4927 11253 4936
rect 11691 4976 11733 4985
rect 11691 4936 11692 4976
rect 11732 4936 11733 4976
rect 11691 4927 11733 4936
rect 12363 4976 12405 4985
rect 12363 4936 12364 4976
rect 12404 4936 12405 4976
rect 12363 4927 12405 4936
rect 12737 4976 12779 4985
rect 12737 4936 12738 4976
rect 12778 4936 12779 4976
rect 12737 4927 12779 4936
rect 12922 4976 12980 4977
rect 12922 4936 12931 4976
rect 12971 4936 12980 4976
rect 12922 4935 12980 4936
rect 13035 4976 13077 4985
rect 13035 4936 13036 4976
rect 13076 4936 13077 4976
rect 13035 4927 13077 4936
rect 13594 4976 13652 4977
rect 13594 4936 13603 4976
rect 13643 4936 13652 4976
rect 13594 4935 13652 4936
rect 16474 4976 16532 4977
rect 16474 4936 16483 4976
rect 16523 4936 16532 4976
rect 16474 4935 16532 4936
rect 18586 4976 18644 4977
rect 20907 4976 20949 4985
rect 18586 4936 18595 4976
rect 18635 4936 18644 4976
rect 18586 4935 18644 4936
rect 20130 4967 20176 4976
rect 20130 4927 20131 4967
rect 20171 4927 20176 4967
rect 20907 4936 20908 4976
rect 20948 4936 20949 4976
rect 20907 4927 20949 4936
rect 21103 4976 21145 4985
rect 21103 4936 21104 4976
rect 21144 4936 21145 4976
rect 21103 4927 21145 4936
rect 21291 4976 21333 4985
rect 21291 4936 21292 4976
rect 21332 4936 21333 4976
rect 21291 4927 21333 4936
rect 21658 4976 21716 4977
rect 21658 4936 21667 4976
rect 21707 4936 21716 4976
rect 21658 4935 21716 4936
rect 21771 4976 21813 4985
rect 21771 4936 21772 4976
rect 21812 4936 21813 4976
rect 21771 4927 21813 4936
rect 22155 4976 22197 4985
rect 22155 4936 22156 4976
rect 22196 4936 22197 4976
rect 22155 4927 22197 4936
rect 22347 4976 22389 4985
rect 22347 4936 22348 4976
rect 22388 4936 22389 4976
rect 22347 4927 22389 4936
rect 7554 4918 7600 4927
rect 20130 4918 20176 4927
rect 7707 4892 7749 4901
rect 7707 4852 7708 4892
rect 7748 4852 7749 4892
rect 7707 4843 7749 4852
rect 8043 4892 8085 4901
rect 8043 4852 8044 4892
rect 8084 4852 8085 4892
rect 8043 4843 8085 4852
rect 11601 4892 11643 4901
rect 11601 4852 11602 4892
rect 11642 4852 11643 4892
rect 11601 4843 11643 4852
rect 15147 4892 15189 4901
rect 15147 4852 15148 4892
rect 15188 4852 15189 4892
rect 15147 4843 15189 4852
rect 16107 4892 16149 4901
rect 16107 4852 16108 4892
rect 16148 4852 16149 4892
rect 16107 4843 16149 4852
rect 18027 4892 18069 4901
rect 18027 4852 18028 4892
rect 18068 4852 18069 4892
rect 18027 4843 18069 4852
rect 20283 4892 20325 4901
rect 20283 4852 20284 4892
rect 20324 4852 20325 4892
rect 20283 4843 20325 4852
rect 7371 4808 7413 4817
rect 7371 4768 7372 4808
rect 7412 4768 7413 4808
rect 7371 4759 7413 4768
rect 10539 4808 10581 4817
rect 10539 4768 10540 4808
rect 10580 4768 10581 4808
rect 10539 4759 10581 4768
rect 6987 4724 7029 4733
rect 6987 4684 6988 4724
rect 7028 4684 7029 4724
rect 6987 4675 7029 4684
rect 9963 4724 10005 4733
rect 9963 4684 9964 4724
rect 10004 4684 10005 4724
rect 9963 4675 10005 4684
rect 10347 4724 10389 4733
rect 10347 4684 10348 4724
rect 10388 4684 10389 4724
rect 10347 4675 10389 4684
rect 18891 4724 18933 4733
rect 18891 4684 18892 4724
rect 18932 4684 18933 4724
rect 18891 4675 18933 4684
rect 21003 4724 21045 4733
rect 21003 4684 21004 4724
rect 21044 4684 21045 4724
rect 21003 4675 21045 4684
rect 576 4556 31392 4580
rect 576 4516 3112 4556
rect 3480 4516 10886 4556
rect 11254 4516 18660 4556
rect 19028 4516 26434 4556
rect 26802 4516 31392 4556
rect 576 4492 31392 4516
rect 7851 4388 7893 4397
rect 7851 4348 7852 4388
rect 7892 4348 7893 4388
rect 7851 4339 7893 4348
rect 13227 4388 13269 4397
rect 13227 4348 13228 4388
rect 13268 4348 13269 4388
rect 13227 4339 13269 4348
rect 16107 4388 16149 4397
rect 16107 4348 16108 4388
rect 16148 4348 16149 4388
rect 16107 4339 16149 4348
rect 6219 4304 6261 4313
rect 6219 4264 6220 4304
rect 6260 4264 6261 4304
rect 6219 4255 6261 4264
rect 8475 4304 8517 4313
rect 8475 4264 8476 4304
rect 8516 4264 8517 4304
rect 8475 4255 8517 4264
rect 11787 4304 11829 4313
rect 11787 4264 11788 4304
rect 11828 4264 11829 4304
rect 11787 4255 11829 4264
rect 13707 4304 13749 4313
rect 13707 4264 13708 4304
rect 13748 4264 13749 4304
rect 13707 4255 13749 4264
rect 14475 4304 14517 4313
rect 14475 4264 14476 4304
rect 14516 4264 14517 4304
rect 14475 4255 14517 4264
rect 17163 4304 17205 4313
rect 17163 4264 17164 4304
rect 17204 4264 17205 4304
rect 17163 4255 17205 4264
rect 8258 4220 8300 4229
rect 8258 4180 8259 4220
rect 8299 4180 8300 4220
rect 8258 4171 8300 4180
rect 9802 4220 9860 4221
rect 9802 4180 9811 4220
rect 9851 4180 9860 4220
rect 9802 4179 9860 4180
rect 10587 4220 10629 4229
rect 10587 4180 10588 4220
rect 10628 4180 10629 4220
rect 10587 4171 10629 4180
rect 15178 4220 15236 4221
rect 15178 4180 15187 4220
rect 15227 4180 15236 4220
rect 15178 4179 15236 4180
rect 7546 4136 7604 4137
rect 7546 4096 7555 4136
rect 7595 4096 7604 4136
rect 7546 4095 7604 4096
rect 8139 4136 8181 4145
rect 8139 4096 8140 4136
rect 8180 4096 8181 4136
rect 8139 4087 8181 4096
rect 8368 4136 8426 4137
rect 8368 4096 8377 4136
rect 8417 4096 8426 4136
rect 8368 4095 8426 4096
rect 8619 4136 8661 4145
rect 8619 4096 8620 4136
rect 8660 4096 8661 4136
rect 8619 4087 8661 4096
rect 9997 4136 10055 4137
rect 9997 4096 10006 4136
rect 10046 4096 10055 4136
rect 9997 4095 10055 4096
rect 10378 4136 10436 4137
rect 10378 4096 10387 4136
rect 10427 4096 10436 4136
rect 10378 4095 10436 4096
rect 11691 4136 11733 4145
rect 11691 4096 11692 4136
rect 11732 4096 11733 4136
rect 11691 4087 11733 4096
rect 11883 4136 11925 4145
rect 11883 4096 11884 4136
rect 11924 4096 11925 4136
rect 11883 4087 11925 4096
rect 13227 4136 13269 4145
rect 13227 4096 13228 4136
rect 13268 4096 13269 4136
rect 13227 4087 13269 4096
rect 13419 4136 13461 4145
rect 13419 4096 13420 4136
rect 13460 4096 13461 4136
rect 13419 4087 13461 4096
rect 13803 4136 13845 4145
rect 13803 4096 13804 4136
rect 13844 4096 13845 4136
rect 13803 4087 13845 4096
rect 14091 4136 14133 4145
rect 14091 4096 14092 4136
rect 14132 4096 14133 4136
rect 14091 4087 14133 4096
rect 15373 4136 15431 4137
rect 15373 4096 15382 4136
rect 15422 4096 15431 4136
rect 15373 4095 15431 4096
rect 15802 4136 15860 4137
rect 15802 4096 15811 4136
rect 15851 4096 15860 4136
rect 15802 4095 15860 4096
rect 16121 4136 16163 4145
rect 16121 4096 16122 4136
rect 16162 4096 16163 4136
rect 16121 4087 16163 4096
rect 7865 4052 7907 4061
rect 7865 4012 7866 4052
rect 7906 4012 7907 4052
rect 7865 4003 7907 4012
rect 8043 4052 8085 4061
rect 8043 4012 8044 4052
rect 8084 4012 8085 4052
rect 8043 4003 8085 4012
rect 15915 4052 15957 4061
rect 15915 4012 15916 4052
rect 15956 4012 15957 4052
rect 15915 4003 15957 4012
rect 7642 3968 7700 3969
rect 7642 3928 7651 3968
rect 7691 3928 7700 3968
rect 7642 3927 7700 3928
rect 13707 3968 13749 3977
rect 13707 3928 13708 3968
rect 13748 3928 13749 3968
rect 13707 3919 13749 3928
rect 13978 3968 14036 3969
rect 13978 3928 13987 3968
rect 14027 3928 14036 3968
rect 13978 3927 14036 3928
rect 14283 3968 14325 3977
rect 14283 3928 14284 3968
rect 14324 3928 14325 3968
rect 14283 3919 14325 3928
rect 576 3800 31392 3824
rect 576 3760 4352 3800
rect 4720 3760 12126 3800
rect 12494 3760 19900 3800
rect 20268 3760 27674 3800
rect 28042 3760 31392 3800
rect 576 3736 31392 3760
rect 576 3044 31392 3068
rect 576 3004 3112 3044
rect 3480 3004 10886 3044
rect 11254 3004 18660 3044
rect 19028 3004 26434 3044
rect 26802 3004 31392 3044
rect 576 2980 31392 3004
rect 576 2288 31392 2312
rect 576 2248 4352 2288
rect 4720 2248 12126 2288
rect 12494 2248 19900 2288
rect 20268 2248 27674 2288
rect 28042 2248 31392 2288
rect 576 2224 31392 2248
rect 576 1532 31392 1556
rect 576 1492 3112 1532
rect 3480 1492 10886 1532
rect 11254 1492 18660 1532
rect 19028 1492 26434 1532
rect 26802 1492 31392 1532
rect 576 1468 31392 1492
rect 576 776 31392 800
rect 576 736 4352 776
rect 4720 736 12126 776
rect 12494 736 19900 776
rect 20268 736 27674 776
rect 28042 736 31392 776
rect 576 712 31392 736
<< via1 >>
rect 4352 27952 4720 27992
rect 12126 27952 12494 27992
rect 19900 27952 20268 27992
rect 27674 27952 28042 27992
rect 844 27784 884 27824
rect 1612 27784 1652 27824
rect 17740 27784 17780 27824
rect 17980 27784 18020 27824
rect 30307 27784 30347 27824
rect 1900 27700 1940 27740
rect 3715 27700 3755 27740
rect 4579 27700 4619 27740
rect 12163 27700 12203 27740
rect 14467 27700 14507 27740
rect 1804 27616 1844 27656
rect 1987 27616 2027 27656
rect 2195 27616 2235 27656
rect 2371 27616 2411 27656
rect 2951 27616 2991 27656
rect 3139 27616 3179 27656
rect 4396 27616 4436 27656
rect 4963 27616 5003 27656
rect 7459 27616 7499 27656
rect 9955 27616 9995 27656
rect 14083 27616 14123 27656
rect 15427 27616 15467 27656
rect 17534 27616 17574 27656
rect 17836 27607 17876 27647
rect 18124 27616 18164 27656
rect 18316 27616 18356 27656
rect 19555 27616 19595 27656
rect 22339 27616 22379 27656
rect 26371 27616 26411 27656
rect 26755 27616 26795 27656
rect 27331 27616 27371 27656
rect 30124 27616 30164 27656
rect 30460 27616 30500 27656
rect 30604 27616 30644 27656
rect 30787 27607 30827 27647
rect 7084 27532 7124 27572
rect 9580 27532 9620 27572
rect 15052 27532 15092 27572
rect 18988 27532 19028 27572
rect 19180 27532 19220 27572
rect 21964 27532 22004 27572
rect 26956 27532 26996 27572
rect 30940 27532 30980 27572
rect 1228 27448 1268 27488
rect 2371 27448 2411 27488
rect 2764 27448 2804 27488
rect 3532 27448 3572 27488
rect 14860 27448 14900 27488
rect 17356 27448 17396 27488
rect 3139 27364 3179 27404
rect 6892 27364 6932 27404
rect 9388 27364 9428 27404
rect 11884 27364 11924 27404
rect 17539 27364 17579 27404
rect 21484 27364 21524 27404
rect 24268 27364 24308 27404
rect 24460 27364 24500 27404
rect 29260 27364 29300 27404
rect 29452 27364 29492 27404
rect 3112 27196 3480 27236
rect 10886 27196 11254 27236
rect 18660 27196 19028 27236
rect 26434 27196 26802 27236
rect 2092 27028 2132 27068
rect 2659 27028 2699 27068
rect 6691 27028 6731 27068
rect 7939 27028 7979 27068
rect 9859 27028 9899 27068
rect 12076 27028 12116 27068
rect 14956 27028 14996 27068
rect 19180 27028 19220 27068
rect 22924 27028 22964 27068
rect 26380 27028 26420 27068
rect 28300 27028 28340 27068
rect 1132 26944 1172 26984
rect 6508 26944 6548 26984
rect 11116 26944 11156 26984
rect 12748 26944 12788 26984
rect 13420 26944 13460 26984
rect 15628 26944 15668 26984
rect 3235 26860 3275 26900
rect 7756 26860 7796 26900
rect 13516 26860 13556 26900
rect 20611 26860 20651 26900
rect 2092 26776 2132 26816
rect 2284 26776 2324 26816
rect 2476 26776 2516 26816
rect 2659 26776 2699 26816
rect 4771 26776 4811 26816
rect 5155 26776 5195 26816
rect 5548 26776 5588 26816
rect 5644 26776 5684 26816
rect 5884 26776 5924 26816
rect 6976 26809 7016 26849
rect 7075 26776 7115 26816
rect 8140 26776 8180 26816
rect 8236 26776 8276 26816
rect 8620 26776 8660 26816
rect 8716 26776 8756 26816
rect 8908 26776 8948 26816
rect 10156 26776 10196 26816
rect 10444 26776 10484 26816
rect 10924 26776 10964 26816
rect 11404 26776 11444 26816
rect 11788 26776 11828 26816
rect 11910 26776 11950 26816
rect 12037 26776 12077 26816
rect 12259 26776 12299 26816
rect 12940 26776 12980 26816
rect 13197 26776 13237 26816
rect 13345 26776 13385 26816
rect 13651 26776 13691 26816
rect 13804 26776 13844 26816
rect 14755 26776 14795 26816
rect 15820 26776 15860 26816
rect 17059 26776 17099 26816
rect 19468 26776 19508 26816
rect 19564 26767 19604 26807
rect 19852 26776 19892 26816
rect 20332 26776 20372 26816
rect 21292 26776 21332 26816
rect 21527 26776 21567 26816
rect 21667 26776 21707 26816
rect 21772 26776 21812 26816
rect 22732 26776 22772 26816
rect 23596 26776 23636 26816
rect 24460 26776 24500 26816
rect 25324 26776 25364 26816
rect 26188 26776 26228 26816
rect 27052 26776 27092 26816
rect 27916 26776 27956 26816
rect 30211 26776 30251 26816
rect 30892 26776 30932 26816
rect 5342 26692 5382 26732
rect 7934 26692 7974 26732
rect 8414 26692 8454 26732
rect 9854 26692 9894 26732
rect 12570 26692 12610 26732
rect 15043 26692 15083 26732
rect 16492 26692 16532 26732
rect 16675 26692 16715 26732
rect 21859 26692 21899 26732
rect 25507 26692 25547 26732
rect 30595 26692 30635 26732
rect 1516 26608 1556 26648
rect 1900 26608 1940 26648
rect 2860 26608 2900 26648
rect 5443 26608 5483 26648
rect 7516 26608 7556 26648
rect 7219 26566 7259 26606
rect 8140 26608 8180 26648
rect 8515 26608 8555 26648
rect 9580 26608 9620 26648
rect 10060 26608 10100 26648
rect 10339 26608 10379 26648
rect 10636 26608 10676 26648
rect 10819 26608 10859 26648
rect 11299 26608 11339 26648
rect 11596 26608 11636 26648
rect 12355 26608 12395 26648
rect 12460 26608 12500 26648
rect 12988 26608 13028 26648
rect 14476 26608 14516 26648
rect 18988 26608 19028 26648
rect 20140 26608 20180 26648
rect 20419 26608 20459 26648
rect 22060 26608 22100 26648
rect 23788 26608 23828 26648
rect 24652 26608 24692 26648
rect 27244 26608 27284 26648
rect 28300 26608 28340 26648
rect 30787 26608 30827 26648
rect 31084 26608 31124 26648
rect 4352 26440 4720 26480
rect 12126 26440 12494 26480
rect 19900 26440 20268 26480
rect 27674 26440 28042 26480
rect 2668 26272 2708 26312
rect 5020 26272 5060 26312
rect 8812 26272 8852 26312
rect 11308 26272 11348 26312
rect 12172 26272 12212 26312
rect 12739 26272 12779 26312
rect 13507 26272 13547 26312
rect 13612 26272 13652 26312
rect 18019 26314 18059 26354
rect 16348 26272 16388 26312
rect 3004 26188 3044 26228
rect 4012 26188 4052 26228
rect 18136 26230 18176 26270
rect 18892 26272 18932 26312
rect 20515 26272 20555 26312
rect 25180 26272 25220 26312
rect 25507 26272 25547 26312
rect 27052 26272 27092 26312
rect 27820 26272 27860 26312
rect 31276 26272 31316 26312
rect 4684 26188 4724 26228
rect 6499 26188 6539 26228
rect 8995 26188 9035 26228
rect 13891 26188 13931 26228
rect 22051 26188 22091 26228
rect 26428 26188 26468 26228
rect 2092 26104 2132 26144
rect 2275 26104 2315 26144
rect 2851 26095 2891 26135
rect 3340 26104 3380 26144
rect 4300 26104 4340 26144
rect 4579 26104 4619 26144
rect 5164 26104 5204 26144
rect 6883 26104 6923 26144
rect 9379 26104 9419 26144
rect 11500 26104 11540 26144
rect 6355 26062 6395 26102
rect 12460 26104 12500 26144
rect 12676 26104 12716 26144
rect 12849 26104 12889 26144
rect 12961 26104 13001 26144
rect 13084 26093 13124 26133
rect 13219 26104 13259 26144
rect 13409 26104 13449 26144
rect 13722 26104 13762 26144
rect 14275 26104 14315 26144
rect 16492 26104 16532 26144
rect 16675 26104 16715 26144
rect 17356 26104 17396 26144
rect 18056 26146 18096 26186
rect 18355 26104 18395 26144
rect 18503 26104 18543 26144
rect 18700 26104 18740 26144
rect 19564 26104 19604 26144
rect 19756 26104 19796 26144
rect 20044 26104 20084 26144
rect 20668 26104 20708 26144
rect 20812 26104 20852 26144
rect 21379 26104 21419 26144
rect 22435 26104 22475 26144
rect 24556 26104 24596 26144
rect 24739 26104 24779 26144
rect 24844 26104 24884 26144
rect 25027 26095 25067 26135
rect 25804 26104 25844 26144
rect 26275 26095 26315 26135
rect 26764 26104 26804 26144
rect 26892 26080 26932 26120
rect 27340 26104 27380 26144
rect 27724 26104 27764 26144
rect 28780 26104 28820 26144
rect 29347 26104 29387 26144
rect 844 26020 884 26060
rect 6163 26020 6203 26060
rect 18220 26020 18260 26060
rect 25714 26020 25754 26060
rect 28972 26020 29012 26060
rect 604 25936 644 25976
rect 1516 25936 1556 25976
rect 1900 25936 1940 25976
rect 2275 25936 2315 25976
rect 16204 25936 16244 25976
rect 17548 25936 17588 25976
rect 18604 25936 18644 25976
rect 20380 25936 20420 25976
rect 24364 25936 24404 25976
rect 24844 25936 24884 25976
rect 28108 25936 28148 25976
rect 5836 25852 5876 25892
rect 21772 25852 21812 25892
rect 3112 25684 3480 25724
rect 10886 25684 11254 25724
rect 18660 25684 19028 25724
rect 26434 25684 26802 25724
rect 5548 25516 5588 25556
rect 7843 25516 7883 25556
rect 8860 25516 8900 25556
rect 21091 25516 21131 25556
rect 26860 25516 26900 25556
rect 28108 25516 28148 25556
rect 1612 25432 1652 25472
rect 2380 25432 2420 25472
rect 7612 25423 7652 25463
rect 9196 25432 9236 25472
rect 10780 25432 10820 25472
rect 11596 25432 11636 25472
rect 14188 25432 14228 25472
rect 14764 25432 14804 25472
rect 18700 25432 18740 25472
rect 25228 25432 25268 25472
rect 25676 25423 25716 25463
rect 26380 25432 26420 25472
rect 30988 25432 31028 25472
rect 652 25348 692 25388
rect 1228 25348 1268 25388
rect 2659 25348 2699 25388
rect 3052 25348 3092 25388
rect 8620 25348 8660 25388
rect 9580 25348 9620 25388
rect 13852 25348 13892 25388
rect 14668 25348 14708 25388
rect 16396 25348 16436 25388
rect 25324 25348 25364 25388
rect 27340 25348 27380 25388
rect 1804 25264 1844 25304
rect 1996 25264 2036 25304
rect 2519 25264 2559 25304
rect 2757 25264 2797 25304
rect 3427 25264 3467 25304
rect 5932 25255 5972 25295
rect 6220 25264 6260 25304
rect 6508 25264 6548 25304
rect 6892 25264 6932 25304
rect 7276 25264 7316 25304
rect 7651 25264 7691 25304
rect 8344 25264 8384 25304
rect 9955 25264 9995 25304
rect 10348 25264 10388 25304
rect 10636 25264 10676 25304
rect 10867 25264 10907 25304
rect 11404 25264 11444 25304
rect 11519 25264 11559 25304
rect 11692 25264 11732 25304
rect 11920 25264 11960 25304
rect 12067 25264 12107 25304
rect 12184 25264 12224 25304
rect 12305 25275 12345 25315
rect 12451 25264 12491 25304
rect 12745 25264 12785 25304
rect 12870 25264 12910 25304
rect 12988 25264 13028 25304
rect 13216 25264 13256 25304
rect 13666 25264 13706 25304
rect 14524 25264 14564 25304
rect 14839 25264 14879 25304
rect 14995 25264 15035 25304
rect 15820 25264 15860 25304
rect 15995 25264 16035 25304
rect 16204 25264 16244 25304
rect 16771 25264 16811 25304
rect 18988 25264 19028 25304
rect 19852 25264 19892 25304
rect 20140 25264 20180 25304
rect 20563 25264 20603 25304
rect 21388 25264 21428 25304
rect 21955 25264 21995 25304
rect 24748 25264 24788 25304
rect 24988 25264 25028 25304
rect 892 25180 932 25220
rect 5836 25180 5876 25220
rect 8179 25180 8219 25220
rect 9340 25180 9380 25220
rect 12451 25180 12491 25220
rect 25160 25222 25200 25262
rect 25445 25264 25485 25304
rect 25699 25264 25739 25304
rect 26092 25264 26132 25304
rect 26275 25264 26315 25304
rect 26380 25264 26420 25304
rect 26563 25264 26603 25304
rect 26999 25264 27039 25304
rect 27139 25264 27179 25304
rect 27244 25264 27284 25304
rect 27523 25264 27563 25304
rect 28780 25264 28820 25304
rect 29644 25264 29684 25304
rect 30508 25264 30548 25304
rect 30796 25264 30836 25304
rect 21086 25180 21126 25220
rect 21571 25180 21611 25220
rect 26668 25180 26708 25220
rect 26871 25180 26911 25220
rect 27831 25180 27871 25220
rect 28963 25180 29003 25220
rect 988 25096 1028 25136
rect 1987 25096 2027 25136
rect 2851 25096 2891 25136
rect 5356 25096 5396 25136
rect 6988 25096 7028 25136
rect 7843 25096 7883 25136
rect 11068 25096 11108 25136
rect 13036 25096 13076 25136
rect 13372 25096 13412 25136
rect 15148 25096 15188 25136
rect 16195 25096 16235 25136
rect 19660 25096 19700 25136
rect 20332 25096 20372 25136
rect 20764 25096 20804 25136
rect 21292 25096 21332 25136
rect 23884 25096 23924 25136
rect 24076 25096 24116 25136
rect 25891 25096 25931 25136
rect 27619 25096 27659 25136
rect 27724 25096 27764 25136
rect 29836 25096 29876 25136
rect 30691 25096 30731 25136
rect 4352 24928 4720 24968
rect 12126 24928 12494 24968
rect 19900 24928 20268 24968
rect 27674 24928 28042 24968
rect 1708 24760 1748 24800
rect 13699 24760 13739 24800
rect 17452 24760 17492 24800
rect 19843 24760 19883 24800
rect 20515 24760 20555 24800
rect 22156 24760 22196 24800
rect 22540 24760 22580 24800
rect 23107 24760 23147 24800
rect 23731 24760 23771 24800
rect 24460 24760 24500 24800
rect 25219 24760 25259 24800
rect 26572 24760 26612 24800
rect 31276 24760 31316 24800
rect 1891 24676 1931 24716
rect 6115 24676 6155 24716
rect 8419 24676 8459 24716
rect 9196 24676 9236 24716
rect 13507 24667 13547 24707
rect 15139 24676 15179 24716
rect 27614 24676 27654 24716
rect 27820 24676 27860 24716
rect 2275 24592 2315 24632
rect 4396 24592 4436 24632
rect 8035 24592 8075 24632
rect 8702 24592 8742 24632
rect 8908 24592 8948 24632
rect 9004 24583 9044 24623
rect 9292 24592 9332 24632
rect 9509 24592 9549 24632
rect 10243 24592 10283 24632
rect 12364 24592 12404 24632
rect 13219 24592 13259 24632
rect 13324 24583 13364 24623
rect 13599 24592 13639 24632
rect 13780 24592 13820 24632
rect 14179 24583 14219 24623
rect 14668 24592 14708 24632
rect 14790 24592 14830 24632
rect 14917 24592 14957 24632
rect 15523 24592 15563 24632
rect 18124 24592 18164 24632
rect 18316 24592 18356 24632
rect 18499 24583 18539 24623
rect 19276 24592 19316 24632
rect 19493 24592 19533 24632
rect 19948 24592 19988 24632
rect 20332 24592 20372 24632
rect 20620 24592 20660 24632
rect 21304 24592 21344 24632
rect 21484 24592 21524 24632
rect 22334 24592 22374 24632
rect 22540 24592 22580 24632
rect 22636 24583 22676 24623
rect 22775 24592 22815 24632
rect 22915 24592 22955 24632
rect 23020 24592 23060 24632
rect 23404 24592 23444 24632
rect 23896 24592 23936 24632
rect 24076 24592 24116 24632
rect 24198 24592 24238 24632
rect 1324 24508 1364 24548
rect 9411 24508 9451 24548
rect 9868 24508 9908 24548
rect 11788 24508 11828 24548
rect 14332 24508 14372 24548
rect 18652 24508 18692 24548
rect 19180 24508 19220 24548
rect 19395 24508 19435 24548
rect 21139 24508 21179 24548
rect 24316 24550 24356 24590
rect 24415 24583 24455 24623
rect 24652 24592 24692 24632
rect 24887 24592 24927 24632
rect 25132 24592 25172 24632
rect 25411 24583 25451 24623
rect 25900 24592 25940 24632
rect 26025 24592 26065 24632
rect 26188 24592 26228 24632
rect 26369 24592 26409 24632
rect 26668 24583 26708 24623
rect 26908 24592 26948 24632
rect 27138 24592 27178 24632
rect 27331 24592 27371 24632
rect 27436 24592 27476 24632
rect 27916 24583 27956 24623
rect 28108 24592 28148 24632
rect 29347 24592 29387 24632
rect 23260 24508 23300 24548
rect 24796 24508 24836 24548
rect 25027 24508 25067 24548
rect 25564 24508 25604 24548
rect 28972 24508 29012 24548
rect 940 24424 980 24464
rect 4204 24424 4244 24464
rect 5548 24424 5588 24464
rect 5932 24424 5972 24464
rect 13036 24424 13076 24464
rect 14956 24424 14996 24464
rect 17644 24424 17684 24464
rect 20812 24424 20852 24464
rect 26092 24424 26132 24464
rect 26812 24424 26852 24464
rect 27436 24424 27476 24464
rect 1084 24340 1124 24380
rect 5068 24340 5108 24380
rect 6508 24340 6548 24380
rect 8707 24340 8747 24380
rect 12172 24340 12212 24380
rect 18220 24340 18260 24380
rect 22339 24340 22379 24380
rect 26371 24340 26411 24380
rect 27619 24340 27659 24380
rect 28780 24340 28820 24380
rect 3112 24172 3480 24212
rect 10886 24172 11254 24212
rect 18660 24172 19028 24212
rect 26434 24172 26802 24212
rect 1036 24004 1076 24044
rect 4588 24004 4628 24044
rect 6172 24004 6212 24044
rect 10819 24004 10859 24044
rect 16876 24004 16916 24044
rect 24364 24004 24404 24044
rect 25468 24004 25508 24044
rect 28108 24004 28148 24044
rect 12652 23920 12692 23960
rect 14668 23920 14708 23960
rect 19516 23920 19556 23960
rect 24499 23920 24539 23960
rect 27244 23920 27284 23960
rect 9292 23836 9332 23876
rect 9628 23836 9668 23876
rect 10444 23836 10484 23876
rect 14956 23836 14996 23876
rect 18403 23836 18443 23876
rect 23596 23836 23636 23876
rect 28972 23836 29012 23876
rect 2563 23752 2603 23792
rect 4108 23752 4148 23792
rect 4396 23752 4436 23792
rect 4972 23743 5012 23783
rect 5260 23752 5300 23792
rect 5548 23752 5588 23792
rect 5932 23752 5972 23792
rect 6646 23752 6686 23792
rect 6979 23752 7019 23792
rect 7660 23752 7700 23792
rect 8716 23752 8756 23792
rect 8812 23752 8852 23792
rect 8971 23752 9011 23792
rect 9091 23752 9131 23792
rect 9196 23752 9236 23792
rect 9484 23752 9524 23792
rect 9772 23752 9812 23792
rect 9964 23752 10004 23792
rect 10103 23752 10143 23792
rect 10243 23752 10283 23792
rect 10348 23752 10388 23792
rect 10631 23752 10671 23792
rect 10819 23752 10859 23792
rect 11008 23752 11048 23792
rect 11164 23752 11204 23792
rect 12364 23752 12404 23792
rect 12652 23752 12692 23792
rect 12767 23752 12807 23792
rect 12940 23752 12980 23792
rect 13132 23752 13172 23792
rect 13516 23752 13556 23792
rect 13996 23752 14036 23792
rect 14275 23752 14315 23792
rect 15331 23752 15371 23792
rect 18124 23752 18164 23792
rect 18796 23752 18836 23792
rect 19027 23752 19067 23792
rect 19660 23752 19700 23792
rect 20035 23752 20075 23792
rect 20140 23752 20180 23792
rect 20764 23752 20804 23792
rect 20908 23752 20948 23792
rect 21724 23752 21764 23792
rect 21868 23752 21908 23792
rect 22339 23752 22379 23792
rect 22457 23752 22497 23792
rect 22617 23752 22657 23792
rect 22723 23752 22763 23792
rect 22857 23752 22897 23792
rect 23416 23752 23456 23792
rect 23692 23752 23732 23792
rect 23811 23752 23851 23792
rect 23932 23752 23972 23792
rect 24067 23752 24107 23792
rect 24708 23752 24748 23792
rect 24844 23752 24884 23792
rect 25079 23752 25119 23792
rect 25219 23743 25259 23783
rect 25324 23752 25364 23792
rect 25612 23752 25652 23792
rect 25847 23752 25887 23792
rect 25987 23743 26027 23783
rect 26092 23752 26132 23792
rect 26467 23752 26507 23792
rect 26775 23752 26815 23792
rect 26947 23752 26987 23792
rect 27244 23752 27284 23792
rect 27628 23752 27668 23792
rect 27772 23752 27812 23792
rect 28780 23752 28820 23792
rect 29347 23752 29387 23792
rect 643 23668 683 23708
rect 2947 23668 2987 23708
rect 3427 23668 3467 23708
rect 4876 23668 4916 23708
rect 6451 23668 6491 23708
rect 7290 23668 7330 23708
rect 8510 23668 8550 23708
rect 14380 23668 14420 23708
rect 17443 23668 17483 23708
rect 19228 23668 19268 23708
rect 23251 23668 23291 23708
rect 24378 23668 24418 23708
rect 27427 23668 27467 23708
rect 4252 23584 4292 23624
rect 7075 23584 7115 23624
rect 7180 23584 7220 23624
rect 8332 23584 8372 23624
rect 8611 23584 8651 23624
rect 9955 23584 9995 23624
rect 11692 23584 11732 23624
rect 13612 23584 13652 23624
rect 17260 23584 17300 23624
rect 20428 23584 20468 23624
rect 20611 23584 20651 23624
rect 21571 23584 21611 23624
rect 22819 23584 22859 23624
rect 24163 23584 24203 23624
rect 25036 23584 25076 23624
rect 25804 23584 25844 23624
rect 26563 23584 26603 23624
rect 26668 23584 26708 23624
rect 27724 23584 27764 23624
rect 31276 23584 31316 23624
rect 4352 23416 4720 23456
rect 12126 23416 12494 23456
rect 19900 23416 20268 23456
rect 27674 23416 28042 23456
rect 1699 23248 1739 23288
rect 3571 23248 3611 23288
rect 4003 23248 4043 23288
rect 4108 23248 4148 23288
rect 4780 23248 4820 23288
rect 5068 23248 5108 23288
rect 5635 23248 5675 23288
rect 11491 23248 11531 23288
rect 12892 23248 12932 23288
rect 15043 23248 15083 23288
rect 18211 23248 18251 23288
rect 18508 23248 18548 23288
rect 19180 23248 19220 23288
rect 20419 23248 20459 23288
rect 20524 23248 20564 23288
rect 21619 23248 21659 23288
rect 28492 23248 28532 23288
rect 2179 23164 2219 23204
rect 2284 23164 2324 23204
rect 3244 23164 3284 23204
rect 4675 23164 4715 23204
rect 5534 23164 5574 23204
rect 6115 23164 6155 23204
rect 10732 23164 10772 23204
rect 15340 23164 15380 23204
rect 16675 23164 16715 23204
rect 17932 23164 17972 23204
rect 19987 23164 20027 23204
rect 20634 23164 20674 23204
rect 20956 23164 20996 23204
rect 25132 23164 25172 23204
rect 25795 23155 25835 23195
rect 26956 23164 26996 23204
rect 844 23080 884 23120
rect 1027 23080 1067 23120
rect 1228 23080 1268 23120
rect 1411 23080 1451 23120
rect 1603 23080 1643 23120
rect 1914 23080 1954 23120
rect 2081 23080 2121 23120
rect 2380 23071 2420 23111
rect 2572 23080 2612 23120
rect 3736 23080 3776 23120
rect 3905 23080 3945 23120
rect 4204 23071 4244 23111
rect 4574 23080 4614 23120
rect 4876 23071 4916 23111
rect 5164 23080 5204 23120
rect 5401 23080 5441 23120
rect 5740 23080 5780 23120
rect 5836 23071 5876 23111
rect 7084 23080 7124 23120
rect 7468 23080 7508 23120
rect 8332 23080 8372 23120
rect 8515 23080 8555 23120
rect 9772 23080 9812 23120
rect 10348 23080 10388 23120
rect 10585 23080 10625 23120
rect 10828 23080 10868 23120
rect 11045 23080 11085 23120
rect 11164 23080 11204 23120
rect 11299 23080 11339 23120
rect 11404 23080 11444 23120
rect 11884 23080 11924 23120
rect 12121 23080 12161 23120
rect 12364 23080 12404 23120
rect 12556 23080 12596 23120
rect 12748 23080 12788 23120
rect 13420 23080 13460 23120
rect 13612 23080 13652 23120
rect 13804 23080 13844 23120
rect 13987 23080 14027 23120
rect 14284 23080 14324 23120
rect 14521 23080 14561 23120
rect 14860 23075 14900 23115
rect 15055 23080 15095 23120
rect 15244 23080 15284 23120
rect 15436 23080 15476 23120
rect 17452 23080 17492 23120
rect 17836 23080 17876 23120
rect 18028 23080 18068 23120
rect 18316 23080 18356 23120
rect 19180 23080 19220 23120
rect 19372 23080 19412 23120
rect 20152 23080 20192 23120
rect 20323 23080 20363 23120
rect 20812 23080 20852 23120
rect 21376 23071 21416 23111
rect 21475 23080 21515 23120
rect 21772 23080 21812 23120
rect 21964 23080 22004 23120
rect 22531 23080 22571 23120
rect 24835 23080 24875 23120
rect 25507 23080 25547 23120
rect 25612 23071 25652 23111
rect 25891 23080 25931 23120
rect 26068 23080 26108 23120
rect 26467 23080 26507 23120
rect 26659 23080 26699 23120
rect 26764 23080 26804 23120
rect 27069 23065 27109 23105
rect 27211 23080 27251 23120
rect 27436 23080 27476 23120
rect 28053 23080 28093 23120
rect 28204 23080 28244 23120
rect 28346 23048 28386 23088
rect 29356 23080 29396 23120
rect 29548 23080 29588 23120
rect 30403 23080 30443 23120
rect 31084 23080 31124 23120
rect 5068 22996 5108 23036
rect 5283 22996 5323 23036
rect 10252 22996 10292 23036
rect 10467 22996 10507 23036
rect 10947 22996 10987 23036
rect 11788 22996 11828 23036
rect 12019 22987 12059 23027
rect 13228 22996 13268 23036
rect 14188 22996 14228 23036
rect 14403 22996 14443 23036
rect 22156 22996 22196 23036
rect 24652 22996 24692 23036
rect 25228 22996 25268 23036
rect 27331 22996 27371 23036
rect 27532 22996 27572 23036
rect 27859 22996 27899 23036
rect 1027 22912 1067 22952
rect 1411 22912 1451 22952
rect 8515 22912 8555 22952
rect 8995 22912 9035 22952
rect 13987 22912 14027 22952
rect 15820 22912 15860 22952
rect 16012 22912 16052 22952
rect 18700 22912 18740 22952
rect 21772 22912 21812 22952
rect 24460 22912 24500 22952
rect 1900 22828 1940 22868
rect 8140 22828 8180 22868
rect 12460 22828 12500 22868
rect 12988 22828 13028 22868
rect 13420 22828 13460 22868
rect 21091 22828 21131 22868
rect 25507 22828 25547 22868
rect 28684 22828 28724 22868
rect 30220 22828 30260 22868
rect 3112 22660 3480 22700
rect 10886 22660 11254 22700
rect 18660 22660 19028 22700
rect 26434 22660 26802 22700
rect 6019 22492 6059 22532
rect 7267 22492 7307 22532
rect 10636 22492 10676 22532
rect 11404 22492 11444 22532
rect 11692 22492 11732 22532
rect 14563 22492 14603 22532
rect 20323 22492 20363 22532
rect 21187 22492 21227 22532
rect 21955 22492 21995 22532
rect 23971 22492 24011 22532
rect 25900 22492 25940 22532
rect 27148 22492 27188 22532
rect 27724 22492 27764 22532
rect 8995 22408 9035 22448
rect 16483 22408 16523 22448
rect 17740 22408 17780 22448
rect 18892 22408 18932 22448
rect 19267 22408 19307 22448
rect 24268 22408 24308 22448
rect 29356 22408 29396 22448
rect 2380 22324 2420 22364
rect 2611 22315 2651 22355
rect 3763 22324 3803 22364
rect 4108 22324 4148 22364
rect 4339 22315 4379 22355
rect 5356 22324 5396 22364
rect 5836 22324 5876 22364
rect 1708 22240 1748 22280
rect 1891 22240 1931 22280
rect 2199 22240 2239 22280
rect 2476 22240 2516 22280
rect 2713 22240 2753 22280
rect 3300 22240 3340 22280
rect 3436 22240 3476 22280
rect 3928 22240 3968 22280
rect 4204 22240 4244 22280
rect 4441 22240 4481 22280
rect 4780 22240 4820 22280
rect 4972 22240 5012 22280
rect 5495 22240 5535 22280
rect 5635 22240 5675 22280
rect 5740 22240 5780 22280
rect 6314 22273 6354 22313
rect 6460 22282 6500 22322
rect 6796 22324 6836 22364
rect 7843 22324 7883 22364
rect 13699 22324 13739 22364
rect 18451 22324 18491 22364
rect 18988 22324 19028 22364
rect 19171 22324 19211 22364
rect 19747 22324 19787 22364
rect 20338 22324 20378 22364
rect 22723 22324 22763 22364
rect 25507 22324 25547 22364
rect 27826 22324 27866 22364
rect 6595 22240 6635 22280
rect 6700 22240 6740 22280
rect 7265 22240 7305 22280
rect 7564 22240 7604 22280
rect 7703 22240 7743 22280
rect 7948 22240 7988 22280
rect 8524 22240 8564 22280
rect 9667 22240 9707 22280
rect 9964 22240 10004 22280
rect 10154 22240 10194 22280
rect 10446 22240 10486 22280
rect 10828 22240 10868 22280
rect 10989 22240 11029 22280
rect 11107 22240 11147 22280
rect 11212 22273 11252 22313
rect 11596 22240 11636 22280
rect 11788 22240 11828 22280
rect 12280 22240 12320 22280
rect 13324 22240 13364 22280
rect 13804 22240 13844 22280
rect 13996 22240 14036 22280
rect 15148 22240 15188 22280
rect 15724 22240 15764 22280
rect 15820 22240 15860 22280
rect 17068 22240 17108 22280
rect 18028 22240 18068 22280
rect 18147 22240 18187 22280
rect 18265 22240 18305 22280
rect 18595 22240 18635 22280
rect 19555 22240 19595 22280
rect 20428 22240 20468 22280
rect 21181 22240 21221 22280
rect 21292 22240 21332 22280
rect 22240 22273 22280 22313
rect 22339 22240 22379 22280
rect 22603 22240 22643 22280
rect 22828 22240 22868 22280
rect 23099 22240 23139 22280
rect 23308 22240 23348 22280
rect 23683 22240 23723 22280
rect 23788 22240 23828 22280
rect 24268 22240 24308 22280
rect 24458 22240 24498 22280
rect 24642 22240 24682 22280
rect 24835 22240 24875 22280
rect 24940 22240 24980 22280
rect 25387 22240 25427 22280
rect 25612 22240 25652 22280
rect 25943 22240 25983 22280
rect 26047 22240 26087 22280
rect 26188 22240 26228 22280
rect 26515 22282 26555 22322
rect 31267 22324 31307 22364
rect 26377 22240 26417 22280
rect 26629 22240 26669 22280
rect 26851 22240 26891 22280
rect 27148 22240 27188 22280
rect 27436 22240 27476 22280
rect 27916 22240 27956 22280
rect 28696 22240 28736 22280
rect 30883 22240 30923 22280
rect 739 22156 779 22196
rect 2092 22156 2132 22196
rect 4876 22156 4916 22196
rect 6017 22156 6057 22196
rect 7468 22156 7508 22196
rect 8222 22156 8262 22196
rect 8428 22156 8468 22196
rect 15518 22156 15558 22196
rect 23212 22156 23252 22196
rect 24739 22156 24779 22196
rect 28531 22156 28571 22196
rect 1987 22072 2027 22112
rect 3139 22072 3179 22112
rect 5116 22072 5156 22112
rect 6220 22072 6260 22112
rect 8035 22072 8075 22112
rect 8323 22072 8363 22112
rect 10060 22072 10100 22112
rect 10339 22072 10379 22112
rect 12115 22072 12155 22112
rect 12739 22072 12779 22112
rect 15619 22072 15659 22112
rect 17932 22072 17972 22112
rect 20131 22072 20171 22112
rect 22459 22072 22499 22112
rect 22915 22072 22955 22112
rect 25699 22072 25739 22112
rect 26668 22072 26708 22112
rect 28972 22072 29012 22112
rect 4352 21904 4720 21944
rect 12126 21904 12494 21944
rect 19900 21904 20268 21944
rect 27674 21904 28042 21944
rect 1315 21736 1355 21776
rect 3532 21736 3572 21776
rect 5347 21736 5387 21776
rect 5923 21736 5963 21776
rect 6316 21736 6356 21776
rect 6883 21736 6923 21776
rect 7372 21736 7412 21776
rect 8620 21736 8660 21776
rect 9763 21736 9803 21776
rect 10435 21736 10475 21776
rect 10723 21736 10763 21776
rect 11203 21736 11243 21776
rect 13603 21736 13643 21776
rect 15907 21736 15947 21776
rect 22156 21736 22196 21776
rect 23596 21736 23636 21776
rect 24172 21736 24212 21776
rect 25564 21736 25604 21776
rect 26380 21736 26420 21776
rect 27259 21736 27299 21776
rect 27580 21736 27620 21776
rect 28636 21736 28676 21776
rect 2846 21652 2886 21692
rect 3639 21652 3679 21692
rect 4771 21652 4811 21692
rect 6028 21652 6068 21692
rect 6782 21652 6822 21692
rect 7852 21652 7892 21692
rect 8092 21652 8132 21692
rect 9388 21652 9428 21692
rect 10938 21652 10978 21692
rect 11418 21652 11458 21692
rect 11740 21652 11780 21692
rect 14764 21652 14804 21692
rect 16723 21652 16763 21692
rect 18307 21652 18347 21692
rect 26284 21652 26324 21692
rect 27998 21652 28038 21692
rect 28963 21652 29003 21692
rect 1132 21568 1172 21608
rect 1327 21568 1367 21608
rect 1516 21568 1556 21608
rect 1621 21568 1661 21608
rect 1843 21568 1883 21608
rect 2044 21568 2084 21608
rect 3052 21568 3092 21608
rect 3148 21559 3188 21599
rect 3331 21568 3371 21608
rect 3436 21568 3476 21608
rect 4003 21559 4043 21599
rect 4439 21568 4479 21608
rect 4684 21568 4724 21608
rect 5500 21568 5540 21608
rect 5644 21568 5684 21608
rect 5822 21568 5862 21608
rect 6124 21559 6164 21599
rect 6412 21568 6452 21608
rect 6629 21568 6669 21608
rect 6988 21568 7028 21608
rect 7084 21559 7124 21599
rect 7372 21568 7412 21608
rect 7564 21568 7604 21608
rect 7756 21568 7796 21608
rect 7948 21568 7988 21608
rect 8284 21568 8324 21608
rect 8428 21568 8468 21608
rect 8716 21568 8756 21608
rect 8953 21568 8993 21608
rect 9292 21568 9332 21608
rect 9484 21568 9524 21608
rect 9667 21568 9707 21608
rect 9975 21568 10015 21608
rect 10131 21568 10171 21608
rect 10348 21568 10388 21608
rect 10627 21568 10667 21608
rect 11107 21568 11147 21608
rect 11587 21559 11627 21599
rect 12211 21568 12251 21608
rect 12643 21568 12683 21608
rect 13516 21568 13556 21608
rect 844 21484 884 21524
rect 1747 21475 1787 21515
rect 4156 21484 4196 21524
rect 4579 21484 4619 21524
rect 4972 21484 5012 21524
rect 6531 21484 6571 21524
rect 12403 21526 12443 21566
rect 13751 21568 13791 21608
rect 13996 21568 14036 21608
rect 14467 21568 14507 21608
rect 15052 21568 15092 21608
rect 8835 21484 8875 21524
rect 10243 21484 10283 21524
rect 13891 21484 13931 21524
rect 14092 21484 14132 21524
rect 14284 21484 14324 21524
rect 14860 21484 14900 21524
rect 15292 21526 15332 21566
rect 15533 21568 15573 21608
rect 16195 21568 16235 21608
rect 16888 21568 16928 21608
rect 17068 21568 17108 21608
rect 17260 21568 17300 21608
rect 18595 21568 18635 21608
rect 18988 21568 19028 21608
rect 19180 21568 19220 21608
rect 19756 21568 19796 21608
rect 19993 21568 20033 21608
rect 20332 21568 20372 21608
rect 20716 21568 20756 21608
rect 21100 21568 21140 21608
rect 21484 21568 21524 21608
rect 21671 21568 21711 21608
rect 21868 21568 21908 21608
rect 22060 21568 22100 21608
rect 22243 21568 22283 21608
rect 22723 21568 22763 21608
rect 22828 21568 22868 21608
rect 23404 21568 23444 21608
rect 23596 21568 23636 21608
rect 24163 21568 24203 21608
rect 24268 21568 24308 21608
rect 24599 21568 24639 21608
rect 24844 21568 24884 21608
rect 25131 21568 25171 21608
rect 25315 21568 25355 21608
rect 25420 21568 25460 21608
rect 25708 21568 25748 21608
rect 26179 21559 26219 21599
rect 26476 21568 26516 21608
rect 27048 21559 27088 21599
rect 27139 21568 27179 21608
rect 27427 21559 27467 21599
rect 28204 21568 28244 21608
rect 28300 21559 28340 21599
rect 28483 21559 28523 21599
rect 29347 21568 29387 21608
rect 15427 21484 15467 21524
rect 15628 21484 15668 21524
rect 15811 21484 15851 21524
rect 16387 21484 16427 21524
rect 18211 21484 18251 21524
rect 18787 21484 18827 21524
rect 19660 21484 19700 21524
rect 19891 21475 19931 21515
rect 24739 21484 24779 21524
rect 24940 21484 24980 21524
rect 5212 21400 5252 21440
rect 12844 21400 12884 21440
rect 17644 21400 17684 21440
rect 18028 21400 18068 21440
rect 20092 21400 20132 21440
rect 20860 21400 20900 21440
rect 23395 21400 23435 21440
rect 25420 21400 25460 21440
rect 604 21316 644 21356
rect 2668 21316 2708 21356
rect 2851 21316 2891 21356
rect 7852 21316 7892 21356
rect 9964 21316 10004 21356
rect 10924 21316 10964 21356
rect 11404 21316 11444 21356
rect 13036 21316 13076 21356
rect 13324 21316 13364 21356
rect 15196 21316 15236 21356
rect 17164 21316 17204 21356
rect 18988 21316 19028 21356
rect 21772 21316 21812 21356
rect 23011 21316 23051 21356
rect 24460 21316 24500 21356
rect 25996 21316 26036 21356
rect 26755 21316 26795 21356
rect 28003 21316 28043 21356
rect 31276 21316 31316 21356
rect 3112 21148 3480 21188
rect 10886 21148 11254 21188
rect 18660 21148 19028 21188
rect 26434 21148 26802 21188
rect 604 20980 644 21020
rect 1228 20980 1268 21020
rect 3532 20980 3572 21020
rect 4963 20980 5003 21020
rect 7372 20980 7412 21020
rect 7948 20980 7988 21020
rect 9052 20980 9092 21020
rect 13084 20980 13124 21020
rect 14371 20980 14411 21020
rect 15628 20980 15668 21020
rect 17155 20980 17195 21020
rect 20515 20980 20555 21020
rect 21292 20980 21332 21020
rect 24451 20980 24491 21020
rect 25804 20980 25844 21020
rect 26380 20980 26420 21020
rect 27715 20980 27755 21020
rect 29836 20980 29876 21020
rect 21868 20896 21908 20936
rect 844 20812 884 20852
rect 3916 20812 3956 20852
rect 4339 20803 4379 20843
rect 5164 20812 5204 20852
rect 6844 20812 6884 20852
rect 7084 20812 7124 20852
rect 8140 20812 8180 20852
rect 8355 20812 8395 20852
rect 8620 20812 8660 20852
rect 9292 20812 9332 20852
rect 14947 20812 14987 20852
rect 19267 20812 19307 20852
rect 19468 20812 19508 20852
rect 1132 20728 1172 20768
rect 1324 20728 1364 20768
rect 1516 20728 1556 20768
rect 1708 20733 1748 20773
rect 1900 20728 1940 20768
rect 2092 20728 2132 20768
rect 2574 20728 2614 20768
rect 3091 20728 3131 20768
rect 3235 20728 3275 20768
rect 4204 20728 4244 20768
rect 4441 20728 4481 20768
rect 4780 20728 4820 20768
rect 4963 20728 5003 20768
rect 5260 20728 5300 20768
rect 5379 20728 5419 20768
rect 5497 20728 5537 20768
rect 5644 20728 5684 20768
rect 5827 20728 5867 20768
rect 6029 20728 6069 20768
rect 6218 20728 6258 20768
rect 6412 20728 6452 20768
rect 6604 20728 6644 20768
rect 7276 20728 7316 20768
rect 7467 20728 7507 20768
rect 7651 20728 7691 20768
rect 8236 20728 8276 20768
rect 8473 20728 8513 20768
rect 8716 20728 8756 20768
rect 8851 20719 8891 20759
rect 8953 20728 8993 20768
rect 11059 20770 11099 20810
rect 19948 20812 19988 20852
rect 24739 20812 24779 20852
rect 25315 20812 25355 20852
rect 28963 20812 29003 20852
rect 9580 20728 9620 20768
rect 9763 20728 9803 20768
rect 10252 20728 10292 20768
rect 11542 20728 11582 20768
rect 11683 20728 11723 20768
rect 12364 20728 12404 20768
rect 12652 20728 12692 20768
rect 12844 20728 12884 20768
rect 13228 20728 13268 20768
rect 13750 20728 13790 20768
rect 14052 20728 14092 20768
rect 14188 20728 14228 20768
rect 14572 20728 14612 20768
rect 14668 20728 14708 20768
rect 14827 20728 14867 20768
rect 15052 20728 15092 20768
rect 15331 20728 15371 20768
rect 16150 20728 16190 20768
rect 16780 20728 16820 20768
rect 17059 20719 17099 20759
rect 17356 20728 17396 20768
rect 17687 20728 17727 20768
rect 17827 20728 17867 20768
rect 17932 20728 17972 20768
rect 18211 20728 18251 20768
rect 18522 20728 18562 20768
rect 18700 20728 18740 20768
rect 18839 20728 18879 20768
rect 19127 20728 19167 20768
rect 19353 20728 19393 20768
rect 19607 20728 19647 20768
rect 19747 20728 19787 20768
rect 19852 20728 19892 20768
rect 20908 20728 20948 20768
rect 21292 20728 21332 20768
rect 21484 20728 21524 20768
rect 22156 20728 22196 20768
rect 23107 20728 23147 20768
rect 24163 20728 24203 20768
rect 24270 20728 24310 20768
rect 25123 20728 25163 20768
rect 25612 20728 25652 20768
rect 26092 20728 26132 20768
rect 26275 20728 26315 20768
rect 26380 20728 26420 20768
rect 26659 20728 26699 20768
rect 26967 20728 27007 20768
rect 27148 20728 27188 20768
rect 27290 20728 27330 20768
rect 27619 20719 27659 20759
rect 27916 20728 27956 20768
rect 28387 20728 28427 20768
rect 28492 20728 28532 20768
rect 29644 20728 29684 20768
rect 30508 20728 30548 20768
rect 30892 20728 30932 20768
rect 31180 20728 31220 20768
rect 1612 20644 1652 20684
rect 2273 20644 2313 20684
rect 3543 20644 3583 20684
rect 4108 20644 4148 20684
rect 6124 20644 6164 20684
rect 7756 20644 7796 20684
rect 7962 20644 8002 20684
rect 9676 20644 9716 20684
rect 9950 20644 9990 20684
rect 12940 20644 12980 20684
rect 14366 20644 14406 20684
rect 15642 20644 15682 20684
rect 16579 20644 16619 20684
rect 18412 20644 18452 20684
rect 23299 20644 23339 20684
rect 27724 20644 27764 20684
rect 30691 20644 30731 20684
rect 1996 20560 2036 20600
rect 2371 20560 2411 20600
rect 2476 20560 2516 20600
rect 2899 20560 2939 20600
rect 3331 20560 3371 20600
rect 3676 20560 3716 20600
rect 5740 20560 5780 20600
rect 6412 20560 6452 20600
rect 10051 20560 10091 20600
rect 10156 20560 10196 20600
rect 10867 20560 10907 20600
rect 11347 20560 11387 20600
rect 13555 20560 13595 20600
rect 13891 20560 13931 20600
rect 15139 20560 15179 20600
rect 15427 20560 15467 20600
rect 15955 20560 15995 20600
rect 18019 20560 18059 20600
rect 18307 20560 18347 20600
rect 18988 20560 19028 20600
rect 20716 20560 20756 20600
rect 22828 20560 22868 20600
rect 24835 20560 24875 20600
rect 25507 20560 25547 20600
rect 25795 20560 25835 20600
rect 26755 20560 26795 20600
rect 26860 20560 26900 20600
rect 27436 20560 27476 20600
rect 28780 20560 28820 20600
rect 30979 20560 31019 20600
rect 4352 20392 4720 20432
rect 12126 20392 12494 20432
rect 19900 20392 20268 20432
rect 27674 20392 28042 20432
rect 2668 20224 2708 20264
rect 3235 20224 3275 20264
rect 5356 20224 5396 20264
rect 6211 20224 6251 20264
rect 6316 20224 6356 20264
rect 7372 20224 7412 20264
rect 8764 20224 8804 20264
rect 11692 20224 11732 20264
rect 12748 20224 12788 20264
rect 12931 20224 12971 20264
rect 13132 20224 13172 20264
rect 14179 20224 14219 20264
rect 14851 20224 14891 20264
rect 14956 20224 14996 20264
rect 16204 20224 16244 20264
rect 16579 20224 16619 20264
rect 17260 20224 17300 20264
rect 18691 20224 18731 20264
rect 18796 20224 18836 20264
rect 19267 20224 19307 20264
rect 19708 20224 19748 20264
rect 24979 20224 25019 20264
rect 28972 20224 29012 20264
rect 4060 20140 4100 20180
rect 4673 20140 4713 20180
rect 4876 20140 4916 20180
rect 13795 20140 13835 20180
rect 17164 20140 17204 20180
rect 17847 20140 17887 20180
rect 20611 20140 20651 20180
rect 24748 20140 24788 20180
rect 25900 20140 25940 20180
rect 27820 20140 27860 20180
rect 28780 20140 28820 20180
rect 31267 20140 31307 20180
rect 1708 20056 1748 20096
rect 2135 20056 2175 20096
rect 2380 20056 2420 20096
rect 2764 20056 2804 20096
rect 3001 20056 3041 20096
rect 3388 20056 3428 20096
rect 3532 20056 3572 20096
rect 4972 20047 5012 20087
rect 5153 20056 5193 20096
rect 5452 20047 5492 20087
rect 5740 20056 5780 20096
rect 5977 20056 6017 20096
rect 6113 20056 6153 20096
rect 6412 20047 6452 20087
rect 6604 20056 6644 20096
rect 6709 20056 6749 20096
rect 6931 20056 6971 20096
rect 7084 20056 7124 20096
rect 7226 20056 7266 20096
rect 7756 20056 7796 20096
rect 8131 20047 8171 20087
rect 8611 20047 8651 20087
rect 9388 20056 9428 20096
rect 9763 20056 9803 20096
rect 12355 20056 12395 20096
rect 13315 20056 13355 20096
rect 13708 20056 13748 20096
rect 13900 20056 13940 20096
rect 14284 20056 14324 20096
rect 14750 20056 14790 20096
rect 15052 20047 15092 20087
rect 15340 20056 15380 20096
rect 15532 20056 15572 20096
rect 15724 20056 15764 20096
rect 15916 20056 15956 20096
rect 16108 20056 16148 20096
rect 16300 20056 16340 20096
rect 16684 20056 16724 20096
rect 17059 20056 17099 20096
rect 17367 20056 17407 20096
rect 17539 20056 17579 20096
rect 17644 20056 17684 20096
rect 18115 20056 18155 20096
rect 18220 20056 18260 20096
rect 18423 20056 18463 20096
rect 18595 20056 18635 20096
rect 18903 20056 18943 20096
rect 19084 20056 19124 20096
rect 19276 20056 19316 20096
rect 19528 20056 19568 20096
rect 20227 20056 20267 20096
rect 22531 20056 22571 20096
rect 23404 20056 23444 20096
rect 23533 20056 23573 20096
rect 23788 20056 23828 20096
rect 24451 20056 24491 20096
rect 25123 20056 25163 20096
rect 25228 20047 25268 20087
rect 25996 20056 26036 20096
rect 26233 20056 26273 20096
rect 26710 20056 26750 20096
rect 27137 20056 27177 20096
rect 27244 20056 27284 20096
rect 27619 20056 27659 20096
rect 27912 20056 27952 20096
rect 28156 20056 28196 20096
rect 30883 20056 30923 20096
rect 2275 19972 2315 20012
rect 2476 19972 2516 20012
rect 2899 19963 2939 20003
rect 3916 19972 3956 20012
rect 4300 19972 4340 20012
rect 5644 19972 5684 20012
rect 5875 19963 5915 20003
rect 6835 19963 6875 20003
rect 8284 19972 8324 20012
rect 12547 19972 12587 20012
rect 22915 19972 22955 20012
rect 24268 19972 24308 20012
rect 24844 19972 24884 20012
rect 26115 19972 26155 20012
rect 26515 19972 26555 20012
rect 11884 19888 11924 19928
rect 14476 19888 14516 19928
rect 20272 19888 20312 19928
rect 23116 19888 23156 19928
rect 931 19804 971 19844
rect 3676 19804 3716 19844
rect 4675 19804 4715 19844
rect 5155 19804 5195 19844
rect 7852 19804 7892 19844
rect 15436 19804 15476 19844
rect 15724 19804 15764 19844
rect 16876 19804 16916 19844
rect 17836 19804 17876 19844
rect 18412 19804 18452 19844
rect 20044 19804 20084 19844
rect 21004 19804 21044 19844
rect 25516 19804 25556 19844
rect 27244 19804 27284 19844
rect 3112 19636 3480 19676
rect 10886 19636 11254 19676
rect 18660 19636 19028 19676
rect 26434 19636 26802 19676
rect 2179 19468 2219 19508
rect 3724 19468 3764 19508
rect 4387 19468 4427 19508
rect 5923 19468 5963 19508
rect 6883 19468 6923 19508
rect 9580 19468 9620 19508
rect 11011 19468 11051 19508
rect 13468 19468 13508 19508
rect 14572 19468 14612 19508
rect 16492 19468 16532 19508
rect 18412 19468 18452 19508
rect 19459 19468 19499 19508
rect 22444 19468 22484 19508
rect 23116 19468 23156 19508
rect 31276 19468 31316 19508
rect 1612 19384 1652 19424
rect 12940 19384 12980 19424
rect 844 19300 884 19340
rect 5452 19300 5492 19340
rect 5667 19300 5707 19340
rect 6700 19300 6740 19340
rect 7756 19300 7796 19340
rect 9772 19300 9812 19340
rect 1804 19216 1844 19256
rect 1996 19216 2036 19256
rect 2177 19216 2217 19256
rect 2476 19216 2516 19256
rect 2947 19216 2987 19256
rect 3052 19216 3092 19256
rect 3427 19216 3467 19256
rect 3738 19216 3778 19256
rect 4012 19216 4052 19256
rect 4131 19216 4171 19256
rect 4249 19216 4289 19256
rect 4382 19216 4422 19256
rect 4684 19216 4724 19256
rect 5068 19216 5108 19256
rect 5260 19216 5300 19256
rect 5548 19216 5588 19256
rect 5785 19216 5825 19256
rect 5921 19216 5961 19256
rect 6220 19216 6260 19256
rect 6359 19216 6399 19256
rect 6499 19216 6539 19256
rect 6604 19216 6644 19256
rect 6881 19216 6921 19256
rect 7178 19249 7218 19289
rect 10444 19300 10484 19340
rect 13228 19300 13268 19340
rect 15939 19300 15979 19340
rect 18700 19300 18740 19340
rect 7852 19216 7892 19256
rect 7971 19216 8011 19256
rect 8089 19216 8129 19256
rect 8716 19216 8756 19256
rect 8908 19216 8948 19256
rect 9187 19216 9227 19256
rect 9304 19249 9344 19289
rect 9868 19216 9908 19256
rect 9987 19216 10027 19256
rect 10099 19216 10139 19256
rect 11308 19216 11348 19256
rect 11680 19216 11720 19256
rect 12643 19207 12683 19247
rect 12940 19216 12980 19256
rect 13912 19216 13952 19256
rect 14083 19216 14123 19256
rect 14394 19216 14434 19256
rect 14764 19216 14804 19256
rect 14883 19216 14923 19256
rect 15052 19216 15092 19256
rect 15191 19216 15231 19256
rect 15331 19216 15371 19256
rect 15436 19216 15476 19256
rect 15820 19216 15860 19256
rect 16060 19258 16100 19298
rect 19747 19300 19787 19340
rect 21868 19300 21908 19340
rect 24047 19300 24087 19340
rect 26572 19300 26612 19340
rect 27052 19300 27092 19340
rect 27267 19300 27307 19340
rect 16300 19216 16340 19256
rect 16984 19216 17024 19256
rect 17164 19216 17204 19256
rect 17303 19216 17343 19256
rect 18019 19216 18059 19256
rect 18136 19249 18176 19289
rect 18604 19216 18644 19256
rect 18796 19216 18836 19256
rect 19276 19216 19316 19256
rect 19445 19216 19485 19256
rect 19607 19216 19647 19256
rect 19852 19216 19892 19256
rect 20403 19216 20443 19256
rect 20803 19216 20843 19256
rect 20995 19216 21035 19256
rect 21292 19216 21332 19256
rect 21484 19216 21524 19256
rect 21772 19216 21812 19256
rect 21964 19216 22004 19256
rect 22147 19216 22187 19256
rect 22627 19216 22667 19256
rect 22924 19216 22964 19256
rect 23116 19216 23156 19256
rect 23241 19216 23281 19256
rect 23404 19216 23444 19256
rect 23945 19216 23985 19256
rect 24163 19216 24203 19256
rect 24268 19216 24308 19256
rect 24652 19216 24692 19256
rect 24835 19216 24875 19256
rect 25324 19216 25364 19256
rect 25612 19216 25652 19256
rect 25996 19216 26036 19256
rect 26659 19216 26699 19256
rect 27148 19216 27188 19256
rect 27385 19216 27425 19256
rect 27624 19216 27664 19256
rect 27820 19216 27860 19256
rect 28108 19216 28148 19256
rect 29347 19216 29387 19256
rect 3258 19132 3298 19172
rect 11006 19132 11046 19172
rect 15523 19132 15563 19172
rect 21388 19132 21428 19172
rect 22458 19132 22498 19172
rect 24748 19132 24788 19172
rect 28963 19132 29003 19172
rect 604 19048 644 19088
rect 1804 19048 1844 19088
rect 2380 19048 2420 19088
rect 3148 19048 3188 19088
rect 3523 19048 3563 19088
rect 3916 19048 3956 19088
rect 4588 19048 4628 19088
rect 5251 19048 5291 19088
rect 6124 19048 6164 19088
rect 7084 19048 7124 19088
rect 8716 19048 8756 19088
rect 9043 19048 9083 19088
rect 10204 19048 10244 19088
rect 11212 19048 11252 19088
rect 11836 19048 11876 19088
rect 13747 19048 13787 19088
rect 14179 19048 14219 19088
rect 14284 19048 14324 19088
rect 15724 19048 15764 19088
rect 16195 19048 16235 19088
rect 16819 19048 16859 19088
rect 17452 19048 17492 19088
rect 17923 19039 17963 19079
rect 19939 19048 19979 19088
rect 20515 19048 20555 19088
rect 22243 19048 22283 19088
rect 22828 19048 22868 19088
rect 23980 19048 24020 19088
rect 25123 19048 25163 19088
rect 25804 19048 25844 19088
rect 26083 19048 26123 19088
rect 26283 19039 26323 19079
rect 27628 19048 27668 19088
rect 28780 19048 28820 19088
rect 4352 18880 4720 18920
rect 12126 18880 12494 18920
rect 19900 18880 20268 18920
rect 27674 18880 28042 18920
rect 748 18712 788 18752
rect 5260 18712 5300 18752
rect 6499 18712 6539 18752
rect 6883 18712 6923 18752
rect 7651 18712 7691 18752
rect 8131 18712 8171 18752
rect 9187 18712 9227 18752
rect 9523 18712 9563 18752
rect 10732 18712 10772 18752
rect 12163 18712 12203 18752
rect 13795 18712 13835 18752
rect 15523 18712 15563 18752
rect 17347 18712 17387 18752
rect 20227 18712 20267 18752
rect 20908 18712 20948 18752
rect 21196 18712 21236 18752
rect 23020 18712 23060 18752
rect 24268 18712 24308 18752
rect 25699 18712 25739 18752
rect 10636 18628 10676 18668
rect 10842 18628 10882 18668
rect 11020 18628 11060 18668
rect 14659 18628 14699 18668
rect 17246 18628 17286 18668
rect 18796 18628 18836 18668
rect 19564 18628 19604 18668
rect 20131 18619 20171 18659
rect 21859 18628 21899 18668
rect 22444 18628 22484 18668
rect 30412 18628 30452 18668
rect 2659 18544 2699 18584
rect 3916 18544 3956 18584
rect 4204 18544 4244 18584
rect 4441 18544 4481 18584
rect 4972 18544 5012 18584
rect 5107 18544 5147 18584
rect 5740 18544 5780 18584
rect 5923 18544 5963 18584
rect 6148 18544 6188 18584
rect 6307 18544 6347 18584
rect 6424 18544 6464 18584
rect 6591 18533 6631 18573
rect 6691 18544 6731 18584
rect 6988 18544 7028 18584
rect 3043 18460 3083 18500
rect 7324 18502 7364 18542
rect 7562 18544 7602 18584
rect 7799 18544 7839 18584
rect 8044 18544 8084 18584
rect 8279 18544 8319 18584
rect 8524 18544 8564 18584
rect 8875 18544 8915 18584
rect 9100 18544 9140 18584
rect 9718 18544 9758 18584
rect 10531 18544 10571 18584
rect 11116 18544 11156 18584
rect 4108 18460 4148 18500
rect 4339 18451 4379 18491
rect 7459 18460 7499 18500
rect 7939 18460 7979 18500
rect 8419 18460 8459 18500
rect 10387 18502 10427 18542
rect 11353 18544 11393 18584
rect 11830 18544 11870 18584
rect 12268 18544 12308 18584
rect 12616 18544 12656 18584
rect 13459 18544 13499 18584
rect 13654 18544 13694 18584
rect 13956 18544 13996 18584
rect 14092 18544 14132 18584
rect 14327 18544 14367 18584
rect 14467 18544 14507 18584
rect 14572 18544 14612 18584
rect 14807 18544 14847 18584
rect 15052 18544 15092 18584
rect 15340 18544 15380 18584
rect 15532 18544 15572 18584
rect 15907 18544 15947 18584
rect 16012 18544 16052 18584
rect 16204 18544 16244 18584
rect 16696 18544 16736 18584
rect 16871 18544 16911 18584
rect 17068 18544 17108 18584
rect 17452 18544 17492 18584
rect 17548 18535 17588 18575
rect 17836 18544 17876 18584
rect 18358 18544 18398 18584
rect 18925 18544 18965 18584
rect 19180 18544 19220 18584
rect 19468 18544 19508 18584
rect 19660 18544 19700 18584
rect 19843 18544 19883 18584
rect 19948 18535 19988 18575
rect 20227 18544 20267 18584
rect 20404 18544 20444 18584
rect 20659 18544 20699 18584
rect 20762 18544 20802 18584
rect 21100 18544 21140 18584
rect 21292 18544 21332 18584
rect 21772 18544 21812 18584
rect 21955 18544 21995 18584
rect 22060 18544 22100 18584
rect 22243 18544 22283 18584
rect 22348 18544 22388 18584
rect 22554 18544 22594 18584
rect 22732 18544 22772 18584
rect 22963 18535 23003 18575
rect 23071 18544 23111 18584
rect 23596 18535 23636 18575
rect 23707 18535 23747 18575
rect 23827 18535 23867 18575
rect 24233 18544 24273 18584
rect 24556 18544 24596 18584
rect 24748 18544 24788 18584
rect 24863 18544 24903 18584
rect 25036 18544 25076 18584
rect 25228 18544 25268 18584
rect 25411 18544 25451 18584
rect 25603 18544 25643 18584
rect 25911 18544 25951 18584
rect 26188 18544 26228 18584
rect 26380 18544 26420 18584
rect 26860 18544 26900 18584
rect 27043 18544 27083 18584
rect 27148 18544 27188 18584
rect 29251 18544 29291 18584
rect 29635 18544 29675 18584
rect 29822 18544 29862 18584
rect 29932 18544 29972 18584
rect 30124 18544 30164 18584
rect 30316 18544 30356 18584
rect 30604 18544 30644 18584
rect 30787 18535 30827 18575
rect 8620 18460 8660 18500
rect 8995 18460 9035 18500
rect 10195 18460 10235 18500
rect 11251 18451 11291 18491
rect 11635 18460 11675 18500
rect 12796 18460 12836 18500
rect 14947 18460 14987 18500
rect 15148 18460 15188 18500
rect 16531 18460 16571 18500
rect 18163 18460 18203 18500
rect 24335 18460 24375 18500
rect 26083 18460 26123 18500
rect 27715 18460 27755 18500
rect 30940 18460 30980 18500
rect 5923 18376 5963 18416
rect 7180 18376 7220 18416
rect 12460 18376 12500 18416
rect 15724 18376 15764 18416
rect 18508 18376 18548 18416
rect 23980 18376 24020 18416
rect 24748 18376 24788 18416
rect 26956 18376 26996 18416
rect 29836 18376 29876 18416
rect 1132 18292 1172 18332
rect 3244 18292 3284 18332
rect 16972 18292 17012 18332
rect 22828 18292 22868 18332
rect 24460 18292 24500 18332
rect 25411 18292 25451 18332
rect 25900 18292 25940 18332
rect 27340 18292 27380 18332
rect 3112 18124 3480 18164
rect 10886 18124 11254 18164
rect 18660 18124 19028 18164
rect 26434 18124 26802 18164
rect 6316 17956 6356 17996
rect 6979 17956 7019 17996
rect 7555 17956 7595 17996
rect 11980 17956 12020 17996
rect 12748 17956 12788 17996
rect 22636 17956 22676 17996
rect 23500 17956 23540 17996
rect 24556 17956 24596 17996
rect 26179 17956 26219 17996
rect 27724 17956 27764 17996
rect 1996 17872 2036 17912
rect 2380 17872 2420 17912
rect 3724 17872 3764 17912
rect 4204 17872 4244 17912
rect 7180 17872 7220 17912
rect 9100 17872 9140 17912
rect 11500 17872 11540 17912
rect 20044 17872 20084 17912
rect 24787 17872 24827 17912
rect 2764 17788 2804 17828
rect 8572 17788 8612 17828
rect 9004 17788 9044 17828
rect 9571 17788 9611 17828
rect 9964 17788 10004 17828
rect 2284 17704 2324 17744
rect 2467 17704 2507 17744
rect 2572 17704 2612 17744
rect 2860 17704 2900 17744
rect 2979 17704 3019 17744
rect 3097 17704 3137 17744
rect 3427 17704 3467 17744
rect 3532 17704 3572 17744
rect 4396 17704 4436 17744
rect 4780 17704 4820 17744
rect 4899 17704 4939 17744
rect 5017 17704 5057 17744
rect 5262 17704 5302 17744
rect 5452 17704 5492 17744
rect 5764 17704 5804 17744
rect 5923 17704 5963 17744
rect 6067 17704 6107 17744
rect 6207 17715 6247 17755
rect 6333 17715 6373 17755
rect 6796 17704 6836 17744
rect 6965 17704 7005 17744
rect 7180 17704 7220 17744
rect 7372 17704 7412 17744
rect 7555 17704 7595 17744
rect 7673 17704 7713 17744
rect 7843 17695 7883 17735
rect 7979 17704 8019 17744
rect 8116 17704 8156 17744
rect 8371 17704 8411 17744
rect 8860 17704 8900 17744
rect 9175 17704 9215 17744
rect 9315 17704 9355 17744
rect 9436 17746 9476 17786
rect 11116 17788 11156 17828
rect 13635 17788 13675 17828
rect 14115 17788 14155 17828
rect 14467 17788 14507 17828
rect 15148 17788 15188 17828
rect 16147 17788 16187 17828
rect 18869 17788 18909 17828
rect 19084 17788 19124 17828
rect 20995 17788 21035 17828
rect 25612 17788 25652 17828
rect 9657 17704 9697 17744
rect 10648 17704 10688 17744
rect 10775 17704 10815 17744
rect 10915 17704 10955 17744
rect 11020 17704 11060 17744
rect 11500 17704 11540 17744
rect 11692 17704 11732 17744
rect 11873 17704 11913 17744
rect 12085 17704 12125 17744
rect 12268 17704 12308 17744
rect 12451 17704 12491 17744
rect 12652 17704 12692 17744
rect 12839 17677 12879 17717
rect 13036 17704 13076 17744
rect 13226 17704 13266 17744
rect 13516 17704 13556 17744
rect 13733 17704 13773 17744
rect 13996 17704 14036 17744
rect 14213 17704 14253 17744
rect 14327 17704 14367 17744
rect 14572 17704 14612 17744
rect 14807 17704 14847 17744
rect 14947 17704 14987 17744
rect 15052 17704 15092 17744
rect 15484 17704 15524 17744
rect 15619 17704 15659 17744
rect 15724 17704 15764 17744
rect 16312 17704 16352 17744
rect 16483 17704 16523 17744
rect 16776 17704 16816 17744
rect 16963 17704 17003 17744
rect 17081 17704 17121 17744
rect 17248 17704 17288 17744
rect 17355 17704 17395 17744
rect 17524 17704 17564 17744
rect 17836 17704 17876 17744
rect 18263 17704 18303 17744
rect 18389 17704 18429 17744
rect 18501 17704 18541 17744
rect 18743 17704 18783 17744
rect 19603 17746 19643 17786
rect 27715 17788 27755 17828
rect 28099 17788 28139 17828
rect 18988 17704 19028 17744
rect 20044 17704 20084 17744
rect 20169 17704 20209 17744
rect 20332 17704 20372 17744
rect 20515 17704 20555 17744
rect 20812 17704 20852 17744
rect 21676 17704 21716 17744
rect 21964 17704 22004 17744
rect 22156 17704 22196 17744
rect 22819 17704 22859 17744
rect 22924 17704 22964 17744
rect 23059 17704 23099 17744
rect 23212 17704 23252 17744
rect 23404 17704 23444 17744
rect 23526 17704 23566 17744
rect 23644 17704 23684 17744
rect 23743 17737 23783 17777
rect 23980 17704 24020 17744
rect 24172 17704 24212 17744
rect 24407 17704 24447 17744
rect 24547 17695 24587 17735
rect 24652 17704 24692 17744
rect 24988 17704 25028 17744
rect 25132 17704 25172 17744
rect 25708 17704 25748 17744
rect 25827 17704 25867 17744
rect 25939 17704 25979 17744
rect 26572 17704 26612 17744
rect 26851 17704 26891 17744
rect 27532 17704 27572 17744
rect 29635 17704 29675 17744
rect 30208 17704 30248 17744
rect 30688 17704 30728 17744
rect 4684 17620 4724 17660
rect 10483 17620 10523 17660
rect 13900 17620 13940 17660
rect 15811 17620 15851 17660
rect 16684 17620 16724 17660
rect 22051 17620 22091 17660
rect 30019 17620 30059 17660
rect 3436 17536 3476 17576
rect 5452 17536 5492 17576
rect 9763 17536 9803 17576
rect 10204 17536 10244 17576
rect 12364 17536 12404 17576
rect 13132 17536 13172 17576
rect 13420 17536 13460 17576
rect 14659 17536 14699 17576
rect 17443 17536 17483 17576
rect 17731 17536 17771 17576
rect 18019 17536 18059 17576
rect 18595 17536 18635 17576
rect 19411 17536 19451 17576
rect 20716 17536 20756 17576
rect 23980 17536 24020 17576
rect 26380 17536 26420 17576
rect 30364 17536 30404 17576
rect 30844 17536 30884 17576
rect 4352 17368 4720 17408
rect 12126 17368 12494 17408
rect 19900 17368 20268 17408
rect 27674 17368 28042 17408
rect 2179 17200 2219 17240
rect 3331 17200 3371 17240
rect 4291 17200 4331 17240
rect 4483 17200 4523 17240
rect 4963 17200 5003 17240
rect 8323 17200 8363 17240
rect 8803 17200 8843 17240
rect 12739 17200 12779 17240
rect 13891 17200 13931 17240
rect 15907 17200 15947 17240
rect 16300 17200 16340 17240
rect 16771 17200 16811 17240
rect 17725 17200 17765 17240
rect 18892 17200 18932 17240
rect 20611 17200 20651 17240
rect 21196 17200 21236 17240
rect 21955 17200 21995 17240
rect 25132 17200 25172 17240
rect 26173 17200 26213 17240
rect 27148 17200 27188 17240
rect 27532 17200 27572 17240
rect 29548 17200 29588 17240
rect 29731 17200 29771 17240
rect 30028 17200 30068 17240
rect 3043 17116 3083 17156
rect 3811 17116 3851 17156
rect 5251 17107 5291 17147
rect 6019 17107 6059 17147
rect 6700 17116 6740 17156
rect 10540 17116 10580 17156
rect 13612 17116 13652 17156
rect 14179 17107 14219 17147
rect 15715 17107 15755 17147
rect 18499 17116 18539 17156
rect 19660 17116 19700 17156
rect 21306 17116 21346 17156
rect 22636 17116 22676 17156
rect 26707 17116 26747 17156
rect 2284 17032 2324 17072
rect 3244 17032 3284 17072
rect 3479 17032 3519 17072
rect 3724 17032 3764 17072
rect 4204 17032 4244 17072
rect 4588 17032 4628 17072
rect 4963 17032 5003 17072
rect 5068 17023 5108 17063
rect 5347 17032 5387 17072
rect 5481 17032 5521 17072
rect 5742 17032 5782 17072
rect 5887 17032 5927 17072
rect 6115 17032 6155 17072
rect 6291 17032 6331 17072
rect 6499 17031 6539 17071
rect 6796 17032 6836 17072
rect 7075 17032 7115 17072
rect 7180 17023 7220 17063
rect 7324 17023 7364 17063
rect 7454 17032 7494 17072
rect 7636 17032 7676 17072
rect 7984 17032 8024 17072
rect 8154 17032 8194 17072
rect 8275 17032 8315 17072
rect 8396 17021 8436 17061
rect 8541 17021 8581 17061
rect 8740 17032 8780 17072
rect 8899 17032 8939 17072
rect 9016 17032 9056 17072
rect 9155 17032 9195 17072
rect 9283 17032 9323 17072
rect 9532 17032 9572 17072
rect 10003 17032 10043 17072
rect 10627 17032 10667 17072
rect 11020 17032 11060 17072
rect 9676 16990 9716 17030
rect 11512 17032 11552 17072
rect 11692 17032 11732 17072
rect 12067 17032 12107 17072
rect 12172 17032 12212 17072
rect 12547 17032 12587 17072
rect 12979 17032 13019 17072
rect 13516 17032 13556 17072
rect 13708 17032 13748 17072
rect 13891 17032 13931 17072
rect 13996 17023 14036 17063
rect 14275 17032 14315 17072
rect 14409 17032 14449 17072
rect 15256 17032 15296 17072
rect 15438 17032 15478 17072
rect 15532 17023 15572 17063
rect 15807 17032 15847 17072
rect 15988 17032 16028 17072
rect 16219 17032 16259 17072
rect 16396 17032 16436 17072
rect 16612 17032 16652 17072
rect 16771 17032 16811 17072
rect 16888 17032 16928 17072
rect 17020 17023 17060 17063
rect 17155 17032 17195 17072
rect 17356 17032 17396 17072
rect 17548 17032 17588 17072
rect 17827 17032 17867 17072
rect 17932 17023 17972 17063
rect 18398 17032 18438 17072
rect 18604 17032 18644 17072
rect 18700 17023 18740 17063
rect 18935 17032 18975 17072
rect 19075 17023 19115 17063
rect 19180 17032 19220 17072
rect 19468 17032 19508 17072
rect 19795 17032 19835 17072
rect 20260 17032 20300 17072
rect 20419 17032 20459 17072
rect 20536 17032 20576 17072
rect 20668 17023 20708 17063
rect 20803 17032 20843 17072
rect 20995 17032 21035 17072
rect 21100 17032 21140 17072
rect 21868 17032 21908 17072
rect 22156 17032 22196 17072
rect 22540 17032 22580 17072
rect 22828 17032 22868 17072
rect 23020 17032 23060 17072
rect 23359 17032 23399 17072
rect 23596 17032 23636 17072
rect 23788 17032 23828 17072
rect 24135 17032 24175 17072
rect 24259 17023 24299 17063
rect 24368 17032 24408 17072
rect 24652 17032 24692 17072
rect 24777 17032 24817 17072
rect 24940 17032 24980 17072
rect 25228 17032 25268 17072
rect 25465 17032 25505 17072
rect 25708 17032 25748 17072
rect 25830 17032 25870 17072
rect 25957 17032 25997 17072
rect 26275 17032 26315 17072
rect 26380 17023 26420 17063
rect 27052 17032 27092 17072
rect 27173 17032 27213 17072
rect 27575 17032 27615 17072
rect 27697 17032 27737 17072
rect 27820 17032 27860 17072
rect 28684 17032 28724 17072
rect 28876 17032 28916 17072
rect 29836 17032 29876 17072
rect 30220 17032 30260 17072
rect 3619 16948 3659 16988
rect 9868 16948 9908 16988
rect 11347 16948 11387 16988
rect 13180 16948 13220 16988
rect 15091 16948 15131 16988
rect 23242 16948 23282 16988
rect 23692 16948 23732 16988
rect 25363 16939 25403 16979
rect 4012 16864 4052 16904
rect 4780 16864 4820 16904
rect 9772 16864 9812 16904
rect 12519 16864 12559 16904
rect 18220 16864 18260 16904
rect 21484 16864 21524 16904
rect 23116 16864 23156 16904
rect 23404 16864 23444 16904
rect 24748 16864 24788 16904
rect 26851 16864 26891 16904
rect 30604 16864 30644 16904
rect 30988 16864 31028 16904
rect 2476 16780 2516 16820
rect 5731 16780 5771 16820
rect 7075 16780 7115 16820
rect 10540 16780 10580 16820
rect 12172 16780 12212 16820
rect 17452 16780 17492 16820
rect 19660 16780 19700 16820
rect 23980 16780 24020 16820
rect 25996 16780 26036 16820
rect 28012 16780 28052 16820
rect 30316 16780 30356 16820
rect 3112 16612 3480 16652
rect 10886 16612 11254 16652
rect 18660 16612 19028 16652
rect 26434 16612 26802 16652
rect 1516 16444 1556 16484
rect 3628 16444 3668 16484
rect 8524 16444 8564 16484
rect 8899 16444 8939 16484
rect 17260 16444 17300 16484
rect 24076 16444 24116 16484
rect 25411 16444 25451 16484
rect 27436 16444 27476 16484
rect 30796 16444 30836 16484
rect 5548 16360 5588 16400
rect 9292 16360 9332 16400
rect 15148 16360 15188 16400
rect 15724 16360 15764 16400
rect 16396 16360 16436 16400
rect 22252 16360 22292 16400
rect 25036 16360 25076 16400
rect 30316 16360 30356 16400
rect 4051 16267 4091 16307
rect 6700 16276 6740 16316
rect 9390 16276 9430 16316
rect 10444 16276 10484 16316
rect 10659 16276 10699 16316
rect 11116 16276 11156 16316
rect 12700 16276 12740 16316
rect 15052 16276 15092 16316
rect 15628 16276 15668 16316
rect 16492 16276 16532 16316
rect 16924 16276 16964 16316
rect 19276 16276 19316 16316
rect 19948 16276 19988 16316
rect 21868 16276 21908 16316
rect 25756 16276 25796 16316
rect 1420 16192 1460 16232
rect 1621 16165 1661 16205
rect 1843 16192 1883 16232
rect 2188 16192 2228 16232
rect 2755 16192 2795 16232
rect 2860 16192 2900 16232
rect 3436 16192 3476 16232
rect 3916 16192 3956 16232
rect 4153 16192 4193 16232
rect 4492 16192 4532 16232
rect 5356 16192 5396 16232
rect 5731 16192 5771 16232
rect 5875 16192 5915 16232
rect 5981 16192 6021 16232
rect 6101 16192 6141 16232
rect 6249 16192 6289 16232
rect 6796 16192 6836 16232
rect 6915 16192 6955 16232
rect 7033 16192 7073 16232
rect 7204 16192 7244 16232
rect 7363 16192 7403 16232
rect 7489 16192 7529 16232
rect 7646 16192 7686 16232
rect 7747 16192 7787 16232
rect 7987 16192 8027 16232
rect 8131 16192 8171 16232
rect 8248 16192 8288 16232
rect 8387 16192 8427 16232
rect 8515 16192 8555 16232
rect 8716 16192 8756 16232
rect 8899 16192 8939 16232
rect 9052 16192 9092 16232
rect 9217 16192 9257 16232
rect 9509 16192 9549 16232
rect 9692 16203 9732 16243
rect 9873 16192 9913 16232
rect 10003 16192 10043 16232
rect 10108 16192 10148 16232
rect 10243 16192 10283 16232
rect 10540 16192 10580 16232
rect 10777 16192 10817 16232
rect 11212 16192 11252 16232
rect 11331 16192 11371 16232
rect 11449 16192 11489 16232
rect 11596 16192 11636 16232
rect 11788 16192 11828 16232
rect 12544 16192 12584 16232
rect 13462 16192 13502 16232
rect 13612 16192 13652 16232
rect 13900 16192 13940 16232
rect 14275 16192 14315 16232
rect 14572 16192 14612 16232
rect 14908 16192 14948 16232
rect 15223 16192 15263 16232
rect 15363 16192 15403 16232
rect 15484 16192 15524 16232
rect 15785 16192 15825 16232
rect 15955 16192 15995 16232
rect 16156 16192 16196 16232
rect 16321 16192 16361 16232
rect 16613 16192 16653 16232
rect 16768 16192 16808 16232
rect 17452 16192 17492 16232
rect 17836 16192 17876 16232
rect 17975 16225 18015 16265
rect 18595 16192 18635 16232
rect 19372 16192 19412 16232
rect 19491 16192 19531 16232
rect 19606 16192 19646 16232
rect 20323 16192 20363 16232
rect 22387 16192 22427 16232
rect 22924 16192 22964 16232
rect 23116 16192 23156 16232
rect 23596 16192 23636 16232
rect 23788 16192 23828 16232
rect 24076 16192 24116 16232
rect 24268 16192 24308 16232
rect 24738 16192 24778 16232
rect 24931 16192 24971 16232
rect 25036 16225 25076 16265
rect 25411 16234 25451 16274
rect 26179 16276 26219 16316
rect 26380 16276 26420 16316
rect 28195 16276 28235 16316
rect 30115 16276 30155 16316
rect 25228 16192 25268 16232
rect 25600 16192 25640 16232
rect 26059 16192 26099 16232
rect 26284 16192 26324 16232
rect 26659 16183 26699 16223
rect 26956 16192 26996 16232
rect 27436 16192 27476 16232
rect 27628 16192 27668 16232
rect 29731 16192 29771 16232
rect 30700 16192 30740 16232
rect 30892 16192 30932 16232
rect 31073 16192 31113 16232
rect 31276 16192 31316 16232
rect 3820 16108 3860 16148
rect 4291 16108 4331 16148
rect 13708 16108 13748 16148
rect 22588 16108 22628 16148
rect 26764 16108 26804 16148
rect 2284 16024 2324 16064
rect 3148 16024 3188 16064
rect 3331 16024 3371 16064
rect 4579 16024 4619 16064
rect 5251 16024 5291 16064
rect 6211 16024 6251 16064
rect 7363 16024 7403 16064
rect 9763 16024 9803 16064
rect 11692 16024 11732 16064
rect 13267 16024 13307 16064
rect 14476 16024 14516 16064
rect 17539 16024 17579 16064
rect 18124 16024 18164 16064
rect 18796 16024 18836 16064
rect 23020 16024 23060 16064
rect 23596 16024 23636 16064
rect 27820 16024 27860 16064
rect 31084 16024 31124 16064
rect 4352 15856 4720 15896
rect 12126 15856 12494 15896
rect 19900 15856 20268 15896
rect 27674 15856 28042 15896
rect 1996 15688 2036 15728
rect 2365 15688 2405 15728
rect 3427 15688 3467 15728
rect 3907 15688 3947 15728
rect 7747 15730 7787 15770
rect 4108 15688 4148 15728
rect 5251 15688 5291 15728
rect 5443 15688 5483 15728
rect 7363 15688 7403 15728
rect 11779 15688 11819 15728
rect 13507 15688 13547 15728
rect 14284 15688 14324 15728
rect 3619 15604 3659 15644
rect 10936 15646 10976 15686
rect 15916 15688 15956 15728
rect 16771 15688 16811 15728
rect 18988 15688 19028 15728
rect 20524 15688 20564 15728
rect 20899 15688 20939 15728
rect 25228 15688 25268 15728
rect 27052 15688 27092 15728
rect 27427 15688 27467 15728
rect 29827 15688 29867 15728
rect 1603 15520 1643 15560
rect 1708 15520 1748 15560
rect 2467 15520 2507 15560
rect 2572 15511 2612 15551
rect 3095 15520 3135 15560
rect 3340 15520 3380 15560
rect 3820 15520 3860 15560
rect 4204 15478 4244 15518
rect 4323 15520 4363 15560
rect 4441 15520 4481 15560
rect 4588 15520 4628 15560
rect 4780 15520 4820 15560
rect 5164 15520 5204 15560
rect 5548 15520 5588 15560
rect 6316 15520 6356 15560
rect 7036 15520 7076 15560
rect 3235 15436 3275 15476
rect 6931 15478 6971 15518
rect 7171 15520 7211 15560
rect 7276 15520 7316 15560
rect 7784 15562 7824 15602
rect 9676 15604 9716 15644
rect 10291 15604 10331 15644
rect 11587 15595 11627 15635
rect 8083 15520 8123 15560
rect 8332 15520 8372 15560
rect 8524 15520 8564 15560
rect 9100 15520 9140 15560
rect 9292 15520 9332 15560
rect 9772 15520 9812 15560
rect 10009 15520 10049 15560
rect 10456 15520 10496 15560
rect 10701 15520 10741 15560
rect 4684 15436 4724 15476
rect 6739 15436 6779 15476
rect 10856 15478 10896 15518
rect 11141 15520 11181 15560
rect 11299 15520 11339 15560
rect 11404 15511 11444 15551
rect 11683 15520 11723 15560
rect 11860 15520 11900 15560
rect 12364 15520 12404 15560
rect 12601 15520 12641 15560
rect 12892 15520 12932 15560
rect 13200 15562 13240 15602
rect 13795 15595 13835 15635
rect 14947 15595 14987 15635
rect 15388 15604 15428 15644
rect 21484 15604 21524 15644
rect 22531 15604 22571 15644
rect 13363 15520 13403 15560
rect 13507 15520 13547 15560
rect 13612 15511 13652 15551
rect 13891 15520 13931 15560
rect 14037 15520 14077 15560
rect 14273 15520 14313 15560
rect 14476 15520 14516 15560
rect 14659 15520 14699 15560
rect 14764 15511 14804 15551
rect 15043 15520 15083 15560
rect 15220 15520 15260 15560
rect 15916 15520 15956 15560
rect 16106 15520 16146 15560
rect 16420 15520 16460 15560
rect 16579 15520 16619 15560
rect 16696 15520 16736 15560
rect 16867 15520 16907 15560
rect 16972 15509 17012 15549
rect 17251 15520 17291 15560
rect 17356 15520 17396 15560
rect 17740 15520 17780 15560
rect 18316 15511 18356 15551
rect 18796 15511 18836 15551
rect 19564 15520 19604 15560
rect 19673 15520 19713 15560
rect 19948 15520 19988 15560
rect 20236 15520 20276 15560
rect 20378 15520 20418 15560
rect 21004 15520 21044 15560
rect 21388 15520 21428 15560
rect 21571 15520 21611 15560
rect 21955 15520 21995 15560
rect 22060 15520 22100 15560
rect 22915 15520 22955 15560
rect 25492 15520 25532 15560
rect 25603 15520 25643 15560
rect 26044 15520 26084 15560
rect 7948 15436 7988 15476
rect 9907 15427 9947 15467
rect 11020 15436 11060 15476
rect 12268 15436 12308 15476
rect 12499 15427 12539 15467
rect 13036 15436 13076 15476
rect 15628 15436 15668 15476
rect 25389 15478 25429 15518
rect 26188 15520 26228 15560
rect 26764 15520 26804 15560
rect 26899 15520 26939 15560
rect 27013 15520 27053 15560
rect 27532 15520 27572 15560
rect 27916 15520 27956 15560
rect 28780 15520 28820 15560
rect 28972 15520 29012 15560
rect 30124 15520 30164 15560
rect 30595 15511 30635 15551
rect 17836 15436 17876 15476
rect 30034 15436 30074 15476
rect 30748 15436 30788 15476
rect 6460 15352 6500 15392
rect 7852 15352 7892 15392
rect 13132 15352 13172 15392
rect 25843 15352 25883 15392
rect 26380 15352 26420 15392
rect 31084 15352 31124 15392
rect 2860 15268 2900 15308
rect 4972 15268 5012 15308
rect 5740 15268 5780 15308
rect 8332 15268 8372 15308
rect 9100 15268 9140 15308
rect 14659 15268 14699 15308
rect 19276 15268 19316 15308
rect 21196 15268 21236 15308
rect 22243 15268 22283 15308
rect 24460 15268 24500 15308
rect 24844 15268 24884 15308
rect 28108 15268 28148 15308
rect 29644 15268 29684 15308
rect 3112 15100 3480 15140
rect 10886 15100 11254 15140
rect 18660 15100 19028 15140
rect 26434 15100 26802 15140
rect 1948 14932 1988 14972
rect 4195 14932 4235 14972
rect 10339 14932 10379 14972
rect 12547 14932 12587 14972
rect 13516 14932 13556 14972
rect 16684 14932 16724 14972
rect 19660 14932 19700 14972
rect 23116 14932 23156 14972
rect 24940 14932 24980 14972
rect 25228 14932 25268 14972
rect 27628 14932 27668 14972
rect 30700 14932 30740 14972
rect 3980 14839 4020 14879
rect 8103 14848 8143 14888
rect 8716 14848 8756 14888
rect 11660 14839 11700 14879
rect 15043 14848 15083 14888
rect 16012 14848 16052 14888
rect 18316 14848 18356 14888
rect 20620 14848 20660 14888
rect 21187 14848 21227 14888
rect 21868 14848 21908 14888
rect 24067 14848 24107 14888
rect 25900 14848 25940 14888
rect 30988 14848 31028 14888
rect 7084 14764 7124 14804
rect 7315 14755 7355 14795
rect 1324 14680 1364 14720
rect 1612 14680 1652 14720
rect 2092 14680 2132 14720
rect 2284 14680 2324 14720
rect 3244 14680 3284 14720
rect 3340 14680 3380 14720
rect 4003 14680 4043 14720
rect 4588 14680 4628 14720
rect 4963 14680 5003 14720
rect 5068 14691 5108 14731
rect 5251 14671 5291 14711
rect 5386 14680 5426 14720
rect 5524 14680 5564 14720
rect 5932 14691 5972 14731
rect 6079 14680 6119 14720
rect 6207 14680 6247 14720
rect 6307 14680 6347 14720
rect 6484 14691 6524 14731
rect 8648 14722 8688 14762
rect 8812 14764 8852 14804
rect 9603 14764 9643 14804
rect 12076 14764 12116 14804
rect 12291 14764 12331 14804
rect 14803 14792 14843 14832
rect 21091 14764 21131 14804
rect 21667 14764 21707 14804
rect 25057 14764 25097 14804
rect 25420 14764 25460 14804
rect 25635 14764 25675 14804
rect 26755 14764 26795 14804
rect 28483 14764 28523 14804
rect 7180 14680 7220 14720
rect 7417 14680 7457 14720
rect 7552 14680 7592 14720
rect 8145 14680 8185 14720
rect 8493 14680 8533 14720
rect 8947 14680 8987 14720
rect 9484 14680 9524 14720
rect 9701 14680 9741 14720
rect 9859 14680 9899 14720
rect 10156 14680 10196 14720
rect 10339 14680 10379 14720
rect 10483 14680 10523 14720
rect 10617 14680 10657 14720
rect 10718 14680 10758 14720
rect 10900 14680 10940 14720
rect 11683 14680 11723 14720
rect 11884 14680 11924 14720
rect 12172 14680 12212 14720
rect 12409 14680 12449 14720
rect 12832 14687 12872 14727
rect 12932 14680 12972 14720
rect 13324 14680 13364 14720
rect 13891 14680 13931 14720
rect 13996 14691 14036 14731
rect 14141 14680 14181 14720
rect 14270 14680 14310 14720
rect 14452 14680 14492 14720
rect 14851 14680 14891 14720
rect 15244 14680 15284 14720
rect 15436 14680 15476 14720
rect 16012 14680 16052 14720
rect 16204 14680 16244 14720
rect 16492 14680 16532 14720
rect 16876 14680 16916 14720
rect 17068 14680 17108 14720
rect 18508 14680 18548 14720
rect 18700 14680 18740 14720
rect 18988 14680 19028 14720
rect 19267 14662 19307 14702
rect 19948 14680 19988 14720
rect 20227 14680 20267 14720
rect 21475 14680 21515 14720
rect 21868 14680 21908 14720
rect 22156 14680 22196 14720
rect 22444 14680 22484 14720
rect 23491 14680 23531 14720
rect 23596 14680 23636 14720
rect 24460 14680 24500 14720
rect 24844 14680 24884 14720
rect 25175 14713 25215 14753
rect 25516 14680 25556 14720
rect 25750 14680 25790 14720
rect 25921 14680 25961 14720
rect 26188 14680 26228 14720
rect 26380 14680 26420 14720
rect 26615 14680 26655 14720
rect 26860 14680 26900 14720
rect 27340 14680 27380 14720
rect 27436 14680 27476 14720
rect 27628 14680 27668 14720
rect 27817 14680 27857 14720
rect 30019 14680 30059 14720
rect 30604 14680 30644 14720
rect 30796 14680 30836 14720
rect 3038 14596 3078 14636
rect 9388 14596 9428 14636
rect 10060 14596 10100 14636
rect 19372 14596 19412 14636
rect 20332 14596 20372 14636
rect 23779 14596 23819 14636
rect 26947 14596 26987 14636
rect 27134 14596 27174 14636
rect 28099 14596 28139 14636
rect 30403 14596 30443 14636
rect 2092 14512 2132 14552
rect 3139 14512 3179 14552
rect 4483 14512 4523 14552
rect 4780 14512 4820 14552
rect 5164 14512 5204 14552
rect 6403 14512 6443 14552
rect 7708 14512 7748 14552
rect 8323 14512 8363 14552
rect 13219 14512 13259 14552
rect 14371 14512 14411 14552
rect 15340 14512 15380 14552
rect 13075 14470 13115 14510
rect 16387 14512 16427 14552
rect 16972 14512 17012 14552
rect 18691 14512 18731 14552
rect 23500 14512 23540 14552
rect 27235 14512 27275 14552
rect 4352 14344 4720 14384
rect 12126 14344 12494 14384
rect 19900 14344 20268 14384
rect 27674 14344 28042 14384
rect 1555 14176 1595 14216
rect 2092 14176 2132 14216
rect 3628 14176 3668 14216
rect 4003 14176 4043 14216
rect 5443 14176 5483 14216
rect 5827 14176 5867 14216
rect 6172 14176 6212 14216
rect 7747 14176 7787 14216
rect 9772 14176 9812 14216
rect 10051 14176 10091 14216
rect 13219 14176 13259 14216
rect 13516 14176 13556 14216
rect 15907 14176 15947 14216
rect 16588 14176 16628 14216
rect 21196 14176 21236 14216
rect 23884 14176 23924 14216
rect 29644 14176 29684 14216
rect 30844 14176 30884 14216
rect 5251 14083 5291 14123
rect 10819 14092 10859 14132
rect 11116 14092 11156 14132
rect 13900 14092 13940 14132
rect 1036 14008 1076 14048
rect 1219 14008 1259 14048
rect 1720 14008 1760 14048
rect 1891 14008 1931 14048
rect 2188 14008 2228 14048
rect 2563 14008 2603 14048
rect 2668 14008 2708 14048
rect 3148 14008 3188 14048
rect 3436 14008 3476 14048
rect 4300 14008 4340 14048
rect 4963 14008 5003 14048
rect 5068 13999 5108 14039
rect 5343 14008 5383 14048
rect 5524 14008 5564 14048
rect 5729 14008 5769 14048
rect 5932 14008 5972 14048
rect 6028 13999 6068 14039
rect 7075 14008 7115 14048
rect 7180 14008 7220 14048
rect 7684 14008 7724 14048
rect 7821 14008 7861 14048
rect 7987 14008 8027 14048
rect 8131 14008 8171 14048
rect 8253 14008 8293 14048
rect 8812 14008 8852 14048
rect 8995 14008 9035 14048
rect 9100 14008 9140 14048
rect 9292 14008 9332 14048
rect 9417 14008 9457 14048
rect 9580 14008 9620 14048
rect 9964 14008 10004 14048
rect 10487 14008 10527 14048
rect 10713 14008 10753 14048
rect 11020 14008 11060 14048
rect 11587 14050 11627 14090
rect 14010 14092 14050 14132
rect 15809 14092 15849 14132
rect 21379 14092 21419 14132
rect 29212 14092 29252 14132
rect 11212 14008 11252 14048
rect 11713 14008 11753 14048
rect 12005 14008 12045 14048
rect 12364 14008 12404 14048
rect 12556 14008 12596 14048
rect 12743 14027 12783 14067
rect 12940 14008 12980 14048
rect 13324 14008 13364 14048
rect 13699 14008 13739 14048
rect 13804 14008 13844 14048
rect 14284 14008 14324 14048
rect 14473 14008 14513 14048
rect 14620 14008 14660 14048
rect 4210 13924 4250 13964
rect 6412 13924 6452 13964
rect 10613 13924 10653 13964
rect 11884 13924 11924 13964
rect 12844 13924 12884 13964
rect 14764 13966 14804 14006
rect 15077 14008 15117 14048
rect 15436 14008 15476 14048
rect 15625 14008 15665 14048
rect 16012 14008 16052 14048
rect 16114 14005 16154 14045
rect 16771 14008 16811 14048
rect 17260 13999 17300 14039
rect 17740 14008 17780 14048
rect 18220 14008 18260 14048
rect 18338 14008 18378 14048
rect 18691 14008 18731 14048
rect 19852 14008 19892 14048
rect 19961 14008 20001 14048
rect 20236 14008 20276 14048
rect 20524 14008 20564 14048
rect 21571 14008 21611 14048
rect 22060 13999 22100 14039
rect 22540 14008 22580 14048
rect 23020 14008 23060 14048
rect 23133 13989 23173 14029
rect 23404 14008 23444 14048
rect 23788 14008 23828 14048
rect 26179 14008 26219 14048
rect 27043 14008 27083 14048
rect 27148 14008 27188 14048
rect 27619 14008 27659 14048
rect 27916 14008 27956 14048
rect 28195 14008 28235 14048
rect 28876 14008 28916 14048
rect 29032 14008 29072 14048
rect 29548 14008 29588 14048
rect 29739 14008 29779 14048
rect 30121 14008 30161 14048
rect 14956 13924 14996 13964
rect 17836 13924 17876 13964
rect 29932 13966 29972 14006
rect 22636 13924 22676 13964
rect 24643 13924 24683 13964
rect 26563 13924 26603 13964
rect 31084 13924 31124 13964
rect 2851 13840 2891 13880
rect 8908 13840 8948 13880
rect 9292 13840 9332 13880
rect 11788 13840 11828 13880
rect 12364 13840 12404 13880
rect 14860 13840 14900 13880
rect 27916 13840 27956 13880
rect 30316 13840 30356 13880
rect 1219 13756 1259 13796
rect 7363 13756 7403 13796
rect 14284 13756 14324 13796
rect 15436 13756 15476 13796
rect 19084 13756 19124 13796
rect 19564 13756 19604 13796
rect 24268 13756 24308 13796
rect 27331 13756 27371 13796
rect 29932 13756 29972 13796
rect 3112 13588 3480 13628
rect 10886 13588 11254 13628
rect 18660 13588 19028 13628
rect 26434 13588 26802 13628
rect 8131 13420 8171 13460
rect 9571 13420 9611 13460
rect 10339 13420 10379 13460
rect 12748 13420 12788 13460
rect 14275 13420 14315 13460
rect 15244 13420 15284 13460
rect 19852 13420 19892 13460
rect 21100 13420 21140 13460
rect 23491 13420 23531 13460
rect 24460 13420 24500 13460
rect 25804 13420 25844 13460
rect 27820 13420 27860 13460
rect 11875 13336 11915 13376
rect 21484 13336 21524 13376
rect 24076 13336 24116 13376
rect 30796 13336 30836 13376
rect 2083 13252 2123 13292
rect 2284 13252 2324 13292
rect 5740 13252 5780 13292
rect 5971 13243 6011 13283
rect 6787 13252 6827 13292
rect 6988 13252 7028 13292
rect 8899 13252 8939 13292
rect 9100 13252 9140 13292
rect 1558 13168 1598 13208
rect 1943 13168 1983 13208
rect 2188 13168 2228 13208
rect 3043 13168 3083 13208
rect 3148 13168 3188 13208
rect 4300 13168 4340 13208
rect 4435 13168 4475 13208
rect 4804 13168 4844 13208
rect 4977 13168 5017 13208
rect 5089 13168 5129 13208
rect 5251 13179 5291 13219
rect 5373 13168 5413 13208
rect 5836 13168 5876 13208
rect 6076 13168 6116 13208
rect 6215 13168 6255 13208
rect 6403 13168 6443 13208
rect 6647 13168 6687 13208
rect 6892 13168 6932 13208
rect 7468 13168 7508 13208
rect 7651 13168 7691 13208
rect 7756 13168 7796 13208
rect 8416 13201 8456 13241
rect 8515 13168 8555 13208
rect 8759 13168 8799 13208
rect 9004 13168 9044 13208
rect 9868 13168 9908 13208
rect 10624 13201 10664 13241
rect 11539 13243 11579 13283
rect 13708 13252 13748 13292
rect 14764 13252 14804 13292
rect 16035 13252 16075 13292
rect 16387 13252 16427 13292
rect 17932 13252 17972 13292
rect 10723 13168 10763 13208
rect 11404 13168 11444 13208
rect 11641 13168 11681 13208
rect 12268 13168 12308 13208
rect 12931 13168 12971 13208
rect 13228 13168 13268 13208
rect 13795 13168 13835 13208
rect 14270 13168 14310 13208
rect 14572 13168 14612 13208
rect 14860 13168 14900 13208
rect 14979 13168 15019 13208
rect 15097 13168 15137 13208
rect 15244 13168 15284 13208
rect 15369 13168 15409 13208
rect 15532 13168 15572 13208
rect 15916 13168 15956 13208
rect 16156 13210 16196 13250
rect 26419 13252 26459 13292
rect 26908 13252 26948 13292
rect 29731 13252 29771 13292
rect 16267 13168 16307 13208
rect 16492 13168 16532 13208
rect 16963 13168 17003 13208
rect 17452 13168 17492 13208
rect 18028 13168 18068 13208
rect 18412 13168 18452 13208
rect 18513 13168 18553 13208
rect 19180 13168 19220 13208
rect 19459 13168 19499 13208
rect 20428 13168 20468 13208
rect 20524 13159 20564 13199
rect 20812 13168 20852 13208
rect 21100 13168 21140 13208
rect 21292 13168 21332 13208
rect 21772 13168 21812 13208
rect 21868 13159 21908 13199
rect 22156 13168 22196 13208
rect 22444 13168 22484 13208
rect 23452 13168 23492 13208
rect 23596 13168 23636 13208
rect 25132 13168 25172 13208
rect 25315 13168 25355 13208
rect 25804 13168 25844 13208
rect 25929 13168 25969 13208
rect 26092 13168 26132 13208
rect 26584 13168 26624 13208
rect 26752 13168 26792 13208
rect 29347 13168 29387 13208
rect 29875 13168 29915 13208
rect 30412 13168 30452 13208
rect 30604 13168 30644 13208
rect 31180 13168 31220 13208
rect 7166 13084 7206 13124
rect 7267 13084 7307 13124
rect 7962 13084 8002 13124
rect 9566 13084 9606 13124
rect 11308 13084 11348 13124
rect 11971 13084 12011 13124
rect 12748 13084 12788 13124
rect 14476 13084 14516 13124
rect 15820 13084 15860 13124
rect 16579 13084 16619 13124
rect 19564 13084 19604 13124
rect 25623 13084 25663 13124
rect 27427 13084 27467 13124
rect 1363 13000 1403 13040
rect 3436 13000 3476 13040
rect 4588 13000 4628 13040
rect 4867 13000 4907 13040
rect 6316 13000 6356 13040
rect 7372 13000 7412 13040
rect 7852 13000 7892 13040
rect 8658 13000 8698 13040
rect 9772 13000 9812 13040
rect 10843 13000 10883 13040
rect 13411 13000 13451 13040
rect 13612 13000 13652 13040
rect 16780 13000 16820 13040
rect 20092 13000 20132 13040
rect 23116 13000 23156 13040
rect 25411 13000 25451 13040
rect 25516 13000 25556 13040
rect 30076 13000 30116 13040
rect 30595 13000 30635 13040
rect 4352 12832 4720 12872
rect 12126 12832 12494 12872
rect 19900 12832 20268 12872
rect 27674 12832 28042 12872
rect 1228 12664 1268 12704
rect 1996 12664 2036 12704
rect 2380 12664 2420 12704
rect 4291 12664 4331 12704
rect 4579 12664 4619 12704
rect 5932 12664 5972 12704
rect 6316 12664 6356 12704
rect 7564 12664 7604 12704
rect 9571 12664 9611 12704
rect 11011 12664 11051 12704
rect 11500 12664 11540 12704
rect 12796 12664 12836 12704
rect 13708 12664 13748 12704
rect 15052 12664 15092 12704
rect 15739 12664 15779 12704
rect 16012 12664 16052 12704
rect 17020 12664 17060 12704
rect 18691 12664 18731 12704
rect 20236 12664 20276 12704
rect 29740 12664 29780 12704
rect 2490 12580 2530 12620
rect 2947 12580 2987 12620
rect 9859 12571 9899 12611
rect 16723 12580 16763 12620
rect 18796 12580 18836 12620
rect 30124 12580 30164 12620
rect 940 12496 980 12536
rect 1075 12496 1115 12536
rect 1603 12496 1643 12536
rect 1708 12496 1748 12536
rect 2179 12496 2219 12536
rect 2284 12496 2324 12536
rect 2615 12496 2655 12536
rect 2860 12496 2900 12536
rect 3959 12496 3999 12536
rect 4099 12496 4139 12536
rect 4204 12496 4244 12536
rect 4780 12496 4820 12536
rect 5068 12496 5108 12536
rect 5260 12496 5300 12536
rect 5452 12496 5492 12536
rect 5836 12496 5876 12536
rect 6019 12496 6059 12536
rect 6231 12496 6271 12536
rect 6403 12496 6443 12536
rect 7084 12496 7124 12536
rect 7468 12496 7508 12536
rect 8323 12496 8363 12536
rect 8668 12496 8708 12536
rect 8969 12496 9009 12536
rect 9139 12496 9179 12536
rect 9571 12496 9611 12536
rect 9676 12487 9716 12527
rect 9951 12496 9991 12536
rect 10132 12485 10172 12525
rect 10348 12496 10388 12536
rect 10463 12496 10503 12536
rect 10636 12496 10676 12536
rect 11164 12496 11204 12536
rect 11308 12496 11348 12536
rect 11596 12496 11636 12536
rect 11833 12496 11873 12536
rect 11980 12496 12020 12536
rect 12172 12496 12212 12536
rect 12616 12496 12656 12536
rect 13084 12496 13124 12536
rect 13420 12496 13460 12536
rect 13804 12496 13844 12536
rect 14041 12496 14081 12536
rect 14659 12496 14699 12536
rect 14764 12496 14804 12536
rect 15520 12487 15560 12527
rect 15916 12496 15956 12536
rect 2755 12412 2795 12452
rect 7939 12412 7979 12452
rect 8515 12412 8555 12452
rect 15619 12454 15659 12494
rect 16108 12496 16148 12536
rect 16918 12496 16958 12536
rect 17164 12496 17204 12536
rect 17879 12496 17919 12536
rect 18124 12496 18164 12536
rect 18590 12496 18630 12536
rect 18892 12487 18932 12527
rect 19660 12496 19700 12536
rect 22147 12496 22187 12536
rect 23062 12496 23102 12536
rect 25411 12496 25451 12536
rect 25996 12496 26036 12536
rect 26188 12496 26228 12536
rect 26755 12496 26795 12536
rect 29644 12496 29684 12536
rect 29817 12496 29857 12536
rect 30028 12496 30068 12536
rect 30220 12496 30260 12536
rect 8812 12412 8852 12452
rect 11731 12403 11771 12443
rect 13923 12412 13963 12452
rect 18019 12412 18059 12452
rect 18220 12412 18260 12452
rect 19570 12412 19610 12452
rect 20611 12412 20651 12452
rect 22531 12412 22571 12452
rect 22867 12412 22907 12452
rect 23875 12412 23915 12452
rect 25795 12412 25835 12452
rect 26380 12412 26420 12452
rect 28300 12412 28340 12452
rect 8035 12328 8075 12368
rect 8908 12328 8948 12368
rect 10348 12328 10388 12368
rect 11980 12328 12020 12368
rect 15235 12328 15275 12368
rect 20236 12328 20276 12368
rect 25996 12328 26036 12368
rect 28876 12328 28916 12368
rect 29260 12328 29300 12368
rect 30508 12328 30548 12368
rect 30892 12328 30932 12368
rect 5260 12244 5300 12284
rect 13219 12244 13259 12284
rect 19468 12244 19508 12284
rect 23500 12244 23540 12284
rect 28684 12244 28724 12284
rect 3112 12076 3480 12116
rect 10886 12076 11254 12116
rect 18660 12076 19028 12116
rect 26434 12076 26802 12116
rect 1420 11908 1460 11948
rect 2284 11908 2324 11948
rect 4780 11908 4820 11948
rect 5644 11908 5684 11948
rect 6604 11908 6644 11948
rect 9475 11908 9515 11948
rect 10060 11908 10100 11948
rect 11779 11908 11819 11948
rect 12931 11908 12971 11948
rect 15340 11908 15380 11948
rect 16099 11908 16139 11948
rect 17356 11908 17396 11948
rect 18115 11908 18155 11948
rect 18595 11908 18635 11948
rect 20428 11908 20468 11948
rect 21676 11908 21716 11948
rect 23491 11908 23531 11948
rect 24076 11908 24116 11948
rect 27148 11908 27188 11948
rect 28588 11908 28628 11948
rect 29155 11908 29195 11948
rect 30316 11908 30356 11948
rect 30700 11908 30740 11948
rect 3340 11824 3380 11864
rect 6124 11824 6164 11864
rect 7267 11824 7307 11864
rect 21964 11824 22004 11864
rect 24316 11815 24356 11855
rect 29356 11824 29396 11864
rect 30988 11824 31028 11864
rect 1996 11740 2036 11780
rect 7762 11740 7802 11780
rect 10588 11740 10628 11780
rect 940 11656 980 11696
rect 1123 11656 1163 11696
rect 1323 11656 1363 11696
rect 1515 11656 1555 11696
rect 1660 11656 1700 11696
rect 1795 11656 1835 11696
rect 1900 11656 1940 11696
rect 2188 11656 2228 11696
rect 2380 11656 2420 11696
rect 2668 11656 2708 11696
rect 3148 11656 3188 11696
rect 3532 11656 3572 11696
rect 3916 11656 3956 11696
rect 4387 11656 4427 11696
rect 4496 11689 4536 11729
rect 4972 11656 5012 11696
rect 5164 11656 5204 11696
rect 5347 11656 5387 11696
rect 5932 11656 5972 11696
rect 6307 11656 6347 11696
rect 6979 11656 7019 11696
rect 7084 11656 7124 11696
rect 8659 11698 8699 11738
rect 12499 11731 12539 11771
rect 12946 11740 12986 11780
rect 13603 11740 13643 11780
rect 15916 11740 15956 11780
rect 19219 11740 19259 11780
rect 19987 11740 20027 11780
rect 20530 11740 20570 11780
rect 7852 11656 7892 11696
rect 8800 11656 8840 11696
rect 9292 11656 9332 11696
rect 9475 11656 9515 11696
rect 9859 11656 9899 11696
rect 9964 11656 10004 11696
rect 10432 11656 10472 11696
rect 11020 11656 11060 11696
rect 11308 11656 11348 11696
rect 12076 11656 12116 11696
rect 12364 11656 12404 11696
rect 12601 11656 12641 11696
rect 13036 11656 13076 11696
rect 13483 11656 13523 11696
rect 13708 11656 13748 11696
rect 14476 11656 14516 11696
rect 14572 11656 14612 11696
rect 14831 11656 14871 11696
rect 14961 11656 15001 11696
rect 15091 11656 15131 11696
rect 15235 11656 15275 11696
rect 15357 11656 15397 11696
rect 15575 11656 15615 11696
rect 15715 11656 15755 11696
rect 15820 11656 15860 11696
rect 16110 11656 16150 11696
rect 16217 11656 16257 11696
rect 16357 11656 16397 11696
rect 16483 11656 16523 11696
rect 16660 11656 16700 11696
rect 16963 11656 17003 11696
rect 17068 11677 17108 11717
rect 17548 11656 17588 11696
rect 17731 11656 17771 11696
rect 18414 11656 18454 11696
rect 20179 11698 20219 11738
rect 21244 11740 21284 11780
rect 25603 11740 25643 11780
rect 27250 11740 27290 11780
rect 18796 11656 18836 11696
rect 18892 11656 18932 11696
rect 19384 11656 19424 11696
rect 20620 11656 20660 11696
rect 21043 11656 21083 11696
rect 21772 11656 21812 11696
rect 22828 11656 22868 11696
rect 23116 11656 23156 11696
rect 23308 11656 23348 11696
rect 23491 11656 23531 11696
rect 24259 11656 24299 11696
rect 25132 11656 25172 11696
rect 25996 11656 26036 11696
rect 26476 11656 26516 11696
rect 26860 11656 26900 11696
rect 27340 11656 27380 11696
rect 27964 11656 28004 11696
rect 28108 11656 28148 11696
rect 28588 11656 28628 11696
rect 28780 11656 28820 11696
rect 28972 11656 29012 11696
rect 29141 11656 29181 11696
rect 29356 11656 29396 11696
rect 29548 11656 29588 11696
rect 29740 11656 29780 11696
rect 29932 11656 29972 11696
rect 30220 11656 30260 11696
rect 30412 11656 30452 11696
rect 30604 11656 30644 11696
rect 30796 11656 30836 11696
rect 2284 11572 2324 11612
rect 5068 11572 5108 11612
rect 5452 11572 5492 11612
rect 5658 11572 5698 11612
rect 6412 11572 6452 11612
rect 6618 11572 6658 11612
rect 11777 11572 11817 11612
rect 13795 11572 13835 11612
rect 14271 11572 14311 11612
rect 14371 11572 14411 11612
rect 17644 11572 17684 11612
rect 18110 11572 18150 11612
rect 18590 11572 18630 11612
rect 22492 11572 22532 11612
rect 29836 11572 29876 11612
rect 1036 11488 1076 11528
rect 2563 11488 2603 11528
rect 2860 11488 2900 11528
rect 3043 11488 3083 11528
rect 4012 11488 4052 11528
rect 4291 11479 4331 11519
rect 5827 11488 5867 11528
rect 7555 11488 7595 11528
rect 8467 11488 8507 11528
rect 8956 11488 8996 11528
rect 11500 11488 11540 11528
rect 11980 11488 12020 11528
rect 12268 11488 12308 11528
rect 16867 11479 16907 11519
rect 18316 11488 18356 11528
rect 24940 11488 24980 11528
rect 26371 11488 26411 11528
rect 27811 11488 27851 11528
rect 4352 11320 4720 11360
rect 12126 11320 12494 11360
rect 19900 11320 20268 11360
rect 27674 11320 28042 11360
rect 1804 11152 1844 11192
rect 3811 11194 3851 11234
rect 2764 11152 2804 11192
rect 5155 11152 5195 11192
rect 5923 11152 5963 11192
rect 7660 11152 7700 11192
rect 8428 11152 8468 11192
rect 9475 11152 9515 11192
rect 10051 11152 10091 11192
rect 10732 11152 10772 11192
rect 11308 11152 11348 11192
rect 11884 11152 11924 11192
rect 13324 11152 13364 11192
rect 13603 11152 13643 11192
rect 14476 11152 14516 11192
rect 15820 11152 15860 11192
rect 18403 11152 18443 11192
rect 18796 11152 18836 11192
rect 21091 11152 21131 11192
rect 22579 11152 22619 11192
rect 24364 11152 24404 11192
rect 25411 11152 25451 11192
rect 26668 11152 26708 11192
rect 27139 11152 27179 11192
rect 29356 11152 29396 11192
rect 29644 11152 29684 11192
rect 30124 11152 30164 11192
rect 940 11068 980 11108
rect 14275 11068 14315 11108
rect 15340 11068 15380 11108
rect 17836 11068 17876 11108
rect 18508 11068 18548 11108
rect 23356 11068 23396 11108
rect 24259 11068 24299 11108
rect 844 10984 884 11024
rect 1036 10984 1076 11024
rect 1411 10984 1451 11024
rect 1516 10984 1556 11024
rect 2476 10984 2516 11024
rect 2611 10984 2651 11024
rect 3139 10984 3179 11024
rect 3244 10984 3284 11024
rect 3841 10984 3881 11024
rect 4147 10984 4187 11024
rect 4843 10984 4883 11024
rect 5068 10984 5108 11024
rect 5591 10984 5631 11024
rect 5836 10984 5876 11024
rect 6700 10984 6740 11024
rect 6883 10984 6923 11024
rect 7036 10984 7076 11024
rect 7201 10984 7241 11024
rect 7493 10984 7533 11024
rect 7756 10984 7796 11024
rect 7973 10984 8013 11024
rect 8524 10984 8564 11024
rect 8761 10984 8801 11024
rect 9580 10984 9620 11024
rect 9955 10984 9995 11024
rect 10266 10984 10306 11024
rect 10444 10984 10484 11024
rect 10583 10984 10623 11024
rect 11404 10984 11444 11024
rect 11539 10975 11579 11015
rect 11641 10984 11681 11024
rect 11788 10984 11828 11024
rect 11980 10984 12020 11024
rect 12211 10984 12251 11024
rect 12931 10984 12971 11024
rect 13036 10984 13076 11024
rect 13505 10984 13545 11024
rect 13708 10984 13748 11024
rect 13804 10975 13844 11015
rect 13943 10984 13983 11024
rect 14188 10984 14228 11024
rect 14476 10984 14516 11024
rect 14668 10984 14708 11024
rect 14860 10984 14900 11024
rect 15043 10984 15083 11024
rect 15235 10984 15275 11024
rect 15543 10984 15583 11024
rect 15724 10984 15764 11024
rect 15916 10984 15956 11024
rect 16771 10984 16811 11024
rect 16876 10984 16916 11024
rect 17452 10984 17492 11024
rect 17731 10984 17771 11024
rect 18302 10984 18342 11024
rect 18604 10975 18644 11015
rect 18979 10984 19019 11024
rect 19948 10984 19988 11024
rect 20716 10984 20756 11024
rect 21196 10984 21236 11024
rect 21580 10984 21620 11024
rect 22339 10975 22379 11015
rect 22444 10984 22484 11024
rect 22828 10984 22868 11024
rect 22947 10984 22987 11024
rect 23068 10984 23108 11024
rect 23203 10975 23243 11015
rect 23639 10984 23679 11024
rect 23884 10984 23924 11024
rect 24161 10984 24201 11024
rect 24460 10975 24500 11015
rect 24638 10984 24678 11024
rect 24748 10984 24788 11024
rect 25099 10984 25139 11024
rect 25324 10984 25364 11024
rect 4012 10900 4052 10940
rect 4963 10900 5003 10940
rect 5731 10900 5771 10940
rect 7372 10900 7412 10940
rect 7875 10900 7915 10940
rect 8643 10900 8683 10940
rect 14083 10900 14123 10940
rect 22732 10900 22772 10940
rect 23779 10900 23819 10940
rect 24945 10942 24985 10982
rect 25612 10984 25652 11024
rect 25900 10984 25940 11024
rect 26275 10984 26315 11024
rect 26380 10984 26420 11024
rect 27436 10984 27476 11024
rect 28588 10984 28628 11024
rect 29260 10984 29300 11024
rect 29443 10984 29483 11024
rect 29644 10984 29684 11024
rect 29829 11003 29869 11043
rect 23980 10900 24020 10940
rect 25219 10900 25259 10940
rect 27346 10900 27386 10940
rect 30028 10942 30068 10982
rect 30220 10984 30260 11024
rect 3916 10816 3956 10856
rect 7276 10816 7316 10856
rect 9772 10816 9812 10856
rect 15043 10816 15083 10856
rect 18124 10816 18164 10856
rect 19024 10816 19064 10856
rect 22051 10816 22091 10856
rect 24844 10816 24884 10856
rect 28876 10816 28916 10856
rect 30412 10816 30452 10856
rect 30796 10816 30836 10856
rect 3427 10732 3467 10772
rect 6883 10732 6923 10772
rect 10252 10732 10292 10772
rect 12316 10732 12356 10772
rect 15532 10732 15572 10772
rect 16972 10732 17012 10772
rect 19555 10732 19595 10772
rect 20323 10732 20363 10772
rect 25612 10732 25652 10772
rect 28195 10732 28235 10772
rect 3112 10564 3480 10604
rect 10886 10564 11254 10604
rect 18660 10564 19028 10604
rect 26434 10564 26802 10604
rect 1660 10396 1700 10436
rect 3340 10396 3380 10436
rect 5251 10396 5291 10436
rect 6412 10396 6452 10436
rect 9052 10396 9092 10436
rect 9484 10396 9524 10436
rect 10147 10396 10187 10436
rect 11404 10396 11444 10436
rect 13315 10396 13355 10436
rect 14908 10396 14948 10436
rect 16636 10396 16676 10436
rect 17251 10396 17291 10436
rect 20668 10396 20708 10436
rect 22051 10396 22091 10436
rect 23980 10396 24020 10436
rect 25036 10396 25076 10436
rect 27811 10396 27851 10436
rect 2275 10312 2315 10352
rect 9916 10286 9956 10326
rect 19363 10312 19403 10352
rect 23155 10312 23195 10352
rect 28492 10312 28532 10352
rect 30412 10312 30452 10352
rect 30796 10312 30836 10352
rect 2659 10228 2699 10268
rect 3619 10228 3659 10268
rect 3820 10228 3860 10268
rect 7171 10228 7211 10268
rect 11506 10228 11546 10268
rect 12019 10228 12059 10268
rect 17548 10228 17588 10268
rect 17763 10228 17803 10268
rect 18028 10228 18068 10268
rect 652 10144 692 10184
rect 844 10144 884 10184
rect 1036 10144 1076 10184
rect 1420 10144 1460 10184
rect 1987 10144 2027 10184
rect 2092 10144 2132 10184
rect 2524 10144 2564 10184
rect 2764 10144 2804 10184
rect 3043 10144 3083 10184
rect 3148 10144 3188 10184
rect 3499 10144 3539 10184
rect 3724 10144 3764 10184
rect 4012 10144 4052 10184
rect 4396 10144 4436 10184
rect 4963 10144 5003 10184
rect 5068 10144 5108 10184
rect 5548 10144 5588 10184
rect 5836 10144 5876 10184
rect 6460 10144 6500 10184
rect 6604 10144 6644 10184
rect 7031 10144 7071 10184
rect 7276 10144 7316 10184
rect 7948 10144 7988 10184
rect 8428 10144 8468 10184
rect 8812 10144 8852 10184
rect 9187 10144 9227 10184
rect 9292 10144 9332 10184
rect 9495 10144 9535 10184
rect 9955 10144 9995 10184
rect 10624 10144 10664 10184
rect 11596 10144 11636 10184
rect 12364 10144 12404 10184
rect 12652 10144 12692 10184
rect 13027 10144 13067 10184
rect 13132 10144 13172 10184
rect 13696 10144 13736 10184
rect 14476 10144 14516 10184
rect 14764 10144 14804 10184
rect 15148 10144 15188 10184
rect 15532 10144 15572 10184
rect 16012 10144 16052 10184
rect 16396 10144 16436 10184
rect 16963 10144 17003 10184
rect 17068 10144 17108 10184
rect 17644 10144 17684 10184
rect 17861 10144 17901 10184
rect 18124 10144 18164 10184
rect 18243 10144 18283 10184
rect 18361 10144 18401 10184
rect 19180 10144 19220 10184
rect 19363 10144 19403 10184
rect 19756 10144 19796 10184
rect 19875 10144 19915 10184
rect 19996 10186 20036 10226
rect 22732 10228 22772 10268
rect 22963 10219 23003 10259
rect 23644 10228 23684 10268
rect 25138 10228 25178 10268
rect 26002 10228 26042 10268
rect 21004 10144 21044 10184
rect 21292 10144 21332 10184
rect 21580 10144 21620 10184
rect 22444 10144 22484 10184
rect 22828 10144 22868 10184
rect 23065 10144 23105 10184
rect 23356 10144 23396 10184
rect 23500 10144 23540 10184
rect 23788 10144 23828 10184
rect 24141 10144 24181 10184
rect 24244 10144 24284 10184
rect 24368 10144 24408 10184
rect 25228 10144 25268 10184
rect 26092 10144 26132 10184
rect 26860 10144 26900 10184
rect 27148 10144 27188 10184
rect 27331 10144 27371 10184
rect 27628 10144 27668 10184
rect 28012 10144 28052 10184
rect 28108 10144 28148 10184
rect 29356 10144 29396 10184
rect 2851 10060 2891 10100
rect 3354 10060 3394 10100
rect 6172 10060 6212 10100
rect 19660 10060 19700 10100
rect 22243 10060 22283 10100
rect 27532 10060 27572 10100
rect 27806 10060 27846 10100
rect 835 9976 875 10016
rect 4492 9976 4532 10016
rect 7363 9976 7403 10016
rect 7843 9976 7883 10016
rect 8140 9976 8180 10016
rect 10780 9976 10820 10016
rect 13852 9976 13892 10016
rect 14275 9976 14315 10016
rect 21676 9976 21716 10016
rect 25795 9976 25835 10016
rect 26659 9976 26699 10016
rect 28012 9976 28052 10016
rect 28684 9976 28724 10016
rect 4352 9808 4720 9848
rect 12126 9808 12494 9848
rect 19900 9808 20268 9848
rect 27674 9808 28042 9848
rect 940 9640 980 9680
rect 1804 9640 1844 9680
rect 4204 9640 4244 9680
rect 4771 9640 4811 9680
rect 6979 9640 7019 9680
rect 7660 9640 7700 9680
rect 8524 9640 8564 9680
rect 9196 9640 9236 9680
rect 9763 9640 9803 9680
rect 10444 9640 10484 9680
rect 10915 9640 10955 9680
rect 12268 9640 12308 9680
rect 13699 9640 13739 9680
rect 13996 9640 14036 9680
rect 14668 9640 14708 9680
rect 15148 9640 15188 9680
rect 15811 9640 15851 9680
rect 17644 9640 17684 9680
rect 17827 9640 17867 9680
rect 18691 9640 18731 9680
rect 20227 9640 20267 9680
rect 20899 9640 20939 9680
rect 21667 9640 21707 9680
rect 23020 9640 23060 9680
rect 23404 9640 23444 9680
rect 24268 9640 24308 9680
rect 24451 9640 24491 9680
rect 25843 9640 25883 9680
rect 27436 9640 27476 9680
rect 2380 9556 2420 9596
rect 6316 9556 6356 9596
rect 13324 9556 13364 9596
rect 15255 9556 15295 9596
rect 15532 9556 15572 9596
rect 25214 9556 25254 9596
rect 25315 9556 25355 9596
rect 26284 9556 26324 9596
rect 26956 9556 26996 9596
rect 940 9472 980 9512
rect 1132 9472 1172 9512
rect 1324 9472 1364 9512
rect 1708 9472 1748 9512
rect 2284 9472 2324 9512
rect 2480 9472 2520 9512
rect 2668 9472 2708 9512
rect 2956 9472 2996 9512
rect 3095 9472 3135 9512
rect 3340 9472 3380 9512
rect 3628 9472 3668 9512
rect 3753 9472 3793 9512
rect 3916 9472 3956 9512
rect 4108 9472 4148 9512
rect 4300 9472 4340 9512
rect 3221 9388 3261 9428
rect 3436 9388 3476 9428
rect 4444 9430 4484 9470
rect 4684 9472 4724 9512
rect 5111 9472 5151 9512
rect 5356 9472 5396 9512
rect 5644 9472 5684 9512
rect 5827 9472 5867 9512
rect 6220 9472 6260 9512
rect 6412 9472 6452 9512
rect 6796 9472 6836 9512
rect 6988 9472 7028 9512
rect 7219 9472 7259 9512
rect 7468 9472 7508 9512
rect 8131 9472 8171 9512
rect 8236 9472 8276 9512
rect 8716 9472 8756 9512
rect 9100 9472 9140 9512
rect 9431 9472 9471 9512
rect 9571 9472 9611 9512
rect 9676 9472 9716 9512
rect 10294 9472 10334 9512
rect 10540 9472 10580 9512
rect 10659 9472 10699 9512
rect 10777 9472 10817 9512
rect 11212 9472 11252 9512
rect 11980 9472 12020 9512
rect 12119 9472 12159 9512
rect 12407 9472 12447 9512
rect 12652 9472 12692 9512
rect 13228 9472 13268 9512
rect 13420 9472 13460 9512
rect 13804 9472 13844 9512
rect 14188 9472 14228 9512
rect 14572 9472 14612 9512
rect 14947 9472 14987 9512
rect 15052 9472 15092 9512
rect 15436 9472 15476 9512
rect 15628 9472 15668 9512
rect 16108 9472 16148 9512
rect 17251 9472 17291 9512
rect 17356 9472 17396 9512
rect 18013 9472 18053 9512
rect 18124 9472 18164 9512
rect 18796 9472 18836 9512
rect 19180 9472 19220 9512
rect 19372 9472 19412 9512
rect 19660 9472 19700 9512
rect 20515 9472 20555 9512
rect 21085 9472 21125 9512
rect 21196 9472 21236 9512
rect 21964 9472 22004 9512
rect 22627 9472 22667 9512
rect 22732 9472 22772 9512
rect 23203 9472 23243 9512
rect 23500 9472 23540 9512
rect 23875 9472 23915 9512
rect 23980 9472 24020 9512
rect 24604 9472 24644 9512
rect 24748 9472 24788 9512
rect 25420 9472 25460 9512
rect 25516 9463 25556 9503
rect 26008 9472 26048 9512
rect 26171 9472 26211 9512
rect 26383 9472 26423 9512
rect 26572 9472 26612 9512
rect 26755 9472 26795 9512
rect 27052 9472 27092 9512
rect 27289 9472 27329 9512
rect 29347 9472 29387 9512
rect 4579 9388 4619 9428
rect 5251 9388 5291 9428
rect 5452 9388 5492 9428
rect 10099 9388 10139 9428
rect 11122 9388 11162 9428
rect 12533 9388 12573 9428
rect 12748 9388 12788 9428
rect 16018 9388 16058 9428
rect 20131 9388 20171 9428
rect 20707 9388 20747 9428
rect 21874 9388 21914 9428
rect 27187 9379 27227 9419
rect 29731 9388 29771 9428
rect 5872 9304 5912 9344
rect 26755 9304 26795 9344
rect 2668 9220 2708 9260
rect 3628 9220 3668 9260
rect 11020 9220 11060 9260
rect 19996 9220 20036 9260
rect 3112 9052 3480 9092
rect 10886 9052 11254 9092
rect 18660 9052 19028 9092
rect 26434 9052 26802 9092
rect 1036 8884 1076 8924
rect 3331 8884 3371 8924
rect 6364 8884 6404 8924
rect 7660 8884 7700 8924
rect 8428 8884 8468 8924
rect 11116 8884 11156 8924
rect 13516 8884 13556 8924
rect 16492 8884 16532 8924
rect 17251 8884 17291 8924
rect 20035 8884 20075 8924
rect 20908 8884 20948 8924
rect 23020 8884 23060 8924
rect 28204 8884 28244 8924
rect 652 8800 692 8840
rect 9244 8791 9284 8831
rect 12220 8791 12260 8831
rect 12451 8800 12491 8840
rect 14188 8800 14228 8840
rect 16867 8800 16907 8840
rect 19747 8800 19787 8840
rect 23404 8800 23444 8840
rect 28396 8800 28436 8840
rect 2947 8716 2987 8756
rect 4786 8716 4826 8756
rect 9964 8716 10004 8756
rect 12652 8716 12692 8756
rect 13228 8716 13268 8756
rect 15532 8716 15572 8756
rect 25138 8716 25178 8756
rect 25948 8716 25988 8756
rect 2563 8632 2603 8672
rect 3329 8632 3369 8672
rect 3628 8632 3668 8672
rect 3820 8632 3860 8672
rect 4204 8632 4244 8672
rect 4876 8632 4916 8672
rect 5452 8632 5492 8672
rect 5683 8632 5723 8672
rect 6028 8632 6068 8672
rect 6604 8632 6644 8672
rect 6988 8632 7028 8672
rect 7267 8632 7307 8672
rect 7376 8639 7416 8679
rect 8131 8632 8171 8672
rect 8236 8632 8276 8672
rect 9283 8632 9323 8672
rect 9643 8632 9683 8672
rect 9763 8632 9803 8672
rect 9868 8632 9908 8672
rect 10336 8632 10376 8672
rect 10819 8632 10859 8672
rect 11788 8632 11828 8672
rect 12259 8632 12299 8672
rect 12835 8632 12875 8672
rect 13564 8632 13604 8672
rect 13708 8632 13748 8672
rect 14188 8632 14228 8672
rect 14380 8632 14420 8672
rect 15043 8632 15083 8672
rect 15148 8632 15188 8672
rect 15628 8632 15668 8672
rect 15747 8632 15787 8672
rect 15865 8632 15905 8672
rect 16195 8632 16235 8672
rect 16492 8632 16532 8672
rect 16684 8632 16724 8672
rect 16867 8632 16907 8672
rect 17068 8632 17108 8672
rect 17251 8632 17291 8672
rect 17878 8632 17918 8672
rect 18508 8632 18548 8672
rect 18650 8632 18690 8672
rect 19459 8632 19499 8672
rect 19564 8632 19604 8672
rect 20236 8632 20276 8672
rect 20332 8632 20372 8672
rect 20611 8632 20651 8672
rect 21475 8632 21515 8672
rect 24172 8632 24212 8672
rect 24556 8632 24596 8672
rect 25228 8632 25268 8672
rect 25804 8632 25844 8672
rect 26764 8632 26804 8672
rect 27148 8632 27188 8672
rect 27244 8632 27284 8672
rect 27532 8632 27572 8672
rect 29068 8632 29108 8672
rect 8439 8548 8479 8588
rect 9484 8548 9524 8588
rect 10492 8548 10532 8588
rect 11130 8548 11170 8588
rect 13132 8548 13172 8588
rect 15244 8548 15284 8588
rect 15351 8548 15391 8588
rect 17683 8548 17723 8588
rect 20030 8548 20070 8588
rect 20919 8548 20959 8588
rect 21091 8548 21131 8588
rect 26942 8548 26982 8588
rect 27043 8548 27083 8588
rect 3532 8464 3572 8504
rect 4300 8464 4340 8504
rect 4579 8464 4619 8504
rect 5308 8464 5348 8504
rect 6124 8464 6164 8504
rect 7171 8455 7211 8495
rect 10915 8464 10955 8504
rect 11683 8464 11723 8504
rect 11980 8464 12020 8504
rect 18796 8464 18836 8504
rect 20707 8464 20747 8504
rect 24652 8464 24692 8504
rect 24931 8464 24971 8504
rect 26092 8464 26132 8504
rect 4352 8296 4720 8336
rect 12126 8296 12494 8336
rect 19900 8296 20268 8336
rect 27674 8296 28042 8336
rect 1468 8128 1508 8168
rect 3043 8128 3083 8168
rect 3340 8128 3380 8168
rect 3811 8128 3851 8168
rect 5827 8128 5867 8168
rect 6307 8128 6347 8168
rect 6604 8128 6644 8168
rect 7660 8128 7700 8168
rect 9091 8128 9131 8168
rect 9859 8128 9899 8168
rect 9964 8128 10004 8168
rect 10732 8128 10772 8168
rect 11404 8128 11444 8168
rect 15820 8128 15860 8168
rect 16195 8128 16235 8168
rect 17539 8128 17579 8168
rect 18211 8128 18251 8168
rect 20131 8128 20171 8168
rect 20332 8128 20372 8168
rect 21100 8128 21140 8168
rect 28108 8128 28148 8168
rect 2764 8044 2804 8084
rect 11980 8044 12020 8084
rect 12184 8044 12224 8084
rect 13027 8044 13067 8084
rect 22147 8044 22187 8084
rect 24067 8035 24107 8075
rect 25132 8044 25172 8084
rect 25795 8044 25835 8084
rect 1315 7951 1355 7991
rect 2668 7960 2708 8000
rect 2851 7960 2891 8000
rect 3148 7960 3188 8000
rect 4108 7960 4148 8000
rect 4845 7960 4885 8000
rect 4993 7960 5033 8000
rect 5285 7960 5325 8000
rect 5932 7960 5972 8000
rect 6412 7960 6452 8000
rect 7267 7960 7307 8000
rect 7372 7960 7412 8000
rect 8035 7960 8075 8000
rect 8140 7960 8180 8000
rect 8620 7960 8660 8000
rect 8812 7960 8852 8000
rect 9292 7960 9332 8000
rect 9580 7960 9620 8000
rect 9763 7960 9803 8000
rect 10074 7960 10114 8000
rect 10252 7960 10292 8000
rect 10636 7960 10676 8000
rect 11500 7960 11540 8000
rect 11717 7960 11757 8000
rect 11875 7960 11915 8000
rect 12695 7960 12735 8000
rect 12931 7960 12971 8000
rect 13276 7960 13316 8000
rect 13577 7960 13617 8000
rect 13731 7960 13771 8000
rect 14476 7960 14516 8000
rect 14611 7960 14651 8000
rect 14956 7960 14996 8000
rect 15148 7960 15188 8000
rect 15379 7960 15419 8000
rect 15724 7960 15764 8000
rect 16396 7960 16436 8000
rect 16684 7960 16724 8000
rect 17207 7960 17247 8000
rect 17452 7960 17492 8000
rect 17740 7960 17780 8000
rect 18028 7960 18068 8000
rect 18364 7960 18404 8000
rect 18508 7960 18548 8000
rect 19267 7960 19307 8000
rect 19372 7960 19412 8000
rect 19799 7960 19839 8000
rect 20044 7960 20084 8000
rect 20428 7960 20468 8000
rect 20659 7960 20699 8000
rect 21772 7960 21812 8000
rect 22828 7960 22868 8000
rect 23308 7960 23348 8000
rect 23779 7960 23819 8000
rect 23884 7951 23924 7991
rect 24171 7960 24211 8000
rect 24340 7949 24380 7989
rect 24542 7960 24582 8000
rect 24652 7960 24692 8000
rect 24844 7960 24884 8000
rect 25031 7960 25071 8000
rect 25216 7960 25256 8000
rect 25420 7960 25460 8000
rect 25612 7960 25652 8000
rect 26179 7960 26219 8000
rect 4018 7876 4058 7916
rect 5164 7876 5204 7916
rect 11619 7876 11659 7916
rect 12835 7876 12875 7916
rect 13420 7876 13460 7916
rect 17347 7876 17387 7916
rect 19939 7876 19979 7916
rect 20563 7867 20603 7907
rect 23218 7876 23258 7916
rect 1996 7792 2036 7832
rect 5068 7792 5108 7832
rect 13516 7792 13556 7832
rect 17740 7792 17780 7832
rect 19555 7792 19595 7832
rect 24556 7792 24596 7832
rect 25219 7792 25259 7832
rect 28300 7792 28340 7832
rect 6124 7708 6164 7748
rect 8323 7708 8363 7748
rect 8620 7708 8660 7748
rect 12172 7708 12212 7748
rect 14659 7708 14699 7748
rect 14956 7708 14996 7748
rect 23116 7708 23156 7748
rect 23779 7708 23819 7748
rect 25420 7708 25460 7748
rect 27724 7708 27764 7748
rect 3112 7540 3480 7580
rect 10886 7540 11254 7580
rect 18660 7540 19028 7580
rect 26434 7540 26802 7580
rect 6028 7372 6068 7412
rect 8035 7372 8075 7412
rect 9388 7372 9428 7412
rect 10252 7372 10292 7412
rect 14476 7372 14516 7412
rect 18979 7372 19019 7412
rect 19660 7372 19700 7412
rect 20812 7372 20852 7412
rect 21187 7372 21227 7412
rect 23356 7372 23396 7412
rect 4204 7288 4244 7328
rect 4652 7279 4692 7319
rect 7180 7288 7220 7328
rect 12892 7288 12932 7328
rect 18499 7288 18539 7328
rect 22380 7279 22420 7319
rect 23500 7288 23540 7328
rect 2131 7204 2171 7244
rect 10354 7204 10394 7244
rect 16204 7204 16244 7244
rect 21676 7204 21716 7244
rect 26476 7204 26516 7244
rect 2326 7120 2366 7160
rect 2572 7120 2612 7160
rect 3244 7120 3284 7160
rect 3436 7120 3476 7160
rect 3820 7120 3860 7160
rect 4675 7120 4715 7160
rect 5068 7120 5108 7160
rect 6109 7120 6149 7160
rect 6223 7120 6263 7160
rect 6787 7120 6827 7160
rect 6892 7153 6932 7193
rect 7747 7120 7787 7160
rect 7852 7120 7892 7160
rect 8323 7120 8363 7160
rect 8631 7120 8671 7160
rect 9187 7120 9227 7160
rect 9298 7120 9338 7160
rect 9772 7120 9812 7160
rect 9964 7120 10004 7160
rect 10444 7120 10484 7160
rect 11116 7120 11156 7160
rect 11500 7120 11540 7160
rect 12268 7120 12308 7160
rect 12652 7120 12692 7160
rect 13219 7120 13259 7160
rect 13324 7120 13364 7160
rect 14179 7120 14219 7160
rect 14851 7120 14891 7160
rect 14956 7120 14996 7160
rect 15628 7120 15668 7160
rect 15724 7120 15764 7160
rect 15863 7120 15903 7160
rect 16003 7120 16043 7160
rect 16108 7120 16148 7160
rect 16396 7120 16436 7160
rect 16588 7120 16628 7160
rect 17443 7120 17483 7160
rect 17548 7120 17588 7160
rect 18211 7120 18251 7160
rect 18316 7120 18356 7160
rect 18940 7120 18980 7160
rect 19084 7120 19124 7160
rect 19708 7120 19748 7160
rect 19852 7120 19892 7160
rect 20611 7120 20651 7160
rect 20716 7120 20756 7160
rect 21182 7120 21222 7160
rect 21484 7120 21524 7160
rect 21772 7120 21812 7160
rect 21891 7120 21931 7160
rect 22009 7120 22049 7160
rect 22339 7120 22379 7160
rect 22732 7120 22772 7160
rect 25075 7162 25115 7202
rect 23020 7120 23060 7160
rect 24064 7120 24104 7160
rect 25228 7120 25268 7160
rect 25420 7120 25460 7160
rect 26135 7120 26175 7160
rect 26275 7120 26315 7160
rect 26380 7120 26420 7160
rect 27235 7120 27275 7160
rect 27543 7120 27583 7160
rect 2942 7036 2982 7076
rect 4876 7036 4916 7076
rect 8524 7036 8564 7076
rect 14284 7036 14324 7076
rect 14490 7036 14530 7076
rect 15425 7036 15465 7076
rect 21388 7036 21428 7076
rect 24220 7036 24260 7076
rect 25324 7036 25364 7076
rect 27436 7036 27476 7076
rect 2467 6952 2507 6992
rect 2764 6952 2804 6992
rect 3043 6952 3083 6992
rect 3148 6952 3188 6992
rect 3916 6952 3956 6992
rect 5740 6952 5780 6992
rect 6691 6943 6731 6983
rect 8419 6952 8459 6992
rect 9955 6952 9995 6992
rect 10147 6952 10187 6992
rect 11596 6952 11636 6992
rect 13612 6952 13652 6992
rect 15244 6952 15284 6992
rect 15523 6952 15563 6992
rect 15628 6952 15668 6992
rect 16396 6952 16436 6992
rect 17836 6952 17876 6992
rect 21004 6952 21044 6992
rect 22156 6952 22196 6992
rect 24883 6952 24923 6992
rect 27331 6952 27371 6992
rect 4352 6784 4720 6824
rect 12126 6784 12494 6824
rect 19900 6784 20268 6824
rect 27674 6784 28042 6824
rect 5068 6616 5108 6656
rect 6220 6616 6260 6656
rect 7660 6616 7700 6656
rect 8812 6616 8852 6656
rect 9676 6616 9716 6656
rect 9859 6616 9899 6656
rect 11788 6616 11828 6656
rect 12259 6616 12299 6656
rect 13324 6616 13364 6656
rect 13699 6616 13739 6656
rect 16108 6616 16148 6656
rect 16780 6616 16820 6656
rect 19171 6616 19211 6656
rect 19939 6616 19979 6656
rect 20995 6616 21035 6656
rect 21763 6616 21803 6656
rect 22243 6616 22283 6656
rect 23875 6616 23915 6656
rect 23980 6616 24020 6656
rect 24364 6616 24404 6656
rect 2755 6532 2795 6572
rect 8131 6532 8171 6572
rect 13914 6532 13954 6572
rect 15244 6532 15284 6572
rect 2380 6448 2420 6488
rect 2597 6448 2637 6488
rect 3139 6448 3179 6488
rect 5590 6448 5630 6488
rect 5932 6448 5972 6488
rect 6071 6448 6111 6488
rect 6412 6448 6452 6488
rect 6527 6448 6567 6488
rect 6700 6448 6740 6488
rect 7267 6448 7307 6488
rect 7378 6450 7418 6490
rect 7819 6448 7859 6488
rect 8044 6448 8084 6488
rect 8332 6448 8372 6488
rect 8716 6448 8756 6488
rect 9388 6448 9428 6488
rect 9523 6448 9563 6488
rect 10012 6448 10052 6488
rect 10156 6448 10196 6488
rect 10583 6448 10623 6488
rect 10828 6448 10868 6488
rect 11395 6448 11435 6488
rect 11500 6448 11540 6488
rect 11927 6448 11967 6488
rect 12172 6448 12212 6488
rect 12844 6448 12884 6488
rect 13132 6448 13172 6488
rect 13603 6448 13643 6488
rect 13708 6448 13748 6488
rect 14039 6448 14079 6488
rect 14284 6448 14324 6488
rect 15038 6448 15078 6488
rect 15340 6439 15380 6479
rect 15715 6448 15755 6488
rect 15820 6448 15860 6488
rect 16300 6448 16340 6488
rect 16684 6448 16724 6488
rect 17164 6448 17204 6488
rect 17401 6448 17441 6488
rect 17932 6448 17972 6488
rect 18316 6448 18356 6488
rect 19468 6448 19508 6488
rect 20125 6448 20165 6488
rect 20236 6448 20276 6488
rect 20663 6448 20703 6488
rect 20908 6448 20948 6488
rect 21196 6448 21236 6488
rect 21379 6448 21419 6488
rect 21484 6448 21524 6488
rect 21924 6448 21964 6488
rect 22060 6448 22100 6488
rect 22348 6448 22388 6488
rect 23596 6448 23636 6488
rect 23777 6448 23817 6488
rect 24076 6439 24116 6479
rect 24263 6448 24303 6488
rect 24451 6448 24491 6488
rect 2284 6364 2324 6404
rect 2515 6355 2555 6395
rect 5395 6364 5435 6404
rect 7939 6364 7979 6404
rect 10723 6364 10763 6404
rect 10924 6364 10964 6404
rect 12067 6364 12107 6404
rect 14179 6364 14219 6404
rect 14380 6364 14420 6404
rect 17068 6364 17108 6404
rect 17283 6364 17323 6404
rect 19378 6364 19418 6404
rect 20803 6364 20843 6404
rect 16003 6280 16043 6320
rect 21292 6280 21332 6320
rect 22540 6280 22580 6320
rect 4684 6196 4724 6236
rect 6412 6196 6452 6236
rect 13900 6196 13940 6236
rect 15043 6196 15083 6236
rect 18556 6196 18596 6236
rect 22924 6196 22964 6236
rect 24451 6196 24491 6236
rect 3112 6028 3480 6068
rect 10886 6028 11254 6068
rect 18660 6028 19028 6068
rect 26434 6028 26802 6068
rect 5740 5860 5780 5900
rect 9676 5860 9716 5900
rect 14380 5860 14420 5900
rect 15043 5860 15083 5900
rect 20611 5860 20651 5900
rect 20908 5860 20948 5900
rect 23212 5860 23252 5900
rect 23596 5860 23636 5900
rect 4876 5776 4916 5816
rect 9004 5776 9044 5816
rect 13420 5776 13460 5816
rect 23788 5776 23828 5816
rect 6700 5692 6740 5732
rect 10659 5692 10699 5732
rect 21292 5692 21332 5732
rect 2462 5608 2502 5648
rect 2764 5608 2804 5648
rect 2947 5608 2987 5648
rect 3628 5608 3668 5648
rect 3907 5608 3947 5648
rect 4563 5608 4603 5648
rect 4683 5608 4723 5648
rect 5068 5608 5108 5648
rect 6115 5608 6155 5648
rect 6220 5608 6260 5648
rect 6604 5608 6644 5648
rect 6796 5608 6836 5648
rect 7123 5608 7163 5648
rect 7318 5608 7358 5648
rect 7459 5608 7499 5648
rect 8140 5608 8180 5648
rect 8620 5608 8660 5648
rect 9379 5608 9419 5648
rect 10060 5608 10100 5648
rect 10540 5608 10580 5648
rect 10777 5608 10817 5648
rect 11107 5608 11147 5648
rect 11212 5608 11252 5648
rect 11644 5608 11684 5648
rect 11834 5608 11874 5648
rect 12172 5608 12212 5648
rect 12556 5608 12596 5648
rect 13027 5608 13067 5648
rect 13144 5615 13184 5655
rect 13804 5608 13844 5648
rect 14083 5608 14123 5648
rect 14380 5608 14420 5648
rect 14755 5608 14795 5648
rect 14860 5608 14900 5648
rect 15484 5608 15524 5648
rect 15628 5608 15668 5648
rect 16204 5608 16244 5648
rect 16323 5608 16363 5648
rect 16441 5608 16481 5648
rect 16684 5608 16724 5648
rect 17068 5608 17108 5648
rect 17635 5608 17675 5648
rect 17740 5608 17780 5648
rect 18412 5608 18452 5648
rect 18796 5608 18836 5648
rect 19180 5608 19220 5648
rect 19564 5608 19604 5648
rect 20428 5608 20468 5648
rect 20611 5608 20651 5648
rect 20812 5608 20852 5648
rect 21004 5608 21044 5648
rect 21667 5608 21707 5648
rect 2563 5524 2603 5564
rect 4108 5524 4148 5564
rect 4218 5524 4258 5564
rect 6403 5524 6443 5564
rect 9484 5524 9524 5564
rect 9690 5524 9730 5564
rect 9859 5524 9899 5564
rect 10444 5524 10484 5564
rect 2668 5440 2708 5480
rect 4003 5440 4043 5480
rect 4588 5440 4628 5480
rect 6124 5440 6164 5480
rect 8515 5440 8555 5480
rect 8812 5440 8852 5480
rect 10147 5440 10187 5480
rect 11500 5440 11540 5480
rect 11980 5440 12020 5480
rect 12652 5440 12692 5480
rect 12931 5431 12971 5471
rect 13612 5440 13652 5480
rect 13891 5440 13931 5480
rect 15331 5440 15371 5480
rect 16108 5440 16148 5480
rect 17164 5440 17204 5480
rect 18028 5440 18068 5480
rect 18307 5440 18347 5480
rect 18988 5440 19028 5480
rect 19267 5440 19307 5480
rect 20236 5440 20276 5480
rect 4352 5272 4720 5312
rect 12126 5272 12494 5312
rect 19900 5272 20268 5312
rect 27674 5272 28042 5312
rect 7372 5104 7412 5144
rect 10348 5104 10388 5144
rect 11395 5104 11435 5144
rect 12259 5104 12299 5144
rect 12556 5104 12596 5144
rect 15532 5104 15572 5144
rect 18412 5104 18452 5144
rect 18691 5104 18731 5144
rect 21436 5104 21476 5144
rect 21868 5104 21908 5144
rect 22252 5104 22292 5144
rect 5059 5020 5099 5060
rect 12835 5020 12875 5060
rect 13219 5020 13259 5060
rect 18906 5020 18946 5060
rect 21978 5020 22018 5060
rect 5443 4936 5483 4976
rect 7555 4927 7595 4967
rect 8419 4936 8459 4976
rect 11212 4936 11252 4976
rect 11692 4936 11732 4976
rect 12364 4936 12404 4976
rect 12738 4936 12778 4976
rect 12931 4936 12971 4976
rect 13036 4936 13076 4976
rect 13603 4936 13643 4976
rect 16483 4936 16523 4976
rect 18595 4936 18635 4976
rect 20131 4927 20171 4967
rect 20908 4936 20948 4976
rect 21104 4936 21144 4976
rect 21292 4936 21332 4976
rect 21667 4936 21707 4976
rect 21772 4936 21812 4976
rect 22156 4936 22196 4976
rect 22348 4936 22388 4976
rect 7708 4852 7748 4892
rect 8044 4852 8084 4892
rect 11602 4852 11642 4892
rect 15148 4852 15188 4892
rect 16108 4852 16148 4892
rect 18028 4852 18068 4892
rect 20284 4852 20324 4892
rect 7372 4768 7412 4808
rect 10540 4768 10580 4808
rect 6988 4684 7028 4724
rect 9964 4684 10004 4724
rect 10348 4684 10388 4724
rect 18892 4684 18932 4724
rect 21004 4684 21044 4724
rect 3112 4516 3480 4556
rect 10886 4516 11254 4556
rect 18660 4516 19028 4556
rect 26434 4516 26802 4556
rect 7852 4348 7892 4388
rect 13228 4348 13268 4388
rect 16108 4348 16148 4388
rect 6220 4264 6260 4304
rect 8476 4264 8516 4304
rect 11788 4264 11828 4304
rect 13708 4264 13748 4304
rect 14476 4264 14516 4304
rect 17164 4264 17204 4304
rect 8259 4180 8299 4220
rect 9811 4180 9851 4220
rect 10588 4180 10628 4220
rect 15187 4180 15227 4220
rect 7555 4096 7595 4136
rect 8140 4096 8180 4136
rect 8377 4096 8417 4136
rect 8620 4096 8660 4136
rect 10006 4096 10046 4136
rect 10387 4096 10427 4136
rect 11692 4096 11732 4136
rect 11884 4096 11924 4136
rect 13228 4096 13268 4136
rect 13420 4096 13460 4136
rect 13804 4096 13844 4136
rect 14092 4096 14132 4136
rect 15382 4096 15422 4136
rect 15811 4096 15851 4136
rect 16122 4096 16162 4136
rect 7866 4012 7906 4052
rect 8044 4012 8084 4052
rect 15916 4012 15956 4052
rect 7651 3928 7691 3968
rect 13708 3928 13748 3968
rect 13987 3928 14027 3968
rect 14284 3928 14324 3968
rect 4352 3760 4720 3800
rect 12126 3760 12494 3800
rect 19900 3760 20268 3800
rect 27674 3760 28042 3800
rect 3112 3004 3480 3044
rect 10886 3004 11254 3044
rect 18660 3004 19028 3044
rect 26434 3004 26802 3044
rect 4352 2248 4720 2288
rect 12126 2248 12494 2288
rect 19900 2248 20268 2288
rect 27674 2248 28042 2288
rect 3112 1492 3480 1532
rect 10886 1492 11254 1532
rect 18660 1492 19028 1532
rect 26434 1492 26802 1532
rect 4352 736 4720 776
rect 12126 736 12494 776
rect 19900 736 20268 776
rect 27674 736 28042 776
<< metal2 >>
rect 16387 28624 16396 28664
rect 16436 28624 30068 28664
rect 30028 28580 30068 28624
rect 9091 28540 9100 28580
rect 9140 28540 29260 28580
rect 29300 28540 29309 28580
rect 30019 28540 30028 28580
rect 30068 28540 30077 28580
rect 2947 28456 2956 28496
rect 2996 28456 9196 28496
rect 9236 28456 9245 28496
rect 13891 28456 13900 28496
rect 13940 28456 25516 28496
rect 25556 28456 25565 28496
rect 1795 28372 1804 28412
rect 1844 28372 7084 28412
rect 7124 28372 7133 28412
rect 3436 28204 6796 28244
rect 6836 28204 6845 28244
rect 3436 28160 3476 28204
rect 2755 28120 2764 28160
rect 2804 28120 3476 28160
rect 3523 28120 3532 28160
rect 3572 28120 8236 28160
rect 8276 28120 8285 28160
rect 27715 28120 27724 28160
rect 27764 28120 30988 28160
rect 31028 28120 31037 28160
rect 1891 28036 1900 28076
rect 1940 28036 5932 28076
rect 5972 28036 5981 28076
rect 2179 27952 2188 27992
rect 2228 27952 2956 27992
rect 2996 27952 3005 27992
rect 4343 27952 4352 27992
rect 4720 27952 4729 27992
rect 12117 27952 12126 27992
rect 12494 27952 12503 27992
rect 14083 27952 14092 27992
rect 14132 27952 14612 27992
rect 19891 27952 19900 27992
rect 20268 27952 20277 27992
rect 25219 27952 25228 27992
rect 25268 27952 27092 27992
rect 27665 27952 27674 27992
rect 28042 27952 28051 27992
rect 14572 27908 14612 27952
rect 27052 27908 27092 27952
rect 844 27868 5452 27908
rect 5492 27868 5501 27908
rect 10627 27868 10636 27908
rect 10676 27868 14516 27908
rect 14572 27868 26956 27908
rect 26996 27868 27005 27908
rect 27052 27868 30356 27908
rect 844 27824 884 27868
rect 835 27784 844 27824
rect 884 27784 893 27824
rect 1603 27784 1612 27824
rect 1652 27784 6988 27824
rect 7028 27784 7037 27824
rect 14476 27740 14516 27868
rect 30316 27824 30356 27868
rect 17731 27784 17740 27824
rect 17780 27784 17980 27824
rect 18020 27784 18029 27824
rect 25411 27784 25420 27824
rect 25460 27784 30164 27824
rect 30298 27784 30307 27824
rect 30347 27784 30356 27824
rect 30124 27740 30164 27784
rect 1769 27700 1900 27740
rect 1940 27700 1949 27740
rect 2467 27700 2476 27740
rect 2516 27700 3715 27740
rect 3755 27700 3764 27740
rect 4570 27700 4579 27740
rect 4619 27700 6700 27740
rect 6740 27700 6749 27740
rect 9283 27700 9292 27740
rect 9332 27700 10060 27740
rect 10100 27700 10109 27740
rect 12154 27700 12163 27740
rect 12203 27700 12940 27740
rect 12980 27700 12989 27740
rect 14458 27700 14467 27740
rect 14507 27700 14516 27740
rect 17059 27700 17068 27740
rect 17108 27700 19604 27740
rect 14188 27656 14420 27661
rect 19564 27656 19604 27700
rect 26380 27700 29260 27740
rect 29300 27700 29309 27740
rect 30124 27700 30836 27740
rect 26380 27656 26420 27700
rect 30796 27656 30836 27700
rect 1673 27616 1804 27656
rect 1844 27616 1853 27656
rect 1978 27616 1987 27656
rect 2027 27616 2036 27656
rect 2186 27616 2195 27656
rect 2235 27616 2275 27656
rect 2362 27616 2371 27656
rect 2411 27616 2668 27656
rect 2708 27616 2717 27656
rect 2909 27616 2951 27656
rect 2991 27616 3000 27656
rect 3130 27616 3139 27656
rect 3188 27616 3319 27656
rect 4265 27616 4396 27656
rect 4436 27616 4445 27656
rect 4954 27616 4963 27656
rect 5003 27616 5740 27656
rect 5780 27616 5789 27656
rect 7363 27616 7372 27656
rect 7412 27616 7459 27656
rect 7499 27616 7543 27656
rect 9946 27616 9955 27656
rect 9995 27616 11308 27656
rect 11348 27616 12172 27656
rect 12212 27616 12221 27656
rect 14074 27616 14083 27656
rect 14123 27621 14420 27656
rect 14123 27616 14228 27621
rect 1996 27488 2036 27616
rect 2188 27572 2228 27616
rect 2956 27572 2996 27616
rect 2179 27532 2188 27572
rect 2228 27532 2237 27572
rect 2947 27532 2956 27572
rect 2996 27532 3005 27572
rect 3244 27532 4800 27572
rect 6499 27532 6508 27572
rect 6548 27532 7084 27572
rect 7124 27532 7133 27572
rect 7459 27532 7468 27572
rect 7508 27532 7517 27572
rect 9449 27532 9580 27572
rect 9620 27532 9629 27572
rect 10531 27532 10540 27572
rect 10580 27532 10589 27572
rect 14179 27532 14188 27572
rect 14228 27532 14237 27572
rect 3244 27488 3284 27532
rect 14380 27488 14420 27621
rect 15331 27616 15340 27656
rect 15380 27616 15427 27656
rect 15467 27616 15511 27656
rect 15619 27616 15628 27656
rect 15668 27616 17534 27656
rect 17574 27616 17583 27656
rect 17836 27647 17876 27656
rect 18115 27616 18124 27656
rect 18164 27616 18173 27656
rect 18307 27616 18316 27656
rect 18356 27616 19180 27656
rect 19220 27616 19229 27656
rect 19546 27616 19555 27656
rect 19595 27616 19604 27656
rect 22330 27616 22339 27656
rect 22388 27616 22519 27656
rect 26362 27616 26371 27656
rect 26411 27616 26420 27656
rect 26746 27616 26755 27656
rect 26795 27616 26860 27656
rect 26900 27616 26935 27656
rect 27322 27616 27331 27656
rect 27371 27616 29356 27656
rect 29396 27616 29405 27656
rect 29993 27616 30124 27656
rect 30164 27616 30173 27656
rect 30329 27616 30412 27656
rect 30452 27616 30460 27656
rect 30500 27616 30509 27656
rect 30595 27616 30604 27656
rect 30644 27616 30691 27656
rect 30778 27647 30836 27656
rect 17836 27572 17876 27607
rect 14921 27532 15052 27572
rect 15092 27532 15101 27572
rect 15715 27532 15724 27572
rect 15764 27532 15773 27572
rect 16780 27532 17876 27572
rect 18124 27572 18164 27616
rect 30604 27572 30644 27616
rect 30778 27607 30787 27647
rect 30827 27607 30836 27647
rect 30778 27606 30836 27607
rect 18124 27532 18932 27572
rect 18979 27532 18988 27572
rect 19028 27532 19180 27572
rect 19220 27532 19229 27572
rect 20832 27532 21100 27572
rect 21140 27532 21149 27572
rect 21833 27532 21964 27572
rect 22004 27532 22013 27572
rect 22531 27532 22540 27572
rect 22580 27532 22589 27572
rect 24931 27532 24940 27572
rect 24980 27532 25152 27572
rect 26825 27532 26956 27572
rect 26996 27532 27005 27572
rect 27331 27532 27340 27572
rect 27380 27532 27389 27572
rect 30595 27532 30604 27572
rect 30644 27532 30653 27572
rect 30883 27532 30892 27572
rect 30932 27532 30940 27572
rect 30980 27532 31063 27572
rect 1219 27448 1228 27488
rect 1268 27448 1277 27488
rect 1996 27448 2092 27488
rect 2132 27448 2141 27488
rect 2249 27448 2371 27488
rect 2420 27448 2429 27488
rect 2633 27448 2764 27488
rect 2804 27448 2813 27488
rect 2860 27448 3284 27488
rect 3401 27448 3532 27488
rect 3572 27448 3581 27488
rect 14380 27448 14612 27488
rect 14729 27448 14860 27488
rect 14900 27448 14909 27488
rect 1228 27404 1268 27448
rect 2860 27404 2900 27448
rect 14572 27404 14612 27448
rect 16780 27404 16820 27532
rect 18892 27488 18932 27532
rect 17347 27448 17356 27488
rect 17396 27448 18836 27488
rect 18892 27448 19084 27488
rect 19124 27448 19133 27488
rect 18796 27404 18836 27448
rect 1228 27364 2900 27404
rect 3130 27364 3139 27404
rect 3179 27364 6836 27404
rect 6883 27364 6892 27404
rect 6932 27364 8620 27404
rect 8660 27364 8669 27404
rect 9379 27364 9388 27404
rect 9428 27364 10732 27404
rect 10772 27364 10781 27404
rect 10828 27364 11884 27404
rect 11924 27364 11933 27404
rect 14572 27364 15820 27404
rect 15860 27364 15869 27404
rect 16099 27364 16108 27404
rect 16148 27364 16820 27404
rect 17530 27364 17539 27404
rect 17588 27364 17719 27404
rect 18796 27364 20428 27404
rect 20468 27364 20477 27404
rect 21187 27364 21196 27404
rect 21236 27364 21484 27404
rect 21524 27364 21533 27404
rect 23395 27364 23404 27404
rect 23444 27364 24268 27404
rect 24308 27364 24317 27404
rect 24451 27364 24460 27404
rect 24500 27364 25900 27404
rect 25940 27364 25949 27404
rect 27907 27364 27916 27404
rect 27956 27364 29164 27404
rect 29204 27364 29260 27404
rect 29300 27364 29309 27404
rect 29443 27364 29452 27404
rect 29492 27364 29644 27404
rect 29684 27364 29693 27404
rect 6796 27320 6836 27364
rect 10828 27320 10868 27364
rect 2860 27280 3916 27320
rect 3956 27280 3965 27320
rect 6796 27280 8524 27320
rect 8564 27280 8573 27320
rect 10339 27280 10348 27320
rect 10388 27280 10868 27320
rect 12067 27280 12076 27320
rect 12116 27280 14764 27320
rect 14804 27280 14813 27320
rect 14947 27280 14956 27320
rect 14996 27280 23308 27320
rect 23348 27280 23357 27320
rect 2860 27152 2900 27280
rect 3103 27196 3112 27236
rect 3480 27196 3489 27236
rect 10877 27196 10886 27236
rect 11254 27196 11263 27236
rect 18651 27196 18660 27236
rect 19028 27196 19037 27236
rect 26425 27196 26434 27236
rect 26802 27196 26811 27236
rect 1132 27112 2900 27152
rect 6316 27112 10444 27152
rect 10484 27112 10493 27152
rect 13507 27112 13516 27152
rect 13556 27112 21004 27152
rect 21044 27112 21053 27152
rect 1132 26984 1172 27112
rect 6316 27068 6356 27112
rect 1961 27028 2092 27068
rect 2132 27028 2141 27068
rect 2650 27028 2659 27068
rect 2699 27028 6356 27068
rect 6569 27028 6691 27068
rect 6740 27028 6749 27068
rect 7930 27028 7939 27068
rect 7979 27028 9580 27068
rect 9620 27028 9629 27068
rect 9850 27028 9859 27068
rect 9899 27028 11212 27068
rect 11252 27028 11261 27068
rect 11945 27028 12076 27068
rect 12116 27028 12125 27068
rect 13411 27028 13420 27068
rect 13460 27028 14956 27068
rect 14996 27028 15005 27068
rect 19049 27028 19180 27068
rect 19220 27028 19229 27068
rect 19363 27028 19372 27068
rect 19412 27028 21812 27068
rect 21955 27028 21964 27068
rect 22004 27028 22924 27068
rect 22964 27028 22973 27068
rect 26371 27028 26380 27068
rect 26420 27028 26860 27068
rect 26900 27028 26909 27068
rect 28291 27028 28300 27068
rect 28340 27028 30124 27068
rect 30164 27028 30173 27068
rect 1123 26944 1132 26984
rect 1172 26944 1181 26984
rect 2092 26944 2860 26984
rect 2900 26944 2909 26984
rect 6377 26944 6508 26984
rect 6548 26944 6557 26984
rect 8515 26944 8524 26984
rect 8564 26944 8852 26984
rect 2092 26816 2132 26944
rect 3113 26860 3235 26900
rect 3284 26860 3293 26900
rect 3523 26860 3532 26900
rect 3572 26860 3581 26900
rect 7747 26860 7756 26900
rect 7796 26860 7948 26900
rect 7988 26860 7997 26900
rect 6976 26851 7016 26858
rect 6946 26849 7016 26851
rect 6946 26837 6976 26849
rect 5644 26816 5684 26825
rect 6782 26816 6892 26837
rect 2083 26776 2092 26816
rect 2132 26776 2141 26816
rect 2275 26776 2284 26816
rect 2324 26776 2476 26816
rect 2516 26776 2525 26816
rect 2650 26776 2659 26816
rect 2708 26776 2860 26816
rect 2900 26776 2909 26816
rect 3148 26776 4588 26816
rect 4628 26776 4637 26816
rect 4762 26776 4771 26816
rect 4811 26776 4820 26816
rect 5059 26776 5068 26816
rect 5108 26776 5155 26816
rect 5195 26776 5239 26816
rect 5417 26776 5548 26816
rect 5588 26776 5597 26816
rect 5684 26776 5731 26816
rect 5875 26776 5884 26816
rect 5924 26776 5932 26816
rect 5972 26776 6055 26816
rect 6499 26776 6508 26816
rect 6548 26797 6892 26816
rect 6932 26809 6976 26837
rect 8236 26816 8276 26825
rect 8716 26816 8756 26825
rect 6932 26800 7016 26809
rect 6932 26797 6986 26800
rect 6548 26776 6822 26797
rect 7066 26776 7075 26816
rect 7115 26776 7124 26816
rect 7171 26776 7180 26816
rect 7220 26776 8140 26816
rect 8180 26776 8189 26816
rect 8489 26776 8620 26816
rect 8660 26776 8669 26816
rect 8812 26816 8852 26944
rect 9292 26944 11057 26984
rect 11107 26944 11116 26984
rect 11156 26944 11692 26984
rect 11732 26944 11741 26984
rect 12739 26944 12748 26984
rect 12788 26944 13268 26984
rect 13315 26944 13324 26984
rect 13364 26944 13420 26984
rect 13460 26944 13495 26984
rect 15593 26944 15628 26984
rect 15668 26944 15724 26984
rect 15764 26944 15773 26984
rect 8812 26776 8908 26816
rect 8948 26776 8957 26816
rect 2476 26732 2516 26776
rect 3148 26732 3188 26776
rect 2476 26692 3188 26732
rect 4780 26648 4820 26776
rect 5644 26732 5684 26776
rect 7084 26732 7124 26776
rect 8236 26732 8276 26776
rect 8716 26732 8756 26776
rect 9292 26732 9332 26944
rect 11017 26900 11057 26944
rect 13228 26900 13268 26944
rect 10156 26860 10924 26900
rect 10964 26860 10973 26900
rect 11017 26860 12172 26900
rect 12212 26860 12221 26900
rect 13228 26860 13516 26900
rect 13556 26860 13565 26900
rect 18307 26860 18316 26900
rect 18356 26860 18365 26900
rect 18499 26860 18508 26900
rect 18548 26860 19372 26900
rect 19412 26860 19421 26900
rect 19468 26860 20611 26900
rect 20651 26860 20660 26900
rect 10156 26816 10196 26860
rect 11788 26816 11828 26860
rect 19468 26816 19508 26860
rect 21772 26816 21812 27028
rect 23395 26860 23404 26900
rect 23444 26860 25364 26900
rect 30115 26860 30124 26900
rect 30164 26860 30173 26900
rect 25324 26816 25364 26860
rect 5211 26692 5260 26732
rect 5300 26692 5342 26732
rect 5382 26692 5391 26732
rect 5635 26692 5644 26732
rect 5684 26692 5693 26732
rect 7037 26692 7084 26732
rect 7124 26692 7133 26732
rect 7180 26692 7934 26732
rect 7974 26692 7983 26732
rect 8131 26692 8140 26732
rect 8180 26692 8276 26732
rect 8323 26692 8332 26732
rect 8372 26692 8414 26732
rect 8454 26692 8660 26732
rect 8716 26692 9332 26732
rect 9388 26776 10156 26816
rect 10313 26776 10444 26816
rect 10484 26776 10924 26816
rect 10964 26776 11404 26816
rect 11444 26776 11453 26816
rect 11779 26776 11788 26816
rect 11828 26776 11837 26816
rect 11884 26776 11910 26816
rect 11950 26776 11959 26816
rect 12028 26776 12037 26816
rect 12077 26776 12116 26816
rect 12250 26776 12259 26816
rect 12299 26776 12556 26816
rect 12596 26776 12605 26816
rect 12931 26776 12940 26816
rect 12980 26776 12989 26816
rect 13188 26776 13197 26816
rect 13237 26776 13268 26816
rect 13315 26776 13324 26816
rect 13385 26776 13495 26816
rect 13642 26776 13651 26816
rect 13691 26776 13700 26816
rect 13795 26776 13804 26816
rect 13844 26776 13975 26816
rect 14746 26776 14755 26816
rect 14795 26776 14804 26816
rect 15811 26776 15820 26816
rect 15860 26776 16820 26816
rect 17050 26776 17059 26816
rect 17108 26776 17239 26816
rect 19459 26776 19468 26816
rect 19508 26776 19517 26816
rect 19564 26807 19604 26816
rect 1385 26608 1516 26648
rect 1556 26608 1565 26648
rect 1769 26608 1900 26648
rect 1940 26608 1949 26648
rect 2851 26608 2860 26648
rect 2900 26608 3340 26648
rect 3380 26608 3389 26648
rect 4675 26608 4684 26648
rect 4724 26608 4820 26648
rect 5321 26608 5443 26648
rect 5492 26608 5501 26648
rect 7180 26606 7220 26692
rect 8620 26648 8660 26692
rect 9388 26648 9428 26776
rect 10156 26767 10196 26776
rect 11404 26732 11444 26776
rect 11884 26732 11924 26776
rect 12076 26732 12116 26776
rect 12940 26732 12980 26776
rect 13228 26732 13268 26776
rect 13660 26732 13700 26776
rect 14764 26732 14804 26776
rect 16780 26732 16820 26776
rect 19651 26776 19660 26816
rect 19700 26776 19852 26816
rect 19892 26776 19901 26816
rect 20201 26776 20332 26816
rect 20372 26776 20381 26816
rect 21161 26776 21196 26816
rect 21236 26776 21292 26816
rect 21332 26776 21341 26816
rect 21396 26776 21484 26816
rect 21524 26776 21527 26816
rect 21567 26776 21576 26816
rect 21658 26776 21667 26816
rect 21707 26776 21716 26816
rect 21763 26776 21772 26816
rect 21812 26776 21821 26816
rect 21868 26776 22732 26816
rect 22772 26776 22781 26816
rect 23107 26776 23116 26816
rect 23156 26776 23596 26816
rect 23636 26776 23645 26816
rect 24067 26776 24076 26816
rect 24116 26776 24460 26816
rect 24500 26776 24509 26816
rect 25315 26776 25324 26816
rect 25364 26776 25373 26816
rect 25891 26776 25900 26816
rect 25940 26776 26188 26816
rect 26228 26776 26237 26816
rect 26921 26776 27052 26816
rect 27092 26776 27101 26816
rect 27148 26776 27916 26816
rect 27956 26776 27965 26816
rect 29347 26776 29356 26816
rect 29396 26776 30211 26816
rect 30251 26776 30260 26816
rect 30883 26776 30892 26816
rect 30932 26776 30941 26816
rect 19564 26732 19604 26767
rect 7433 26608 7516 26648
rect 7556 26608 7564 26648
rect 7604 26608 7613 26648
rect 8131 26608 8140 26648
rect 8180 26608 8189 26648
rect 8506 26608 8515 26648
rect 8555 26608 8564 26648
rect 8620 26608 9428 26648
rect 9484 26692 9854 26732
rect 9894 26692 9903 26732
rect 10723 26692 10732 26732
rect 10772 26692 10781 26732
rect 11404 26692 11924 26732
rect 11980 26692 12116 26732
rect 12521 26692 12570 26732
rect 12610 26692 12652 26732
rect 12692 26692 12701 26732
rect 12940 26692 13124 26732
rect 13228 26692 13516 26732
rect 13556 26692 13565 26732
rect 13660 26692 13996 26732
rect 14036 26692 14804 26732
rect 14921 26692 15043 26732
rect 15092 26692 15101 26732
rect 16483 26692 16492 26732
rect 16532 26692 16675 26732
rect 16715 26692 16724 26732
rect 16780 26692 17548 26732
rect 17588 26692 17597 26732
rect 17731 26692 17740 26732
rect 17780 26692 19604 26732
rect 19660 26692 20564 26732
rect 7180 26566 7219 26606
rect 7259 26566 7268 26606
rect 7180 26564 7220 26566
rect 4204 26524 7220 26564
rect 8140 26564 8180 26608
rect 8524 26564 8564 26608
rect 9484 26564 9524 26692
rect 10732 26648 10772 26692
rect 9571 26608 9580 26648
rect 9620 26608 9751 26648
rect 10051 26608 10060 26648
rect 10100 26608 10156 26648
rect 10196 26608 10231 26648
rect 10330 26608 10339 26648
rect 10388 26608 10519 26648
rect 10627 26608 10636 26648
rect 10676 26608 10685 26648
rect 10732 26608 10819 26648
rect 10859 26608 10868 26648
rect 11107 26608 11116 26648
rect 11156 26608 11299 26648
rect 11339 26608 11348 26648
rect 11465 26608 11596 26648
rect 11636 26608 11645 26648
rect 8140 26524 8428 26564
rect 8468 26524 8477 26564
rect 8524 26524 9524 26564
rect 10636 26564 10676 26608
rect 10636 26524 11788 26564
rect 11828 26524 11837 26564
rect 4204 26480 4244 26524
rect 2083 26440 2092 26480
rect 2132 26440 4244 26480
rect 4343 26440 4352 26480
rect 4720 26440 4729 26480
rect 4876 26440 7756 26480
rect 7796 26440 7805 26480
rect 7939 26440 7948 26480
rect 7988 26440 10444 26480
rect 10484 26440 10493 26480
rect 4876 26312 4916 26440
rect 5155 26356 5164 26396
rect 5204 26356 5300 26396
rect 5347 26356 5356 26396
rect 5396 26356 11884 26396
rect 11924 26356 11933 26396
rect 5260 26312 5300 26356
rect 11980 26312 12020 26692
rect 13084 26648 13124 26692
rect 14764 26648 14804 26692
rect 19660 26648 19700 26692
rect 12346 26608 12355 26648
rect 12395 26608 12404 26648
rect 12451 26608 12460 26648
rect 12500 26608 12631 26648
rect 12857 26608 12940 26648
rect 12980 26608 12988 26648
rect 13028 26608 13037 26648
rect 13084 26608 13708 26648
rect 13748 26608 13757 26648
rect 13891 26608 13900 26648
rect 13940 26608 14476 26648
rect 14516 26608 14525 26648
rect 14764 26608 18412 26648
rect 18452 26608 18461 26648
rect 18883 26608 18892 26648
rect 18932 26608 18988 26648
rect 19028 26608 19063 26648
rect 19468 26608 19700 26648
rect 20009 26608 20140 26648
rect 20180 26608 20189 26648
rect 20297 26608 20419 26648
rect 20468 26608 20477 26648
rect 12364 26564 12404 26608
rect 12364 26524 12844 26564
rect 12884 26524 12893 26564
rect 17347 26524 17356 26564
rect 17396 26524 18508 26564
rect 18548 26524 18557 26564
rect 12117 26440 12126 26480
rect 12494 26440 12503 26480
rect 18028 26440 18988 26480
rect 19028 26440 19037 26480
rect 12643 26356 12652 26396
rect 12692 26356 12788 26396
rect 12748 26312 12788 26356
rect 18028 26354 18068 26440
rect 19468 26396 19508 26608
rect 20524 26564 20564 26692
rect 21676 26564 21716 26776
rect 21868 26732 21908 26776
rect 27148 26732 27188 26776
rect 21850 26692 21859 26732
rect 21899 26692 21908 26732
rect 24739 26692 24748 26732
rect 24788 26692 25507 26732
rect 25547 26692 25556 26732
rect 26275 26692 26284 26732
rect 26324 26692 27188 26732
rect 30586 26692 30595 26732
rect 30635 26692 30700 26732
rect 30740 26692 30775 26732
rect 22051 26608 22060 26648
rect 22100 26608 22109 26648
rect 23587 26608 23596 26648
rect 23636 26608 23788 26648
rect 23828 26608 23837 26648
rect 24521 26608 24556 26648
rect 24596 26608 24652 26648
rect 24692 26608 24701 26648
rect 25795 26608 25804 26648
rect 25844 26608 27244 26648
rect 27284 26608 27293 26648
rect 28169 26608 28300 26648
rect 28340 26608 28349 26648
rect 29155 26608 29164 26648
rect 29204 26608 30028 26648
rect 30068 26608 30787 26648
rect 30827 26608 30836 26648
rect 20524 26524 21716 26564
rect 19891 26440 19900 26480
rect 20268 26440 20277 26480
rect 18010 26314 18019 26354
rect 18059 26314 18068 26354
rect 18136 26356 19508 26396
rect 19564 26356 20660 26396
rect 2659 26272 2668 26312
rect 2708 26272 4916 26312
rect 5011 26272 5020 26312
rect 5060 26272 5068 26312
rect 5108 26272 5191 26312
rect 5260 26272 8140 26312
rect 8180 26272 8189 26312
rect 8803 26272 8812 26312
rect 8852 26272 10196 26312
rect 11107 26272 11116 26312
rect 11156 26272 11308 26312
rect 11348 26272 11357 26312
rect 11980 26272 12172 26312
rect 12212 26272 12221 26312
rect 12730 26272 12739 26312
rect 12779 26272 12788 26312
rect 12844 26272 13507 26312
rect 13547 26272 13556 26312
rect 13603 26272 13612 26312
rect 13652 26272 14668 26312
rect 14708 26272 14717 26312
rect 16291 26272 16300 26312
rect 16340 26272 16348 26312
rect 16388 26272 16471 26312
rect 2092 26188 2476 26228
rect 2516 26188 2525 26228
rect 2844 26188 2956 26228
rect 2996 26188 3004 26228
rect 3044 26188 3956 26228
rect 4003 26188 4012 26228
rect 4052 26188 4684 26228
rect 4724 26188 4733 26228
rect 4924 26188 5548 26228
rect 5588 26188 5597 26228
rect 6377 26188 6499 26228
rect 6548 26188 6557 26228
rect 8986 26188 8995 26228
rect 9035 26188 9580 26228
rect 9620 26188 9629 26228
rect 2092 26144 2132 26188
rect 3916 26144 3956 26188
rect 4924 26144 4964 26188
rect 10156 26144 10196 26272
rect 12844 26228 12884 26272
rect 18136 26270 18176 26356
rect 18883 26272 18892 26312
rect 18932 26272 19084 26312
rect 19124 26272 19133 26312
rect 18127 26230 18136 26270
rect 18176 26230 18185 26270
rect 19564 26228 19604 26356
rect 20506 26272 20515 26312
rect 20555 26272 20564 26312
rect 20524 26228 20564 26272
rect 12802 26188 12844 26228
rect 12884 26188 12893 26228
rect 12956 26188 13324 26228
rect 13364 26188 13516 26228
rect 13556 26188 13565 26228
rect 13769 26188 13891 26228
rect 13940 26188 13949 26228
rect 16963 26188 16972 26228
rect 17012 26188 18067 26228
rect 18403 26188 18412 26228
rect 18452 26188 18461 26228
rect 18883 26188 18892 26228
rect 18932 26188 19604 26228
rect 12844 26144 12884 26188
rect 12956 26144 12996 26188
rect 18027 26186 18067 26188
rect 18027 26146 18056 26186
rect 18096 26146 18105 26186
rect 18412 26144 18452 26188
rect 19564 26144 19604 26188
rect 20044 26188 20564 26228
rect 20044 26144 20084 26188
rect 20620 26144 20660 26356
rect 22060 26228 22100 26608
rect 30892 26564 30932 26776
rect 31075 26608 31084 26648
rect 31124 26608 31255 26648
rect 28195 26524 28204 26564
rect 28244 26524 30932 26564
rect 27665 26440 27674 26480
rect 28042 26440 28051 26480
rect 23875 26356 23884 26396
rect 23924 26356 25940 26396
rect 22627 26272 22636 26312
rect 22676 26272 25180 26312
rect 25220 26272 25229 26312
rect 25385 26272 25507 26312
rect 25556 26272 25565 26312
rect 22042 26188 22051 26228
rect 22091 26188 22100 26228
rect 24844 26188 25228 26228
rect 25268 26188 25420 26228
rect 25460 26188 25469 26228
rect 24844 26144 24884 26188
rect 25900 26144 25940 26356
rect 28588 26356 30124 26396
rect 30164 26356 30173 26396
rect 25987 26272 25996 26312
rect 26036 26272 27052 26312
rect 27092 26272 27101 26312
rect 27689 26272 27820 26312
rect 27860 26272 27869 26312
rect 26179 26188 26188 26228
rect 26228 26188 26428 26228
rect 26468 26188 26477 26228
rect 28588 26144 28628 26356
rect 2083 26104 2092 26144
rect 2132 26104 2141 26144
rect 2266 26104 2275 26144
rect 2315 26104 2324 26144
rect 2284 26060 2324 26104
rect 2842 26135 2860 26144
rect 2842 26095 2851 26135
rect 2900 26104 3031 26144
rect 3209 26104 3340 26144
rect 3380 26104 3389 26144
rect 3916 26104 4012 26144
rect 4052 26104 4300 26144
rect 4340 26104 4349 26144
rect 4570 26104 4579 26144
rect 4619 26104 4780 26144
rect 4820 26104 4964 26144
rect 5033 26104 5164 26144
rect 5204 26104 5213 26144
rect 6874 26104 6883 26144
rect 6932 26104 7063 26144
rect 9370 26104 9379 26144
rect 9428 26104 9559 26144
rect 10156 26104 11500 26144
rect 11540 26104 11549 26144
rect 12329 26104 12460 26144
rect 12500 26104 12509 26144
rect 12556 26104 12676 26144
rect 12716 26104 12725 26144
rect 12840 26104 12849 26144
rect 12889 26104 12898 26144
rect 12952 26104 12961 26144
rect 13001 26104 13010 26144
rect 2891 26095 2900 26104
rect 2842 26094 2900 26095
rect 3340 26060 3380 26104
rect 6346 26062 6355 26102
rect 6395 26062 6404 26102
rect 835 26020 844 26060
rect 884 26020 2188 26060
rect 2228 26020 2237 26060
rect 2284 26020 2476 26060
rect 2516 26020 2525 26060
rect 3340 26020 5356 26060
rect 5396 26020 5405 26060
rect 5731 26020 5740 26060
rect 5780 26020 6163 26060
rect 6203 26020 6212 26060
rect 595 25936 604 25976
rect 644 25936 1132 25976
rect 1172 25936 1181 25976
rect 1385 25936 1516 25976
rect 1556 25936 1565 25976
rect 1769 25936 1900 25976
rect 1940 25936 1949 25976
rect 2266 25936 2275 25976
rect 2315 25936 5260 25976
rect 5300 25936 5309 25976
rect 6364 25892 6404 26062
rect 12556 26060 12596 26104
rect 13075 26093 13084 26133
rect 13124 26093 13133 26133
rect 13210 26104 13219 26144
rect 13259 26104 13268 26144
rect 13400 26104 13409 26144
rect 13460 26104 13589 26144
rect 13673 26104 13722 26144
rect 13762 26104 13804 26144
rect 13844 26104 13853 26144
rect 14266 26104 14275 26144
rect 14315 26104 15340 26144
rect 15380 26104 15389 26144
rect 16483 26104 16492 26144
rect 16532 26104 16675 26144
rect 16715 26104 16724 26144
rect 17347 26104 17356 26144
rect 17396 26104 17972 26144
rect 18346 26104 18355 26144
rect 18395 26104 18452 26144
rect 18494 26104 18503 26144
rect 18543 26104 18552 26144
rect 18691 26104 18700 26144
rect 18740 26104 19084 26144
rect 19124 26104 19133 26144
rect 19555 26104 19564 26144
rect 19604 26104 19613 26144
rect 19660 26104 19756 26144
rect 19796 26104 19805 26144
rect 20035 26104 20044 26144
rect 20084 26104 20093 26144
rect 20620 26104 20668 26144
rect 20708 26104 20717 26144
rect 20803 26104 20812 26144
rect 20852 26104 20983 26144
rect 21370 26104 21379 26144
rect 21419 26104 21428 26144
rect 22339 26104 22348 26144
rect 22388 26104 22435 26144
rect 22475 26104 22519 26144
rect 24355 26104 24364 26144
rect 24404 26104 24556 26144
rect 24596 26104 24605 26144
rect 24730 26104 24739 26144
rect 24779 26104 24788 26144
rect 24835 26104 24844 26144
rect 24884 26104 24893 26144
rect 25018 26135 25036 26144
rect 6787 26020 6796 26060
rect 6836 26020 6845 26060
rect 8227 26020 8236 26060
rect 8276 26020 9216 26060
rect 11395 26020 11404 26060
rect 11444 26020 12596 26060
rect 13084 25976 13124 26093
rect 11779 25936 11788 25976
rect 11828 25936 13124 25976
rect 13228 25976 13268 26104
rect 17356 26060 17396 26104
rect 14851 26020 14860 26060
rect 14900 26020 14909 26060
rect 16204 26020 17396 26060
rect 16204 25976 16244 26020
rect 17932 25976 17972 26104
rect 18508 26060 18548 26104
rect 18089 26020 18220 26060
rect 18260 26020 18269 26060
rect 18499 26020 18508 26060
rect 18548 26020 18590 26060
rect 19660 25976 19700 26104
rect 20044 26060 20084 26104
rect 21388 26060 21428 26104
rect 24748 26060 24788 26104
rect 25018 26095 25027 26135
rect 25076 26104 25207 26144
rect 25673 26104 25708 26144
rect 25748 26104 25804 26144
rect 25844 26104 25853 26144
rect 25900 26135 26324 26144
rect 25900 26104 26275 26135
rect 25067 26095 25076 26104
rect 25018 26094 25076 26095
rect 26266 26095 26275 26104
rect 26315 26095 26324 26135
rect 26633 26104 26764 26144
rect 26804 26104 26813 26144
rect 26266 26094 26324 26095
rect 26858 26080 26892 26120
rect 26932 26080 26941 26120
rect 27209 26104 27340 26144
rect 27380 26104 27389 26144
rect 27715 26104 27724 26144
rect 27764 26104 28628 26144
rect 28684 26272 30604 26312
rect 30644 26272 31276 26312
rect 31316 26272 31325 26312
rect 28684 26144 28724 26272
rect 28771 26188 28780 26228
rect 28820 26188 29356 26228
rect 29396 26188 29405 26228
rect 29356 26144 29396 26188
rect 28684 26104 28780 26144
rect 28820 26104 28829 26144
rect 29338 26104 29347 26144
rect 29387 26104 29396 26144
rect 26858 26060 26898 26080
rect 19747 26020 19756 26060
rect 19796 26020 20084 26060
rect 20131 26020 20140 26060
rect 20180 26020 21428 26060
rect 21484 26020 22272 26060
rect 24748 26020 24844 26060
rect 24884 26020 24893 26060
rect 25705 26020 25714 26060
rect 25754 26020 25900 26060
rect 25940 26020 25949 26060
rect 26371 26020 26380 26060
rect 26420 26020 26898 26060
rect 28841 26020 28972 26060
rect 29012 26020 29021 26060
rect 29155 26020 29164 26060
rect 29204 26020 29213 26060
rect 13228 25936 13804 25976
rect 13844 25936 13853 25976
rect 16195 25936 16204 25976
rect 16244 25936 16253 25976
rect 17417 25936 17548 25976
rect 17588 25936 17597 25976
rect 17932 25936 18412 25976
rect 18452 25936 18461 25976
rect 18595 25936 18604 25976
rect 18644 25936 19468 25976
rect 19508 25936 19700 25976
rect 20371 25936 20380 25976
rect 20420 25936 21388 25976
rect 21428 25936 21437 25976
rect 21484 25892 21524 26020
rect 24067 25936 24076 25976
rect 24116 25936 24364 25976
rect 24404 25936 24413 25976
rect 24835 25936 24844 25976
rect 24884 25936 26956 25976
rect 26996 25936 27005 25976
rect 27977 25936 28108 25976
rect 28148 25936 28157 25976
rect 3043 25852 3052 25892
rect 3092 25852 5452 25892
rect 5492 25852 5501 25892
rect 5827 25852 5836 25892
rect 5876 25852 5932 25892
rect 5972 25852 6007 25892
rect 6364 25852 8332 25892
rect 8372 25852 8381 25892
rect 8611 25852 8620 25892
rect 8660 25852 12652 25892
rect 12692 25852 12701 25892
rect 20269 25852 21524 25892
rect 21763 25852 21772 25892
rect 21812 25852 22828 25892
rect 22868 25852 22877 25892
rect 23779 25852 23788 25892
rect 23828 25852 30892 25892
rect 30932 25852 30941 25892
rect 20269 25808 20309 25852
rect 1516 25768 2860 25808
rect 2900 25768 2909 25808
rect 6883 25768 6892 25808
rect 6932 25768 15244 25808
rect 15284 25768 15293 25808
rect 17635 25768 17644 25808
rect 17684 25768 20309 25808
rect 643 25348 652 25388
rect 692 25348 844 25388
rect 884 25348 893 25388
rect 1097 25348 1228 25388
rect 1268 25348 1277 25388
rect 1516 25304 1556 25768
rect 3103 25684 3112 25724
rect 3480 25684 3489 25724
rect 3715 25684 3724 25724
rect 3764 25684 7564 25724
rect 7604 25684 9004 25724
rect 9044 25684 9053 25724
rect 10877 25684 10886 25724
rect 11254 25684 11263 25724
rect 18651 25684 18660 25724
rect 19028 25684 19037 25724
rect 21283 25684 21292 25724
rect 21332 25684 26092 25724
rect 26132 25684 26141 25724
rect 26425 25684 26434 25724
rect 26802 25684 26811 25724
rect 2380 25600 7468 25640
rect 7508 25600 7517 25640
rect 10060 25600 16876 25640
rect 16916 25600 16925 25640
rect 18115 25600 18124 25640
rect 18164 25600 21772 25640
rect 21812 25600 21821 25640
rect 23875 25600 23884 25640
rect 23924 25600 28148 25640
rect 2380 25472 2420 25600
rect 10060 25556 10100 25600
rect 28108 25556 28148 25600
rect 3052 25516 5548 25556
rect 5588 25516 5597 25556
rect 7834 25516 7843 25556
rect 7883 25516 8140 25556
rect 8180 25516 8189 25556
rect 8851 25516 8860 25556
rect 8900 25516 10100 25556
rect 11683 25516 11692 25556
rect 11732 25516 12308 25556
rect 1603 25432 1612 25472
rect 1652 25432 1783 25472
rect 2371 25432 2380 25472
rect 2420 25432 2429 25472
rect 3052 25388 3092 25516
rect 5443 25432 5452 25472
rect 5492 25463 7652 25472
rect 5492 25432 7612 25463
rect 9187 25432 9196 25472
rect 9236 25432 10060 25472
rect 10100 25432 10109 25472
rect 10627 25432 10636 25472
rect 10676 25432 10780 25472
rect 10820 25432 10829 25472
rect 11587 25432 11596 25472
rect 11636 25432 11788 25472
rect 11828 25432 11837 25472
rect 7612 25414 7652 25423
rect 12268 25388 12308 25516
rect 14530 25516 16108 25556
rect 16148 25516 16157 25556
rect 21082 25516 21091 25556
rect 21131 25516 21580 25556
rect 21620 25516 21629 25556
rect 21676 25516 23980 25556
rect 24020 25516 24029 25556
rect 25396 25516 26860 25556
rect 26900 25516 26909 25556
rect 28099 25516 28108 25556
rect 28148 25516 28157 25556
rect 14530 25472 14570 25516
rect 21676 25472 21716 25516
rect 14057 25432 14188 25472
rect 14228 25432 14237 25472
rect 14428 25432 14570 25472
rect 14755 25432 14764 25472
rect 14804 25432 16436 25472
rect 18691 25432 18700 25472
rect 18740 25432 18749 25472
rect 19075 25432 19084 25472
rect 19124 25432 21716 25472
rect 25097 25432 25228 25472
rect 25268 25432 25277 25472
rect 14428 25388 14468 25432
rect 16396 25388 16436 25432
rect 2563 25348 2572 25388
rect 2612 25348 2659 25388
rect 2699 25348 2743 25388
rect 3043 25348 3052 25388
rect 3092 25348 3101 25388
rect 3235 25348 3244 25388
rect 3284 25348 3293 25388
rect 5251 25348 5260 25388
rect 5300 25348 5644 25388
rect 5684 25348 6258 25388
rect 6979 25348 6988 25388
rect 7028 25348 7037 25388
rect 7171 25348 7180 25388
rect 7220 25348 7412 25388
rect 8611 25348 8620 25388
rect 8660 25348 9100 25388
rect 9140 25348 9149 25388
rect 9571 25348 9580 25388
rect 9620 25348 10732 25388
rect 10772 25348 10781 25388
rect 12268 25348 12329 25388
rect 12425 25348 12556 25388
rect 12596 25348 13324 25388
rect 13364 25348 13804 25388
rect 13844 25348 13852 25388
rect 13892 25348 14468 25388
rect 14537 25348 14668 25388
rect 14708 25348 14717 25388
rect 15964 25348 16108 25388
rect 16148 25348 16157 25388
rect 16387 25348 16396 25388
rect 16436 25348 16445 25388
rect 17539 25348 17548 25388
rect 17588 25348 17597 25388
rect 6218 25304 6258 25348
rect 6988 25304 7028 25348
rect 7372 25304 7412 25348
rect 12289 25315 12329 25348
rect 1516 25264 1804 25304
rect 1844 25264 1853 25304
rect 1987 25264 1996 25304
rect 2036 25264 2380 25304
rect 2420 25264 2429 25304
rect 2510 25264 2519 25304
rect 2559 25264 2568 25304
rect 2748 25264 2757 25304
rect 2797 25264 2956 25304
rect 2996 25264 3005 25304
rect 3340 25264 3427 25304
rect 3467 25264 5740 25304
rect 5780 25264 5789 25304
rect 5923 25264 5932 25304
rect 5972 25264 6103 25304
rect 6211 25264 6220 25304
rect 6260 25264 6269 25304
rect 6377 25264 6508 25304
rect 6548 25264 6557 25304
rect 6761 25264 6892 25304
rect 6932 25264 6941 25304
rect 6988 25264 7276 25304
rect 7316 25264 7325 25304
rect 7372 25264 7651 25304
rect 7691 25264 7700 25304
rect 8323 25264 8332 25304
rect 8384 25264 8503 25304
rect 9283 25264 9292 25304
rect 9332 25264 9955 25304
rect 9995 25264 10004 25304
rect 10313 25264 10348 25304
rect 10388 25264 10444 25304
rect 10484 25264 10493 25304
rect 10627 25264 10636 25304
rect 10676 25264 10685 25304
rect 10819 25264 10828 25304
rect 10907 25264 10999 25304
rect 11273 25264 11404 25304
rect 11444 25264 11453 25304
rect 11500 25264 11519 25304
rect 11559 25264 11568 25304
rect 11683 25264 11692 25304
rect 11732 25264 11863 25304
rect 11911 25264 11920 25304
rect 11960 25264 11969 25304
rect 12046 25264 12067 25304
rect 12107 25264 12116 25304
rect 12172 25264 12184 25304
rect 12224 25264 12233 25304
rect 12289 25275 12305 25315
rect 12345 25275 12354 25315
rect 12460 25304 12500 25348
rect 14428 25304 14468 25348
rect 15964 25304 16004 25348
rect 18700 25304 18740 25432
rect 20044 25304 20084 25432
rect 25396 25388 25436 25516
rect 25577 25463 25708 25472
rect 25577 25432 25676 25463
rect 25748 25432 26324 25472
rect 26371 25432 26380 25472
rect 26420 25432 26516 25472
rect 26947 25432 26956 25472
rect 26996 25432 27005 25472
rect 30979 25432 30988 25472
rect 31028 25432 31037 25472
rect 25676 25414 25716 25423
rect 26284 25388 26324 25432
rect 21763 25348 21772 25388
rect 21812 25348 21821 25388
rect 23683 25348 23692 25388
rect 23732 25348 25028 25388
rect 25315 25348 25324 25388
rect 25364 25348 25436 25388
rect 26153 25348 26284 25388
rect 26324 25348 26333 25388
rect 21388 25304 21428 25313
rect 24988 25304 25028 25348
rect 26284 25304 26324 25348
rect 26476 25304 26516 25432
rect 26851 25348 26860 25388
rect 26900 25348 26911 25388
rect 12442 25264 12451 25304
rect 12491 25264 12500 25304
rect 12701 25264 12745 25304
rect 12785 25264 12794 25304
rect 12861 25264 12870 25304
rect 12910 25264 12919 25304
rect 12979 25264 12988 25304
rect 13028 25264 13037 25304
rect 13097 25264 13216 25304
rect 13268 25264 13666 25304
rect 13706 25264 13715 25304
rect 14428 25264 14524 25304
rect 14564 25264 14573 25304
rect 14729 25264 14839 25304
rect 14900 25264 14909 25304
rect 14986 25264 14995 25304
rect 15035 25264 15092 25304
rect 15139 25264 15148 25304
rect 15188 25264 15820 25304
rect 15860 25264 15869 25304
rect 15964 25264 15995 25304
rect 16035 25264 16044 25304
rect 16195 25264 16204 25304
rect 16244 25264 16375 25304
rect 16762 25264 16771 25304
rect 16811 25264 17068 25304
rect 17108 25264 17117 25304
rect 18700 25264 18988 25304
rect 19028 25264 19037 25304
rect 19843 25264 19852 25304
rect 19892 25264 20084 25304
rect 20131 25264 20140 25304
rect 20180 25264 20189 25304
rect 20332 25264 20563 25304
rect 20603 25264 20612 25304
rect 21353 25264 21388 25304
rect 21428 25264 21484 25304
rect 21524 25264 21676 25304
rect 21716 25264 21725 25304
rect 21946 25264 21955 25304
rect 21995 25264 22348 25304
rect 22388 25264 22397 25304
rect 23884 25264 24748 25304
rect 24788 25264 24797 25304
rect 24979 25264 24988 25304
rect 25028 25264 25037 25304
rect 25314 25264 25420 25304
rect 25485 25264 25494 25304
rect 25690 25264 25699 25304
rect 25739 25264 25748 25304
rect 26083 25264 26092 25304
rect 26132 25264 26141 25304
rect 26266 25264 26275 25304
rect 26315 25264 26324 25304
rect 26371 25264 26380 25304
rect 26420 25264 26429 25304
rect 26476 25264 26563 25304
rect 26603 25264 26612 25304
rect 2519 25220 2559 25264
rect 883 25180 892 25220
rect 932 25180 1324 25220
rect 1364 25180 1373 25220
rect 1603 25180 1612 25220
rect 1652 25180 2559 25220
rect 643 25096 652 25136
rect 692 25096 988 25136
rect 1028 25096 1037 25136
rect 1865 25096 1987 25136
rect 2036 25096 2045 25136
rect 2842 25096 2851 25136
rect 2891 25096 3148 25136
rect 3188 25096 3197 25136
rect 3340 25052 3380 25264
rect 5932 25246 5972 25255
rect 5443 25180 5452 25220
rect 5492 25180 5836 25220
rect 5876 25180 5885 25220
rect 5836 25136 5876 25180
rect 6892 25136 6932 25264
rect 7276 25220 7316 25264
rect 7276 25180 8179 25220
rect 8219 25180 8228 25220
rect 8515 25180 8524 25220
rect 8564 25180 9340 25220
rect 9380 25180 9389 25220
rect 10636 25136 10676 25264
rect 11500 25220 11540 25264
rect 11919 25220 11959 25264
rect 11500 25180 11959 25220
rect 5225 25096 5356 25136
rect 5396 25096 5405 25136
rect 5836 25096 6932 25136
rect 6979 25096 6988 25136
rect 7028 25096 7037 25136
rect 7834 25096 7843 25136
rect 7883 25096 10676 25136
rect 11011 25096 11020 25136
rect 11060 25096 11068 25136
rect 11108 25096 11191 25136
rect 2275 25012 2284 25052
rect 2324 25012 3380 25052
rect 6988 25052 7028 25096
rect 6988 25012 11404 25052
rect 11444 25012 11453 25052
rect 11500 24968 11540 25180
rect 12046 25136 12086 25264
rect 12172 25220 12212 25264
rect 12748 25220 12788 25264
rect 12137 25180 12172 25220
rect 12212 25180 12221 25220
rect 12329 25180 12451 25220
rect 12500 25180 12509 25220
rect 12739 25180 12748 25220
rect 12788 25180 12797 25220
rect 12879 25136 12919 25264
rect 12988 25220 13028 25264
rect 15052 25220 15092 25264
rect 20140 25220 20180 25264
rect 12988 25180 13036 25220
rect 13076 25180 13085 25220
rect 15052 25180 17260 25220
rect 17300 25180 17309 25220
rect 18499 25180 18508 25220
rect 18548 25180 20180 25220
rect 20332 25136 20372 25264
rect 21388 25255 21428 25264
rect 20611 25180 20620 25220
rect 20660 25180 21086 25220
rect 21126 25180 21135 25220
rect 21562 25180 21571 25220
rect 21611 25180 21868 25220
rect 21908 25180 21917 25220
rect 22444 25180 22924 25220
rect 22964 25180 22973 25220
rect 22444 25136 22484 25180
rect 23884 25136 23924 25264
rect 25151 25222 25160 25262
rect 25200 25222 25220 25262
rect 25180 25220 25220 25222
rect 25708 25220 25748 25264
rect 25180 25180 25268 25220
rect 12046 25096 12844 25136
rect 12884 25096 12919 25136
rect 13027 25096 13036 25136
rect 13076 25096 13085 25136
rect 13363 25096 13372 25136
rect 13412 25096 14380 25136
rect 14420 25096 14429 25136
rect 15139 25096 15148 25136
rect 15188 25096 15197 25136
rect 15331 25096 15340 25136
rect 15380 25096 16195 25136
rect 16235 25096 16244 25136
rect 19529 25096 19660 25136
rect 19700 25096 19709 25136
rect 20323 25096 20332 25136
rect 20372 25096 20381 25136
rect 20633 25096 20716 25136
rect 20756 25096 20764 25136
rect 20804 25096 20813 25136
rect 21283 25096 21292 25136
rect 21332 25096 22484 25136
rect 22723 25096 22732 25136
rect 22772 25096 23884 25136
rect 23924 25096 23933 25136
rect 24067 25096 24076 25136
rect 24116 25096 24125 25136
rect 12046 25052 12086 25096
rect 11587 25012 11596 25052
rect 11636 25012 12086 25052
rect 4343 24928 4352 24968
rect 4720 24928 4729 24968
rect 8803 24928 8812 24968
rect 8852 24928 11540 24968
rect 12117 24928 12126 24968
rect 12494 24928 12503 24968
rect 13036 24884 13076 25096
rect 10435 24844 10444 24884
rect 10484 24844 10636 24884
rect 10676 24844 11020 24884
rect 11060 24844 11069 24884
rect 13036 24844 14406 24884
rect 1577 24760 1708 24800
rect 1748 24760 1757 24800
rect 8044 24760 11308 24800
rect 11348 24760 11357 24800
rect 13690 24760 13699 24800
rect 13739 24760 13900 24800
rect 13940 24760 13949 24800
rect 1882 24676 1891 24716
rect 1931 24676 4588 24716
rect 4628 24676 4637 24716
rect 6106 24676 6115 24716
rect 6155 24676 7468 24716
rect 7508 24676 7517 24716
rect 8044 24632 8084 24760
rect 14366 24716 14406 24844
rect 15148 24716 15188 25096
rect 15235 25012 15244 25052
rect 15284 25012 23788 25052
rect 23828 25012 23837 25052
rect 17452 24928 19372 24968
rect 19412 24928 19421 24968
rect 19891 24928 19900 24968
rect 20268 24928 20277 24968
rect 17452 24800 17492 24928
rect 17539 24844 17548 24884
rect 17588 24844 20620 24884
rect 20660 24844 20669 24884
rect 22540 24844 23780 24884
rect 22540 24800 22580 24844
rect 23740 24800 23780 24844
rect 16195 24760 16204 24800
rect 16244 24760 17452 24800
rect 17492 24760 17501 24800
rect 18124 24760 19843 24800
rect 19892 24760 19901 24800
rect 20393 24760 20515 24800
rect 20564 24760 20573 24800
rect 21667 24760 21676 24800
rect 21716 24760 21725 24800
rect 21859 24760 21868 24800
rect 21908 24760 22156 24800
rect 22196 24760 22205 24800
rect 22531 24760 22540 24800
rect 22580 24760 22589 24800
rect 23098 24760 23107 24800
rect 23156 24760 23287 24800
rect 23722 24760 23731 24800
rect 23771 24760 23788 24800
rect 23828 24760 23940 24800
rect 8410 24676 8419 24716
rect 8459 24676 9196 24716
rect 9236 24676 9245 24716
rect 9379 24676 9388 24716
rect 9428 24676 9772 24716
rect 9812 24676 10292 24716
rect 10252 24632 10292 24676
rect 13228 24676 13324 24716
rect 13364 24676 13373 24716
rect 13498 24707 13516 24716
rect 13228 24632 13268 24676
rect 13498 24667 13507 24707
rect 13556 24676 13687 24716
rect 13789 24676 13996 24716
rect 14036 24676 14045 24716
rect 14366 24676 14708 24716
rect 14755 24676 14764 24716
rect 14804 24676 14813 24716
rect 15130 24676 15139 24716
rect 15179 24676 15188 24716
rect 15265 24676 17068 24716
rect 17108 24676 17117 24716
rect 13547 24667 13556 24676
rect 13498 24666 13556 24667
rect 13789 24632 13829 24676
rect 14668 24632 14708 24676
rect 14764 24632 14804 24676
rect 15265 24632 15305 24676
rect 18124 24632 18164 24760
rect 21676 24716 21716 24760
rect 24076 24716 24116 25096
rect 25228 25052 25268 25180
rect 25420 25180 25748 25220
rect 25420 25136 25460 25180
rect 25411 25096 25420 25136
rect 25460 25096 25469 25136
rect 25699 25096 25708 25136
rect 25748 25096 25891 25136
rect 25931 25096 25940 25136
rect 25228 25012 25996 25052
rect 26036 25012 26045 25052
rect 26092 24968 26132 25264
rect 26380 25220 26420 25264
rect 26871 25220 26911 25348
rect 26956 25304 26996 25432
rect 30988 25388 31028 25432
rect 27043 25348 27052 25388
rect 27092 25348 27340 25388
rect 27380 25348 27389 25388
rect 27497 25348 27628 25388
rect 27668 25348 31028 25388
rect 27532 25304 27572 25348
rect 26956 25264 26999 25304
rect 27039 25264 27048 25304
rect 27130 25264 27139 25304
rect 27179 25264 27188 25304
rect 27235 25264 27244 25304
rect 27284 25264 27415 25304
rect 27514 25264 27523 25304
rect 27563 25264 27572 25304
rect 28745 25264 28780 25304
rect 28820 25264 28876 25304
rect 28916 25264 28925 25304
rect 29635 25264 29644 25304
rect 29684 25264 29932 25304
rect 29972 25264 29981 25304
rect 30499 25264 30508 25304
rect 30548 25264 30557 25304
rect 30787 25264 30796 25304
rect 30836 25264 30845 25304
rect 27148 25220 27188 25264
rect 30508 25220 30548 25264
rect 26333 25180 26380 25220
rect 26420 25180 26429 25220
rect 26537 25180 26668 25220
rect 26708 25180 26717 25220
rect 26862 25180 26871 25220
rect 26911 25180 26920 25220
rect 27043 25180 27052 25220
rect 27092 25180 27188 25220
rect 27244 25180 27831 25220
rect 27871 25180 28108 25220
rect 28148 25180 28157 25220
rect 28579 25180 28588 25220
rect 28628 25180 28963 25220
rect 29003 25180 29012 25220
rect 29068 25180 30548 25220
rect 27244 25136 27284 25180
rect 29068 25136 29108 25180
rect 26467 25096 26476 25136
rect 26516 25096 27284 25136
rect 27331 25096 27340 25136
rect 27380 25096 27619 25136
rect 27659 25096 27668 25136
rect 27715 25096 27724 25136
rect 27764 25096 29108 25136
rect 29705 25096 29836 25136
rect 29876 25096 29885 25136
rect 29932 25096 30691 25136
rect 30731 25096 30740 25136
rect 18220 24676 18836 24716
rect 18979 24676 18988 24716
rect 19028 24676 20660 24716
rect 2266 24592 2275 24632
rect 2324 24592 2455 24632
rect 2755 24592 2764 24632
rect 2804 24592 4108 24632
rect 4148 24592 4157 24632
rect 4387 24592 4396 24632
rect 4436 24592 5740 24632
rect 5780 24592 5789 24632
rect 8026 24592 8035 24632
rect 8075 24592 8084 24632
rect 8515 24592 8524 24632
rect 8564 24592 8702 24632
rect 8742 24592 8751 24632
rect 8899 24592 8908 24632
rect 8948 24592 8957 24632
rect 9004 24623 9091 24632
rect 4396 24548 4436 24592
rect 8908 24548 8948 24592
rect 9044 24592 9091 24623
rect 9161 24592 9292 24632
rect 9332 24592 9341 24632
rect 9475 24592 9484 24632
rect 9549 24592 9655 24632
rect 10234 24592 10243 24632
rect 10283 24592 10292 24632
rect 11788 24592 12364 24632
rect 12404 24592 12413 24632
rect 13210 24592 13219 24632
rect 13259 24592 13268 24632
rect 13324 24623 13364 24632
rect 9004 24548 9044 24583
rect 11788 24548 11828 24592
rect 13590 24592 13599 24632
rect 13639 24592 13652 24632
rect 13771 24592 13780 24632
rect 13820 24592 13829 24632
rect 14057 24623 14188 24632
rect 14057 24592 14179 24623
rect 14228 24592 14237 24632
rect 14659 24592 14668 24632
rect 14708 24592 14717 24632
rect 14764 24592 14790 24632
rect 14830 24592 14851 24632
rect 14908 24592 14917 24632
rect 14996 24592 15097 24632
rect 15244 24592 15305 24632
rect 15514 24592 15523 24632
rect 15563 24592 15820 24632
rect 15860 24592 15869 24632
rect 18115 24592 18124 24632
rect 18164 24592 18173 24632
rect 13324 24548 13364 24583
rect 13612 24548 13652 24592
rect 14170 24583 14179 24592
rect 14219 24583 14228 24592
rect 14170 24582 14228 24583
rect 15244 24548 15284 24592
rect 18220 24548 18260 24676
rect 18796 24632 18836 24676
rect 19948 24632 19988 24676
rect 20620 24632 20660 24676
rect 21484 24676 21580 24716
rect 21620 24676 21629 24716
rect 21676 24676 22815 24716
rect 21484 24632 21524 24676
rect 22775 24632 22815 24676
rect 22924 24676 23308 24716
rect 23348 24676 23357 24716
rect 23404 24676 24116 24716
rect 24172 24928 26764 24968
rect 26804 24928 26813 24968
rect 22924 24632 22964 24676
rect 23404 24632 23444 24676
rect 24172 24632 24212 24928
rect 27340 24884 27380 25096
rect 29932 25052 29972 25096
rect 30796 25052 30836 25264
rect 28291 25012 28300 25052
rect 28340 25012 29972 25052
rect 30019 25012 30028 25052
rect 30068 25012 30836 25052
rect 27665 24928 27674 24968
rect 28042 24928 28051 24968
rect 28099 24928 28108 24968
rect 28148 24928 30412 24968
rect 30452 24928 31468 24968
rect 31508 24928 31517 24968
rect 24643 24844 24652 24884
rect 24692 24844 25748 24884
rect 24451 24760 24460 24800
rect 24500 24760 25119 24800
rect 25193 24760 25219 24800
rect 25259 24760 25324 24800
rect 25364 24760 25373 24800
rect 25079 24716 25119 24760
rect 25708 24716 25748 24844
rect 26092 24844 27380 24884
rect 28675 24844 28684 24884
rect 28724 24844 30796 24884
rect 30836 24844 30845 24884
rect 26092 24800 26132 24844
rect 24259 24676 24268 24716
rect 24308 24676 24692 24716
rect 24835 24676 24844 24716
rect 24884 24676 24893 24716
rect 25079 24676 25172 24716
rect 24652 24632 24692 24676
rect 24844 24632 24884 24676
rect 25132 24632 25172 24676
rect 25228 24676 25516 24716
rect 25556 24676 25565 24716
rect 25612 24676 25748 24716
rect 26034 24760 26092 24800
rect 26132 24760 26141 24800
rect 26537 24760 26572 24800
rect 26612 24760 26668 24800
rect 26708 24760 26717 24800
rect 28003 24760 28012 24800
rect 28052 24760 28492 24800
rect 28532 24760 28541 24800
rect 28867 24760 28876 24800
rect 28916 24760 30028 24800
rect 30068 24760 31276 24800
rect 31316 24760 31325 24800
rect 18307 24592 18316 24632
rect 18356 24592 18365 24632
rect 18490 24623 18508 24632
rect 1027 24508 1036 24548
rect 1076 24508 1324 24548
rect 1364 24508 1373 24548
rect 1420 24508 2112 24548
rect 4204 24508 4436 24548
rect 1420 24464 1460 24508
rect 4204 24464 4244 24508
rect 6796 24464 6836 24528
rect 8707 24508 8716 24548
rect 8756 24508 8948 24548
rect 8995 24508 9004 24548
rect 9044 24508 9411 24548
rect 9451 24508 9460 24548
rect 9859 24508 9868 24548
rect 9908 24508 10004 24548
rect 10051 24508 10060 24548
rect 10100 24508 10109 24548
rect 11779 24508 11788 24548
rect 11828 24508 11837 24548
rect 13123 24508 13132 24548
rect 13172 24508 13364 24548
rect 13603 24508 13612 24548
rect 13652 24508 13695 24548
rect 14323 24508 14332 24548
rect 14372 24508 14476 24548
rect 14516 24508 15284 24548
rect 931 24424 940 24464
rect 980 24424 1460 24464
rect 4195 24424 4204 24464
rect 4244 24424 4253 24464
rect 5539 24424 5548 24464
rect 5588 24424 5597 24464
rect 5923 24424 5932 24464
rect 5972 24424 6836 24464
rect 5548 24380 5588 24424
rect 9964 24380 10004 24508
rect 16780 24464 16820 24528
rect 17731 24508 17740 24548
rect 17780 24508 18260 24548
rect 18316 24548 18356 24592
rect 18490 24583 18499 24623
rect 18548 24592 18679 24632
rect 18796 24592 19276 24632
rect 19316 24592 19325 24632
rect 19459 24592 19468 24632
rect 19533 24592 19639 24632
rect 19939 24592 19948 24632
rect 19988 24592 19997 24632
rect 20297 24592 20332 24632
rect 20372 24592 20428 24632
rect 20468 24592 20477 24632
rect 20611 24592 20620 24632
rect 20660 24592 20669 24632
rect 21182 24592 21292 24632
rect 21344 24592 21362 24632
rect 21475 24592 21484 24632
rect 21524 24592 21533 24632
rect 21580 24592 22334 24632
rect 22374 24592 22383 24632
rect 22531 24592 22540 24632
rect 22580 24592 22589 24632
rect 22636 24623 22676 24632
rect 18539 24583 18548 24592
rect 18490 24582 18548 24583
rect 18316 24508 18452 24548
rect 18595 24508 18604 24548
rect 18644 24508 18652 24548
rect 18692 24508 18775 24548
rect 19171 24508 19180 24548
rect 19220 24508 19229 24548
rect 19386 24508 19395 24548
rect 19435 24508 19756 24548
rect 19796 24508 19805 24548
rect 20995 24508 21004 24548
rect 21044 24508 21139 24548
rect 21179 24508 21188 24548
rect 18412 24464 18452 24508
rect 19180 24464 19220 24508
rect 21580 24464 21620 24592
rect 22540 24548 22580 24592
rect 21955 24508 21964 24548
rect 22004 24508 22580 24548
rect 22766 24592 22775 24632
rect 22815 24592 22824 24632
rect 22906 24592 22915 24632
rect 22955 24592 22964 24632
rect 23011 24592 23020 24632
rect 23060 24592 23116 24632
rect 23156 24592 23191 24632
rect 23395 24592 23404 24632
rect 23444 24592 23453 24632
rect 23774 24592 23884 24632
rect 23936 24592 23954 24632
rect 24067 24592 24076 24632
rect 24116 24592 24125 24632
rect 24172 24592 24198 24632
rect 24238 24592 24247 24632
rect 24415 24623 24460 24632
rect 22636 24548 22676 24583
rect 24076 24548 24116 24592
rect 24316 24590 24356 24599
rect 24313 24550 24316 24590
rect 24455 24592 24460 24623
rect 24500 24592 24586 24632
rect 24643 24592 24652 24632
rect 24692 24592 24701 24632
rect 24844 24592 24887 24632
rect 24927 24592 24936 24632
rect 25123 24592 25132 24632
rect 25172 24592 25181 24632
rect 24415 24574 24455 24583
rect 24313 24548 24356 24550
rect 25228 24548 25268 24676
rect 25612 24632 25652 24676
rect 26034 24632 26074 24760
rect 26141 24676 26188 24716
rect 26228 24676 26237 24716
rect 26915 24676 26956 24716
rect 26996 24676 27005 24716
rect 27483 24676 27532 24716
rect 27572 24676 27614 24716
rect 27654 24676 27663 24716
rect 27811 24676 27820 24716
rect 27860 24676 28300 24716
rect 28340 24676 28349 24716
rect 28972 24676 29836 24716
rect 29876 24676 29885 24716
rect 26188 24632 26228 24676
rect 26915 24632 26955 24676
rect 28972 24632 29012 24676
rect 25402 24623 25652 24632
rect 25402 24583 25411 24623
rect 25451 24592 25652 24623
rect 25699 24592 25708 24632
rect 25748 24592 25900 24632
rect 25940 24592 25949 24632
rect 26016 24592 26025 24632
rect 26065 24592 26074 24632
rect 26179 24592 26188 24632
rect 26228 24592 26237 24632
rect 26360 24592 26369 24632
rect 26420 24592 26540 24632
rect 26668 24623 26708 24632
rect 25451 24583 25460 24592
rect 25402 24582 25460 24583
rect 26899 24592 26908 24632
rect 26948 24592 26957 24632
rect 27052 24592 27138 24632
rect 27178 24592 27187 24632
rect 27322 24592 27331 24632
rect 27371 24592 27380 24632
rect 27427 24592 27436 24632
rect 27476 24592 27820 24632
rect 27860 24592 27869 24632
rect 27916 24623 27956 24632
rect 26668 24548 26708 24583
rect 27052 24548 27092 24592
rect 27340 24548 27380 24592
rect 28099 24592 28108 24632
rect 28148 24592 29012 24632
rect 29338 24592 29347 24632
rect 29396 24592 29527 24632
rect 27916 24548 27956 24583
rect 22636 24508 22732 24548
rect 22772 24508 22836 24548
rect 23011 24508 23020 24548
rect 23060 24508 23260 24548
rect 23300 24508 23309 24548
rect 23971 24508 23980 24548
rect 24020 24508 24116 24548
rect 24163 24508 24172 24548
rect 24212 24541 24356 24548
rect 24212 24508 24353 24541
rect 24713 24508 24796 24548
rect 24836 24508 24844 24548
rect 24884 24508 24893 24548
rect 25018 24508 25027 24548
rect 25067 24508 25268 24548
rect 25555 24508 25564 24548
rect 25604 24508 25613 24548
rect 26668 24508 26860 24548
rect 26900 24508 26909 24548
rect 27043 24508 27052 24548
rect 27092 24508 27101 24548
rect 27331 24508 27340 24548
rect 27380 24508 27427 24548
rect 27916 24508 28684 24548
rect 28724 24508 28733 24548
rect 28841 24508 28972 24548
rect 29012 24508 29021 24548
rect 29731 24508 29740 24548
rect 29780 24508 29789 24548
rect 22636 24464 22676 24508
rect 23020 24464 23060 24508
rect 25564 24464 25604 24508
rect 11779 24424 11788 24464
rect 11828 24424 12556 24464
rect 12596 24424 12605 24464
rect 13027 24424 13036 24464
rect 13076 24424 13516 24464
rect 13556 24424 13565 24464
rect 14947 24424 14956 24464
rect 14996 24424 15148 24464
rect 15188 24424 15197 24464
rect 16780 24424 17644 24464
rect 17684 24424 17693 24464
rect 18124 24424 18220 24464
rect 18260 24424 18269 24464
rect 18412 24424 20236 24464
rect 20276 24424 20285 24464
rect 20803 24424 20812 24464
rect 20852 24424 21292 24464
rect 21332 24424 21620 24464
rect 21667 24424 21676 24464
rect 21716 24424 22676 24464
rect 22819 24424 22828 24464
rect 22868 24424 23060 24464
rect 23299 24424 23308 24464
rect 23348 24424 25604 24464
rect 25961 24424 26092 24464
rect 26132 24424 26141 24464
rect 26755 24424 26764 24464
rect 26804 24424 26812 24464
rect 26852 24424 26935 24464
rect 27427 24424 27436 24464
rect 27476 24424 28396 24464
rect 28436 24424 28445 24464
rect 18124 24380 18164 24424
rect 355 24340 364 24380
rect 404 24340 1084 24380
rect 1124 24340 1133 24380
rect 4937 24340 4972 24380
rect 5012 24340 5068 24380
rect 5108 24340 5117 24380
rect 5548 24340 5972 24380
rect 6499 24340 6508 24380
rect 6548 24340 7660 24380
rect 7700 24340 7709 24380
rect 8419 24340 8428 24380
rect 8468 24340 8707 24380
rect 8747 24340 8756 24380
rect 9964 24340 10444 24380
rect 10484 24340 10493 24380
rect 12041 24340 12172 24380
rect 12212 24340 12221 24380
rect 13987 24340 13996 24380
rect 14036 24340 18164 24380
rect 18211 24340 18220 24380
rect 18260 24340 21484 24380
rect 21524 24340 21533 24380
rect 21763 24340 21772 24380
rect 21812 24340 22339 24380
rect 22379 24340 22444 24380
rect 22484 24340 22548 24380
rect 25987 24340 25996 24380
rect 26036 24340 26371 24380
rect 26411 24340 26420 24380
rect 27610 24340 27619 24380
rect 27659 24340 27668 24380
rect 28771 24340 28780 24380
rect 28820 24340 28972 24380
rect 29012 24340 29021 24380
rect 5932 24296 5972 24340
rect 27628 24296 27668 24340
rect 5932 24256 10540 24296
rect 10580 24256 10589 24296
rect 19459 24256 19468 24296
rect 19508 24256 23116 24296
rect 23156 24256 23165 24296
rect 27619 24256 27628 24296
rect 27668 24256 27715 24296
rect 3103 24172 3112 24212
rect 3480 24172 3489 24212
rect 6019 24172 6028 24212
rect 6068 24172 10100 24212
rect 10877 24172 10886 24212
rect 11254 24172 11263 24212
rect 13315 24172 13324 24212
rect 13364 24172 14188 24212
rect 14228 24172 15724 24212
rect 15764 24172 15773 24212
rect 16195 24172 16204 24212
rect 16244 24172 18548 24212
rect 18651 24172 18660 24212
rect 19028 24172 19037 24212
rect 19171 24172 19180 24212
rect 19220 24172 25036 24212
rect 25076 24172 25085 24212
rect 26425 24172 26434 24212
rect 26802 24172 26811 24212
rect 10060 24128 10100 24172
rect 18508 24128 18548 24172
rect 1219 24088 1228 24128
rect 1268 24088 5548 24128
rect 5588 24088 5597 24128
rect 5731 24088 5740 24128
rect 5780 24088 8756 24128
rect 10060 24088 17012 24128
rect 18508 24088 21868 24128
rect 21908 24088 21917 24128
rect 24599 24088 28588 24128
rect 28628 24088 28637 24128
rect 8716 24044 8756 24088
rect 16972 24044 17012 24088
rect 1027 24004 1036 24044
rect 1076 24004 2380 24044
rect 2420 24004 2429 24044
rect 4457 24004 4588 24044
rect 4628 24004 4637 24044
rect 6163 24004 6172 24044
rect 6212 24004 8620 24044
rect 8660 24004 8669 24044
rect 8716 24004 9964 24044
rect 10004 24004 10013 24044
rect 10810 24004 10819 24044
rect 10859 24004 13228 24044
rect 13268 24004 13277 24044
rect 13516 24004 14668 24044
rect 14708 24004 14717 24044
rect 16387 24004 16396 24044
rect 16436 24004 16876 24044
rect 16916 24004 16925 24044
rect 16972 24004 23308 24044
rect 23348 24004 23357 24044
rect 24355 24004 24364 24044
rect 24404 24004 24460 24044
rect 24500 24004 24535 24044
rect 6988 23920 10540 23960
rect 10580 23920 10589 23960
rect 12643 23920 12652 23960
rect 12692 23920 12748 23960
rect 12788 23920 12852 23960
rect 12940 23920 13420 23960
rect 13460 23920 13469 23960
rect 1507 23836 1516 23876
rect 1556 23836 1565 23876
rect 3235 23836 3244 23876
rect 3284 23836 4436 23876
rect 4396 23792 4436 23836
rect 4684 23836 5972 23876
rect 2275 23752 2284 23792
rect 2324 23752 2563 23792
rect 2603 23752 2612 23792
rect 3811 23752 3820 23792
rect 3860 23752 4108 23792
rect 4148 23752 4157 23792
rect 4387 23752 4396 23792
rect 4436 23752 4445 23792
rect 4684 23708 4724 23836
rect 5932 23792 5972 23836
rect 6988 23792 7028 23920
rect 12652 23876 12692 23920
rect 12940 23876 12980 23920
rect 7363 23836 7372 23876
rect 7412 23836 8852 23876
rect 9091 23836 9100 23876
rect 9140 23836 9292 23876
rect 9332 23836 9341 23876
rect 9619 23836 9628 23876
rect 9668 23836 10156 23876
rect 10196 23836 10205 23876
rect 10313 23836 10444 23876
rect 10484 23836 10493 23876
rect 10828 23836 12692 23876
rect 12748 23836 12980 23876
rect 13036 23836 13132 23876
rect 13172 23836 13181 23876
rect 8812 23817 8852 23836
rect 8812 23792 8859 23817
rect 10060 23792 10100 23836
rect 10828 23792 10868 23836
rect 12748 23792 12788 23836
rect 13036 23792 13076 23836
rect 13516 23792 13556 24004
rect 14659 23920 14668 23960
rect 14708 23920 14996 23960
rect 17251 23920 17260 23960
rect 17300 23920 19516 23960
rect 19556 23920 19565 23960
rect 19939 23920 19948 23960
rect 19988 23920 22156 23960
rect 22196 23920 22205 23960
rect 22349 23920 22676 23960
rect 24355 23920 24364 23960
rect 24404 23920 24499 23960
rect 24539 23920 24548 23960
rect 14956 23876 14996 23920
rect 22349 23876 22389 23920
rect 22636 23876 22676 23920
rect 13996 23836 14188 23876
rect 14228 23836 14237 23876
rect 14947 23836 14956 23876
rect 14996 23836 15005 23876
rect 16003 23836 16012 23876
rect 16052 23836 16061 23876
rect 16675 23836 16684 23876
rect 16724 23836 18403 23876
rect 18443 23836 18452 23876
rect 20227 23836 20236 23876
rect 20276 23836 20285 23876
rect 21475 23836 21484 23876
rect 21524 23836 22389 23876
rect 22612 23836 22676 23876
rect 22732 23836 23212 23876
rect 23252 23836 23261 23876
rect 23491 23836 23500 23876
rect 23540 23836 23596 23876
rect 23636 23836 23671 23876
rect 23932 23836 23980 23876
rect 24020 23836 24029 23876
rect 24076 23836 24172 23876
rect 24212 23836 24221 23876
rect 13996 23792 14036 23836
rect 20236 23792 20276 23836
rect 22612 23792 22652 23836
rect 22732 23792 22772 23836
rect 23932 23792 23972 23836
rect 24076 23792 24116 23836
rect 4841 23752 4972 23792
rect 5012 23752 5021 23792
rect 5129 23752 5260 23792
rect 5300 23752 5309 23792
rect 5539 23752 5548 23792
rect 5588 23752 5740 23792
rect 5780 23752 5789 23792
rect 5897 23752 5932 23792
rect 5972 23752 6028 23792
rect 6068 23752 6077 23792
rect 6637 23752 6646 23792
rect 6686 23752 6836 23792
rect 6970 23752 6979 23792
rect 7019 23752 7028 23792
rect 7529 23752 7660 23792
rect 7700 23752 7709 23792
rect 8585 23752 8620 23792
rect 8660 23752 8716 23792
rect 8756 23752 8765 23792
rect 8852 23752 8859 23792
rect 8962 23752 8971 23792
rect 9011 23752 9020 23792
rect 9082 23752 9091 23792
rect 9131 23752 9140 23792
rect 9187 23752 9196 23792
rect 9236 23752 9292 23792
rect 9332 23752 9367 23792
rect 9411 23752 9484 23792
rect 9524 23752 9533 23792
rect 9641 23752 9676 23792
rect 9716 23752 9772 23792
rect 9812 23752 9821 23792
rect 9955 23752 9964 23792
rect 10004 23752 10013 23792
rect 10060 23752 10103 23792
rect 10143 23752 10152 23792
rect 10234 23752 10243 23792
rect 10283 23752 10292 23792
rect 10339 23752 10348 23792
rect 10388 23752 10397 23792
rect 10622 23752 10631 23792
rect 10671 23752 10680 23792
rect 10810 23752 10819 23792
rect 10859 23752 10868 23792
rect 10999 23752 11008 23792
rect 11048 23752 11060 23792
rect 11155 23752 11164 23792
rect 11204 23752 11308 23792
rect 11348 23752 11357 23792
rect 12163 23752 12172 23792
rect 12212 23752 12364 23792
rect 12404 23752 12413 23792
rect 12521 23752 12556 23792
rect 12596 23752 12652 23792
rect 12692 23752 12701 23792
rect 12748 23752 12767 23792
rect 12807 23752 12816 23792
rect 12876 23752 12940 23792
rect 12980 23752 13076 23792
rect 13123 23752 13132 23792
rect 13172 23752 13460 23792
rect 13507 23752 13516 23792
rect 13556 23752 13565 23792
rect 13987 23752 13996 23792
rect 14036 23752 14045 23792
rect 14266 23752 14275 23792
rect 14315 23752 15092 23792
rect 15322 23752 15331 23792
rect 15380 23752 15511 23792
rect 17251 23752 17260 23792
rect 17300 23752 17740 23792
rect 17780 23752 17789 23792
rect 18115 23752 18124 23792
rect 18164 23752 18173 23792
rect 18787 23752 18796 23792
rect 18836 23752 19027 23792
rect 19067 23752 19180 23792
rect 19220 23752 19229 23792
rect 19529 23752 19660 23792
rect 19700 23752 19709 23792
rect 19843 23752 19852 23792
rect 19892 23752 20035 23792
rect 20075 23752 20084 23792
rect 20131 23752 20140 23792
rect 20180 23752 20276 23792
rect 20515 23752 20524 23792
rect 20564 23752 20764 23792
rect 20804 23752 20813 23792
rect 20899 23752 20908 23792
rect 20948 23752 21044 23792
rect 21593 23752 21676 23792
rect 21716 23752 21724 23792
rect 21764 23752 21773 23792
rect 21859 23752 21868 23792
rect 21908 23752 21964 23792
rect 22004 23752 22039 23792
rect 22156 23752 22339 23792
rect 22379 23752 22388 23792
rect 22448 23752 22457 23792
rect 22497 23752 22508 23792
rect 22608 23752 22617 23792
rect 22657 23752 22666 23792
rect 22714 23752 22723 23792
rect 22763 23752 22772 23792
rect 22819 23752 22828 23792
rect 22897 23752 22999 23792
rect 23299 23752 23308 23792
rect 23348 23752 23416 23792
rect 23456 23752 23479 23792
rect 23596 23752 23692 23792
rect 23732 23752 23741 23792
rect 23802 23752 23811 23792
rect 23851 23752 23860 23792
rect 23923 23752 23932 23792
rect 23972 23752 23981 23792
rect 24058 23752 24067 23792
rect 24107 23752 24116 23792
rect 4972 23734 5012 23743
rect 6796 23708 6836 23752
rect 8812 23743 8852 23752
rect 634 23668 643 23708
rect 683 23668 1612 23708
rect 1652 23668 1996 23708
rect 2036 23668 2045 23708
rect 2938 23668 2947 23708
rect 2987 23668 3427 23708
rect 3467 23668 3476 23708
rect 4012 23668 4532 23708
rect 4684 23668 4876 23708
rect 4916 23668 4925 23708
rect 5923 23668 5932 23708
rect 5972 23668 6451 23708
rect 6491 23668 6500 23708
rect 6796 23668 7180 23708
rect 7220 23668 7229 23708
rect 7281 23668 7290 23708
rect 7330 23668 7852 23708
rect 7892 23668 7901 23708
rect 8035 23668 8044 23708
rect 8084 23668 8510 23708
rect 8550 23668 8559 23708
rect 4012 23624 4052 23668
rect 1228 23584 4052 23624
rect 4108 23584 4252 23624
rect 4292 23584 4301 23624
rect 1228 23456 1268 23584
rect 1132 23416 1268 23456
rect 1132 23204 1172 23416
rect 1411 23332 1420 23372
rect 1460 23332 2900 23372
rect 2860 23288 2900 23332
rect 4108 23288 4148 23584
rect 4492 23540 4532 23668
rect 6691 23584 6700 23624
rect 6740 23584 7075 23624
rect 7115 23584 7124 23624
rect 7171 23584 7180 23624
rect 7220 23584 7276 23624
rect 7316 23584 7351 23624
rect 8201 23584 8236 23624
rect 8276 23584 8332 23624
rect 8372 23584 8381 23624
rect 8602 23584 8611 23624
rect 8651 23584 8660 23624
rect 4492 23500 6124 23540
rect 6164 23500 6173 23540
rect 7084 23456 7124 23584
rect 8620 23540 8660 23584
rect 8976 23540 9016 23752
rect 9100 23708 9140 23752
rect 9100 23668 9196 23708
rect 9236 23668 9245 23708
rect 7555 23500 7564 23540
rect 7604 23500 8660 23540
rect 8803 23500 8812 23540
rect 8852 23500 9016 23540
rect 9411 23456 9451 23752
rect 9964 23708 10004 23752
rect 9964 23668 10060 23708
rect 10100 23668 10164 23708
rect 9946 23584 9955 23624
rect 9995 23584 10004 23624
rect 4343 23416 4352 23456
rect 4720 23416 4729 23456
rect 7084 23416 9484 23456
rect 9524 23416 9611 23456
rect 4780 23332 5740 23372
rect 5780 23332 5789 23372
rect 4780 23288 4820 23332
rect 9964 23288 10004 23584
rect 10252 23456 10292 23752
rect 10347 23540 10387 23752
rect 10636 23708 10676 23752
rect 11020 23708 11060 23752
rect 13420 23708 13460 23752
rect 15052 23708 15092 23752
rect 10627 23668 10636 23708
rect 10676 23668 10718 23708
rect 11011 23668 11020 23708
rect 11060 23668 13324 23708
rect 13364 23668 13373 23708
rect 13420 23668 14036 23708
rect 14371 23668 14380 23708
rect 14420 23668 14668 23708
rect 14708 23668 14717 23708
rect 15052 23668 17443 23708
rect 17483 23668 17492 23708
rect 13996 23624 14036 23668
rect 18124 23624 18164 23752
rect 19219 23668 19228 23708
rect 19268 23668 20908 23708
rect 20948 23668 20957 23708
rect 21004 23624 21044 23752
rect 22156 23708 22196 23752
rect 22468 23708 22508 23752
rect 22147 23668 22156 23708
rect 22196 23668 22205 23708
rect 22423 23668 22444 23708
rect 22484 23668 22508 23708
rect 23203 23668 23212 23708
rect 23291 23668 23383 23708
rect 23596 23624 23636 23752
rect 23811 23708 23851 23752
rect 24599 23708 24639 24088
rect 25411 24004 25420 24044
rect 25460 24004 25468 24044
rect 25508 24004 25591 24044
rect 27331 24004 27340 24044
rect 27380 24004 28108 24044
rect 28148 24004 28157 24044
rect 25315 23920 25324 23960
rect 25364 23920 25373 23960
rect 25507 23920 25516 23960
rect 25556 23920 27244 23960
rect 27284 23920 29108 23960
rect 25324 23876 25364 23920
rect 24739 23836 24748 23876
rect 24788 23836 24797 23876
rect 24940 23836 25228 23876
rect 25268 23836 25277 23876
rect 25324 23836 25652 23876
rect 24699 23752 24708 23792
rect 24748 23752 24788 23836
rect 24940 23792 24980 23836
rect 25612 23792 25652 23836
rect 25996 23836 26764 23876
rect 26804 23836 26813 23876
rect 25996 23792 26036 23836
rect 27628 23792 27668 23920
rect 28841 23836 28972 23876
rect 29012 23836 29021 23876
rect 29068 23792 29108 23920
rect 30211 23836 30220 23876
rect 30260 23836 30269 23876
rect 24835 23752 24844 23792
rect 24884 23752 24980 23792
rect 25070 23752 25079 23792
rect 25119 23752 25128 23792
rect 25210 23783 25268 23792
rect 23811 23668 23980 23708
rect 24020 23668 24029 23708
rect 24369 23668 24378 23708
rect 24418 23668 24639 23708
rect 25079 23708 25119 23752
rect 25210 23743 25219 23783
rect 25259 23743 25268 23783
rect 25315 23752 25324 23792
rect 25364 23752 25495 23792
rect 25603 23752 25612 23792
rect 25652 23752 25661 23792
rect 25838 23752 25847 23792
rect 25887 23752 25896 23792
rect 25978 23783 26036 23792
rect 25210 23742 25268 23743
rect 25228 23708 25268 23742
rect 25847 23708 25887 23752
rect 25978 23743 25987 23783
rect 26027 23743 26036 23783
rect 26083 23752 26092 23792
rect 26132 23752 26141 23792
rect 26345 23752 26467 23792
rect 26516 23752 26525 23792
rect 26644 23752 26668 23792
rect 26708 23752 26775 23792
rect 26815 23752 26824 23792
rect 26938 23752 26947 23792
rect 26987 23752 26996 23792
rect 27043 23752 27052 23792
rect 27092 23787 27188 23792
rect 27235 23787 27244 23792
rect 27092 23752 27244 23787
rect 27284 23752 27293 23792
rect 27619 23752 27628 23792
rect 27668 23752 27677 23792
rect 27763 23752 27772 23792
rect 27812 23752 28204 23792
rect 28244 23752 28253 23792
rect 28771 23752 28780 23792
rect 28820 23752 28876 23792
rect 28916 23752 28951 23792
rect 29059 23752 29068 23792
rect 29108 23752 29117 23792
rect 29251 23752 29260 23792
rect 29300 23752 29347 23792
rect 29387 23752 29431 23792
rect 25978 23742 26036 23743
rect 25079 23668 25171 23708
rect 25228 23668 25420 23708
rect 25460 23668 25887 23708
rect 26092 23708 26132 23752
rect 26956 23708 26996 23752
rect 27148 23747 27284 23752
rect 27772 23708 27812 23752
rect 26092 23668 27010 23708
rect 27305 23668 27340 23708
rect 27380 23668 27427 23708
rect 27467 23668 27485 23708
rect 27619 23668 27628 23708
rect 27668 23668 27812 23708
rect 28204 23708 28244 23752
rect 28204 23668 29548 23708
rect 29588 23668 29597 23708
rect 25131 23624 25171 23668
rect 26970 23624 27010 23668
rect 11561 23584 11596 23624
rect 11636 23584 11692 23624
rect 11732 23584 11741 23624
rect 13603 23584 13612 23624
rect 13652 23584 13708 23624
rect 13748 23584 13783 23624
rect 13996 23584 17260 23624
rect 17300 23584 17644 23624
rect 17684 23584 18164 23624
rect 18211 23584 18220 23624
rect 18260 23584 19948 23624
rect 19988 23584 19997 23624
rect 20297 23584 20428 23624
rect 20468 23584 20477 23624
rect 20602 23584 20611 23624
rect 20660 23584 20791 23624
rect 21004 23584 21571 23624
rect 21611 23584 21620 23624
rect 22810 23584 22819 23624
rect 22859 23584 22868 23624
rect 22915 23584 22924 23624
rect 22964 23584 23500 23624
rect 23540 23584 23636 23624
rect 24154 23584 24163 23624
rect 24203 23584 24364 23624
rect 24404 23584 24413 23624
rect 25027 23584 25036 23624
rect 25076 23584 25085 23624
rect 25131 23584 25516 23624
rect 25556 23584 25565 23624
rect 25673 23584 25804 23624
rect 25844 23584 25853 23624
rect 26275 23584 26284 23624
rect 26324 23584 26563 23624
rect 26603 23584 26612 23624
rect 26659 23584 26668 23624
rect 26708 23584 26839 23624
rect 26970 23584 27436 23624
rect 27476 23584 27485 23624
rect 27593 23584 27724 23624
rect 27764 23584 29932 23624
rect 29972 23584 29981 23624
rect 31171 23584 31180 23624
rect 31220 23584 31276 23624
rect 31316 23584 31351 23624
rect 22828 23540 22868 23584
rect 10347 23500 11692 23540
rect 11732 23500 11741 23540
rect 12835 23500 12844 23540
rect 12884 23500 20756 23540
rect 22828 23500 24460 23540
rect 24500 23500 24509 23540
rect 20716 23456 20756 23500
rect 10252 23416 10444 23456
rect 10484 23416 11500 23456
rect 11540 23416 11549 23456
rect 12117 23416 12126 23456
rect 12494 23416 12503 23456
rect 15052 23416 19468 23456
rect 19508 23416 19517 23456
rect 19891 23416 19900 23456
rect 20268 23416 20277 23456
rect 20428 23416 20674 23456
rect 20716 23416 24748 23456
rect 24788 23416 24797 23456
rect 10627 23332 10636 23372
rect 10676 23332 13460 23372
rect 1690 23248 1699 23288
rect 1739 23248 2324 23288
rect 2371 23248 2380 23288
rect 2420 23248 2804 23288
rect 2860 23248 3571 23288
rect 3611 23248 3620 23288
rect 3811 23248 3820 23288
rect 3860 23248 4003 23288
rect 4043 23248 4052 23288
rect 4099 23248 4108 23288
rect 4148 23248 4157 23288
rect 4483 23248 4492 23288
rect 4532 23248 4780 23288
rect 4820 23248 4829 23288
rect 5059 23248 5068 23288
rect 5108 23248 5323 23288
rect 5539 23248 5548 23288
rect 5588 23248 5635 23288
rect 5675 23248 5719 23288
rect 7459 23248 7468 23288
rect 7508 23248 8140 23288
rect 8180 23248 8189 23288
rect 9964 23248 10388 23288
rect 2284 23204 2324 23248
rect 844 23164 940 23204
rect 980 23164 989 23204
rect 1036 23164 1172 23204
rect 2170 23164 2179 23204
rect 2219 23164 2228 23204
rect 2275 23164 2284 23204
rect 2324 23164 2668 23204
rect 2708 23164 2717 23204
rect 844 23120 884 23164
rect 1036 23120 1076 23164
rect 2188 23120 2228 23164
rect 2764 23120 2804 23248
rect 5283 23204 5323 23248
rect 3113 23164 3244 23204
rect 3284 23164 3293 23204
rect 3724 23164 4675 23204
rect 4715 23164 4724 23204
rect 4924 23164 5068 23204
rect 5108 23164 5117 23204
rect 5283 23164 5534 23204
rect 5574 23164 5583 23204
rect 5635 23164 5644 23204
rect 5684 23164 6115 23204
rect 6155 23164 6164 23204
rect 7084 23164 7564 23204
rect 7604 23164 7613 23204
rect 8995 23164 9004 23204
rect 9044 23164 9676 23204
rect 9716 23164 9725 23204
rect 9772 23164 10252 23204
rect 10292 23164 10301 23204
rect 835 23080 844 23120
rect 884 23080 893 23120
rect 1018 23080 1027 23120
rect 1067 23080 1076 23120
rect 1219 23080 1228 23120
rect 1268 23080 1277 23120
rect 1402 23080 1411 23120
rect 1451 23080 1460 23120
rect 1594 23080 1603 23120
rect 1652 23080 1783 23120
rect 1905 23080 1914 23120
rect 1954 23080 2081 23120
rect 2132 23080 2141 23120
rect 2188 23080 2284 23120
rect 2324 23080 2333 23120
rect 2380 23111 2420 23120
rect 905 22912 1027 22952
rect 1076 22912 1085 22952
rect 1228 22784 1268 23080
rect 1420 23036 1460 23080
rect 2563 23080 2572 23120
rect 2612 23080 2804 23120
rect 3724 23120 3764 23164
rect 4924 23120 4964 23164
rect 7084 23120 7124 23164
rect 9772 23120 9812 23164
rect 10348 23120 10388 23248
rect 10594 23248 10987 23288
rect 11107 23248 11116 23288
rect 11156 23248 11491 23288
rect 11531 23248 11540 23288
rect 11779 23248 11788 23288
rect 11828 23248 12596 23288
rect 12883 23248 12892 23288
rect 12932 23248 13132 23288
rect 13172 23248 13181 23288
rect 10594 23120 10634 23248
rect 10947 23204 10987 23248
rect 10723 23164 10732 23204
rect 10772 23164 10903 23204
rect 10947 23164 11085 23204
rect 11045 23123 11085 23164
rect 11308 23164 11404 23204
rect 11444 23164 11453 23204
rect 11875 23164 11884 23204
rect 11924 23164 12404 23204
rect 11045 23120 11199 23123
rect 11308 23120 11348 23164
rect 12364 23120 12404 23164
rect 12556 23120 12596 23248
rect 13420 23120 13460 23332
rect 15052 23288 15092 23416
rect 20428 23372 20468 23416
rect 20634 23372 20674 23416
rect 25036 23372 25076 23584
rect 27665 23416 27674 23456
rect 28042 23416 28051 23456
rect 14371 23248 14380 23288
rect 14420 23248 14900 23288
rect 15034 23248 15043 23288
rect 15083 23248 15092 23288
rect 15148 23332 15244 23372
rect 15284 23332 15293 23372
rect 15715 23332 15724 23372
rect 15764 23332 20468 23372
rect 20515 23332 20524 23372
rect 20564 23332 20573 23372
rect 20634 23332 23308 23372
rect 23348 23332 23357 23372
rect 24355 23332 24364 23372
rect 24404 23332 25076 23372
rect 29923 23332 29932 23372
rect 29972 23332 31180 23372
rect 31220 23332 31229 23372
rect 13507 23164 13516 23204
rect 13556 23164 13652 23204
rect 13795 23164 13804 23204
rect 13844 23164 13891 23204
rect 13987 23164 13996 23204
rect 14036 23164 14083 23204
rect 14530 23164 14668 23204
rect 14708 23164 14717 23204
rect 13612 23120 13652 23164
rect 13804 23120 13844 23164
rect 13996 23120 14036 23164
rect 14530 23120 14570 23164
rect 3724 23080 3736 23120
rect 3776 23080 3785 23120
rect 3896 23080 3905 23120
rect 3945 23080 4108 23120
rect 4148 23080 4157 23120
rect 4204 23111 4291 23120
rect 2380 23060 2420 23071
rect 4244 23080 4291 23111
rect 4387 23080 4396 23120
rect 4436 23080 4574 23120
rect 4614 23080 4628 23120
rect 2380 23036 2496 23060
rect 4204 23036 4244 23071
rect 1420 22996 1900 23036
rect 1940 22996 1949 23036
rect 2179 22996 2188 23036
rect 2228 23020 2496 23036
rect 2228 22996 2420 23020
rect 4195 22996 4204 23036
rect 4244 22996 4253 23036
rect 4588 22952 4628 23080
rect 4876 23111 4964 23120
rect 4916 23080 4964 23111
rect 5033 23080 5164 23120
rect 5204 23080 5213 23120
rect 5321 23080 5401 23120
rect 5441 23080 5452 23120
rect 5492 23080 5501 23120
rect 5609 23080 5740 23120
rect 5780 23080 5789 23120
rect 5836 23111 5876 23120
rect 4876 23062 4916 23071
rect 7075 23080 7084 23120
rect 7124 23080 7133 23120
rect 7337 23080 7468 23120
rect 7508 23080 7517 23120
rect 8227 23080 8236 23120
rect 8276 23080 8332 23120
rect 8372 23080 8407 23120
rect 8506 23080 8515 23120
rect 8555 23080 8908 23120
rect 8948 23080 8957 23120
rect 9763 23080 9772 23120
rect 9812 23080 9821 23120
rect 10339 23080 10348 23120
rect 10388 23080 10397 23120
rect 10576 23080 10585 23120
rect 10625 23080 10634 23120
rect 10819 23080 10828 23120
rect 10868 23080 10915 23120
rect 11010 23080 11045 23120
rect 11085 23083 11164 23120
rect 11085 23080 11094 23083
rect 11155 23080 11164 23083
rect 11204 23080 11213 23120
rect 11290 23080 11299 23120
rect 11339 23080 11348 23120
rect 11395 23080 11404 23120
rect 11444 23080 11540 23120
rect 11875 23080 11884 23120
rect 11924 23080 11933 23120
rect 12112 23080 12121 23120
rect 12161 23080 12308 23120
rect 12355 23080 12364 23120
rect 12404 23080 12413 23120
rect 12547 23080 12556 23120
rect 12596 23080 12605 23120
rect 12713 23080 12748 23120
rect 12788 23080 12844 23120
rect 12884 23080 12893 23120
rect 13411 23080 13420 23120
rect 13460 23080 13469 23120
rect 13603 23080 13612 23120
rect 13652 23080 13661 23120
rect 13795 23080 13804 23120
rect 13844 23080 13853 23120
rect 13978 23080 13987 23120
rect 14027 23080 14036 23120
rect 14153 23080 14188 23120
rect 14228 23080 14284 23120
rect 14324 23080 14333 23120
rect 14512 23080 14521 23120
rect 14561 23080 14570 23120
rect 14860 23115 14900 23248
rect 15148 23120 15188 23332
rect 20524 23288 20564 23332
rect 23308 23288 23348 23332
rect 15244 23248 17836 23288
rect 17876 23248 17885 23288
rect 18089 23248 18211 23288
rect 18260 23248 18269 23288
rect 18377 23248 18508 23288
rect 18548 23248 18557 23288
rect 19049 23248 19180 23288
rect 19220 23248 19229 23288
rect 20227 23248 20236 23288
rect 20276 23248 20419 23288
rect 20459 23248 20468 23288
rect 20515 23248 20524 23288
rect 20564 23248 20611 23288
rect 20716 23248 21292 23288
rect 21332 23248 21341 23288
rect 21610 23248 21619 23288
rect 21659 23248 21772 23288
rect 21812 23248 21821 23288
rect 23308 23248 28103 23288
rect 28483 23248 28492 23288
rect 28532 23248 28916 23288
rect 15244 23120 15284 23248
rect 20716 23204 20756 23248
rect 15331 23164 15340 23204
rect 15380 23164 16204 23204
rect 16244 23164 16253 23204
rect 16553 23164 16675 23204
rect 16724 23164 16733 23204
rect 17251 23164 17260 23204
rect 17300 23164 17932 23204
rect 17972 23164 17981 23204
rect 18316 23164 19412 23204
rect 19651 23164 19660 23204
rect 19700 23164 19987 23204
rect 20027 23164 20036 23204
rect 20140 23164 20428 23204
rect 20468 23164 20477 23204
rect 20625 23164 20634 23204
rect 20674 23164 20756 23204
rect 20947 23164 20956 23204
rect 20996 23164 22156 23204
rect 22196 23164 22205 23204
rect 22339 23164 22348 23204
rect 22388 23164 23212 23204
rect 23252 23164 23261 23204
rect 25027 23164 25036 23204
rect 25076 23164 25132 23204
rect 25172 23164 25207 23204
rect 25756 23195 25844 23204
rect 18316 23120 18356 23164
rect 19372 23120 19412 23164
rect 20140 23120 20180 23164
rect 22540 23120 22580 23164
rect 25756 23155 25795 23195
rect 25835 23155 25844 23195
rect 26179 23164 26188 23204
rect 26228 23164 26708 23204
rect 26825 23164 26956 23204
rect 26996 23164 27005 23204
rect 27139 23164 27148 23204
rect 27188 23164 27260 23204
rect 25756 23154 25844 23155
rect 5836 23036 5876 23071
rect 5059 22996 5068 23036
rect 5108 22996 5117 23036
rect 5251 22996 5260 23036
rect 5323 22996 5431 23036
rect 5827 22996 5836 23036
rect 5876 22996 5923 23036
rect 10121 22996 10252 23036
rect 10292 22996 10301 23036
rect 5068 22952 5108 22996
rect 1402 22912 1411 22952
rect 1451 22912 3436 22952
rect 3476 22912 3485 22952
rect 4588 22912 5108 22952
rect 8393 22912 8515 22952
rect 8564 22912 8573 22952
rect 8803 22912 8812 22952
rect 8852 22912 8995 22952
rect 9035 22912 9044 22952
rect 10348 22868 10388 23080
rect 10828 23036 10868 23080
rect 11164 23036 11204 23080
rect 10458 22996 10467 23036
rect 10507 22996 10540 23036
rect 10580 22996 10638 23036
rect 10819 22996 10828 23036
rect 10868 22996 10877 23036
rect 10938 22996 10947 23036
rect 10987 22996 10996 23036
rect 11164 22996 11308 23036
rect 11348 22996 11357 23036
rect 10947 22952 10987 22996
rect 10627 22912 10636 22952
rect 10676 22912 10987 22952
rect 11500 22868 11540 23080
rect 11657 22996 11788 23036
rect 11828 22996 11837 23036
rect 1699 22828 1708 22868
rect 1748 22828 1900 22868
rect 1940 22828 1949 22868
rect 2947 22828 2956 22868
rect 2996 22828 7948 22868
rect 7988 22828 7997 22868
rect 8131 22828 8140 22868
rect 8180 22828 8716 22868
rect 8756 22828 8765 22868
rect 8899 22828 8908 22868
rect 8948 22828 10060 22868
rect 10100 22828 10109 22868
rect 10348 22828 10828 22868
rect 10868 22828 11540 22868
rect 11884 22784 11924 23080
rect 12268 23036 12308 23080
rect 12748 23036 12788 23080
rect 14729 23075 14860 23115
rect 14900 23075 14909 23115
rect 15046 23080 15055 23120
rect 15095 23080 15188 23120
rect 15235 23080 15244 23120
rect 15284 23080 15293 23120
rect 15360 23080 15436 23120
rect 15476 23080 15485 23120
rect 17321 23080 17452 23120
rect 17492 23080 17501 23120
rect 17705 23080 17740 23120
rect 17780 23080 17836 23120
rect 17876 23080 17885 23120
rect 18019 23080 18028 23120
rect 18068 23080 18199 23120
rect 18307 23080 18316 23120
rect 18356 23080 18365 23120
rect 19171 23080 19180 23120
rect 19220 23080 19229 23120
rect 19363 23080 19372 23120
rect 19412 23080 19564 23120
rect 19604 23080 19613 23120
rect 19747 23080 19756 23120
rect 19796 23080 19988 23120
rect 20140 23080 20152 23120
rect 20192 23080 20201 23120
rect 20269 23080 20323 23120
rect 20363 23080 20385 23120
rect 20803 23080 20812 23120
rect 20852 23080 21140 23120
rect 21245 23080 21292 23120
rect 21332 23111 21416 23120
rect 21332 23080 21376 23111
rect 12010 23027 12076 23036
rect 12010 22987 12019 23027
rect 12059 22996 12076 23027
rect 12116 22996 12199 23036
rect 12259 22996 12268 23036
rect 12308 22996 12788 23036
rect 13219 22996 13228 23036
rect 13268 22996 13612 23036
rect 13652 22996 13661 23036
rect 14179 22996 14188 23036
rect 14228 22996 14237 23036
rect 14371 22996 14380 23036
rect 14443 22996 14551 23036
rect 12059 22987 12068 22996
rect 12010 22986 12068 22987
rect 13865 22912 13987 22952
rect 14036 22912 14045 22952
rect 14188 22868 14228 22996
rect 14860 22952 14900 23075
rect 15436 23036 15476 23080
rect 19180 23036 19220 23080
rect 15427 22996 15436 23036
rect 15476 22996 15485 23036
rect 15724 22996 15956 23036
rect 18211 22996 18220 23036
rect 18260 22996 19220 23036
rect 19948 23036 19988 23080
rect 20269 23036 20309 23080
rect 19948 22996 20309 23036
rect 15724 22952 15764 22996
rect 14860 22912 15764 22952
rect 15811 22912 15820 22952
rect 15860 22912 15869 22952
rect 12329 22828 12364 22868
rect 12404 22828 12460 22868
rect 12500 22828 12509 22868
rect 12979 22828 12988 22868
rect 13028 22828 13036 22868
rect 13076 22828 13159 22868
rect 13289 22828 13324 22868
rect 13364 22828 13420 22868
rect 13460 22828 13469 22868
rect 14083 22828 14092 22868
rect 14132 22828 14228 22868
rect 15820 22784 15860 22912
rect 15916 22868 15956 22996
rect 21100 22952 21140 23080
rect 21466 23080 21475 23120
rect 21524 23080 21655 23120
rect 21763 23080 21772 23120
rect 21812 23080 21821 23120
rect 21955 23080 21964 23120
rect 22004 23080 22060 23120
rect 22100 23080 22135 23120
rect 22522 23080 22531 23120
rect 22571 23080 22580 23120
rect 24826 23080 24835 23120
rect 24875 23080 25132 23120
rect 25172 23080 25181 23120
rect 25315 23080 25324 23120
rect 25364 23080 25507 23120
rect 25556 23080 25565 23120
rect 25612 23111 25652 23120
rect 21376 23062 21416 23071
rect 21772 23036 21812 23080
rect 21763 22996 21772 23036
rect 21812 22996 21859 23036
rect 22025 22996 22156 23036
rect 22196 22996 22205 23036
rect 16003 22912 16012 22952
rect 16052 22912 16183 22952
rect 18307 22912 18316 22952
rect 18356 22912 18700 22952
rect 18740 22912 18749 22952
rect 19267 22912 19276 22952
rect 19316 22912 20908 22952
rect 20948 22912 20957 22952
rect 21100 22912 21772 22952
rect 21812 22912 21821 22952
rect 15916 22828 18220 22868
rect 18260 22828 18269 22868
rect 20707 22828 20716 22868
rect 20756 22828 21091 22868
rect 21131 22828 21140 22868
rect 1228 22744 2572 22784
rect 2612 22744 2621 22784
rect 7747 22744 7756 22784
rect 7796 22744 10444 22784
rect 10484 22744 10493 22784
rect 10780 22744 11788 22784
rect 11828 22744 11924 22784
rect 12163 22744 12172 22784
rect 12212 22744 14612 22784
rect 15820 22744 22540 22784
rect 22580 22744 22589 22784
rect 10780 22700 10820 22744
rect 1027 22660 1036 22700
rect 1076 22660 2764 22700
rect 2804 22660 2813 22700
rect 3103 22660 3112 22700
rect 3480 22660 3489 22700
rect 7843 22660 7852 22700
rect 7892 22660 10820 22700
rect 10877 22660 10886 22700
rect 11254 22660 11263 22700
rect 8419 22576 8428 22616
rect 8468 22576 13246 22616
rect 451 22492 460 22532
rect 500 22492 5396 22532
rect 5993 22492 6019 22532
rect 6059 22492 6124 22532
rect 6164 22492 6173 22532
rect 6307 22492 6316 22532
rect 6356 22492 6365 22532
rect 7171 22492 7180 22532
rect 7220 22492 7267 22532
rect 7307 22492 7351 22532
rect 7468 22492 7948 22532
rect 7988 22492 7997 22532
rect 8332 22492 8524 22532
rect 8564 22492 8573 22532
rect 9667 22492 9676 22532
rect 9716 22492 10388 22532
rect 10505 22492 10636 22532
rect 10676 22492 10685 22532
rect 11273 22492 11308 22532
rect 11348 22492 11404 22532
rect 11444 22492 11453 22532
rect 11561 22492 11692 22532
rect 11732 22492 11741 22532
rect 5356 22448 5396 22492
rect 2083 22408 2092 22448
rect 2132 22408 4148 22448
rect 0 22364 400 22384
rect 4108 22364 4148 22408
rect 4204 22408 4300 22448
rect 4340 22408 4349 22448
rect 4684 22408 4780 22448
rect 4820 22408 4829 22448
rect 5356 22408 5452 22448
rect 5492 22408 5501 22448
rect 0 22324 556 22364
rect 596 22324 605 22364
rect 1219 22324 1228 22364
rect 1268 22324 1940 22364
rect 2179 22324 2188 22364
rect 2228 22324 2380 22364
rect 2420 22324 2429 22364
rect 2602 22355 3532 22364
rect 0 22304 400 22324
rect 1900 22280 1940 22324
rect 2602 22315 2611 22355
rect 2651 22324 3532 22355
rect 3572 22324 3581 22364
rect 3754 22324 3763 22364
rect 3803 22324 3916 22364
rect 3956 22324 3965 22364
rect 4099 22324 4108 22364
rect 4148 22324 4157 22364
rect 2651 22315 2660 22324
rect 2602 22314 2660 22315
rect 4204 22280 4244 22408
rect 4330 22355 4396 22364
rect 4330 22315 4339 22355
rect 4379 22324 4396 22355
rect 4436 22324 4519 22364
rect 4379 22315 4388 22324
rect 4330 22314 4388 22315
rect 4684 22280 4724 22408
rect 4780 22324 5068 22364
rect 5108 22324 5117 22364
rect 5347 22324 5356 22364
rect 5396 22324 5548 22364
rect 5588 22324 5597 22364
rect 5827 22324 5836 22364
rect 5876 22324 6007 22364
rect 4780 22280 4820 22324
rect 6316 22313 6356 22492
rect 6665 22324 6796 22364
rect 6836 22324 6845 22364
rect 1577 22240 1708 22280
rect 1748 22240 1757 22280
rect 1882 22240 1891 22280
rect 1931 22240 1940 22280
rect 2083 22240 2092 22280
rect 2132 22240 2199 22280
rect 2239 22240 2263 22280
rect 2467 22240 2476 22280
rect 2516 22240 2525 22280
rect 2704 22240 2713 22280
rect 2753 22240 2762 22280
rect 3291 22240 3300 22280
rect 259 22156 268 22196
rect 308 22156 739 22196
rect 779 22156 788 22196
rect 1411 22156 1420 22196
rect 1460 22156 2092 22196
rect 2132 22156 2141 22196
rect 1315 22072 1324 22112
rect 1364 22072 1987 22112
rect 2027 22072 2284 22112
rect 2324 22072 2333 22112
rect 2476 22028 2516 22240
rect 2722 22196 2762 22240
rect 3340 22196 3380 22280
rect 3427 22240 3436 22280
rect 3476 22240 3607 22280
rect 3715 22240 3724 22280
rect 3764 22240 3928 22280
rect 3968 22240 3977 22280
rect 4195 22240 4204 22280
rect 4244 22240 4253 22280
rect 4432 22240 4441 22280
rect 4481 22240 4724 22280
rect 4771 22240 4780 22280
rect 4820 22240 4829 22280
rect 4963 22240 4972 22280
rect 5012 22240 5143 22280
rect 5364 22240 5452 22280
rect 5492 22240 5495 22280
rect 5535 22240 5544 22280
rect 5626 22240 5635 22280
rect 5675 22240 5684 22280
rect 5731 22240 5740 22280
rect 5780 22240 5911 22280
rect 6305 22273 6314 22313
rect 6354 22273 6363 22313
rect 6451 22282 6460 22322
rect 6500 22282 6509 22322
rect 4450 22196 4490 22240
rect 2659 22156 2668 22196
rect 2708 22156 2762 22196
rect 3331 22156 3340 22196
rect 3380 22156 3389 22196
rect 4195 22156 4204 22196
rect 4244 22156 4490 22196
rect 4745 22156 4876 22196
rect 4916 22156 4925 22196
rect 3017 22072 3139 22112
rect 3188 22072 3197 22112
rect 4876 22072 5116 22112
rect 5156 22072 5165 22112
rect 4876 22028 4916 22072
rect 451 21988 460 22028
rect 500 21988 1036 22028
rect 1076 21988 1085 22028
rect 1603 21988 1612 22028
rect 1652 21988 2516 22028
rect 2860 21988 4916 22028
rect 0 21944 400 21964
rect 2860 21944 2900 21988
rect 5644 21944 5684 22240
rect 6460 22196 6500 22282
rect 7468 22280 7508 22492
rect 7843 22408 7852 22448
rect 7892 22408 7901 22448
rect 7852 22364 7892 22408
rect 8332 22364 8372 22492
rect 8419 22408 8428 22448
rect 8468 22408 8995 22448
rect 9035 22408 9044 22448
rect 9676 22408 10252 22448
rect 10292 22408 10301 22448
rect 7555 22324 7564 22364
rect 7604 22324 7651 22364
rect 7834 22324 7843 22364
rect 7883 22324 7939 22364
rect 8044 22324 8372 22364
rect 6586 22240 6595 22280
rect 6635 22240 6644 22280
rect 6691 22240 6700 22280
rect 6740 22240 6822 22280
rect 7256 22240 7265 22280
rect 7305 22240 7508 22280
rect 7564 22280 7604 22324
rect 8044 22280 8084 22324
rect 8524 22280 8564 22289
rect 9676 22280 9716 22408
rect 10348 22364 10388 22492
rect 13206 22448 13246 22576
rect 14572 22532 14612 22744
rect 22636 22700 22676 23016
rect 24521 22996 24652 23036
rect 24692 22996 24701 23036
rect 24844 22952 24884 23080
rect 25612 23036 25652 23071
rect 25219 22996 25228 23036
rect 25268 22996 25277 23036
rect 25516 22996 25652 23036
rect 24451 22912 24460 22952
rect 24500 22912 24884 22952
rect 25228 22868 25268 22996
rect 25516 22952 25556 22996
rect 25756 22952 25796 23154
rect 26668 23120 26708 23164
rect 27220 23120 27260 23164
rect 28063 23120 28103 23248
rect 28204 23164 28588 23204
rect 28628 23164 28637 23204
rect 28204 23120 28244 23164
rect 25882 23080 25891 23120
rect 25931 23080 25940 23120
rect 26059 23080 26068 23120
rect 26132 23080 26248 23120
rect 26371 23080 26380 23120
rect 26420 23080 26467 23120
rect 26507 23080 26551 23120
rect 26650 23080 26659 23120
rect 26699 23080 26708 23120
rect 26755 23080 26764 23120
rect 26804 23080 26813 23120
rect 25900 23036 25940 23080
rect 26764 23036 26804 23080
rect 25900 22996 26804 23036
rect 27052 23065 27069 23105
rect 27109 23065 27118 23105
rect 27202 23080 27211 23120
rect 27251 23080 27260 23120
rect 27427 23080 27436 23120
rect 27476 23080 27607 23120
rect 28044 23080 28053 23120
rect 28093 23080 28103 23120
rect 28195 23080 28204 23120
rect 28244 23080 28253 23120
rect 27052 22952 27092 23065
rect 28063 23036 28103 23080
rect 28337 23048 28346 23088
rect 28386 23048 28395 23088
rect 27209 22996 27244 23036
rect 27284 22996 27331 23036
rect 27371 22996 27389 23036
rect 27523 22996 27532 23036
rect 27572 22996 27628 23036
rect 27668 22996 27703 23036
rect 27811 22996 27820 23036
rect 27899 22996 27991 23036
rect 28063 22996 28204 23036
rect 28244 22996 28253 23036
rect 28355 22952 28395 23048
rect 28876 23036 28916 23248
rect 29155 23080 29164 23120
rect 29204 23080 29356 23120
rect 29396 23080 29405 23120
rect 29539 23080 29548 23120
rect 29588 23080 29719 23120
rect 30281 23080 30316 23120
rect 30356 23080 30403 23120
rect 30443 23080 30461 23120
rect 30953 23080 31084 23120
rect 31124 23080 31133 23120
rect 25507 22912 25516 22952
rect 25556 22912 25652 22952
rect 25756 22912 26284 22952
rect 26324 22912 26333 22952
rect 27052 22912 27148 22952
rect 27188 22912 27197 22952
rect 27820 22912 28395 22952
rect 28780 22996 28916 23036
rect 25612 22868 25652 22912
rect 27820 22868 27860 22912
rect 25228 22828 25507 22868
rect 25547 22828 25556 22868
rect 25612 22828 27860 22868
rect 27907 22828 27916 22868
rect 27956 22828 28684 22868
rect 28724 22828 28733 22868
rect 28780 22784 28820 22996
rect 30211 22828 30220 22868
rect 30260 22828 31276 22868
rect 31316 22828 31325 22868
rect 27619 22744 27628 22784
rect 27668 22744 28820 22784
rect 18651 22660 18660 22700
rect 19028 22660 19037 22700
rect 19267 22660 19276 22700
rect 19316 22660 22676 22700
rect 26425 22660 26434 22700
rect 26802 22660 26811 22700
rect 14755 22576 14764 22616
rect 14804 22576 16876 22616
rect 16916 22576 16925 22616
rect 20332 22576 22060 22616
rect 22100 22576 22109 22616
rect 23011 22576 23020 22616
rect 23060 22576 23828 22616
rect 26851 22576 26860 22616
rect 26900 22576 30124 22616
rect 30164 22576 30173 22616
rect 20332 22532 20372 22576
rect 14554 22492 14563 22532
rect 14603 22492 14612 22532
rect 17443 22492 17452 22532
rect 17492 22492 19316 22532
rect 20314 22492 20323 22532
rect 20363 22492 20372 22532
rect 21178 22492 21187 22532
rect 21227 22492 21772 22532
rect 21812 22492 21821 22532
rect 21946 22492 21955 22532
rect 21995 22492 22156 22532
rect 22196 22492 22205 22532
rect 22252 22492 23692 22532
rect 23732 22492 23741 22532
rect 19276 22448 19316 22492
rect 22252 22448 22292 22492
rect 23788 22448 23828 22576
rect 23962 22492 23971 22532
rect 24011 22492 24268 22532
rect 24308 22492 24317 22532
rect 25699 22492 25708 22532
rect 25748 22492 25900 22532
rect 25940 22492 25949 22532
rect 26275 22492 26284 22532
rect 26324 22492 27148 22532
rect 27188 22492 27197 22532
rect 27593 22492 27724 22532
rect 27764 22492 27773 22532
rect 10435 22408 10444 22448
rect 10484 22408 11156 22448
rect 10348 22324 10964 22364
rect 10924 22280 10964 22324
rect 11116 22280 11156 22408
rect 7651 22240 7660 22280
rect 7700 22240 7703 22280
rect 7743 22240 7831 22280
rect 7939 22240 7948 22280
rect 7988 22240 8084 22280
rect 8393 22240 8524 22280
rect 8564 22240 8573 22280
rect 9658 22240 9667 22280
rect 9707 22240 9716 22280
rect 9833 22240 9964 22280
rect 10004 22240 10013 22280
rect 10109 22240 10154 22280
rect 10194 22240 10203 22280
rect 10437 22240 10446 22280
rect 10486 22240 10495 22280
rect 10627 22240 10636 22280
rect 10676 22240 10828 22280
rect 10868 22240 10877 22280
rect 10924 22240 10989 22280
rect 11029 22240 11038 22280
rect 11098 22240 11107 22280
rect 11147 22240 11156 22280
rect 11212 22408 12268 22448
rect 12308 22408 12317 22448
rect 13206 22408 16483 22448
rect 16523 22408 16532 22448
rect 17731 22408 17740 22448
rect 17780 22408 18124 22448
rect 18164 22408 18173 22448
rect 18220 22408 18892 22448
rect 18932 22408 18941 22448
rect 19258 22408 19267 22448
rect 19307 22408 19316 22448
rect 19363 22408 19372 22448
rect 19412 22408 20309 22448
rect 11212 22313 11252 22408
rect 18220 22364 18260 22408
rect 20269 22364 20309 22408
rect 22156 22408 22292 22448
rect 22349 22408 22636 22448
rect 22676 22408 22685 22448
rect 23788 22408 24268 22448
rect 24308 22408 24317 22448
rect 26524 22408 26668 22448
rect 26708 22408 26717 22448
rect 27148 22408 29164 22448
rect 29204 22408 29356 22448
rect 29396 22408 29405 22448
rect 11491 22324 11500 22364
rect 11540 22324 11828 22364
rect 11788 22280 11828 22324
rect 13324 22324 13699 22364
rect 13739 22324 13748 22364
rect 14275 22324 14284 22364
rect 14324 22324 15188 22364
rect 13324 22280 13364 22324
rect 15148 22280 15188 22324
rect 17068 22324 18260 22364
rect 18442 22324 18451 22364
rect 18491 22324 18604 22364
rect 18644 22324 18653 22364
rect 18857 22324 18988 22364
rect 19028 22324 19171 22364
rect 19211 22324 19220 22364
rect 19625 22324 19747 22364
rect 19796 22324 19805 22364
rect 20269 22324 20338 22364
rect 20378 22324 21676 22364
rect 21716 22324 21725 22364
rect 15820 22280 15860 22289
rect 17068 22280 17108 22324
rect 22156 22322 22196 22408
rect 22156 22313 22280 22322
rect 22156 22282 22240 22313
rect 11212 22264 11252 22273
rect 11465 22240 11596 22280
rect 11636 22240 11645 22280
rect 11779 22240 11788 22280
rect 11828 22240 11837 22280
rect 11971 22240 11980 22280
rect 12020 22240 12280 22280
rect 12320 22240 12329 22280
rect 12931 22240 12940 22280
rect 12980 22240 13324 22280
rect 13364 22240 13373 22280
rect 13699 22240 13708 22280
rect 13748 22240 13804 22280
rect 13844 22240 13879 22280
rect 13987 22240 13996 22280
rect 14036 22240 14092 22280
rect 14132 22240 14167 22280
rect 15017 22240 15148 22280
rect 15188 22240 15197 22280
rect 15523 22240 15532 22280
rect 15572 22240 15724 22280
rect 15764 22240 15773 22280
rect 15860 22240 15916 22280
rect 15956 22240 15991 22280
rect 16937 22240 17068 22280
rect 17108 22240 17117 22280
rect 17897 22240 18028 22280
rect 18068 22240 18077 22280
rect 18138 22240 18147 22280
rect 18187 22240 18196 22280
rect 18256 22240 18265 22280
rect 18305 22240 18452 22280
rect 18499 22240 18508 22280
rect 18548 22240 18595 22280
rect 18635 22240 19555 22280
rect 19595 22240 19604 22280
rect 20419 22240 20428 22280
rect 20468 22240 20908 22280
rect 20948 22240 20957 22280
rect 21149 22240 21181 22280
rect 21221 22240 21236 22280
rect 21283 22240 21292 22280
rect 21332 22240 22060 22280
rect 22100 22240 22109 22280
rect 22349 22280 22389 22408
rect 22601 22324 22723 22364
rect 22772 22324 22781 22364
rect 23107 22324 23116 22364
rect 23156 22324 23186 22364
rect 23395 22324 23404 22364
rect 23444 22324 23732 22364
rect 23116 22280 23156 22324
rect 23692 22280 23732 22324
rect 24079 22324 24884 22364
rect 25498 22324 25507 22364
rect 25547 22324 25804 22364
rect 25844 22324 25853 22364
rect 25911 22324 26092 22364
rect 26132 22324 26141 22364
rect 22240 22264 22280 22273
rect 22330 22240 22339 22280
rect 22379 22240 22389 22280
rect 22594 22240 22603 22280
rect 22643 22240 22676 22280
rect 22819 22240 22828 22280
rect 22868 22240 22999 22280
rect 23090 22240 23099 22280
rect 23139 22240 23156 22280
rect 23299 22240 23308 22280
rect 23348 22240 23582 22280
rect 23674 22240 23683 22280
rect 23723 22240 23732 22280
rect 23779 22240 23788 22280
rect 23828 22240 23959 22280
rect 6604 22196 6644 22240
rect 5993 22156 6017 22196
rect 6057 22156 6124 22196
rect 6164 22156 6173 22196
rect 6403 22156 6412 22196
rect 6452 22156 6500 22196
rect 6595 22156 6604 22196
rect 6644 22156 6691 22196
rect 6782 22112 6822 22240
rect 7564 22231 7604 22240
rect 8524 22231 8564 22240
rect 10156 22196 10196 22240
rect 10444 22196 10484 22240
rect 10938 22238 11012 22240
rect 10938 22196 10978 22238
rect 15820 22231 15860 22240
rect 18147 22196 18187 22240
rect 18412 22196 18452 22240
rect 21196 22196 21236 22240
rect 7337 22156 7468 22196
rect 7508 22156 7517 22196
rect 8044 22156 8222 22196
rect 8262 22156 8271 22196
rect 8419 22156 8428 22196
rect 8468 22156 8477 22196
rect 9484 22156 9676 22196
rect 9716 22156 9725 22196
rect 10147 22156 10156 22196
rect 10196 22156 10205 22196
rect 10399 22156 10444 22196
rect 10484 22156 10493 22196
rect 10938 22156 13804 22196
rect 13844 22156 15518 22196
rect 15558 22156 15567 22196
rect 16099 22156 16108 22196
rect 16148 22156 18316 22196
rect 18356 22156 18365 22196
rect 18412 22156 19180 22196
rect 19220 22156 19229 22196
rect 21187 22156 21196 22196
rect 21236 22156 22252 22196
rect 22292 22156 22301 22196
rect 8044 22112 8084 22156
rect 8428 22112 8468 22156
rect 9484 22112 9524 22156
rect 5731 22072 5740 22112
rect 5780 22072 6220 22112
rect 6260 22072 6822 22112
rect 7913 22072 8035 22112
rect 8084 22072 8093 22112
rect 8201 22072 8236 22112
rect 8276 22072 8323 22112
rect 8363 22072 8381 22112
rect 8428 22072 9524 22112
rect 9929 22072 10060 22112
rect 10100 22072 10109 22112
rect 10243 22072 10252 22112
rect 10292 22072 10339 22112
rect 10379 22072 10423 22112
rect 10732 22072 12115 22112
rect 12155 22072 12164 22112
rect 12617 22072 12739 22112
rect 12788 22072 12797 22112
rect 13699 22072 13708 22112
rect 13748 22072 15619 22112
rect 15659 22072 15668 22112
rect 17923 22072 17932 22112
rect 17972 22072 18220 22112
rect 18260 22072 18988 22112
rect 19028 22072 19037 22112
rect 20122 22072 20131 22112
rect 20171 22072 20332 22112
rect 20372 22072 20381 22112
rect 20803 22072 20812 22112
rect 20852 22072 22459 22112
rect 22499 22072 22540 22112
rect 22580 22072 22589 22112
rect 7075 21988 7084 22028
rect 7124 21988 10348 22028
rect 10388 21988 10397 22028
rect 10732 21944 10772 22072
rect 22636 22028 22676 22240
rect 23542 22196 23582 22240
rect 24079 22196 24119 22324
rect 24844 22280 24884 22324
rect 25911 22280 25951 22324
rect 26524 22322 26564 22408
rect 26506 22282 26515 22322
rect 26555 22282 26564 22322
rect 26034 22280 26084 22281
rect 27148 22280 27188 22408
rect 27817 22324 27826 22364
rect 27866 22324 28588 22364
rect 28628 22324 28637 22364
rect 30403 22324 30412 22364
rect 30452 22324 30461 22364
rect 31258 22324 31267 22364
rect 31316 22324 31447 22364
rect 23203 22156 23212 22196
rect 23252 22156 23383 22196
rect 23542 22156 24119 22196
rect 24172 22240 24268 22280
rect 24308 22240 24317 22280
rect 24449 22240 24458 22280
rect 24498 22240 24507 22280
rect 24599 22240 24642 22280
rect 24682 22240 24691 22280
rect 24826 22240 24835 22280
rect 24875 22240 24884 22280
rect 24931 22240 24940 22280
rect 24980 22240 25036 22280
rect 25076 22240 25111 22280
rect 25289 22240 25387 22280
rect 25460 22240 25469 22280
rect 25577 22240 25612 22280
rect 25652 22240 25708 22280
rect 25748 22240 25757 22280
rect 25911 22240 25943 22280
rect 25983 22240 25992 22280
rect 26034 22240 26047 22280
rect 26087 22240 26096 22280
rect 26179 22240 26188 22280
rect 26228 22240 26237 22280
rect 26368 22240 26377 22280
rect 26417 22240 26426 22280
rect 26620 22240 26629 22280
rect 26669 22240 26708 22280
rect 26842 22240 26851 22280
rect 26891 22240 26947 22280
rect 27139 22240 27148 22280
rect 27188 22240 27197 22280
rect 27427 22240 27436 22280
rect 27476 22240 27724 22280
rect 27764 22240 27773 22280
rect 27907 22240 27916 22280
rect 27956 22240 28087 22280
rect 28195 22240 28204 22280
rect 28244 22240 28684 22280
rect 28736 22240 28745 22280
rect 29443 22240 29452 22280
rect 29492 22240 30883 22280
rect 30923 22240 30932 22280
rect 24172 22196 24212 22240
rect 24172 22156 24364 22196
rect 24404 22156 24413 22196
rect 24460 22112 24500 22240
rect 22906 22072 22915 22112
rect 22955 22072 23060 22112
rect 24451 22072 24460 22112
rect 24500 22072 24509 22112
rect 21475 21988 21484 22028
rect 21524 21988 22676 22028
rect 23020 21944 23060 22072
rect 24599 22028 24639 22240
rect 24844 22196 24884 22240
rect 26034 22196 26074 22240
rect 24730 22156 24739 22196
rect 24779 22156 24788 22196
rect 24844 22156 25132 22196
rect 25172 22156 25181 22196
rect 25507 22156 25516 22196
rect 25556 22156 25804 22196
rect 25844 22156 26074 22196
rect 23779 21988 23788 22028
rect 23828 21988 24639 22028
rect 24748 22028 24788 22156
rect 25690 22072 25699 22112
rect 25739 22072 26092 22112
rect 26132 22072 26141 22112
rect 26188 22028 26228 22240
rect 26380 22196 26420 22240
rect 26668 22196 26708 22240
rect 26860 22196 26900 22240
rect 26371 22156 26380 22196
rect 26420 22156 26464 22196
rect 26659 22156 26668 22196
rect 26708 22156 26725 22196
rect 26851 22156 26860 22196
rect 26900 22156 26909 22196
rect 28522 22156 28531 22196
rect 28571 22156 29356 22196
rect 29396 22156 29405 22196
rect 26275 22072 26284 22112
rect 26324 22072 26668 22112
rect 26708 22072 26717 22112
rect 27427 22072 27436 22112
rect 27476 22072 28972 22112
rect 29012 22072 29021 22112
rect 24748 21988 29260 22028
rect 29300 21988 29309 22028
rect 24599 21944 24639 21988
rect 0 21904 2900 21944
rect 4343 21904 4352 21944
rect 4720 21904 4729 21944
rect 5644 21904 6739 21944
rect 7555 21904 7564 21944
rect 7604 21904 7988 21944
rect 8803 21904 8812 21944
rect 8852 21904 10772 21944
rect 12117 21904 12126 21944
rect 12494 21904 12503 21944
rect 19891 21904 19900 21944
rect 20268 21904 20277 21944
rect 23020 21904 24364 21944
rect 24404 21904 24413 21944
rect 24599 21904 25132 21944
rect 25172 21904 26860 21944
rect 26900 21904 26909 21944
rect 27665 21904 27674 21944
rect 28042 21904 28051 21944
rect 0 21884 400 21904
rect 1132 21820 3148 21860
rect 3188 21820 3197 21860
rect 3331 21820 3340 21860
rect 3380 21820 5540 21860
rect 1132 21608 1172 21820
rect 1306 21736 1315 21776
rect 1355 21736 1612 21776
rect 1652 21736 1661 21776
rect 1987 21736 1996 21776
rect 2036 21736 2084 21776
rect 3401 21736 3532 21776
rect 3572 21736 3581 21776
rect 4963 21736 4972 21776
rect 5012 21736 5347 21776
rect 5387 21736 5396 21776
rect 2044 21608 2084 21736
rect 2179 21652 2188 21692
rect 2228 21652 2846 21692
rect 2886 21652 3436 21692
rect 3476 21652 3639 21692
rect 3679 21652 4148 21692
rect 4483 21652 4492 21692
rect 4532 21652 4771 21692
rect 4811 21652 4820 21692
rect 4108 21608 4148 21652
rect 5500 21608 5540 21820
rect 5932 21820 6604 21860
rect 6644 21820 6653 21860
rect 5932 21776 5972 21820
rect 6699 21776 6739 21904
rect 7948 21860 7988 21904
rect 7948 21820 8660 21860
rect 8620 21776 8660 21820
rect 9772 21820 9868 21860
rect 9908 21820 9917 21860
rect 10060 21820 11252 21860
rect 13603 21820 13612 21860
rect 13652 21820 17260 21860
rect 17300 21820 17309 21860
rect 21929 21820 22060 21860
rect 22100 21820 23308 21860
rect 23348 21820 23357 21860
rect 25699 21820 25708 21860
rect 25748 21820 27148 21860
rect 27188 21820 27620 21860
rect 9772 21776 9812 21820
rect 5914 21736 5923 21776
rect 5963 21736 5972 21776
rect 6019 21736 6028 21776
rect 6068 21736 6164 21776
rect 6307 21736 6316 21776
rect 6356 21736 6487 21776
rect 6699 21736 6883 21776
rect 6923 21736 6932 21776
rect 7363 21736 7372 21776
rect 7412 21736 7660 21776
rect 7700 21736 7709 21776
rect 8611 21736 8620 21776
rect 8660 21736 8669 21776
rect 8962 21736 9580 21776
rect 9620 21736 9629 21776
rect 9754 21736 9763 21776
rect 9803 21736 9812 21776
rect 6019 21652 6028 21692
rect 6068 21652 6077 21692
rect 1123 21568 1132 21608
rect 1172 21568 1181 21608
rect 1318 21568 1327 21608
rect 1367 21568 1376 21608
rect 1507 21575 1516 21608
rect 0 21524 400 21544
rect 1324 21524 1364 21568
rect 1418 21535 1516 21575
rect 1556 21535 1565 21608
rect 1612 21568 1621 21608
rect 1661 21568 1670 21608
rect 1795 21568 1804 21608
rect 1883 21568 1975 21608
rect 2035 21568 2044 21608
rect 2084 21568 2093 21608
rect 2921 21568 3052 21608
rect 3092 21568 3101 21608
rect 3148 21599 3188 21608
rect 0 21484 460 21524
rect 500 21484 509 21524
rect 835 21484 844 21524
rect 884 21484 893 21524
rect 1289 21484 1324 21524
rect 1364 21484 1373 21524
rect 0 21464 400 21484
rect 844 21440 884 21484
rect 1612 21440 1652 21568
rect 3322 21584 3331 21608
rect 1738 21515 2900 21524
rect 1738 21475 1747 21515
rect 1787 21484 2900 21515
rect 1787 21475 1796 21484
rect 1738 21474 1796 21475
rect 844 21400 1420 21440
rect 1460 21400 1469 21440
rect 1603 21400 1612 21440
rect 1652 21400 1661 21440
rect 2860 21356 2900 21484
rect 460 21316 604 21356
rect 644 21316 653 21356
rect 2659 21316 2668 21356
rect 2708 21316 2717 21356
rect 2842 21316 2851 21356
rect 2891 21316 2900 21356
rect 0 21104 400 21124
rect 460 21104 500 21316
rect 2668 21188 2708 21316
rect 3148 21272 3188 21559
rect 3292 21568 3331 21584
rect 3371 21568 3380 21608
rect 3427 21568 3436 21608
rect 3476 21568 3532 21608
rect 3572 21568 3607 21608
rect 3881 21568 3916 21608
rect 3956 21599 4052 21608
rect 3956 21568 4003 21599
rect 3292 21544 3380 21568
rect 3994 21559 4003 21568
rect 4043 21559 4052 21599
rect 4108 21568 4439 21608
rect 4479 21568 4488 21608
rect 4675 21568 4684 21608
rect 4724 21568 4876 21608
rect 4916 21568 4925 21608
rect 5340 21568 5452 21608
rect 5492 21568 5500 21608
rect 5540 21568 5549 21608
rect 5635 21568 5644 21608
rect 5684 21568 5822 21608
rect 5862 21568 5871 21608
rect 3994 21558 4052 21559
rect 3292 21524 3332 21544
rect 3235 21484 3244 21524
rect 3284 21484 3332 21524
rect 4012 21440 4052 21558
rect 5644 21524 5684 21568
rect 4099 21484 4108 21524
rect 4148 21484 4156 21524
rect 4196 21484 4279 21524
rect 4570 21484 4579 21524
rect 4619 21484 4780 21524
rect 4820 21484 4829 21524
rect 4963 21484 4972 21524
rect 5012 21484 5143 21524
rect 5539 21484 5548 21524
rect 5588 21484 5684 21524
rect 6028 21440 6068 21652
rect 6124 21599 6164 21736
rect 8962 21692 9002 21736
rect 10060 21692 10100 21820
rect 10732 21776 10772 21820
rect 11212 21776 11252 21820
rect 10313 21736 10435 21776
rect 10484 21736 10493 21776
rect 10714 21736 10723 21776
rect 10763 21736 10772 21776
rect 10862 21736 10924 21776
rect 10964 21736 10978 21776
rect 11194 21736 11203 21776
rect 11243 21736 11252 21776
rect 11418 21736 12940 21776
rect 12980 21736 12989 21776
rect 13577 21736 13603 21776
rect 13643 21736 13708 21776
rect 13748 21736 13757 21776
rect 10732 21692 10772 21736
rect 10938 21692 10978 21736
rect 11418 21692 11458 21736
rect 15052 21692 15092 21820
rect 15139 21736 15148 21776
rect 15188 21736 15907 21776
rect 15947 21736 15956 21776
rect 18019 21736 18028 21776
rect 18068 21736 18604 21776
rect 18644 21736 18653 21776
rect 20899 21736 20908 21776
rect 20948 21736 21908 21776
rect 6629 21652 6782 21692
rect 6822 21652 6831 21692
rect 7337 21652 7468 21692
rect 7508 21652 7852 21692
rect 7892 21652 7901 21692
rect 7948 21652 8092 21692
rect 8132 21652 8141 21692
rect 8227 21652 8236 21692
rect 8276 21652 9002 21692
rect 9379 21652 9388 21692
rect 9428 21652 10100 21692
rect 10147 21652 10156 21692
rect 10196 21652 10218 21692
rect 10348 21652 10772 21692
rect 10929 21652 10938 21692
rect 10978 21652 11418 21692
rect 11458 21652 11467 21692
rect 11657 21652 11740 21692
rect 11780 21652 11788 21692
rect 11828 21652 11837 21692
rect 11971 21652 11980 21692
rect 12020 21652 14764 21692
rect 14804 21652 14813 21692
rect 15052 21652 15327 21692
rect 15486 21652 15532 21692
rect 15572 21652 15581 21692
rect 16003 21652 16012 21692
rect 16052 21652 16723 21692
rect 16763 21652 16772 21692
rect 16972 21652 18307 21692
rect 18347 21652 18356 21692
rect 18412 21652 19276 21692
rect 19316 21652 19325 21692
rect 20236 21652 20756 21692
rect 6629 21608 6669 21652
rect 7372 21608 7412 21652
rect 7948 21608 7988 21652
rect 8962 21608 9002 21652
rect 9676 21608 9716 21652
rect 10156 21608 10196 21652
rect 10348 21608 10388 21652
rect 6307 21568 6316 21608
rect 6356 21568 6412 21608
rect 6452 21568 6487 21608
rect 6595 21568 6604 21608
rect 6669 21568 6775 21608
rect 6857 21568 6988 21608
rect 7028 21568 7037 21608
rect 7084 21599 7124 21608
rect 6124 21550 6164 21559
rect 7363 21568 7372 21608
rect 7412 21568 7421 21608
rect 7555 21568 7564 21608
rect 7604 21568 7613 21608
rect 7747 21568 7756 21608
rect 7796 21568 7805 21608
rect 7939 21568 7948 21608
rect 7988 21568 7997 21608
rect 8044 21568 8284 21608
rect 8324 21568 8333 21608
rect 8419 21568 8428 21608
rect 8468 21568 8599 21608
rect 8702 21568 8716 21608
rect 8756 21568 8765 21608
rect 8944 21568 8953 21608
rect 8993 21568 9002 21608
rect 9283 21568 9292 21608
rect 9332 21568 9341 21608
rect 9475 21568 9484 21608
rect 9524 21568 9533 21608
rect 9658 21568 9667 21608
rect 9707 21568 9716 21608
rect 9966 21575 9975 21608
rect 9868 21568 9975 21575
rect 10015 21568 10024 21608
rect 10122 21568 10131 21608
rect 10171 21568 10196 21608
rect 10339 21568 10348 21608
rect 10388 21568 10397 21608
rect 10618 21568 10627 21608
rect 10667 21568 10732 21608
rect 10772 21568 10807 21608
rect 11036 21568 11045 21608
rect 11085 21568 11107 21608
rect 11147 21568 11216 21608
rect 11465 21599 11596 21608
rect 11465 21568 11587 21599
rect 11636 21568 11645 21608
rect 11875 21568 11884 21608
rect 11924 21568 12211 21608
rect 12251 21568 12260 21608
rect 12634 21568 12643 21608
rect 12692 21568 12823 21608
rect 13385 21568 13516 21608
rect 13556 21568 13565 21608
rect 13612 21568 13751 21608
rect 13791 21568 13800 21608
rect 13987 21568 13996 21608
rect 14036 21568 14188 21608
rect 14228 21568 14237 21608
rect 14458 21568 14467 21608
rect 14516 21568 14647 21608
rect 14921 21568 15052 21608
rect 15092 21568 15101 21608
rect 6522 21484 6531 21524
rect 6571 21484 6796 21524
rect 6836 21484 6845 21524
rect 4012 21400 5212 21440
rect 5252 21400 5740 21440
rect 5780 21400 5789 21440
rect 6028 21400 6988 21440
rect 7028 21400 7037 21440
rect 7084 21356 7124 21559
rect 7564 21524 7604 21568
rect 7555 21484 7564 21524
rect 7604 21484 7651 21524
rect 7756 21440 7796 21568
rect 8044 21524 8084 21568
rect 8702 21524 8742 21568
rect 9292 21524 9332 21568
rect 8035 21484 8044 21524
rect 8084 21484 8093 21524
rect 8702 21484 8756 21524
rect 8826 21484 8835 21524
rect 8875 21484 8884 21524
rect 9292 21484 9388 21524
rect 9428 21484 9437 21524
rect 7267 21400 7276 21440
rect 7316 21400 8236 21440
rect 8276 21400 8285 21440
rect 8716 21356 8756 21484
rect 7084 21316 7796 21356
rect 7843 21316 7852 21356
rect 7892 21316 8756 21356
rect 7756 21272 7796 21316
rect 3148 21232 4780 21272
rect 4820 21232 4829 21272
rect 7756 21232 8428 21272
rect 8468 21232 8477 21272
rect 8835 21188 8875 21484
rect 2668 21148 2956 21188
rect 2996 21148 3005 21188
rect 3103 21148 3112 21188
rect 3480 21148 3489 21188
rect 7939 21148 7948 21188
rect 7988 21148 8875 21188
rect 9484 21104 9524 21568
rect 9868 21535 10015 21568
rect 11578 21559 11587 21568
rect 11627 21559 11636 21568
rect 11578 21558 11636 21559
rect 9868 21440 9908 21535
rect 12394 21526 12403 21566
rect 12443 21526 12500 21566
rect 12460 21524 12500 21526
rect 13612 21524 13652 21568
rect 15287 21566 15327 21652
rect 15532 21608 15572 21652
rect 16972 21608 17012 21652
rect 18412 21608 18452 21652
rect 20236 21608 20276 21652
rect 20716 21608 20756 21652
rect 21484 21652 21772 21692
rect 21812 21652 21821 21692
rect 21484 21608 21524 21652
rect 21868 21608 21908 21736
rect 22060 21608 22100 21820
rect 27580 21776 27620 21820
rect 22147 21736 22156 21776
rect 22196 21736 22732 21776
rect 22772 21736 22781 21776
rect 23561 21736 23596 21776
rect 23636 21736 23692 21776
rect 23732 21736 23741 21776
rect 24163 21736 24172 21776
rect 24212 21736 24556 21776
rect 24596 21736 24605 21776
rect 24652 21736 25420 21776
rect 25460 21736 25564 21776
rect 25604 21736 25613 21776
rect 26371 21736 26380 21776
rect 26420 21736 26668 21776
rect 26708 21736 26717 21776
rect 26851 21736 26860 21776
rect 26900 21736 27259 21776
rect 27299 21736 27308 21776
rect 27571 21736 27580 21776
rect 27620 21736 27629 21776
rect 28099 21736 28108 21776
rect 28148 21736 28157 21776
rect 28627 21736 28636 21776
rect 28676 21736 29452 21776
rect 29492 21736 29501 21776
rect 24652 21692 24692 21736
rect 28108 21692 28148 21736
rect 22531 21652 22540 21692
rect 22580 21652 23156 21692
rect 23116 21608 23156 21652
rect 23980 21652 24652 21692
rect 24692 21652 24701 21692
rect 25123 21652 25132 21692
rect 25172 21652 25218 21692
rect 25603 21652 25612 21692
rect 25652 21652 25748 21692
rect 23980 21608 24020 21652
rect 25131 21608 25171 21652
rect 25708 21608 25748 21652
rect 25996 21652 26284 21692
rect 26324 21652 26572 21692
rect 26612 21652 26621 21692
rect 27048 21652 27436 21692
rect 27476 21652 27485 21692
rect 27867 21652 27916 21692
rect 27956 21652 27998 21692
rect 28038 21652 28047 21692
rect 28108 21652 28340 21692
rect 28954 21652 28963 21692
rect 29012 21652 29143 21692
rect 15524 21568 15533 21608
rect 15573 21568 15582 21608
rect 15628 21568 16052 21608
rect 16099 21568 16108 21608
rect 16148 21568 16195 21608
rect 16235 21568 16279 21608
rect 16766 21568 16876 21608
rect 16928 21568 17012 21608
rect 17059 21568 17068 21608
rect 17108 21568 17117 21608
rect 17251 21568 17260 21608
rect 17300 21568 17644 21608
rect 17684 21568 17693 21608
rect 17932 21568 18452 21608
rect 18499 21568 18508 21608
rect 18548 21568 18595 21608
rect 18635 21568 18679 21608
rect 18857 21568 18988 21608
rect 19028 21568 19037 21608
rect 19171 21568 19180 21608
rect 19220 21568 19351 21608
rect 19564 21568 19756 21608
rect 19796 21568 19805 21608
rect 19984 21568 19993 21608
rect 20033 21568 20276 21608
rect 20323 21568 20332 21608
rect 20372 21568 20503 21608
rect 20585 21568 20716 21608
rect 20756 21568 20765 21608
rect 21091 21568 21100 21608
rect 21140 21568 21149 21608
rect 21475 21568 21484 21608
rect 21524 21568 21533 21608
rect 21629 21568 21671 21608
rect 21711 21568 21720 21608
rect 21859 21568 21868 21608
rect 21908 21568 21917 21608
rect 22051 21568 22060 21608
rect 22100 21568 22109 21608
rect 22234 21568 22243 21608
rect 22292 21568 22423 21608
rect 22714 21568 22723 21608
rect 22763 21568 22772 21608
rect 22819 21568 22828 21608
rect 22868 21568 22999 21608
rect 23116 21568 23404 21608
rect 23444 21568 23453 21608
rect 23587 21568 23596 21608
rect 23636 21568 24020 21608
rect 24154 21568 24163 21608
rect 24203 21568 24212 21608
rect 24259 21568 24268 21608
rect 24308 21568 24317 21608
rect 24451 21568 24460 21608
rect 24500 21568 24599 21608
rect 24639 21568 24648 21608
rect 24835 21568 24844 21608
rect 24884 21568 25015 21608
rect 25122 21568 25131 21608
rect 25171 21568 25180 21608
rect 25306 21568 25315 21608
rect 25355 21568 25364 21608
rect 25411 21568 25420 21608
rect 25460 21568 25591 21608
rect 25699 21568 25708 21608
rect 25748 21568 25757 21608
rect 15283 21526 15292 21566
rect 15332 21526 15341 21566
rect 15628 21524 15668 21568
rect 16012 21524 16052 21568
rect 17068 21524 17108 21568
rect 10234 21484 10243 21524
rect 10283 21484 10484 21524
rect 12460 21484 13268 21524
rect 13603 21484 13612 21524
rect 13652 21484 13661 21524
rect 13853 21484 13891 21524
rect 13931 21484 13940 21524
rect 14083 21484 14092 21524
rect 14132 21484 14284 21524
rect 14324 21484 14333 21524
rect 14851 21484 14860 21524
rect 14900 21484 14909 21524
rect 15389 21484 15427 21524
rect 15467 21484 15476 21524
rect 15619 21484 15628 21524
rect 15668 21484 15677 21524
rect 15724 21484 15811 21524
rect 15851 21484 15860 21524
rect 16012 21484 16387 21524
rect 16427 21484 16436 21524
rect 16675 21484 16684 21524
rect 16724 21484 17108 21524
rect 9868 21400 10252 21440
rect 10292 21400 10301 21440
rect 9955 21316 9964 21356
rect 10004 21316 10060 21356
rect 10100 21316 10164 21356
rect 10444 21272 10484 21484
rect 10924 21400 11404 21440
rect 11444 21400 11453 21440
rect 11587 21400 11596 21440
rect 11636 21400 12844 21440
rect 12884 21400 12893 21440
rect 10924 21356 10964 21400
rect 13228 21356 13268 21484
rect 13900 21440 13940 21484
rect 14860 21440 14900 21484
rect 15436 21440 15476 21484
rect 13891 21400 13900 21440
rect 13940 21400 13949 21440
rect 14083 21400 14092 21440
rect 14132 21400 15380 21440
rect 15427 21400 15436 21440
rect 15476 21400 15485 21440
rect 10915 21316 10924 21356
rect 10964 21316 10973 21356
rect 11395 21316 11404 21356
rect 11444 21316 11453 21356
rect 13027 21316 13036 21356
rect 13076 21316 13085 21356
rect 13219 21316 13228 21356
rect 13268 21316 13324 21356
rect 13364 21316 13399 21356
rect 15187 21316 15196 21356
rect 15236 21316 15245 21356
rect 11404 21272 11444 21316
rect 9955 21232 9964 21272
rect 10004 21232 10484 21272
rect 10531 21232 10540 21272
rect 10580 21232 11444 21272
rect 13036 21272 13076 21316
rect 13036 21232 14380 21272
rect 14420 21232 14429 21272
rect 15196 21188 15236 21316
rect 15340 21272 15380 21400
rect 15724 21272 15764 21484
rect 17932 21440 17972 21568
rect 18089 21484 18211 21524
rect 18260 21484 18269 21524
rect 18778 21484 18787 21524
rect 18827 21484 19468 21524
rect 19508 21484 19517 21524
rect 17635 21400 17644 21440
rect 17684 21400 17972 21440
rect 18019 21400 18028 21440
rect 18068 21400 18077 21440
rect 17033 21316 17164 21356
rect 17204 21316 17213 21356
rect 15340 21232 15764 21272
rect 18028 21272 18068 21400
rect 18499 21316 18508 21356
rect 18548 21316 18988 21356
rect 19028 21316 19037 21356
rect 19564 21272 19604 21568
rect 20332 21524 20372 21568
rect 19651 21484 19660 21524
rect 19700 21484 19709 21524
rect 19882 21515 20372 21524
rect 19660 21356 19700 21484
rect 19882 21475 19891 21515
rect 19931 21484 20372 21515
rect 19931 21475 19940 21484
rect 19882 21474 19940 21475
rect 20035 21400 20044 21440
rect 20084 21400 20092 21440
rect 20132 21400 20215 21440
rect 20777 21400 20860 21440
rect 20900 21400 20908 21440
rect 20948 21400 20957 21440
rect 21100 21356 21140 21568
rect 21676 21524 21716 21568
rect 21868 21524 21908 21568
rect 22732 21524 22772 21568
rect 24172 21524 24212 21568
rect 21667 21484 21676 21524
rect 21716 21484 21725 21524
rect 21868 21484 22060 21524
rect 22100 21484 22109 21524
rect 22732 21484 22924 21524
rect 22964 21484 22973 21524
rect 23020 21484 24172 21524
rect 24212 21484 24221 21524
rect 23020 21440 23060 21484
rect 24268 21440 24308 21568
rect 25324 21524 25364 21568
rect 25996 21524 26036 21652
rect 26083 21568 26092 21608
rect 26132 21599 26263 21608
rect 26132 21568 26179 21599
rect 26170 21559 26179 21568
rect 26219 21568 26263 21599
rect 26467 21568 26476 21608
rect 26516 21568 26525 21608
rect 27048 21599 27088 21652
rect 27436 21608 27476 21652
rect 26219 21559 26228 21568
rect 26170 21558 26228 21559
rect 24355 21484 24364 21524
rect 24404 21484 24739 21524
rect 24779 21484 24788 21524
rect 24931 21484 24940 21524
rect 24980 21484 24989 21524
rect 25123 21484 25132 21524
rect 25172 21484 25364 21524
rect 25420 21484 26036 21524
rect 24940 21440 24980 21484
rect 25420 21440 25460 21484
rect 26476 21440 26516 21568
rect 27130 21568 27139 21608
rect 27179 21568 27244 21608
rect 27284 21568 27319 21608
rect 27418 21599 27523 21608
rect 27048 21550 27088 21559
rect 27418 21559 27427 21599
rect 27467 21568 27523 21599
rect 27619 21568 27628 21608
rect 27668 21568 28204 21608
rect 28244 21568 28253 21608
rect 28300 21599 28340 21652
rect 27467 21559 27476 21568
rect 27418 21558 27476 21559
rect 28300 21550 28340 21559
rect 28474 21599 28684 21608
rect 28474 21559 28483 21599
rect 28523 21568 28684 21599
rect 28724 21568 28733 21608
rect 29338 21568 29347 21608
rect 29396 21568 29527 21608
rect 28523 21559 28532 21568
rect 28474 21558 28532 21559
rect 30403 21484 30412 21524
rect 30452 21484 30461 21524
rect 21859 21400 21868 21440
rect 21908 21400 23060 21440
rect 23273 21400 23308 21440
rect 23348 21400 23395 21440
rect 23435 21400 23453 21440
rect 24268 21400 24980 21440
rect 25411 21400 25420 21440
rect 25460 21400 25469 21440
rect 26476 21400 27532 21440
rect 27572 21400 27581 21440
rect 24940 21356 24980 21400
rect 19660 21316 21140 21356
rect 21353 21316 21484 21356
rect 21524 21316 21772 21356
rect 21812 21316 21821 21356
rect 23002 21316 23011 21356
rect 23051 21316 23116 21356
rect 23156 21316 23191 21356
rect 24329 21316 24460 21356
rect 24500 21316 24509 21356
rect 24940 21316 25324 21356
rect 25364 21316 25373 21356
rect 25987 21316 25996 21356
rect 26036 21316 26045 21356
rect 26659 21316 26668 21356
rect 26708 21316 26755 21356
rect 26795 21316 26839 21356
rect 27619 21316 27628 21356
rect 27668 21316 28003 21356
rect 28043 21316 28052 21356
rect 29539 21316 29548 21356
rect 29588 21316 30988 21356
rect 31028 21316 31276 21356
rect 31316 21316 31325 21356
rect 21388 21272 21428 21316
rect 18028 21232 19508 21272
rect 19564 21232 21428 21272
rect 22819 21232 22828 21272
rect 22868 21232 24844 21272
rect 24884 21232 24893 21272
rect 19468 21188 19508 21232
rect 9667 21148 9676 21188
rect 9716 21148 10143 21188
rect 10877 21148 10886 21188
rect 11254 21148 11263 21188
rect 15196 21148 15628 21188
rect 15668 21148 15677 21188
rect 18651 21148 18660 21188
rect 19028 21148 19037 21188
rect 19468 21148 21004 21188
rect 21044 21148 21053 21188
rect 10103 21104 10143 21148
rect 25996 21104 26036 21316
rect 26425 21148 26434 21188
rect 26802 21148 26811 21188
rect 0 21064 500 21104
rect 844 21064 3572 21104
rect 0 21044 400 21064
rect 451 20980 460 21020
rect 500 20980 604 21020
rect 644 20980 653 21020
rect 844 20852 884 21064
rect 3532 21020 3572 21064
rect 3628 21064 5068 21104
rect 5108 21064 6452 21104
rect 9091 21064 9100 21104
rect 9140 21064 9327 21104
rect 9484 21064 9812 21104
rect 10103 21064 11596 21104
rect 11636 21064 11645 21104
rect 14851 21064 14860 21104
rect 14900 21064 27088 21104
rect 28675 21064 28684 21104
rect 28724 21064 30316 21104
rect 30356 21064 30365 21104
rect 1097 20980 1228 21020
rect 1268 20980 1277 21020
rect 1356 20980 1420 21020
rect 1460 20980 3380 21020
rect 3523 20980 3532 21020
rect 3572 20980 3581 21020
rect 835 20812 844 20852
rect 884 20812 893 20852
rect 1411 20812 1420 20852
rect 1460 20812 1469 20852
rect 1420 20768 1460 20812
rect 1516 20768 1556 20980
rect 1708 20896 3244 20936
rect 3284 20896 3293 20936
rect 1708 20773 1748 20896
rect 3340 20852 3380 20980
rect 3628 20852 3668 21064
rect 4954 20980 4963 21020
rect 5003 20980 5548 21020
rect 5588 20980 5597 21020
rect 3916 20896 5068 20936
rect 5108 20896 5117 20936
rect 5164 20896 5684 20936
rect 5731 20896 5740 20936
rect 5780 20896 6057 20936
rect 3916 20852 3956 20896
rect 5164 20852 5204 20896
rect 1843 20812 1900 20852
rect 1940 20812 1949 20852
rect 3100 20812 3668 20852
rect 3907 20812 3916 20852
rect 3956 20812 3965 20852
rect 4265 20843 4396 20852
rect 4265 20812 4339 20843
rect 1123 20728 1132 20768
rect 1172 20728 1181 20768
rect 1315 20728 1324 20768
rect 1364 20728 1460 20768
rect 1507 20728 1516 20768
rect 1556 20728 1565 20768
rect 1699 20733 1708 20773
rect 1748 20733 1757 20773
rect 1843 20768 1883 20812
rect 2574 20768 2614 20777
rect 3100 20768 3140 20812
rect 4330 20803 4339 20812
rect 4379 20812 4396 20843
rect 4436 20812 4445 20852
rect 5033 20812 5164 20852
rect 5204 20812 5213 20852
rect 5260 20812 5548 20852
rect 5588 20812 5597 20852
rect 4379 20803 4388 20812
rect 4330 20802 4388 20803
rect 5260 20768 5300 20812
rect 5644 20768 5684 20896
rect 5812 20812 5836 20852
rect 5876 20812 5885 20852
rect 5812 20768 5853 20812
rect 6017 20768 6057 20896
rect 6412 20852 6452 21064
rect 7241 20980 7372 21020
rect 7412 20980 7421 21020
rect 7817 20980 7948 21020
rect 7988 20980 7997 21020
rect 9043 20980 9052 21020
rect 9092 20980 9196 21020
rect 9236 20980 9245 21020
rect 9287 20936 9327 21064
rect 9379 20980 9388 21020
rect 9428 20980 9676 21020
rect 9716 20980 9725 21020
rect 9772 20936 9812 21064
rect 11875 20980 11884 21020
rect 11924 20980 13084 21020
rect 13124 20980 13133 21020
rect 13891 20980 13900 21020
rect 13940 20980 14371 21020
rect 14411 20980 14420 21020
rect 14476 20980 15188 21020
rect 15427 20980 15436 21020
rect 15476 20980 15628 21020
rect 15668 20980 15677 21020
rect 16963 20980 16972 21020
rect 17012 20980 17155 21020
rect 17195 20980 17204 21020
rect 18883 20980 18892 21020
rect 18932 20980 19412 21020
rect 20419 20980 20428 21020
rect 20468 20980 20515 21020
rect 20555 20980 20599 21020
rect 21161 20980 21292 21020
rect 21332 20980 21341 21020
rect 24425 20980 24451 21020
rect 24491 20980 24556 21020
rect 24596 20980 24605 21020
rect 25673 20980 25804 21020
rect 25844 20980 25853 21020
rect 26371 20980 26380 21020
rect 26420 20980 26860 21020
rect 26900 20980 26909 21020
rect 14476 20936 14516 20980
rect 7084 20896 7276 20936
rect 7316 20896 7325 20936
rect 7555 20896 7564 20936
rect 7604 20896 8180 20936
rect 8227 20896 8236 20936
rect 8276 20896 8285 20936
rect 9287 20896 9716 20936
rect 9772 20896 10387 20936
rect 7084 20852 7124 20896
rect 8140 20852 8180 20896
rect 8236 20852 8276 20896
rect 6211 20812 6220 20852
rect 6260 20812 6305 20852
rect 6412 20812 6844 20852
rect 6884 20812 6893 20852
rect 7075 20812 7084 20852
rect 7124 20812 7133 20852
rect 7459 20812 7468 20852
rect 7508 20812 7517 20852
rect 7651 20812 7660 20852
rect 7700 20812 7743 20852
rect 8131 20812 8140 20852
rect 8180 20812 8189 20852
rect 8236 20812 8355 20852
rect 8395 20812 8404 20852
rect 8489 20812 8620 20852
rect 8660 20812 8669 20852
rect 9283 20812 9292 20852
rect 9332 20812 9580 20852
rect 9620 20812 9629 20852
rect 6220 20768 6260 20812
rect 6412 20768 6452 20812
rect 7468 20768 7508 20812
rect 7703 20768 7743 20812
rect 9676 20768 9716 20896
rect 10252 20768 10292 20777
rect 1843 20728 1900 20768
rect 1940 20728 1949 20768
rect 2057 20728 2092 20768
rect 2132 20728 2188 20768
rect 2228 20728 2237 20768
rect 2443 20728 2572 20768
rect 2614 20728 2621 20768
rect 3082 20728 3091 20768
rect 3131 20728 3140 20768
rect 3226 20728 3235 20768
rect 3275 20728 3532 20768
rect 3572 20728 3581 20768
rect 4003 20728 4012 20768
rect 4052 20728 4204 20768
rect 4244 20728 4253 20768
rect 4432 20728 4441 20768
rect 4481 20728 4588 20768
rect 4628 20728 4637 20768
rect 4771 20728 4780 20768
rect 4820 20728 4829 20768
rect 4954 20728 4963 20768
rect 5012 20728 5143 20768
rect 5251 20728 5260 20768
rect 5300 20728 5309 20768
rect 5370 20728 5379 20768
rect 5419 20728 5428 20768
rect 5488 20728 5497 20768
rect 5537 20728 5588 20768
rect 5635 20728 5644 20768
rect 5684 20728 5693 20768
rect 5812 20728 5827 20768
rect 5867 20728 5876 20768
rect 6017 20728 6029 20768
rect 6069 20728 6078 20768
rect 6209 20728 6218 20768
rect 6258 20728 6267 20768
rect 6403 20728 6412 20768
rect 6452 20728 6461 20768
rect 6595 20728 6604 20768
rect 6644 20728 6796 20768
rect 6836 20728 6845 20768
rect 7145 20728 7276 20768
rect 7316 20728 7325 20768
rect 7421 20728 7467 20768
rect 7507 20728 7516 20768
rect 7642 20728 7651 20768
rect 7691 20728 7743 20768
rect 8105 20728 8236 20768
rect 8276 20728 8285 20768
rect 8393 20728 8473 20768
rect 8513 20728 8524 20768
rect 8564 20728 8573 20768
rect 8702 20728 8716 20768
rect 8756 20728 8765 20768
rect 8842 20759 8900 20768
rect 8842 20757 8851 20759
rect 0 20684 400 20704
rect 0 20644 460 20684
rect 500 20644 509 20684
rect 0 20624 400 20644
rect 1132 20600 1172 20728
rect 2574 20719 2614 20728
rect 4780 20684 4820 20728
rect 1603 20644 1612 20684
rect 1652 20644 2132 20684
rect 2249 20644 2273 20684
rect 2313 20644 2380 20684
rect 2420 20644 2429 20684
rect 2851 20644 2860 20684
rect 2900 20644 3543 20684
rect 3583 20644 4108 20684
rect 4148 20644 4157 20684
rect 4780 20644 5260 20684
rect 5300 20644 5309 20684
rect 2092 20600 2132 20644
rect 5379 20600 5419 20728
rect 5548 20684 5588 20728
rect 8476 20684 8516 20728
rect 5548 20644 5876 20684
rect 6115 20644 6124 20684
rect 6164 20644 6508 20684
rect 6548 20644 6557 20684
rect 7721 20644 7756 20684
rect 7796 20644 7852 20684
rect 7892 20644 7901 20684
rect 7953 20644 7962 20684
rect 8002 20644 8516 20684
rect 5836 20600 5876 20644
rect 8702 20600 8742 20728
rect 1132 20560 1612 20600
rect 1652 20560 1661 20600
rect 1865 20560 1996 20600
rect 2036 20560 2045 20600
rect 2092 20560 2188 20600
rect 2228 20560 2237 20600
rect 2362 20560 2371 20600
rect 2411 20560 2420 20600
rect 2467 20560 2476 20600
rect 2516 20560 2764 20600
rect 2804 20560 2813 20600
rect 2890 20560 2899 20600
rect 2939 20560 3052 20600
rect 3092 20560 3101 20600
rect 3209 20560 3331 20600
rect 3380 20560 3389 20600
rect 3667 20560 3676 20600
rect 3716 20560 3916 20600
rect 3956 20560 3965 20600
rect 4387 20560 4396 20600
rect 4436 20560 5419 20600
rect 5609 20560 5740 20600
rect 5780 20560 5789 20600
rect 5836 20560 6220 20600
rect 6260 20560 6269 20600
rect 6403 20560 6412 20600
rect 6452 20560 6604 20600
rect 6644 20560 6653 20600
rect 8227 20560 8236 20600
rect 8276 20560 8742 20600
rect 8835 20719 8851 20757
rect 8891 20719 8900 20759
rect 8944 20728 8953 20768
rect 8993 20728 9004 20768
rect 9044 20728 9133 20768
rect 9379 20728 9388 20768
rect 9428 20728 9580 20768
rect 9620 20728 9629 20768
rect 9676 20728 9763 20768
rect 9803 20728 10252 20768
rect 10252 20719 10292 20728
rect 8835 20717 8900 20719
rect 2380 20516 2420 20560
rect 8835 20516 8875 20717
rect 9667 20644 9676 20684
rect 9716 20644 9950 20684
rect 9990 20644 9999 20684
rect 10347 20600 10387 20896
rect 11068 20896 14516 20936
rect 15148 20936 15188 20980
rect 15148 20896 15916 20936
rect 15956 20896 15965 20936
rect 11068 20810 11108 20896
rect 14083 20812 14092 20852
rect 14132 20812 14141 20852
rect 14825 20812 14860 20852
rect 14900 20812 14947 20852
rect 14987 20812 15005 20852
rect 11050 20770 11059 20810
rect 11099 20770 11108 20810
rect 11533 20728 11542 20768
rect 11582 20728 11683 20768
rect 11723 20728 11732 20768
rect 11779 20728 11788 20768
rect 11828 20728 12364 20768
rect 12404 20728 12413 20768
rect 12547 20728 12556 20768
rect 12596 20728 12652 20768
rect 12692 20728 12727 20768
rect 12835 20728 12844 20768
rect 12884 20728 13015 20768
rect 13123 20728 13132 20768
rect 13172 20728 13228 20768
rect 13268 20728 13652 20768
rect 13741 20728 13750 20768
rect 13790 20728 13900 20768
rect 13940 20728 13949 20768
rect 14043 20728 14052 20768
rect 14092 20728 14132 20812
rect 14668 20768 14708 20777
rect 15148 20768 15188 20896
rect 19372 20852 19412 20980
rect 19459 20896 19468 20936
rect 19508 20896 19988 20936
rect 21737 20896 21868 20936
rect 21908 20896 21917 20936
rect 19948 20852 19988 20896
rect 24556 20852 24596 20980
rect 27048 20936 27088 21064
rect 27593 20980 27715 21020
rect 27764 20980 27773 21020
rect 28195 20980 28204 21020
rect 28244 20980 29836 21020
rect 29876 20980 29885 21020
rect 25699 20896 25708 20936
rect 25748 20896 26420 20936
rect 27048 20896 27177 20936
rect 17059 20812 17068 20852
rect 17108 20812 17260 20852
rect 17300 20812 17492 20852
rect 17452 20768 17492 20812
rect 17932 20812 18412 20852
rect 18452 20812 18461 20852
rect 18691 20812 18700 20852
rect 18740 20812 18836 20852
rect 19075 20812 19084 20852
rect 19124 20812 19133 20852
rect 19258 20812 19267 20852
rect 19307 20812 19412 20852
rect 19459 20812 19468 20852
rect 19508 20812 19756 20852
rect 19796 20812 19805 20852
rect 19939 20812 19948 20852
rect 19988 20812 19997 20852
rect 21292 20812 21580 20852
rect 21620 20812 21629 20852
rect 21868 20812 21964 20852
rect 22004 20812 22013 20852
rect 24163 20812 24172 20852
rect 24212 20812 24404 20852
rect 24556 20812 24739 20852
rect 24779 20812 24788 20852
rect 25193 20812 25315 20852
rect 25364 20812 25373 20852
rect 25603 20812 25612 20852
rect 25652 20812 26132 20852
rect 17932 20768 17972 20812
rect 18796 20768 18836 20812
rect 19084 20768 19124 20812
rect 21292 20768 21332 20812
rect 21868 20768 21908 20812
rect 24364 20768 24404 20812
rect 26092 20768 26132 20812
rect 26380 20768 26420 20896
rect 27137 20768 27177 20896
rect 28291 20812 28300 20852
rect 28340 20812 28963 20852
rect 29003 20812 29012 20852
rect 29347 20812 29356 20852
rect 29396 20812 31220 20852
rect 28492 20768 28532 20812
rect 31180 20768 31220 20812
rect 14179 20728 14188 20768
rect 14228 20728 14372 20768
rect 14441 20728 14572 20768
rect 14612 20728 14621 20768
rect 14818 20728 14827 20768
rect 14867 20728 14876 20768
rect 15043 20728 15052 20768
rect 15092 20728 15188 20768
rect 15322 20728 15331 20768
rect 15371 20728 15628 20768
rect 15668 20728 15677 20768
rect 16141 20728 16150 20768
rect 16190 20728 16396 20768
rect 16436 20728 16445 20768
rect 16771 20728 16780 20768
rect 16820 20759 17164 20768
rect 16820 20728 17059 20759
rect 13612 20684 13652 20728
rect 14332 20684 14372 20728
rect 14668 20684 14708 20728
rect 14836 20684 14876 20728
rect 17050 20719 17059 20728
rect 17099 20728 17164 20759
rect 17204 20728 17213 20768
rect 17347 20728 17356 20768
rect 17396 20728 17405 20768
rect 17452 20728 17687 20768
rect 17727 20728 17736 20768
rect 17818 20728 17827 20768
rect 17867 20728 17876 20768
rect 17923 20728 17932 20768
rect 17972 20728 17981 20768
rect 18089 20728 18211 20768
rect 18260 20728 18269 20768
rect 18391 20728 18508 20768
rect 18562 20728 18700 20768
rect 18740 20728 18749 20768
rect 18796 20728 18839 20768
rect 18879 20728 18888 20768
rect 19084 20728 19127 20768
rect 19167 20728 19176 20768
rect 19228 20728 19353 20768
rect 19393 20728 19402 20768
rect 19598 20728 19607 20768
rect 19647 20728 19656 20768
rect 19738 20728 19747 20768
rect 19787 20728 19796 20768
rect 19843 20728 19852 20768
rect 19892 20728 20180 20768
rect 20611 20728 20620 20768
rect 20660 20728 20812 20768
rect 20852 20728 20908 20768
rect 20948 20728 20957 20768
rect 21283 20728 21292 20768
rect 21332 20728 21341 20768
rect 21475 20728 21484 20768
rect 21524 20728 21908 20768
rect 22025 20728 22156 20768
rect 22196 20728 22205 20768
rect 23098 20728 23107 20768
rect 23156 20728 23287 20768
rect 24154 20728 24163 20768
rect 24203 20728 24212 20768
rect 24261 20728 24270 20768
rect 24310 20728 24319 20768
rect 24364 20728 25123 20768
rect 25163 20728 25172 20768
rect 25603 20728 25612 20768
rect 25652 20728 25661 20768
rect 26083 20728 26092 20768
rect 26132 20728 26141 20768
rect 26266 20728 26275 20768
rect 26315 20728 26324 20768
rect 26371 20728 26380 20768
rect 26420 20728 26551 20768
rect 26650 20728 26659 20768
rect 26699 20728 26708 20768
rect 26836 20728 26860 20768
rect 26900 20728 26967 20768
rect 27007 20728 27016 20768
rect 27137 20728 27148 20768
rect 27188 20728 27197 20768
rect 27281 20728 27290 20768
rect 27330 20759 27668 20768
rect 27330 20728 27619 20759
rect 17099 20719 17108 20728
rect 17050 20718 17108 20719
rect 17356 20684 17396 20728
rect 17836 20684 17876 20728
rect 10732 20644 11884 20684
rect 11924 20644 11933 20684
rect 12931 20644 12940 20684
rect 12980 20644 13111 20684
rect 13603 20644 13612 20684
rect 13652 20644 13661 20684
rect 14332 20644 14366 20684
rect 14406 20644 14532 20684
rect 14659 20644 14668 20684
rect 14708 20644 14755 20684
rect 14836 20644 15642 20684
rect 15682 20644 15916 20684
rect 15956 20644 15965 20684
rect 16570 20644 16579 20684
rect 16619 20644 16972 20684
rect 17012 20644 17021 20684
rect 17356 20644 17740 20684
rect 17780 20644 17789 20684
rect 17836 20644 18412 20684
rect 18452 20644 18461 20684
rect 10732 20600 10772 20644
rect 14332 20600 14372 20644
rect 14836 20600 14876 20644
rect 9379 20560 9388 20600
rect 9428 20560 10051 20600
rect 10091 20560 10100 20600
rect 10147 20560 10156 20600
rect 10196 20560 10772 20600
rect 10858 20560 10867 20600
rect 10907 20560 10916 20600
rect 11273 20560 11347 20600
rect 11387 20560 11404 20600
rect 11444 20560 11453 20600
rect 13546 20560 13555 20600
rect 13595 20560 13829 20600
rect 13882 20560 13891 20600
rect 13931 20560 13940 20600
rect 14332 20560 14876 20600
rect 15017 20560 15139 20600
rect 15188 20560 15197 20600
rect 15418 20560 15427 20600
rect 15467 20560 15628 20600
rect 15668 20560 15677 20600
rect 15881 20560 15955 20600
rect 15995 20560 16012 20600
rect 16052 20560 16061 20600
rect 17897 20560 18019 20600
rect 18068 20560 18077 20600
rect 18185 20560 18307 20600
rect 18356 20560 18365 20600
rect 18979 20560 18988 20600
rect 19028 20560 19084 20600
rect 19124 20560 19159 20600
rect 10876 20516 10916 20560
rect 931 20476 940 20516
rect 980 20476 2420 20516
rect 7939 20476 7948 20516
rect 7988 20476 8875 20516
rect 9187 20476 9196 20516
rect 9236 20476 10252 20516
rect 10292 20476 10916 20516
rect 13789 20432 13829 20560
rect 13900 20516 13940 20560
rect 19228 20516 19268 20728
rect 19607 20684 19647 20728
rect 19756 20684 19796 20728
rect 19363 20644 19372 20684
rect 19412 20644 19647 20684
rect 19747 20644 19756 20684
rect 19796 20644 19843 20684
rect 19459 20560 19468 20600
rect 19508 20560 20044 20600
rect 20084 20560 20093 20600
rect 20140 20516 20180 20728
rect 24172 20684 24212 20728
rect 24279 20684 24319 20728
rect 25612 20684 25652 20728
rect 26284 20684 26324 20728
rect 26668 20684 26708 20728
rect 20995 20644 21004 20684
rect 21044 20644 23299 20684
rect 23339 20644 23348 20684
rect 24125 20644 24172 20684
rect 24212 20644 24221 20684
rect 24279 20644 25132 20684
rect 25172 20644 26572 20684
rect 26612 20644 26621 20684
rect 26668 20644 27244 20684
rect 27284 20644 27293 20684
rect 20707 20560 20716 20600
rect 20756 20560 20765 20600
rect 22819 20560 22828 20600
rect 22868 20560 23596 20600
rect 23636 20560 23645 20600
rect 24826 20560 24835 20600
rect 24875 20560 25324 20600
rect 25364 20560 25373 20600
rect 25481 20560 25507 20600
rect 25547 20560 25612 20600
rect 25652 20560 25661 20600
rect 25786 20560 25795 20600
rect 25835 20560 25844 20600
rect 26746 20560 26755 20600
rect 26795 20560 26804 20600
rect 26851 20560 26860 20600
rect 26900 20560 27031 20600
rect 13900 20476 16876 20516
rect 16916 20476 16925 20516
rect 18403 20476 18412 20516
rect 18452 20476 20180 20516
rect 20716 20516 20756 20560
rect 25804 20516 25844 20560
rect 20716 20476 23404 20516
rect 23444 20476 23453 20516
rect 25699 20476 25708 20516
rect 25748 20476 25844 20516
rect 26764 20516 26804 20560
rect 27340 20516 27380 20728
rect 27610 20719 27619 20728
rect 27659 20719 27668 20759
rect 27785 20728 27916 20768
rect 27956 20728 27965 20768
rect 28378 20728 28387 20768
rect 28427 20728 28436 20768
rect 28483 20728 28492 20768
rect 28532 20728 28541 20768
rect 28963 20728 28972 20768
rect 29012 20728 29644 20768
rect 29684 20728 29693 20768
rect 30377 20728 30508 20768
rect 30548 20728 30557 20768
rect 30787 20728 30796 20768
rect 30836 20728 30892 20768
rect 30932 20728 30967 20768
rect 31171 20728 31180 20768
rect 31220 20728 31229 20768
rect 27610 20718 27668 20719
rect 28396 20684 28436 20728
rect 27715 20644 27724 20684
rect 27764 20644 28204 20684
rect 28244 20644 28253 20684
rect 28396 20644 28492 20684
rect 28532 20644 30691 20684
rect 30731 20644 30740 20684
rect 30796 20644 31660 20684
rect 31700 20644 31709 20684
rect 27427 20560 27436 20600
rect 27476 20560 28580 20600
rect 28649 20560 28684 20600
rect 28724 20560 28780 20600
rect 28820 20560 28829 20600
rect 26764 20476 26815 20516
rect 27235 20476 27244 20516
rect 27284 20476 27380 20516
rect 28540 20516 28580 20560
rect 30796 20516 30836 20644
rect 28540 20476 30836 20516
rect 30892 20560 30979 20600
rect 31019 20560 31028 20600
rect 4343 20392 4352 20432
rect 4720 20392 4729 20432
rect 8419 20392 8428 20432
rect 8468 20392 11884 20432
rect 11924 20392 11933 20432
rect 12117 20392 12126 20432
rect 12494 20392 12503 20432
rect 13789 20392 14476 20432
rect 14516 20392 14525 20432
rect 18691 20392 18700 20432
rect 18740 20392 18749 20432
rect 1795 20308 1804 20348
rect 1844 20308 3052 20348
rect 3092 20308 6028 20348
rect 6068 20308 6077 20348
rect 9667 20308 9676 20348
rect 9716 20308 11404 20348
rect 11444 20308 11453 20348
rect 12748 20308 13385 20348
rect 0 20264 400 20284
rect 12748 20264 12788 20308
rect 0 20224 980 20264
rect 2563 20224 2572 20264
rect 2612 20224 2668 20264
rect 2708 20224 2743 20264
rect 3113 20224 3235 20264
rect 3284 20224 3293 20264
rect 4684 20224 5164 20264
rect 5204 20224 5213 20264
rect 5347 20224 5356 20264
rect 5396 20224 5527 20264
rect 5827 20224 5836 20264
rect 5876 20224 6211 20264
rect 6251 20224 6260 20264
rect 6307 20224 6316 20264
rect 6356 20224 6604 20264
rect 6644 20224 6653 20264
rect 6787 20224 6796 20264
rect 6836 20224 7372 20264
rect 7412 20224 7421 20264
rect 8524 20224 8764 20264
rect 8804 20224 9908 20264
rect 11657 20224 11692 20264
rect 11732 20224 11788 20264
rect 11828 20224 11837 20264
rect 12547 20224 12556 20264
rect 12596 20224 12748 20264
rect 12835 20224 12844 20264
rect 12884 20224 12931 20264
rect 12971 20224 13015 20264
rect 13123 20224 13132 20264
rect 13172 20224 13303 20264
rect 0 20204 400 20224
rect 940 20180 980 20224
rect 4684 20180 4724 20224
rect 6316 20180 6356 20224
rect 8524 20180 8564 20224
rect 9868 20180 9908 20224
rect 12748 20215 12788 20224
rect 13345 20180 13385 20308
rect 16876 20308 17644 20348
rect 17684 20308 17693 20348
rect 16876 20264 16916 20308
rect 18700 20264 18740 20392
rect 19276 20264 19316 20476
rect 19891 20392 19900 20432
rect 20268 20392 20277 20432
rect 26775 20348 26815 20476
rect 30892 20432 30932 20560
rect 27665 20392 27674 20432
rect 28042 20392 28051 20432
rect 29923 20392 29932 20432
rect 29972 20392 30932 20432
rect 23491 20308 23500 20348
rect 23540 20308 26668 20348
rect 26708 20308 26717 20348
rect 26775 20308 27148 20348
rect 27188 20308 28052 20348
rect 14057 20224 14179 20264
rect 14228 20224 14237 20264
rect 14659 20224 14668 20264
rect 14708 20224 14851 20264
rect 14891 20224 14900 20264
rect 14947 20224 14956 20264
rect 14996 20224 15148 20264
rect 15188 20224 15197 20264
rect 15244 20224 15572 20264
rect 15907 20224 15916 20264
rect 15956 20224 16204 20264
rect 16244 20224 16253 20264
rect 16457 20224 16579 20264
rect 16628 20224 16916 20264
rect 17251 20224 17260 20264
rect 17300 20224 18068 20264
rect 18682 20224 18691 20264
rect 18731 20224 18740 20264
rect 18787 20224 18796 20264
rect 18836 20224 18892 20264
rect 18932 20224 18967 20264
rect 19258 20224 19267 20264
rect 19307 20224 19316 20264
rect 19372 20224 19708 20264
rect 19748 20224 19757 20264
rect 24163 20224 24172 20264
rect 24212 20224 24979 20264
rect 25019 20224 25028 20264
rect 15244 20180 15284 20224
rect 940 20140 4060 20180
rect 4100 20140 4109 20180
rect 4608 20140 4673 20180
rect 4713 20140 4724 20180
rect 4867 20140 4876 20180
rect 4916 20140 4925 20180
rect 5836 20140 6356 20180
rect 6691 20140 6700 20180
rect 6740 20140 6776 20180
rect 7200 20140 7276 20180
rect 7316 20140 7325 20180
rect 7875 20140 8276 20180
rect 4876 20096 4916 20140
rect 5836 20096 5876 20140
rect 6699 20096 6739 20140
rect 7276 20096 7316 20140
rect 7875 20096 7915 20140
rect 8236 20096 8276 20140
rect 8502 20140 8564 20180
rect 8611 20140 8620 20180
rect 8660 20140 9772 20180
rect 9812 20140 9821 20180
rect 9868 20140 12020 20180
rect 8502 20096 8542 20140
rect 9772 20096 9812 20140
rect 1699 20056 1708 20096
rect 1748 20056 1757 20096
rect 1891 20056 1900 20096
rect 1940 20056 2135 20096
rect 2175 20056 2184 20096
rect 2275 20056 2284 20096
rect 2324 20056 2380 20096
rect 2420 20056 2764 20096
rect 2804 20056 2813 20096
rect 2992 20056 3001 20096
rect 3041 20056 3052 20096
rect 3092 20056 3181 20096
rect 3257 20056 3340 20096
rect 3380 20056 3388 20096
rect 3428 20056 3437 20096
rect 3523 20056 3532 20096
rect 3572 20056 3820 20096
rect 3860 20056 3869 20096
rect 4675 20056 4684 20096
rect 4724 20056 4916 20096
rect 4972 20087 5012 20096
rect 0 19844 400 19864
rect 0 19804 460 19844
rect 500 19804 509 19844
rect 809 19804 844 19844
rect 884 19804 931 19844
rect 971 19804 989 19844
rect 0 19784 400 19804
rect 1708 19508 1748 20056
rect 5144 20056 5153 20096
rect 5204 20056 5324 20096
rect 5452 20087 5492 20096
rect 4972 20012 5012 20047
rect 5705 20056 5740 20096
rect 5780 20056 5836 20096
rect 5876 20056 5885 20096
rect 5968 20056 5977 20096
rect 6017 20056 6026 20096
rect 6104 20056 6113 20096
rect 6164 20056 6284 20096
rect 6412 20087 6604 20096
rect 5452 20012 5492 20047
rect 5986 20012 6026 20056
rect 6452 20056 6604 20087
rect 6644 20056 6653 20096
rect 6699 20056 6709 20096
rect 6749 20056 6758 20096
rect 6883 20056 6892 20096
rect 6971 20056 7084 20096
rect 7124 20056 7133 20096
rect 7217 20056 7226 20096
rect 7266 20056 7316 20096
rect 7363 20056 7372 20096
rect 7412 20056 7756 20096
rect 7796 20056 7915 20096
rect 8009 20087 8140 20096
rect 8009 20056 8131 20087
rect 8180 20056 8189 20096
rect 8236 20056 8542 20096
rect 8585 20087 8716 20096
rect 8585 20056 8611 20087
rect 6412 20038 6452 20047
rect 8122 20047 8131 20056
rect 8171 20047 8180 20056
rect 8122 20046 8180 20047
rect 8602 20047 8611 20056
rect 8651 20056 8716 20087
rect 8756 20056 8765 20096
rect 9257 20056 9388 20096
rect 9428 20056 9437 20096
rect 9754 20056 9763 20096
rect 9803 20056 9812 20096
rect 8651 20047 8660 20056
rect 8602 20046 8660 20047
rect 2266 19972 2275 20012
rect 2315 19972 2324 20012
rect 2467 19972 2476 20012
rect 2516 19972 2525 20012
rect 2890 20003 3860 20012
rect 2284 19508 2324 19972
rect 2476 19760 2516 19972
rect 2890 19963 2899 20003
rect 2939 19972 3860 20003
rect 3907 19972 3916 20012
rect 3956 19972 3965 20012
rect 4169 19972 4300 20012
rect 4340 19972 4349 20012
rect 4972 19972 5260 20012
rect 5300 19972 5309 20012
rect 5452 19972 5644 20012
rect 5684 19972 5693 20012
rect 5866 20003 5924 20012
rect 2939 19963 2948 19972
rect 2890 19962 2948 19963
rect 3820 19844 3860 19972
rect 3916 19928 3956 19972
rect 5866 19963 5875 20003
rect 5915 19963 5924 20003
rect 5986 19972 6028 20012
rect 6068 19972 6077 20012
rect 6826 20003 6884 20012
rect 5866 19962 5924 19963
rect 6826 19963 6835 20003
rect 6875 19963 6884 20003
rect 8275 19972 8284 20012
rect 8324 19972 8333 20012
rect 6826 19962 6884 19963
rect 5884 19928 5924 19962
rect 6844 19928 6884 19962
rect 8284 19928 8324 19972
rect 3916 19888 4724 19928
rect 5884 19888 6604 19928
rect 6644 19888 6653 19928
rect 6844 19888 8084 19928
rect 8131 19888 8140 19928
rect 8180 19888 8324 19928
rect 11020 19928 11060 19992
rect 11980 19928 12020 20140
rect 13324 20140 13385 20180
rect 13673 20140 13795 20180
rect 13844 20140 13853 20180
rect 15148 20140 15284 20180
rect 15532 20180 15572 20224
rect 18028 20180 18068 20224
rect 19372 20180 19412 20224
rect 15532 20140 15764 20180
rect 16675 20140 16684 20180
rect 16724 20140 16771 20180
rect 17033 20140 17164 20180
rect 17204 20140 17213 20180
rect 17356 20140 17847 20180
rect 17887 20140 17896 20180
rect 18028 20140 18644 20180
rect 19296 20140 19372 20180
rect 19412 20140 19421 20180
rect 20602 20140 20611 20180
rect 20651 20140 20660 20180
rect 20803 20140 20812 20180
rect 20852 20140 22580 20180
rect 24617 20140 24748 20180
rect 24788 20140 24797 20180
rect 13324 20096 13364 20140
rect 15148 20096 15188 20140
rect 15724 20096 15764 20140
rect 16684 20096 16724 20140
rect 17356 20096 17396 20140
rect 18604 20096 18644 20140
rect 19372 20096 19412 20140
rect 20620 20096 20660 20140
rect 22540 20096 22580 20140
rect 25756 20096 25796 20308
rect 28012 20264 28052 20308
rect 26563 20224 26572 20264
rect 26612 20224 26996 20264
rect 28003 20224 28012 20264
rect 28052 20224 28061 20264
rect 28841 20224 28972 20264
rect 29012 20224 29021 20264
rect 25891 20140 25900 20180
rect 25940 20140 26668 20180
rect 26708 20140 26717 20180
rect 26956 20096 26996 20224
rect 27811 20140 27820 20180
rect 27860 20140 28108 20180
rect 28148 20140 28157 20180
rect 28771 20140 28780 20180
rect 28820 20140 29548 20180
rect 29588 20140 29597 20180
rect 29923 20140 29932 20180
rect 29972 20140 31267 20180
rect 31307 20140 31316 20180
rect 12346 20056 12355 20096
rect 12395 20056 12844 20096
rect 12884 20056 12893 20096
rect 13306 20056 13315 20096
rect 13355 20056 13364 20096
rect 13699 20056 13708 20096
rect 13748 20056 13757 20096
rect 13891 20056 13900 20096
rect 13940 20056 14071 20096
rect 14153 20056 14284 20096
rect 14324 20056 14333 20096
rect 14380 20056 14750 20096
rect 14790 20056 14799 20096
rect 15052 20087 15188 20096
rect 13708 20012 13748 20056
rect 14380 20012 14420 20056
rect 15092 20056 15188 20087
rect 15244 20056 15340 20096
rect 15380 20056 15389 20096
rect 15520 20093 15532 20096
rect 15052 20012 15092 20047
rect 15244 20012 15284 20056
rect 15499 20031 15532 20093
rect 15572 20056 15630 20096
rect 15715 20056 15724 20096
rect 15764 20056 15773 20096
rect 15907 20056 15916 20096
rect 15956 20056 15965 20096
rect 16099 20056 16108 20096
rect 16148 20056 16157 20096
rect 16204 20056 16300 20096
rect 16340 20056 16349 20096
rect 16675 20056 16684 20096
rect 16724 20056 16733 20096
rect 17050 20056 17059 20096
rect 17099 20056 17108 20096
rect 15572 20031 15581 20056
rect 12538 19972 12547 20012
rect 12587 19972 12748 20012
rect 12788 19972 12797 20012
rect 13324 19972 13748 20012
rect 14371 19972 14380 20012
rect 14420 19972 14551 20012
rect 14659 19972 14668 20012
rect 14708 19972 15092 20012
rect 15235 19972 15244 20012
rect 15284 19972 15293 20012
rect 13324 19928 13364 19972
rect 14380 19928 14420 19972
rect 15916 19928 15956 20056
rect 11020 19888 11884 19928
rect 11924 19888 11933 19928
rect 11980 19888 13324 19928
rect 13364 19888 13373 19928
rect 13507 19888 13516 19928
rect 13556 19888 14420 19928
rect 14467 19888 14476 19928
rect 14516 19888 15956 19928
rect 16108 19928 16148 20056
rect 16204 20012 16244 20056
rect 17068 20012 17108 20056
rect 17260 20056 17367 20096
rect 17407 20056 17416 20096
rect 17530 20056 17539 20096
rect 17579 20056 17588 20096
rect 17635 20056 17644 20096
rect 17684 20056 17693 20096
rect 18106 20056 18115 20096
rect 18155 20056 18164 20096
rect 18211 20056 18220 20096
rect 18260 20056 18356 20096
rect 17260 20012 17300 20056
rect 17548 20012 17588 20056
rect 16195 19972 16204 20012
rect 16244 19972 16253 20012
rect 16771 19972 16780 20012
rect 16820 19972 17108 20012
rect 17251 19972 17260 20012
rect 17300 19972 17309 20012
rect 17443 19972 17452 20012
rect 17492 19972 17588 20012
rect 17644 19928 17684 20056
rect 18124 20012 18164 20056
rect 16108 19888 16492 19928
rect 16532 19888 16541 19928
rect 17155 19888 17164 19928
rect 17204 19888 17684 19928
rect 17836 19972 18164 20012
rect 4684 19844 4724 19888
rect 8044 19844 8084 19888
rect 14476 19844 14516 19888
rect 17836 19844 17876 19972
rect 2563 19804 2572 19844
rect 2612 19804 3676 19844
rect 3716 19804 3725 19844
rect 3820 19804 4396 19844
rect 4436 19804 4445 19844
rect 4666 19804 4675 19844
rect 4715 19804 4724 19844
rect 5059 19804 5068 19844
rect 5108 19804 5155 19844
rect 5195 19804 5239 19844
rect 7459 19804 7468 19844
rect 7508 19804 7852 19844
rect 7892 19804 7901 19844
rect 8044 19804 13036 19844
rect 13076 19804 13085 19844
rect 13891 19804 13900 19844
rect 13940 19804 14516 19844
rect 14851 19804 14860 19844
rect 14900 19804 15436 19844
rect 15476 19804 15485 19844
rect 15715 19804 15724 19844
rect 15764 19804 15916 19844
rect 15956 19804 15965 19844
rect 16867 19804 16876 19844
rect 16916 19804 17644 19844
rect 17684 19804 17693 19844
rect 17827 19804 17836 19844
rect 17876 19804 17885 19844
rect 18316 19760 18356 20056
rect 18412 20056 18423 20096
rect 18463 20056 18472 20096
rect 18586 20056 18595 20096
rect 18635 20056 18644 20096
rect 18700 20056 18903 20096
rect 18943 20056 18952 20096
rect 19075 20056 19084 20096
rect 19124 20056 19171 20096
rect 19267 20056 19276 20096
rect 19316 20056 19412 20096
rect 19519 20056 19528 20096
rect 19604 20056 19708 20096
rect 20218 20056 20227 20096
rect 20267 20056 20276 20096
rect 20620 20056 22156 20096
rect 22196 20056 22205 20096
rect 22522 20056 22531 20096
rect 22571 20056 22580 20096
rect 23395 20056 23404 20096
rect 23444 20056 23453 20096
rect 23524 20056 23533 20096
rect 23573 20056 23596 20096
rect 23636 20056 23713 20096
rect 23779 20056 23788 20096
rect 23828 20056 23837 20096
rect 24442 20056 24451 20096
rect 24491 20056 24652 20096
rect 24692 20056 24701 20096
rect 25001 20056 25123 20096
rect 25172 20056 25181 20096
rect 25228 20087 25324 20096
rect 18412 20012 18452 20056
rect 18700 20012 18740 20056
rect 19084 20012 19124 20056
rect 20236 20012 20276 20056
rect 18412 19972 18508 20012
rect 18548 19972 18740 20012
rect 19075 19972 19084 20012
rect 19124 19972 19133 20012
rect 19363 19972 19372 20012
rect 19412 19972 21236 20012
rect 21859 19972 21868 20012
rect 21908 19972 21917 20012
rect 22906 19972 22915 20012
rect 22955 19972 23060 20012
rect 18412 19888 19180 19928
rect 19220 19888 19229 19928
rect 19651 19888 19660 19928
rect 19700 19888 20272 19928
rect 20312 19888 21140 19928
rect 18412 19844 18452 19888
rect 18403 19804 18412 19844
rect 18452 19804 18461 19844
rect 18595 19804 18604 19844
rect 18644 19804 20044 19844
rect 20084 19804 20093 19844
rect 20995 19804 21004 19844
rect 21044 19804 21053 19844
rect 2476 19720 2956 19760
rect 2996 19720 3005 19760
rect 6211 19720 6220 19760
rect 6260 19720 11692 19760
rect 11732 19720 11741 19760
rect 14371 19720 14380 19760
rect 14420 19720 17260 19760
rect 17300 19720 17309 19760
rect 18316 19720 18452 19760
rect 18499 19720 18508 19760
rect 18548 19720 20812 19760
rect 20852 19720 20861 19760
rect 3103 19636 3112 19676
rect 3480 19636 3489 19676
rect 7084 19636 10156 19676
rect 10196 19636 10205 19676
rect 10877 19636 10886 19676
rect 11254 19636 11263 19676
rect 11491 19636 11500 19676
rect 11540 19636 17972 19676
rect 1708 19468 2179 19508
rect 2219 19468 2228 19508
rect 2284 19468 3724 19508
rect 3764 19468 3773 19508
rect 4265 19468 4387 19508
rect 4436 19468 4445 19508
rect 5914 19468 5923 19508
rect 5963 19468 5972 19508
rect 6595 19468 6604 19508
rect 6644 19468 6883 19508
rect 6923 19468 6932 19508
rect 0 19424 400 19444
rect 0 19384 652 19424
rect 692 19384 701 19424
rect 1603 19384 1612 19424
rect 1652 19384 3628 19424
rect 3668 19384 3677 19424
rect 5548 19384 5836 19424
rect 5876 19384 5885 19424
rect 0 19364 400 19384
rect 809 19300 844 19340
rect 884 19300 940 19340
rect 980 19300 989 19340
rect 1804 19300 2188 19340
rect 2228 19300 2237 19340
rect 2956 19300 3724 19340
rect 3764 19300 3773 19340
rect 4012 19300 4588 19340
rect 4628 19300 4637 19340
rect 5251 19300 5260 19340
rect 5300 19300 5452 19340
rect 5492 19300 5501 19340
rect 1804 19256 1844 19300
rect 2476 19256 2516 19265
rect 2956 19256 2996 19300
rect 4012 19256 4052 19300
rect 4684 19256 4724 19265
rect 5548 19256 5588 19384
rect 5932 19340 5972 19468
rect 7084 19340 7124 19636
rect 7171 19552 7180 19592
rect 7220 19552 11060 19592
rect 11020 19508 11060 19552
rect 9571 19468 9580 19508
rect 9620 19468 10732 19508
rect 10772 19468 10781 19508
rect 11002 19468 11011 19508
rect 11051 19468 11060 19508
rect 13411 19468 13420 19508
rect 13460 19468 13468 19508
rect 13508 19468 13591 19508
rect 14441 19468 14572 19508
rect 14612 19468 14621 19508
rect 15139 19468 15148 19508
rect 15188 19468 16492 19508
rect 16532 19468 16541 19508
rect 5658 19300 5667 19340
rect 5707 19300 5972 19340
rect 6211 19300 6220 19340
rect 6260 19300 6307 19340
rect 6691 19300 6700 19340
rect 6740 19300 7124 19340
rect 7180 19384 12652 19424
rect 12692 19384 12701 19424
rect 12809 19384 12940 19424
rect 12980 19384 12989 19424
rect 6220 19256 6260 19300
rect 7180 19289 7220 19384
rect 7651 19300 7660 19340
rect 7700 19300 7756 19340
rect 7796 19300 7831 19340
rect 8098 19300 9196 19340
rect 9236 19300 9245 19340
rect 9484 19300 9772 19340
rect 9812 19300 9821 19340
rect 10435 19300 10444 19340
rect 10484 19300 10636 19340
rect 10676 19300 10685 19340
rect 12739 19300 12748 19340
rect 12788 19300 12980 19340
rect 13097 19300 13228 19340
rect 13268 19300 13277 19340
rect 14092 19300 14668 19340
rect 14708 19300 14717 19340
rect 15139 19300 15148 19340
rect 15188 19300 15764 19340
rect 15808 19300 15916 19340
rect 15979 19300 15988 19340
rect 1795 19216 1804 19256
rect 1844 19216 1853 19256
rect 1987 19216 1996 19256
rect 2036 19216 2045 19256
rect 2168 19216 2177 19256
rect 2217 19216 2380 19256
rect 2420 19216 2429 19256
rect 2516 19216 2764 19256
rect 2804 19216 2813 19256
rect 2938 19216 2947 19256
rect 2987 19216 2996 19256
rect 3043 19216 3052 19256
rect 3092 19216 3223 19256
rect 3418 19216 3427 19256
rect 3467 19216 3532 19256
rect 3572 19216 3607 19256
rect 3689 19216 3738 19256
rect 3778 19216 3820 19256
rect 3860 19216 3869 19256
rect 4003 19216 4012 19256
rect 4052 19216 4061 19256
rect 4108 19216 4131 19256
rect 4171 19216 4180 19256
rect 4240 19216 4249 19256
rect 4289 19216 4300 19256
rect 4340 19216 4382 19256
rect 4422 19216 4500 19256
rect 4937 19216 5068 19256
rect 5108 19216 5117 19256
rect 5251 19216 5260 19256
rect 5300 19216 5309 19256
rect 5539 19216 5548 19256
rect 5588 19216 5597 19256
rect 5776 19216 5785 19256
rect 5825 19216 5856 19256
rect 5912 19216 5921 19256
rect 5961 19216 6124 19256
rect 6164 19216 6173 19256
rect 6350 19216 6359 19256
rect 6399 19216 6408 19256
rect 6490 19216 6499 19256
rect 6539 19216 6548 19256
rect 6595 19216 6604 19256
rect 6644 19216 6775 19256
rect 6872 19216 6881 19256
rect 6932 19216 7052 19256
rect 7169 19249 7178 19289
rect 7218 19249 7227 19289
rect 8098 19256 8138 19300
rect 9484 19298 9524 19300
rect 9304 19289 9524 19298
rect 7721 19216 7756 19256
rect 7796 19216 7852 19256
rect 7892 19216 7901 19256
rect 7948 19216 7971 19256
rect 8011 19216 8020 19256
rect 8080 19216 8089 19256
rect 8129 19216 8138 19256
rect 8707 19216 8716 19256
rect 8756 19216 8765 19256
rect 8899 19216 8908 19256
rect 8948 19216 9004 19256
rect 9044 19216 9079 19256
rect 9178 19216 9187 19256
rect 9227 19216 9236 19256
rect 9344 19258 9524 19289
rect 11308 19256 11348 19265
rect 12940 19256 12980 19300
rect 14092 19256 14132 19300
rect 15724 19256 15764 19300
rect 16035 19298 16075 19468
rect 16035 19258 16060 19298
rect 16100 19258 16109 19298
rect 16492 19256 16532 19468
rect 17932 19424 17972 19636
rect 18412 19508 18452 19720
rect 18651 19636 18660 19676
rect 19028 19636 19037 19676
rect 18403 19468 18412 19508
rect 18452 19468 18461 19508
rect 19433 19468 19459 19508
rect 19499 19468 19564 19508
rect 19604 19468 19613 19508
rect 21004 19424 21044 19804
rect 21100 19760 21140 19888
rect 21196 19844 21236 19972
rect 23020 19928 23060 19972
rect 23020 19888 23116 19928
rect 23156 19888 23165 19928
rect 21196 19804 22828 19844
rect 22868 19804 22877 19844
rect 21100 19720 23020 19760
rect 23060 19720 23069 19760
rect 22627 19552 22636 19592
rect 22676 19552 23308 19592
rect 23348 19552 23357 19592
rect 23404 19508 23444 20056
rect 22435 19468 22444 19508
rect 22484 19468 22493 19508
rect 23107 19468 23116 19508
rect 23156 19468 23444 19508
rect 22444 19424 22484 19468
rect 23788 19424 23828 20056
rect 25268 20056 25324 20087
rect 25364 20056 25399 20096
rect 25507 20056 25516 20096
rect 25556 20056 25996 20096
rect 26036 20056 26045 20096
rect 26224 20056 26233 20096
rect 26273 20056 26572 20096
rect 26612 20056 26621 20096
rect 26701 20056 26710 20096
rect 26750 20056 26860 20096
rect 26900 20056 26909 20096
rect 26956 20056 27137 20096
rect 27177 20056 27186 20096
rect 27235 20056 27244 20096
rect 27284 20056 27532 20096
rect 27572 20056 27619 20096
rect 27659 20056 27703 20096
rect 27903 20056 27912 20096
rect 27952 20056 28052 20096
rect 28147 20056 28156 20096
rect 28196 20056 28244 20096
rect 29443 20056 29452 20096
rect 29492 20056 30883 20096
rect 30923 20056 30932 20096
rect 25228 20038 25268 20047
rect 28012 20012 28052 20056
rect 24259 19972 24268 20012
rect 24308 19972 24317 20012
rect 24713 19972 24748 20012
rect 24788 19972 24844 20012
rect 24884 19972 24893 20012
rect 25795 19972 25804 20012
rect 25844 19972 26115 20012
rect 26155 19972 26164 20012
rect 26506 19972 26515 20012
rect 26555 19972 26956 20012
rect 26996 19972 27244 20012
rect 27284 19972 27293 20012
rect 28012 19972 28108 20012
rect 28148 19972 28157 20012
rect 24268 19928 24308 19972
rect 28204 19928 28244 20056
rect 31104 19972 31372 20012
rect 31412 19972 31421 20012
rect 24268 19888 25132 19928
rect 25172 19888 25181 19928
rect 26371 19888 26380 19928
rect 26420 19888 26900 19928
rect 27139 19888 27148 19928
rect 27188 19888 28244 19928
rect 25507 19804 25516 19844
rect 25556 19804 25565 19844
rect 17932 19384 21044 19424
rect 21388 19384 22348 19424
rect 22388 19384 22397 19424
rect 22444 19384 23828 19424
rect 21388 19340 21428 19384
rect 25516 19340 25556 19804
rect 26860 19760 26900 19888
rect 27235 19804 27244 19844
rect 27284 19804 27293 19844
rect 27619 19804 27628 19844
rect 27668 19804 29644 19844
rect 29684 19804 29693 19844
rect 26851 19720 26860 19760
rect 26900 19720 26909 19760
rect 26425 19636 26434 19676
rect 26802 19636 26811 19676
rect 27052 19384 27148 19424
rect 27188 19384 27197 19424
rect 27052 19340 27092 19384
rect 27244 19340 27284 19804
rect 27715 19552 27724 19592
rect 27764 19552 30316 19592
rect 30356 19552 30365 19592
rect 27532 19468 28204 19508
rect 28244 19468 28492 19508
rect 28532 19468 28541 19508
rect 30499 19468 30508 19508
rect 30548 19468 31276 19508
rect 31316 19468 31325 19508
rect 17164 19300 17452 19340
rect 17492 19300 17501 19340
rect 18316 19300 18700 19340
rect 18740 19300 18749 19340
rect 19738 19300 19747 19340
rect 19787 19300 20140 19340
rect 20180 19300 20716 19340
rect 20756 19300 20765 19340
rect 21004 19300 21428 19340
rect 21484 19300 21868 19340
rect 21908 19300 23116 19340
rect 23156 19300 23165 19340
rect 23308 19300 24047 19340
rect 24087 19300 24556 19340
rect 24596 19300 24605 19340
rect 25516 19300 26036 19340
rect 26441 19300 26572 19340
rect 26612 19300 26621 19340
rect 27043 19300 27052 19340
rect 27092 19300 27101 19340
rect 27244 19300 27267 19340
rect 27307 19300 27316 19340
rect 17164 19256 17204 19300
rect 18316 19298 18356 19300
rect 18136 19289 18356 19298
rect 9304 19240 9344 19249
rect 9737 19216 9772 19256
rect 9812 19216 9868 19256
rect 9908 19216 9917 19256
rect 9964 19216 9987 19256
rect 10027 19216 10036 19256
rect 10090 19216 10099 19256
rect 10139 19216 10156 19256
rect 10196 19216 10270 19256
rect 11177 19216 11308 19256
rect 11348 19216 11357 19256
rect 11657 19216 11680 19256
rect 11720 19216 11788 19256
rect 11828 19216 11837 19256
rect 12547 19216 12556 19256
rect 12596 19247 12727 19256
rect 12596 19216 12643 19247
rect 595 19048 604 19088
rect 644 19048 652 19088
rect 692 19048 775 19088
rect 1795 19048 1804 19088
rect 1844 19048 1853 19088
rect 1804 18920 1844 19048
rect 1996 19004 2036 19216
rect 2476 19207 2516 19216
rect 3249 19132 3258 19172
rect 3298 19132 3628 19172
rect 3668 19132 3677 19172
rect 3820 19132 4012 19172
rect 4052 19132 4061 19172
rect 3820 19088 3860 19132
rect 2371 19048 2380 19088
rect 2420 19048 2572 19088
rect 2612 19048 2621 19088
rect 3139 19048 3148 19088
rect 3188 19048 3319 19088
rect 3514 19048 3523 19088
rect 3563 19048 3860 19088
rect 3907 19048 3916 19088
rect 3956 19048 3965 19088
rect 3916 19004 3956 19048
rect 1996 18964 3956 19004
rect 1804 18880 3436 18920
rect 3476 18880 3485 18920
rect 4108 18836 4148 19216
rect 4684 19172 4724 19216
rect 5260 19172 5300 19216
rect 5816 19172 5856 19216
rect 6220 19207 6260 19216
rect 6359 19172 6399 19216
rect 6508 19172 6548 19216
rect 7948 19172 7988 19216
rect 4684 19132 5164 19172
rect 5204 19132 5213 19172
rect 5260 19132 5548 19172
rect 5588 19132 5597 19172
rect 5816 19132 6028 19172
rect 6068 19132 6077 19172
rect 6307 19132 6316 19172
rect 6356 19132 6399 19172
rect 6499 19132 6508 19172
rect 6548 19132 7220 19172
rect 7267 19132 7276 19172
rect 7316 19132 7988 19172
rect 7180 19088 7220 19132
rect 8098 19088 8138 19216
rect 8716 19172 8756 19216
rect 8716 19132 8908 19172
rect 8948 19132 8957 19172
rect 9196 19088 9236 19216
rect 9964 19172 10004 19216
rect 11308 19207 11348 19216
rect 12634 19207 12643 19216
rect 12683 19216 12727 19247
rect 12931 19216 12940 19256
rect 12980 19216 12989 19256
rect 13790 19216 13900 19256
rect 13952 19216 13970 19256
rect 14074 19216 14083 19256
rect 14132 19216 14263 19256
rect 14345 19216 14394 19256
rect 14434 19216 14476 19256
rect 14516 19216 14525 19256
rect 14633 19216 14764 19256
rect 14804 19216 14813 19256
rect 14860 19216 14883 19256
rect 14923 19216 14932 19256
rect 15043 19216 15052 19256
rect 15092 19216 15101 19256
rect 15148 19216 15191 19256
rect 15231 19216 15240 19256
rect 15322 19216 15331 19256
rect 15371 19216 15380 19256
rect 15427 19216 15436 19256
rect 15476 19216 15607 19256
rect 15724 19216 15820 19256
rect 15860 19216 15869 19256
rect 16195 19216 16204 19256
rect 16244 19216 16300 19256
rect 16340 19216 16375 19256
rect 16492 19216 16972 19256
rect 17024 19216 17033 19256
rect 17155 19216 17164 19256
rect 17204 19216 17213 19256
rect 17294 19216 17303 19256
rect 17343 19216 17352 19256
rect 17827 19216 17836 19256
rect 17876 19216 18019 19256
rect 18059 19216 18068 19256
rect 18176 19258 18356 19289
rect 21004 19256 21044 19300
rect 21484 19256 21524 19300
rect 23308 19256 23348 19300
rect 25516 19256 25556 19300
rect 25996 19256 26036 19300
rect 27532 19256 27572 19468
rect 27628 19384 28876 19424
rect 28916 19384 28925 19424
rect 27628 19256 27668 19384
rect 27811 19300 27820 19340
rect 27860 19300 28204 19340
rect 28244 19300 28253 19340
rect 30595 19300 30604 19340
rect 30644 19300 30653 19340
rect 27820 19256 27860 19300
rect 18136 19240 18176 19249
rect 18473 19216 18604 19256
rect 18644 19216 18653 19256
rect 18787 19216 18796 19256
rect 18836 19216 18845 19256
rect 19145 19216 19276 19256
rect 19316 19216 19325 19256
rect 19436 19216 19445 19256
rect 19485 19216 19494 19256
rect 19561 19216 19570 19256
rect 19647 19216 19741 19256
rect 19843 19216 19852 19256
rect 19892 19216 19901 19256
rect 20394 19216 20403 19256
rect 20443 19216 20671 19256
rect 20794 19216 20803 19256
rect 20843 19216 20852 19256
rect 20986 19216 20995 19256
rect 21035 19216 21044 19256
rect 21161 19216 21292 19256
rect 21332 19216 21341 19256
rect 21475 19216 21484 19256
rect 21524 19216 21533 19256
rect 21641 19216 21772 19256
rect 21812 19216 21821 19256
rect 21955 19216 21964 19256
rect 22004 19216 22013 19256
rect 22138 19216 22147 19256
rect 22196 19216 22327 19256
rect 22505 19216 22627 19256
rect 22676 19216 22685 19256
rect 22793 19216 22924 19256
rect 22964 19216 23116 19256
rect 23156 19216 23165 19256
rect 23232 19216 23241 19256
rect 23281 19216 23348 19256
rect 23395 19216 23404 19256
rect 23444 19216 23575 19256
rect 23849 19216 23945 19256
rect 24020 19216 24029 19256
rect 24154 19216 24163 19256
rect 24203 19216 24212 19256
rect 24259 19216 24268 19256
rect 24308 19216 24364 19256
rect 24404 19216 24439 19256
rect 24643 19216 24652 19256
rect 24692 19216 24701 19256
rect 24826 19216 24835 19256
rect 24884 19216 25015 19256
rect 25315 19216 25324 19256
rect 25364 19216 25556 19256
rect 25603 19216 25612 19256
rect 25652 19216 25783 19256
rect 25987 19216 25996 19256
rect 26036 19216 26045 19256
rect 26371 19216 26380 19256
rect 26420 19216 26659 19256
rect 26699 19216 26708 19256
rect 27017 19216 27148 19256
rect 27188 19216 27197 19256
rect 27376 19216 27385 19256
rect 27425 19216 27572 19256
rect 27615 19216 27624 19256
rect 27664 19216 27673 19256
rect 27811 19216 27820 19256
rect 27860 19216 27869 19256
rect 28099 19216 28108 19256
rect 28148 19216 28396 19256
rect 28436 19216 28445 19256
rect 29321 19216 29347 19256
rect 29387 19216 29452 19256
rect 29492 19216 29501 19256
rect 12683 19207 12692 19216
rect 12634 19206 12692 19207
rect 12652 19172 12692 19206
rect 14860 19172 14900 19216
rect 9379 19132 9388 19172
rect 9428 19132 10004 19172
rect 10723 19132 10732 19172
rect 10772 19132 11006 19172
rect 11046 19132 11055 19172
rect 12652 19132 13708 19172
rect 13748 19132 13757 19172
rect 14836 19132 14860 19172
rect 14900 19132 14909 19172
rect 15051 19088 15091 19216
rect 4291 19048 4300 19088
rect 4340 19048 4588 19088
rect 4628 19048 5012 19088
rect 5242 19048 5251 19088
rect 5291 19048 5300 19088
rect 6115 19048 6124 19088
rect 6164 19048 6988 19088
rect 7028 19048 7084 19088
rect 7124 19048 7133 19088
rect 7180 19048 8138 19088
rect 8585 19048 8716 19088
rect 8756 19048 8765 19088
rect 8860 19048 9043 19088
rect 9083 19048 9092 19088
rect 9196 19048 9964 19088
rect 10004 19048 10204 19088
rect 10244 19048 10253 19088
rect 11203 19048 11212 19088
rect 11252 19048 11261 19088
rect 11827 19048 11836 19088
rect 11876 19048 11980 19088
rect 12020 19048 12029 19088
rect 13738 19048 13747 19088
rect 13787 19048 13796 19088
rect 13891 19048 13900 19088
rect 13940 19048 14179 19088
rect 14219 19048 14228 19088
rect 14275 19048 14284 19088
rect 14324 19048 15091 19088
rect 4972 18920 5012 19048
rect 5260 19004 5300 19048
rect 5260 18964 6412 19004
rect 6452 18964 6461 19004
rect 6508 18920 6548 19048
rect 8860 19004 8900 19048
rect 11212 19004 11252 19048
rect 13756 19004 13796 19048
rect 15148 19004 15188 19216
rect 15340 19172 15380 19216
rect 17303 19172 17343 19216
rect 18796 19172 18836 19216
rect 15235 19132 15244 19172
rect 15284 19132 15380 19172
rect 15514 19132 15523 19172
rect 15563 19132 15956 19172
rect 16483 19132 16492 19172
rect 16532 19132 17343 19172
rect 17452 19132 18836 19172
rect 19445 19172 19485 19216
rect 19852 19172 19892 19216
rect 20631 19172 20671 19216
rect 20812 19172 20852 19216
rect 21964 19172 22004 19216
rect 23404 19172 23444 19216
rect 24172 19172 24212 19216
rect 19445 19132 19660 19172
rect 19700 19132 19709 19172
rect 19852 19132 20332 19172
rect 20372 19132 20381 19172
rect 20631 19132 20716 19172
rect 20756 19132 20765 19172
rect 20812 19132 21388 19172
rect 21428 19132 21437 19172
rect 21964 19132 22252 19172
rect 22292 19132 22301 19172
rect 22449 19132 22458 19172
rect 22498 19132 23060 19172
rect 23404 19132 24500 19172
rect 4343 18880 4352 18920
rect 4720 18880 4729 18920
rect 4972 18880 6548 18920
rect 8620 18964 8900 19004
rect 9187 18964 9196 19004
rect 9236 18964 10156 19004
rect 10196 18964 10205 19004
rect 11212 18964 13516 19004
rect 13556 18964 13565 19004
rect 13756 18964 14476 19004
rect 14516 18964 14525 19004
rect 15051 18964 15188 19004
rect 15436 19048 15724 19088
rect 15764 19048 15773 19088
rect 4108 18796 8524 18836
rect 8564 18796 8573 18836
rect 8620 18752 8660 18964
rect 15051 18920 15091 18964
rect 15436 18920 15476 19048
rect 8899 18880 8908 18920
rect 8948 18880 9572 18920
rect 12117 18880 12126 18920
rect 12494 18880 12503 18920
rect 13891 18880 13900 18920
rect 13940 18880 15091 18920
rect 15139 18880 15148 18920
rect 15188 18880 15476 18920
rect 9196 18796 9388 18836
rect 9428 18796 9437 18836
rect 9196 18752 9236 18796
rect 9532 18752 9572 18880
rect 15916 18836 15956 19132
rect 17452 19088 17492 19132
rect 23020 19088 23060 19132
rect 16003 19048 16012 19088
rect 16052 19048 16195 19088
rect 16235 19048 16244 19088
rect 16300 19048 16819 19088
rect 16859 19048 17164 19088
rect 17204 19048 17213 19088
rect 17443 19048 17452 19088
rect 17492 19048 17501 19088
rect 17914 19079 18028 19088
rect 14476 18796 15244 18836
rect 15284 18796 15293 18836
rect 15916 18796 16204 18836
rect 16244 18796 16253 18836
rect 739 18712 748 18752
rect 788 18712 3628 18752
rect 3668 18712 3677 18752
rect 5059 18712 5068 18752
rect 5108 18712 5260 18752
rect 5300 18712 5309 18752
rect 6490 18712 6499 18752
rect 6539 18712 6604 18752
rect 6644 18712 6679 18752
rect 6761 18712 6883 18752
rect 6932 18712 6941 18752
rect 7625 18712 7651 18752
rect 7691 18712 7756 18752
rect 7796 18712 7805 18752
rect 8122 18712 8131 18752
rect 8171 18712 8660 18752
rect 9178 18712 9187 18752
rect 9227 18712 9236 18752
rect 9514 18712 9523 18752
rect 9563 18712 9572 18752
rect 10723 18712 10732 18752
rect 10772 18712 11308 18752
rect 11348 18712 11357 18752
rect 11875 18712 11884 18752
rect 11924 18712 12163 18752
rect 12203 18712 12556 18752
rect 12596 18712 12605 18752
rect 13673 18712 13708 18752
rect 13748 18712 13795 18752
rect 13835 18712 13853 18752
rect 13965 18712 14188 18752
rect 14228 18712 14237 18752
rect 13965 18668 14005 18712
rect 2668 18628 8620 18668
rect 8660 18628 8669 18668
rect 8716 18628 8908 18668
rect 8948 18628 8957 18668
rect 9004 18628 9676 18668
rect 9716 18628 9725 18668
rect 10339 18628 10348 18668
rect 10388 18628 10436 18668
rect 10531 18628 10540 18668
rect 10580 18628 10636 18668
rect 10676 18628 10711 18668
rect 10833 18628 10842 18668
rect 10882 18628 11020 18668
rect 11060 18628 11069 18668
rect 11116 18628 11540 18668
rect 2668 18584 2708 18628
rect 8716 18584 8756 18628
rect 9004 18584 9044 18628
rect 2650 18544 2659 18584
rect 2699 18544 2708 18584
rect 3139 18544 3148 18584
rect 3188 18544 3916 18584
rect 3956 18544 3965 18584
rect 4073 18544 4108 18584
rect 4148 18544 4204 18584
rect 4244 18544 4253 18584
rect 4432 18544 4441 18584
rect 4481 18544 4684 18584
rect 4724 18544 4733 18584
rect 4841 18544 4972 18584
rect 5012 18544 5021 18584
rect 5098 18544 5107 18584
rect 5147 18544 5156 18584
rect 5443 18544 5452 18584
rect 5492 18544 5740 18584
rect 5780 18544 5789 18584
rect 5836 18544 5923 18584
rect 5963 18544 5972 18584
rect 6026 18544 6124 18584
rect 6188 18544 6206 18584
rect 6298 18544 6307 18584
rect 6347 18544 6356 18584
rect 6415 18544 6424 18584
rect 6464 18544 6499 18584
rect 5116 18500 5156 18544
rect 5836 18500 5876 18544
rect 6316 18500 6356 18544
rect 6424 18500 6464 18544
rect 6582 18533 6591 18573
rect 6631 18533 6640 18573
rect 6682 18544 6691 18584
rect 6740 18544 6871 18584
rect 6979 18544 6988 18584
rect 7028 18544 7180 18584
rect 7220 18544 7229 18584
rect 7517 18544 7562 18584
rect 7602 18544 7611 18584
rect 7747 18544 7756 18584
rect 7796 18544 7799 18584
rect 7839 18544 7927 18584
rect 8035 18544 8044 18584
rect 8084 18544 8093 18584
rect 8227 18544 8236 18584
rect 8276 18544 8279 18584
rect 8319 18544 8407 18584
rect 8515 18544 8524 18584
rect 8564 18544 8756 18584
rect 8866 18544 8875 18584
rect 8915 18544 9044 18584
rect 9091 18544 9100 18584
rect 9140 18544 9271 18584
rect 9709 18544 9718 18584
rect 9758 18544 10156 18584
rect 10196 18544 10205 18584
rect 1987 18460 1996 18500
rect 2036 18460 2045 18500
rect 3034 18460 3043 18500
rect 3083 18460 3092 18500
rect 3715 18460 3724 18500
rect 3764 18460 4108 18500
rect 4148 18460 4157 18500
rect 4330 18491 4876 18500
rect 3052 18332 3092 18460
rect 4330 18451 4339 18491
rect 4379 18460 4876 18491
rect 4916 18460 4925 18500
rect 5059 18460 5068 18500
rect 5108 18460 5156 18500
rect 5816 18460 5876 18500
rect 6211 18460 6220 18500
rect 6260 18460 6356 18500
rect 6403 18460 6412 18500
rect 6452 18460 6464 18500
rect 4379 18451 4388 18460
rect 4330 18450 4388 18451
rect 5816 18332 5856 18460
rect 6600 18416 6640 18533
rect 7276 18502 7324 18542
rect 7364 18502 7373 18542
rect 7276 18500 7316 18502
rect 7564 18500 7604 18544
rect 7180 18460 7316 18500
rect 7450 18460 7459 18500
rect 7499 18460 7508 18500
rect 7555 18460 7564 18500
rect 7604 18460 7613 18500
rect 7930 18460 7939 18500
rect 7979 18460 7988 18500
rect 7180 18416 7220 18460
rect 5914 18376 5923 18416
rect 5963 18376 6640 18416
rect 7171 18376 7180 18416
rect 7220 18376 7229 18416
rect 7468 18332 7508 18460
rect 7948 18332 7988 18460
rect 8044 18416 8084 18544
rect 10396 18542 10436 18628
rect 11116 18584 11156 18628
rect 11500 18584 11540 18628
rect 12625 18628 14005 18668
rect 12625 18584 12665 18628
rect 13965 18584 14005 18628
rect 14092 18628 14284 18668
rect 14324 18628 14333 18668
rect 14092 18584 14132 18628
rect 14476 18584 14516 18796
rect 16300 18752 16340 19048
rect 17914 19039 17923 19079
rect 17963 19048 18028 19079
rect 18068 19048 18103 19088
rect 19930 19048 19939 19088
rect 19979 19048 19988 19088
rect 20035 19048 20044 19088
rect 20084 19048 20515 19088
rect 20555 19048 20564 19088
rect 22234 19048 22243 19088
rect 22283 19048 22292 19088
rect 22819 19048 22828 19088
rect 22868 19048 22877 19088
rect 23020 19048 23980 19088
rect 24020 19048 24029 19088
rect 17963 19039 17972 19048
rect 17914 19038 17972 19039
rect 19948 19004 19988 19048
rect 19804 18964 19988 19004
rect 22252 19004 22292 19048
rect 22828 19004 22868 19048
rect 22252 18964 22868 19004
rect 14755 18712 14764 18752
rect 14804 18712 15305 18752
rect 15401 18712 15436 18752
rect 15476 18712 15523 18752
rect 15563 18712 15581 18752
rect 15907 18712 16340 18752
rect 16963 18712 16972 18752
rect 17012 18712 17286 18752
rect 17338 18712 17347 18752
rect 17387 18712 18604 18752
rect 18644 18712 18653 18752
rect 18700 18712 18932 18752
rect 19267 18712 19276 18752
rect 19316 18712 19700 18752
rect 15265 18668 15305 18712
rect 15907 18668 15947 18712
rect 17246 18668 17286 18712
rect 18700 18668 18740 18712
rect 18892 18668 18932 18712
rect 14650 18628 14659 18668
rect 14699 18628 15052 18668
rect 15092 18628 15101 18668
rect 15265 18628 15947 18668
rect 16195 18628 16204 18668
rect 16244 18628 16253 18668
rect 16867 18628 16876 18668
rect 16916 18628 16925 18668
rect 17237 18628 17246 18668
rect 17286 18628 17295 18668
rect 17356 18628 17876 18668
rect 15907 18584 15947 18628
rect 16204 18584 16244 18628
rect 16876 18584 16916 18628
rect 10522 18544 10531 18584
rect 10571 18544 10580 18584
rect 11107 18544 11116 18584
rect 11156 18544 11165 18584
rect 11273 18544 11353 18584
rect 11393 18544 11404 18584
rect 11444 18544 11453 18584
rect 11500 18544 11830 18584
rect 11870 18544 12212 18584
rect 12259 18544 12268 18584
rect 12308 18544 12460 18584
rect 12500 18544 12509 18584
rect 12556 18544 12616 18584
rect 12656 18544 12665 18584
rect 12835 18544 12844 18584
rect 12884 18544 13459 18584
rect 13499 18544 13508 18584
rect 13645 18544 13654 18584
rect 13694 18544 13708 18584
rect 13748 18544 13834 18584
rect 13947 18544 13956 18584
rect 13996 18544 14005 18584
rect 14083 18544 14092 18584
rect 14132 18544 14141 18584
rect 14284 18544 14327 18584
rect 14367 18544 14376 18584
rect 14458 18544 14467 18584
rect 14507 18544 14516 18584
rect 14563 18544 14572 18584
rect 14612 18544 14743 18584
rect 14798 18544 14807 18584
rect 14847 18544 14856 18584
rect 15043 18544 15052 18584
rect 15092 18544 15101 18584
rect 15235 18544 15244 18584
rect 15284 18544 15340 18584
rect 15380 18544 15415 18584
rect 15523 18544 15532 18584
rect 15572 18544 15581 18584
rect 15898 18544 15907 18584
rect 15947 18544 15956 18584
rect 16003 18544 16012 18584
rect 16052 18544 16061 18584
rect 16195 18544 16204 18584
rect 16244 18544 16291 18584
rect 16579 18544 16588 18584
rect 16628 18544 16696 18584
rect 16736 18544 16759 18584
rect 16829 18544 16871 18584
rect 16911 18544 16920 18584
rect 17059 18544 17068 18584
rect 17108 18544 17239 18584
rect 10378 18502 10387 18542
rect 10427 18502 10436 18542
rect 10540 18500 10580 18544
rect 12172 18500 12212 18544
rect 8297 18460 8419 18500
rect 8468 18460 8477 18500
rect 8611 18460 8620 18500
rect 8660 18460 8924 18500
rect 8986 18460 8995 18500
rect 9035 18460 9044 18500
rect 9571 18460 9580 18500
rect 9620 18460 10195 18500
rect 10235 18460 10244 18500
rect 10540 18491 11308 18500
rect 10540 18460 11251 18491
rect 8044 18376 8716 18416
rect 8756 18376 8765 18416
rect 8884 18332 8924 18460
rect 9004 18416 9044 18460
rect 11242 18451 11251 18460
rect 11291 18460 11308 18491
rect 11348 18460 11357 18500
rect 11626 18460 11635 18500
rect 11675 18460 12116 18500
rect 12163 18460 12172 18500
rect 12212 18460 12221 18500
rect 11291 18451 11300 18460
rect 11242 18450 11300 18451
rect 9004 18376 9140 18416
rect 1123 18292 1132 18332
rect 1172 18292 2284 18332
rect 2324 18292 2333 18332
rect 2380 18292 3092 18332
rect 3235 18292 3244 18332
rect 3284 18292 3293 18332
rect 5816 18292 6892 18332
rect 6932 18292 6941 18332
rect 7468 18292 7756 18332
rect 7796 18292 7805 18332
rect 7948 18292 8524 18332
rect 8564 18292 8573 18332
rect 8884 18292 9004 18332
rect 9044 18292 9053 18332
rect 2380 17912 2420 18292
rect 3244 18248 3284 18292
rect 9100 18248 9140 18376
rect 12076 18332 12116 18460
rect 12556 18416 12596 18544
rect 13468 18500 13508 18544
rect 14284 18500 14324 18544
rect 14807 18500 14847 18544
rect 12748 18460 12796 18500
rect 12836 18460 12845 18500
rect 13468 18460 13900 18500
rect 13940 18460 13949 18500
rect 14275 18460 14284 18500
rect 14324 18460 14333 18500
rect 14668 18460 14847 18500
rect 14938 18460 14947 18500
rect 14987 18460 14996 18500
rect 12748 18416 12788 18460
rect 14668 18416 14708 18460
rect 12451 18376 12460 18416
rect 12500 18376 12596 18416
rect 12643 18376 12652 18416
rect 12692 18376 12788 18416
rect 13987 18376 13996 18416
rect 14036 18376 14380 18416
rect 14420 18376 14429 18416
rect 14659 18376 14668 18416
rect 14708 18376 14717 18416
rect 10627 18292 10636 18332
rect 10676 18292 13556 18332
rect 2476 18208 3284 18248
rect 6595 18208 6604 18248
rect 6644 18208 9196 18248
rect 9236 18208 9300 18248
rect 1865 17872 1996 17912
rect 2036 17872 2045 17912
rect 2371 17872 2380 17912
rect 2420 17872 2429 17912
rect 2284 17788 2380 17828
rect 2420 17788 2429 17828
rect 2284 17744 2324 17788
rect 2476 17744 2516 18208
rect 3103 18124 3112 18164
rect 3480 18124 3489 18164
rect 9004 18124 9257 18164
rect 10877 18124 10886 18164
rect 11254 18124 11263 18164
rect 11308 18124 11500 18164
rect 11540 18124 12460 18164
rect 12500 18124 12509 18164
rect 9004 18080 9044 18124
rect 9217 18080 9257 18124
rect 11308 18080 11348 18124
rect 6211 18040 6220 18080
rect 6260 18040 6356 18080
rect 6316 17996 6356 18040
rect 6988 18040 7695 18080
rect 6988 17996 7028 18040
rect 2860 17956 3724 17996
rect 3764 17956 3773 17996
rect 6307 17956 6316 17996
rect 6356 17956 6365 17996
rect 6970 17956 6979 17996
rect 7019 17956 7028 17996
rect 7171 17956 7180 17996
rect 7220 17956 7555 17996
rect 7595 17956 7604 17996
rect 2633 17788 2668 17828
rect 2708 17788 2764 17828
rect 2804 17788 2813 17828
rect 2860 17744 2900 17956
rect 3715 17872 3724 17912
rect 3764 17872 3820 17912
rect 3860 17872 3895 17912
rect 4073 17872 4204 17912
rect 4244 17872 4253 17912
rect 4963 17872 4972 17912
rect 5012 17872 5932 17912
rect 5972 17872 5981 17912
rect 6211 17872 6220 17912
rect 6260 17872 6269 17912
rect 6364 17872 7180 17912
rect 7220 17872 7229 17912
rect 2947 17788 2956 17828
rect 2996 17788 3476 17828
rect 3436 17744 3476 17788
rect 5068 17788 5356 17828
rect 5396 17788 5405 17828
rect 5068 17779 5108 17788
rect 5026 17744 5108 17779
rect 6216 17755 6256 17872
rect 6364 17755 6404 17872
rect 7655 17828 7695 18040
rect 8620 18040 9044 18080
rect 9091 18040 9100 18080
rect 9140 18040 9149 18080
rect 9217 18040 11348 18080
rect 11395 18040 11404 18080
rect 11444 18040 12364 18080
rect 12404 18040 12413 18080
rect 8620 17912 8660 18040
rect 9100 17912 9140 18040
rect 6595 17788 6604 17828
rect 6644 17788 6932 17828
rect 2275 17704 2284 17744
rect 2324 17704 2333 17744
rect 2458 17704 2467 17744
rect 2507 17704 2516 17744
rect 2563 17704 2572 17744
rect 2612 17704 2743 17744
rect 2851 17704 2860 17744
rect 2900 17704 2909 17744
rect 2956 17704 2979 17744
rect 3019 17704 3028 17744
rect 3088 17704 3097 17744
rect 3137 17704 3148 17744
rect 3188 17704 3277 17744
rect 3418 17704 3427 17744
rect 3467 17704 3476 17744
rect 3523 17704 3532 17744
rect 3572 17704 4204 17744
rect 4244 17704 4253 17744
rect 4387 17704 4396 17744
rect 4436 17704 4567 17744
rect 4649 17704 4780 17744
rect 4820 17704 4829 17744
rect 4890 17704 4899 17744
rect 4939 17704 4964 17744
rect 5008 17704 5017 17744
rect 5057 17739 5108 17744
rect 5057 17704 5066 17739
rect 5253 17704 5262 17744
rect 5302 17704 5347 17744
rect 5443 17704 5452 17744
rect 5492 17704 5501 17744
rect 5642 17704 5740 17744
rect 5804 17704 5822 17744
rect 5914 17704 5923 17744
rect 5963 17704 5972 17744
rect 6058 17704 6067 17744
rect 6107 17704 6116 17744
rect 6198 17715 6207 17755
rect 6247 17715 6256 17755
rect 6324 17715 6333 17755
rect 6373 17715 6404 17755
rect 6892 17744 6932 17788
rect 7372 17788 7468 17828
rect 7508 17788 7517 17828
rect 7561 17788 7695 17828
rect 7996 17872 8660 17912
rect 8707 17872 8716 17912
rect 8756 17872 8765 17912
rect 9091 17872 9100 17912
rect 9140 17872 9149 17912
rect 7996 17828 8036 17872
rect 8716 17828 8756 17872
rect 9217 17828 9257 18040
rect 11212 17996 11252 18040
rect 9763 17956 9772 17996
rect 9812 17956 11020 17996
rect 11060 17956 11069 17996
rect 11203 17956 11212 17996
rect 11252 17956 11261 17996
rect 9426 17872 9676 17912
rect 9716 17872 9725 17912
rect 9964 17872 11500 17912
rect 11540 17872 11549 17912
rect 7996 17788 8044 17828
rect 8084 17788 8196 17828
rect 8489 17788 8572 17828
rect 8612 17788 8620 17828
rect 8660 17788 8669 17828
rect 8716 17788 9004 17828
rect 9044 17788 9053 17828
rect 9217 17788 9332 17828
rect 7372 17744 7412 17788
rect 7561 17744 7601 17788
rect 7996 17744 8036 17788
rect 9292 17744 9332 17788
rect 9426 17786 9466 17872
rect 9964 17828 10004 17872
rect 9562 17788 9571 17828
rect 9611 17788 9908 17828
rect 9955 17788 9964 17828
rect 10004 17788 10013 17828
rect 10444 17788 10540 17828
rect 10580 17788 10589 17828
rect 10723 17788 10732 17828
rect 10772 17788 11116 17828
rect 11156 17788 11165 17828
rect 9426 17746 9436 17786
rect 9476 17746 9485 17786
rect 9868 17744 9908 17788
rect 10444 17744 10484 17788
rect 11692 17744 11732 18040
rect 13516 17996 13556 18292
rect 14668 18164 14708 18376
rect 14956 18332 14996 18460
rect 15052 18416 15092 18544
rect 15139 18460 15148 18500
rect 15188 18460 15319 18500
rect 15052 18376 15244 18416
rect 15284 18376 15293 18416
rect 15363 18332 15403 18544
rect 15532 18500 15572 18544
rect 15532 18460 15947 18500
rect 15619 18376 15628 18416
rect 15668 18376 15724 18416
rect 15764 18376 15799 18416
rect 14755 18292 14764 18332
rect 14804 18292 14996 18332
rect 15191 18292 15403 18332
rect 15907 18332 15947 18460
rect 16012 18416 16052 18544
rect 17356 18500 17396 18628
rect 17836 18584 17876 18628
rect 18367 18628 18740 18668
rect 18787 18628 18796 18668
rect 18836 18628 18845 18668
rect 18892 18628 19564 18668
rect 19604 18628 19613 18668
rect 18367 18584 18407 18628
rect 18796 18584 18836 18628
rect 19660 18584 19700 18712
rect 19804 18584 19844 18964
rect 19891 18880 19900 18920
rect 20268 18880 20277 18920
rect 23203 18880 23212 18920
rect 23252 18880 23404 18920
rect 23444 18880 24404 18920
rect 20236 18796 21292 18836
rect 21332 18796 21341 18836
rect 20236 18752 20276 18796
rect 24364 18752 24404 18880
rect 24460 18836 24500 19132
rect 24652 19004 24692 19216
rect 24739 19132 24748 19172
rect 24788 19132 28963 19172
rect 29003 19132 29012 19172
rect 24835 19048 24844 19088
rect 24884 19048 25123 19088
rect 25163 19048 25172 19088
rect 25673 19048 25804 19088
rect 25844 19048 25853 19088
rect 26074 19048 26083 19088
rect 26123 19048 26228 19088
rect 26275 19079 26284 19088
rect 26275 19048 26283 19079
rect 26324 19048 26454 19088
rect 27497 19048 27628 19088
rect 27668 19048 27677 19088
rect 28771 19048 28780 19088
rect 28820 19048 31084 19088
rect 31124 19048 31133 19088
rect 24652 18964 26092 19004
rect 26132 18964 26141 19004
rect 26188 18920 26228 19048
rect 26283 19030 26323 19039
rect 26380 18964 30508 19004
rect 30548 18964 30557 19004
rect 26380 18920 26420 18964
rect 25603 18880 25612 18920
rect 25652 18880 26420 18920
rect 27665 18880 27674 18920
rect 28042 18880 28051 18920
rect 28867 18880 28876 18920
rect 28916 18880 30164 18920
rect 28876 18836 28916 18880
rect 24460 18796 28916 18836
rect 29443 18796 29452 18836
rect 29492 18796 29932 18836
rect 29972 18796 29981 18836
rect 20218 18712 20227 18752
rect 20267 18712 20276 18752
rect 20323 18712 20332 18752
rect 20372 18712 20908 18752
rect 20948 18712 20957 18752
rect 21187 18712 21196 18752
rect 21236 18712 21245 18752
rect 23011 18712 23020 18752
rect 23060 18712 23191 18752
rect 23971 18712 23980 18752
rect 24020 18712 24268 18752
rect 24308 18712 24317 18752
rect 24364 18712 24692 18752
rect 24931 18712 24940 18752
rect 24980 18712 25268 18752
rect 25411 18712 25420 18752
rect 25460 18712 25699 18752
rect 25739 18712 27380 18752
rect 27427 18712 27436 18752
rect 27476 18712 27860 18752
rect 21196 18668 21236 18712
rect 24652 18668 24692 18712
rect 20122 18659 20524 18668
rect 20122 18619 20131 18659
rect 20171 18628 20524 18659
rect 20564 18628 21236 18668
rect 21850 18628 21859 18668
rect 21899 18628 22292 18668
rect 22339 18628 22348 18668
rect 22388 18628 22444 18668
rect 22484 18628 22519 18668
rect 22924 18628 23212 18668
rect 23252 18628 23261 18668
rect 23692 18628 23788 18668
rect 23828 18628 23837 18668
rect 24067 18628 24076 18668
rect 24116 18628 24596 18668
rect 24652 18628 25076 18668
rect 20171 18619 20180 18628
rect 20122 18618 20180 18619
rect 22252 18584 22292 18628
rect 22924 18584 22964 18628
rect 23692 18584 23732 18628
rect 24556 18584 24596 18628
rect 25036 18584 25076 18628
rect 25228 18584 25268 18712
rect 27340 18668 27380 18712
rect 27820 18668 27860 18712
rect 29164 18712 29780 18752
rect 29164 18668 29204 18712
rect 29740 18668 29780 18712
rect 25612 18628 25804 18668
rect 25844 18628 25853 18668
rect 26275 18628 26284 18668
rect 26324 18628 26333 18668
rect 26467 18628 26476 18668
rect 26516 18628 27092 18668
rect 27340 18628 27764 18668
rect 27820 18628 29204 18668
rect 29260 18628 29644 18668
rect 29684 18628 29693 18668
rect 29740 18628 29876 18668
rect 30019 18628 30028 18668
rect 30068 18628 30077 18668
rect 25612 18584 25652 18628
rect 26284 18584 26324 18628
rect 27052 18584 27092 18628
rect 17443 18544 17452 18584
rect 17492 18544 17501 18584
rect 17548 18575 17684 18584
rect 16195 18460 16204 18500
rect 16244 18460 16531 18500
rect 16571 18460 17396 18500
rect 17452 18416 17492 18544
rect 17588 18544 17684 18575
rect 17827 18544 17836 18584
rect 17876 18544 18007 18584
rect 18349 18544 18358 18584
rect 18398 18544 18407 18584
rect 18595 18544 18604 18584
rect 18644 18544 18836 18584
rect 18916 18544 18925 18584
rect 18965 18544 19028 18584
rect 19145 18544 19180 18584
rect 19220 18544 19276 18584
rect 19316 18544 19325 18584
rect 19459 18544 19468 18584
rect 19508 18544 19517 18584
rect 19651 18544 19660 18584
rect 19700 18544 19709 18584
rect 19804 18544 19843 18584
rect 19883 18544 19892 18584
rect 19948 18575 19988 18584
rect 17548 18526 17588 18535
rect 16012 18376 16588 18416
rect 16628 18376 16637 18416
rect 17251 18376 17260 18416
rect 17300 18376 17492 18416
rect 17644 18332 17684 18544
rect 18988 18500 19028 18544
rect 18154 18460 18163 18500
rect 18203 18460 18212 18500
rect 18979 18460 18988 18500
rect 19028 18460 19037 18500
rect 15907 18292 16492 18332
rect 16532 18292 16541 18332
rect 16963 18292 16972 18332
rect 17012 18292 17021 18332
rect 17443 18292 17452 18332
rect 17492 18292 17684 18332
rect 14668 18124 14847 18164
rect 11971 17956 11980 17996
rect 12020 17956 12172 17996
rect 12212 17956 12221 17996
rect 12547 17956 12556 17996
rect 12596 17956 12748 17996
rect 12788 17956 12797 17996
rect 13516 17956 14284 17996
rect 14324 17956 14668 17996
rect 14708 17956 14717 17996
rect 13123 17872 13132 17912
rect 13172 17872 13181 17912
rect 13132 17828 13172 17872
rect 12124 17788 13172 17828
rect 13219 17788 13228 17828
rect 13268 17788 13277 17828
rect 12124 17744 12164 17788
rect 12652 17744 12692 17788
rect 13228 17744 13268 17788
rect 13516 17744 13556 17956
rect 14807 17912 14847 18124
rect 13891 17872 13900 17912
rect 13940 17872 14324 17912
rect 14371 17872 14380 17912
rect 14420 17872 14847 17912
rect 14284 17828 14324 17872
rect 13626 17788 13635 17828
rect 13675 17788 13996 17828
rect 14036 17788 14115 17828
rect 14155 17788 14196 17828
rect 14284 17788 14367 17828
rect 14441 17788 14467 17828
rect 14507 17788 14572 17828
rect 14612 17788 14621 17828
rect 14327 17744 14367 17788
rect 14807 17744 14847 17872
rect 15191 17828 15231 18292
rect 16972 18248 17012 18292
rect 18172 18248 18212 18460
rect 19468 18416 19508 18544
rect 20218 18544 20227 18584
rect 20267 18544 20276 18584
rect 20395 18544 20404 18584
rect 20468 18544 20584 18584
rect 20631 18544 20659 18584
rect 20699 18544 20708 18584
rect 20753 18544 20762 18584
rect 20802 18544 20812 18584
rect 20852 18544 20942 18584
rect 21091 18544 21100 18584
rect 21140 18544 21236 18584
rect 21283 18544 21292 18584
rect 21332 18544 21463 18584
rect 21667 18544 21676 18584
rect 21716 18544 21772 18584
rect 21812 18544 21847 18584
rect 21946 18544 21955 18584
rect 21995 18544 22004 18584
rect 22051 18544 22060 18584
rect 22100 18544 22109 18584
rect 22234 18544 22243 18584
rect 22283 18544 22292 18584
rect 22339 18544 22348 18584
rect 22388 18544 22397 18584
rect 22444 18544 22554 18584
rect 22594 18544 22732 18584
rect 22772 18544 22781 18584
rect 22924 18575 23012 18584
rect 22924 18544 22963 18575
rect 19948 18500 19988 18535
rect 19651 18460 19660 18500
rect 19700 18460 19988 18500
rect 20236 18500 20276 18544
rect 20631 18500 20671 18544
rect 21196 18500 21236 18544
rect 21964 18500 22004 18544
rect 20236 18460 20332 18500
rect 20372 18460 20381 18500
rect 20536 18460 20671 18500
rect 21187 18460 21196 18500
rect 21236 18460 21245 18500
rect 21859 18460 21868 18500
rect 21908 18460 22004 18500
rect 18307 18376 18316 18416
rect 18356 18376 18508 18416
rect 18548 18376 19508 18416
rect 20536 18416 20576 18460
rect 20536 18376 21388 18416
rect 21428 18376 21437 18416
rect 20536 18332 20576 18376
rect 18403 18292 18412 18332
rect 18452 18292 20576 18332
rect 22060 18248 22100 18544
rect 22348 18416 22388 18544
rect 22444 18500 22484 18544
rect 22954 18535 22963 18544
rect 23003 18535 23012 18575
rect 23062 18544 23071 18584
rect 23111 18544 23408 18584
rect 23465 18544 23596 18584
rect 23636 18544 23645 18584
rect 23692 18575 23747 18584
rect 23692 18544 23707 18575
rect 22954 18534 23012 18535
rect 23368 18500 23408 18544
rect 23596 18526 23636 18535
rect 23707 18526 23747 18535
rect 23818 18575 23980 18584
rect 23818 18535 23827 18575
rect 23867 18544 23980 18575
rect 24020 18544 24029 18584
rect 24224 18544 24233 18584
rect 24273 18544 24364 18584
rect 24404 18544 24413 18584
rect 24547 18544 24556 18584
rect 24596 18544 24605 18584
rect 24739 18544 24748 18584
rect 24788 18544 24797 18584
rect 24844 18544 24863 18584
rect 24903 18544 24931 18584
rect 25027 18544 25036 18584
rect 25076 18544 25085 18584
rect 25219 18544 25228 18584
rect 25268 18544 25277 18584
rect 25402 18544 25411 18584
rect 25451 18544 25460 18584
rect 25594 18544 25603 18584
rect 25643 18544 25652 18584
rect 25804 18544 25911 18584
rect 25951 18544 25960 18584
rect 26179 18544 26188 18584
rect 26228 18544 26324 18584
rect 26371 18544 26380 18584
rect 26420 18544 26551 18584
rect 26755 18544 26764 18584
rect 26804 18544 26860 18584
rect 26900 18544 26935 18584
rect 27034 18544 27043 18584
rect 27083 18544 27092 18584
rect 27139 18544 27148 18584
rect 27188 18544 27572 18584
rect 23867 18535 23876 18544
rect 23818 18534 23876 18535
rect 24748 18500 24788 18544
rect 24844 18500 24884 18544
rect 22435 18460 22444 18500
rect 22484 18460 22493 18500
rect 23368 18460 23500 18500
rect 23540 18460 23549 18500
rect 24326 18460 24335 18500
rect 24375 18460 24788 18500
rect 24835 18460 24844 18500
rect 24884 18460 24893 18500
rect 24364 18416 24404 18460
rect 22348 18376 23252 18416
rect 23971 18376 23980 18416
rect 24020 18376 24404 18416
rect 24547 18376 24556 18416
rect 24596 18376 24748 18416
rect 24788 18376 24797 18416
rect 23212 18332 23252 18376
rect 25036 18332 25076 18544
rect 25420 18500 25460 18544
rect 25420 18460 25612 18500
rect 25652 18460 25661 18500
rect 25804 18416 25844 18544
rect 26380 18500 26420 18544
rect 25961 18460 26083 18500
rect 26132 18460 26141 18500
rect 26380 18460 27340 18500
rect 27380 18460 27389 18500
rect 27532 18416 27572 18544
rect 27724 18500 27764 18628
rect 29260 18584 29300 18628
rect 29836 18584 29876 18628
rect 30028 18584 30068 18628
rect 30124 18584 30164 18880
rect 30307 18712 30316 18752
rect 30356 18712 30365 18752
rect 30316 18584 30356 18712
rect 30403 18628 30412 18668
rect 30452 18628 30700 18668
rect 30740 18628 30749 18668
rect 29242 18544 29251 18584
rect 29291 18544 29300 18584
rect 29539 18544 29548 18584
rect 29588 18544 29635 18584
rect 29675 18544 29719 18584
rect 29813 18544 29822 18584
rect 29862 18544 29876 18584
rect 29923 18544 29932 18584
rect 29972 18544 30068 18584
rect 30115 18544 30124 18584
rect 30164 18544 30173 18584
rect 30307 18544 30316 18584
rect 30356 18544 30365 18584
rect 30595 18544 30604 18584
rect 30644 18544 30653 18584
rect 30778 18575 31124 18584
rect 27706 18460 27715 18500
rect 27755 18460 27764 18500
rect 29472 18460 30316 18500
rect 30356 18460 30365 18500
rect 25804 18376 26228 18416
rect 26825 18376 26956 18416
rect 26996 18376 27005 18416
rect 27532 18376 27724 18416
rect 27764 18376 27773 18416
rect 29705 18376 29836 18416
rect 29876 18376 29885 18416
rect 22243 18292 22252 18332
rect 22292 18292 22636 18332
rect 22676 18292 22828 18332
rect 22868 18292 22877 18332
rect 23212 18292 24268 18332
rect 24308 18292 24317 18332
rect 24451 18292 24460 18332
rect 24500 18292 25076 18332
rect 25402 18292 25411 18332
rect 25451 18292 25460 18332
rect 25891 18292 25900 18332
rect 25940 18292 25949 18332
rect 15427 18208 15436 18248
rect 15476 18208 17012 18248
rect 17251 18208 17260 18248
rect 17300 18208 18212 18248
rect 19084 18208 21964 18248
rect 22004 18208 22013 18248
rect 22060 18208 23020 18248
rect 23060 18208 23069 18248
rect 23203 18208 23212 18248
rect 23252 18208 24364 18248
rect 24404 18208 24413 18248
rect 18651 18124 18660 18164
rect 19028 18124 19037 18164
rect 19084 18080 19124 18208
rect 25420 18164 25460 18292
rect 25900 18248 25940 18292
rect 19267 18124 19276 18164
rect 19316 18124 25460 18164
rect 25708 18208 25940 18248
rect 17827 18040 17836 18080
rect 17876 18040 19124 18080
rect 20227 18040 20236 18080
rect 20276 18040 20620 18080
rect 20660 18040 20669 18080
rect 20803 18040 20812 18080
rect 20852 18040 21580 18080
rect 21620 18040 23444 18080
rect 23587 18040 23596 18080
rect 23636 18040 23876 18080
rect 15427 17956 15436 17996
rect 15476 17956 20564 17996
rect 22147 17956 22156 17996
rect 22196 17956 22636 17996
rect 22676 17956 22685 17996
rect 20524 17912 20564 17956
rect 16387 17872 16396 17912
rect 16436 17872 17396 17912
rect 15139 17788 15148 17828
rect 15188 17788 15231 17828
rect 15715 17788 15724 17828
rect 15764 17788 16147 17828
rect 16187 17788 16196 17828
rect 16771 17788 16780 17828
rect 16820 17788 17130 17828
rect 16780 17744 16820 17788
rect 17090 17744 17130 17788
rect 17356 17744 17396 17872
rect 18028 17872 18988 17912
rect 19028 17872 19037 17912
rect 19747 17872 19756 17912
rect 19796 17872 20044 17912
rect 20084 17872 20093 17912
rect 20140 17872 20428 17912
rect 20468 17872 20477 17912
rect 20524 17872 22292 17912
rect 6665 17704 6796 17744
rect 6836 17704 6845 17744
rect 6892 17704 6965 17744
rect 7005 17704 7014 17744
rect 7171 17704 7180 17744
rect 7220 17704 7229 17744
rect 7363 17704 7372 17744
rect 7412 17704 7421 17744
rect 7546 17704 7555 17744
rect 7595 17704 7604 17744
rect 7664 17704 7673 17744
rect 7713 17704 7722 17744
rect 2956 17660 2996 17704
rect 4924 17660 4964 17704
rect 5260 17660 5300 17704
rect 5452 17660 5492 17704
rect 5932 17660 5972 17704
rect 6076 17660 6116 17704
rect 7180 17660 7220 17704
rect 2956 17620 3724 17660
rect 3764 17620 3773 17660
rect 4579 17620 4588 17660
rect 4628 17620 4684 17660
rect 4724 17620 4759 17660
rect 4924 17620 4972 17660
rect 5012 17620 5021 17660
rect 5251 17620 5260 17660
rect 5300 17620 5309 17660
rect 5417 17620 5548 17660
rect 5588 17620 5597 17660
rect 5885 17620 5932 17660
rect 5972 17620 5981 17660
rect 6076 17620 6508 17660
rect 6548 17620 6557 17660
rect 7180 17620 7276 17660
rect 7316 17620 7325 17660
rect 5548 17576 5588 17620
rect 2083 17536 2092 17576
rect 2132 17536 3436 17576
rect 3476 17536 3628 17576
rect 3668 17536 3677 17576
rect 5321 17536 5452 17576
rect 5492 17536 5501 17576
rect 5548 17536 6412 17576
rect 6452 17536 6461 17576
rect 7372 17408 7412 17704
rect 7682 17660 7722 17704
rect 7834 17735 7915 17744
rect 7834 17695 7843 17735
rect 7883 17695 7915 17735
rect 7970 17704 7979 17744
rect 8019 17704 8036 17744
rect 8107 17704 8116 17744
rect 8156 17704 8276 17744
rect 8323 17704 8332 17744
rect 8411 17704 8503 17744
rect 8620 17704 8860 17744
rect 8900 17704 8909 17744
rect 9065 17704 9175 17744
rect 9236 17704 9245 17744
rect 9292 17704 9315 17744
rect 9355 17704 9364 17744
rect 9648 17704 9657 17744
rect 9697 17704 9706 17744
rect 9868 17704 10484 17744
rect 10526 17704 10636 17744
rect 10688 17704 10706 17744
rect 10766 17704 10775 17744
rect 10815 17704 10824 17744
rect 10906 17704 10915 17744
rect 10955 17704 10964 17744
rect 11011 17704 11020 17744
rect 11060 17704 11191 17744
rect 11491 17704 11500 17744
rect 11540 17704 11549 17744
rect 11683 17704 11692 17744
rect 11732 17704 11741 17744
rect 11837 17704 11873 17744
rect 11913 17704 11924 17744
rect 12076 17704 12085 17744
rect 12125 17704 12164 17744
rect 12220 17704 12268 17744
rect 12308 17704 12317 17744
rect 12442 17704 12451 17744
rect 12491 17704 12547 17744
rect 12643 17704 12652 17744
rect 12692 17704 12701 17744
rect 7834 17694 7915 17695
rect 7459 17620 7468 17660
rect 7508 17620 7722 17660
rect 7875 17576 7915 17694
rect 8236 17660 8276 17704
rect 8620 17660 8660 17704
rect 8227 17620 8236 17660
rect 8276 17620 8285 17660
rect 8611 17620 8620 17660
rect 8660 17620 8669 17660
rect 7651 17536 7660 17576
rect 7700 17536 9196 17576
rect 9236 17536 9245 17576
rect 9652 17492 9692 17704
rect 10775 17660 10815 17704
rect 10243 17620 10252 17660
rect 10292 17620 10483 17660
rect 10523 17620 10815 17660
rect 10924 17660 10964 17704
rect 11500 17660 11540 17704
rect 11884 17660 11924 17704
rect 10924 17620 11308 17660
rect 11348 17620 11357 17660
rect 11500 17620 11596 17660
rect 11636 17620 11645 17660
rect 11875 17620 11884 17660
rect 11924 17620 11933 17660
rect 12220 17576 12260 17704
rect 12460 17660 12500 17704
rect 12830 17677 12839 17717
rect 12879 17677 12888 17717
rect 13027 17704 13036 17744
rect 13076 17704 13085 17744
rect 13181 17704 13226 17744
rect 13266 17704 13275 17744
rect 13507 17704 13516 17744
rect 13556 17704 13565 17744
rect 13699 17704 13708 17744
rect 13773 17704 13879 17744
rect 13987 17704 13996 17744
rect 14036 17704 14045 17744
rect 14204 17704 14213 17744
rect 14253 17704 14262 17744
rect 14318 17704 14327 17744
rect 14367 17704 14376 17744
rect 14537 17704 14572 17744
rect 14612 17704 14668 17744
rect 14708 17704 14717 17744
rect 14798 17704 14807 17744
rect 14847 17704 14856 17744
rect 14938 17704 14947 17744
rect 14987 17704 14996 17744
rect 15043 17704 15052 17744
rect 15092 17704 15139 17744
rect 15475 17704 15484 17744
rect 15524 17704 15533 17744
rect 15610 17704 15619 17744
rect 15659 17704 15668 17744
rect 15715 17704 15724 17744
rect 15764 17704 15820 17744
rect 15860 17704 15895 17744
rect 16190 17704 16300 17744
rect 16352 17704 16370 17744
rect 16474 17704 16483 17744
rect 16532 17704 16663 17744
rect 16733 17704 16776 17744
rect 16816 17704 16825 17744
rect 16954 17704 16963 17744
rect 17003 17704 17012 17744
rect 17072 17704 17081 17744
rect 17121 17704 17130 17744
rect 17239 17704 17248 17744
rect 17288 17704 17297 17744
rect 17346 17704 17355 17744
rect 17395 17704 17404 17744
rect 17515 17704 17524 17744
rect 17564 17704 17836 17744
rect 17876 17704 17885 17744
rect 12451 17620 12460 17660
rect 12500 17620 12509 17660
rect 12844 17576 12884 17677
rect 13036 17660 13076 17704
rect 13036 17620 13900 17660
rect 13940 17620 13949 17660
rect 13996 17576 14036 17704
rect 14213 17660 14253 17704
rect 14572 17660 14612 17704
rect 14213 17620 14612 17660
rect 9754 17536 9763 17576
rect 9803 17536 10060 17576
rect 10100 17536 10109 17576
rect 10195 17536 10204 17576
rect 10244 17536 10348 17576
rect 10388 17536 10397 17576
rect 11331 17536 12260 17576
rect 12355 17536 12364 17576
rect 12404 17536 12652 17576
rect 12692 17536 12701 17576
rect 12835 17536 12844 17576
rect 12884 17536 12893 17576
rect 13001 17536 13132 17576
rect 13172 17536 13181 17576
rect 13411 17536 13420 17576
rect 13460 17536 13900 17576
rect 13940 17536 13949 17576
rect 13996 17536 14188 17576
rect 14228 17536 14237 17576
rect 14650 17536 14659 17576
rect 14699 17536 14708 17576
rect 9652 17452 9676 17492
rect 9716 17452 9725 17492
rect 11331 17408 11371 17536
rect 13996 17492 14036 17536
rect 4343 17368 4352 17408
rect 4720 17368 4729 17408
rect 7372 17368 11371 17408
rect 12028 17452 14036 17492
rect 12028 17324 12068 17452
rect 14668 17408 14708 17536
rect 12117 17368 12126 17408
rect 12494 17368 12503 17408
rect 14659 17368 14668 17408
rect 14708 17368 14717 17408
rect 14956 17324 14996 17704
rect 15052 17660 15092 17704
rect 15043 17620 15052 17660
rect 15092 17620 15101 17660
rect 15484 17576 15524 17704
rect 15628 17660 15668 17704
rect 16972 17660 17012 17704
rect 17246 17660 17286 17704
rect 18028 17660 18068 17872
rect 20140 17828 20180 17872
rect 18595 17788 18604 17828
rect 18644 17788 18653 17828
rect 18787 17788 18796 17828
rect 18836 17788 18869 17828
rect 18909 17788 18967 17828
rect 19075 17788 19084 17828
rect 19124 17788 19255 17828
rect 19660 17788 20180 17828
rect 20227 17788 20236 17828
rect 20276 17788 20285 17828
rect 20332 17788 20995 17828
rect 21035 17788 21044 17828
rect 21187 17788 21196 17828
rect 21236 17788 22060 17828
rect 22100 17788 22196 17828
rect 18604 17744 18644 17788
rect 19660 17786 19700 17788
rect 19594 17746 19603 17786
rect 19643 17746 19700 17786
rect 20236 17744 20276 17788
rect 20332 17744 20372 17788
rect 22156 17744 22196 17788
rect 18115 17704 18124 17744
rect 18164 17704 18263 17744
rect 18303 17704 18312 17744
rect 18367 17704 18389 17744
rect 18429 17704 18438 17744
rect 18492 17704 18501 17744
rect 18541 17704 18644 17744
rect 18691 17704 18700 17744
rect 18740 17704 18743 17744
rect 18783 17704 18871 17744
rect 18979 17704 18988 17744
rect 19028 17704 19159 17744
rect 20035 17704 20044 17744
rect 20084 17704 20093 17744
rect 20160 17704 20169 17744
rect 20209 17704 20276 17744
rect 20323 17704 20332 17744
rect 20372 17704 20381 17744
rect 20506 17704 20515 17744
rect 20564 17704 20695 17744
rect 20803 17704 20812 17744
rect 20852 17704 21004 17744
rect 21044 17704 21053 17744
rect 21667 17704 21676 17744
rect 21716 17704 21725 17744
rect 21833 17704 21964 17744
rect 22004 17704 22013 17744
rect 22147 17704 22156 17744
rect 22196 17704 22205 17744
rect 18367 17660 18407 17704
rect 15581 17620 15628 17660
rect 15668 17620 15677 17660
rect 15802 17620 15811 17660
rect 15851 17620 16204 17660
rect 16244 17620 16253 17660
rect 16675 17620 16684 17660
rect 16724 17620 17012 17660
rect 17100 17620 17260 17660
rect 17300 17620 17309 17660
rect 17452 17620 18068 17660
rect 18307 17620 18316 17660
rect 18356 17620 18407 17660
rect 17246 17576 17286 17620
rect 17452 17576 17492 17620
rect 20044 17576 20084 17704
rect 21676 17660 21716 17704
rect 20323 17620 20332 17660
rect 20372 17620 22051 17660
rect 22091 17620 22100 17660
rect 15324 17536 15436 17576
rect 15476 17536 15524 17576
rect 16867 17536 16876 17576
rect 16916 17536 17286 17576
rect 17434 17536 17443 17576
rect 17483 17536 17492 17576
rect 17722 17536 17731 17576
rect 17771 17536 17780 17576
rect 17827 17536 17836 17576
rect 17876 17536 18019 17576
rect 18059 17536 18068 17576
rect 18403 17536 18412 17576
rect 18452 17536 18595 17576
rect 18635 17536 18644 17576
rect 19180 17536 19411 17576
rect 19451 17536 19460 17576
rect 20044 17536 20524 17576
rect 20564 17536 20573 17576
rect 20707 17536 20716 17576
rect 20756 17536 20812 17576
rect 20852 17536 20887 17576
rect 15484 17408 15524 17536
rect 17740 17492 17780 17536
rect 19180 17492 19220 17536
rect 16675 17452 16684 17492
rect 16724 17452 17780 17492
rect 19171 17452 19180 17492
rect 19220 17452 19229 17492
rect 19468 17452 21772 17492
rect 21812 17452 21821 17492
rect 19468 17408 19508 17452
rect 22060 17408 22100 17620
rect 22252 17492 22292 17872
rect 22819 17788 22828 17828
rect 22868 17788 22964 17828
rect 23107 17788 23116 17828
rect 23156 17788 23308 17828
rect 23348 17788 23357 17828
rect 22924 17744 22964 17788
rect 23212 17744 23252 17788
rect 23404 17744 23444 18040
rect 23491 17956 23500 17996
rect 23540 17956 23671 17996
rect 23587 17788 23596 17828
rect 23636 17788 23780 17828
rect 23740 17786 23780 17788
rect 23740 17777 23783 17786
rect 23740 17746 23743 17777
rect 22339 17704 22348 17744
rect 22388 17704 22819 17744
rect 22859 17704 22868 17744
rect 23050 17704 23059 17744
rect 23099 17704 23156 17744
rect 23203 17704 23212 17744
rect 23252 17704 23261 17744
rect 23395 17704 23404 17744
rect 23444 17704 23453 17744
rect 23500 17704 23526 17744
rect 23566 17704 23575 17744
rect 23635 17704 23644 17744
rect 23684 17704 23693 17744
rect 23743 17728 23783 17737
rect 23836 17744 23876 18040
rect 24547 17956 24556 17996
rect 24596 17956 24844 17996
rect 24884 17956 24893 17996
rect 24355 17872 24364 17912
rect 24404 17872 24787 17912
rect 24827 17872 24836 17912
rect 24067 17788 24076 17828
rect 24116 17788 24125 17828
rect 24259 17788 24268 17828
rect 24308 17788 25612 17828
rect 25652 17788 25661 17828
rect 24076 17744 24116 17788
rect 25708 17744 25748 18208
rect 26188 17996 26228 18376
rect 30604 18332 30644 18544
rect 30778 18535 30787 18575
rect 30827 18544 31124 18575
rect 30827 18535 30836 18544
rect 30778 18534 30836 18535
rect 27331 18292 27340 18332
rect 27380 18292 27436 18332
rect 27476 18292 27511 18332
rect 28963 18292 28972 18332
rect 29012 18292 30220 18332
rect 30260 18292 30644 18332
rect 30892 18460 30940 18500
rect 30980 18460 30989 18500
rect 30892 18248 30932 18460
rect 26275 18208 26284 18248
rect 26324 18208 30932 18248
rect 31084 18164 31124 18544
rect 26425 18124 26434 18164
rect 26802 18124 26811 18164
rect 27619 18124 27628 18164
rect 27668 18124 31124 18164
rect 25795 17956 25804 17996
rect 25844 17956 25853 17996
rect 26170 17956 26179 17996
rect 26219 17956 26228 17996
rect 27715 17956 27724 17996
rect 27764 17956 30220 17996
rect 30260 17956 30269 17996
rect 25804 17744 25844 17956
rect 27532 17788 27715 17828
rect 27755 17788 27764 17828
rect 27977 17788 28099 17828
rect 28148 17788 28157 17828
rect 29856 17788 30988 17828
rect 31028 17788 31037 17828
rect 27532 17744 27572 17788
rect 23836 17704 23980 17744
rect 24020 17704 24029 17744
rect 24076 17704 24172 17744
rect 24212 17704 24221 17744
rect 24276 17704 24364 17744
rect 24404 17704 24407 17744
rect 24447 17704 24456 17744
rect 24538 17735 24596 17744
rect 22732 17576 22772 17704
rect 22924 17695 22964 17704
rect 23116 17660 23156 17704
rect 23500 17660 23540 17704
rect 23107 17620 23116 17660
rect 23156 17620 23165 17660
rect 23395 17620 23404 17660
rect 23444 17620 23540 17660
rect 23644 17576 23684 17704
rect 24161 17702 24212 17704
rect 24538 17695 24547 17735
rect 24587 17695 24596 17735
rect 24643 17704 24652 17744
rect 24692 17704 24988 17744
rect 25028 17704 25037 17744
rect 25123 17704 25132 17744
rect 25172 17704 25516 17744
rect 25556 17704 25565 17744
rect 25699 17704 25708 17744
rect 25748 17704 25757 17744
rect 25804 17704 25827 17744
rect 25867 17704 25876 17744
rect 25930 17704 25939 17744
rect 25979 17704 25988 17744
rect 26563 17704 26572 17744
rect 26612 17704 26851 17744
rect 26891 17704 26900 17744
rect 27523 17704 27532 17744
rect 27572 17704 27581 17744
rect 29513 17704 29635 17744
rect 29684 17704 29693 17744
rect 30199 17704 30208 17744
rect 30248 17704 30548 17744
rect 30679 17704 30688 17744
rect 30740 17704 30868 17744
rect 24538 17694 24596 17695
rect 24556 17660 24596 17694
rect 25132 17660 25172 17704
rect 25940 17660 25980 17704
rect 30508 17660 30548 17704
rect 23875 17620 23884 17660
rect 23924 17620 24500 17660
rect 24556 17620 25172 17660
rect 25411 17620 25420 17660
rect 25460 17620 25980 17660
rect 29897 17620 30019 17660
rect 30068 17620 30077 17660
rect 30508 17620 30892 17660
rect 30932 17620 30941 17660
rect 24460 17576 24500 17620
rect 22732 17536 23684 17576
rect 23971 17536 23980 17576
rect 24020 17536 24268 17576
rect 24308 17536 24317 17576
rect 24460 17536 26380 17576
rect 26420 17536 26429 17576
rect 26668 17536 30364 17576
rect 30404 17536 30413 17576
rect 30508 17536 30844 17576
rect 30884 17536 30893 17576
rect 22252 17452 23020 17492
rect 23060 17452 23069 17492
rect 23203 17452 23212 17492
rect 23252 17452 26572 17492
rect 26612 17452 26621 17492
rect 26668 17408 26708 17536
rect 30508 17492 30548 17536
rect 26755 17452 26764 17492
rect 26804 17452 30548 17492
rect 15484 17368 16911 17408
rect 4300 17284 5068 17324
rect 5108 17284 5117 17324
rect 6019 17284 6028 17324
rect 6068 17284 6153 17324
rect 7267 17284 7276 17324
rect 7316 17284 8948 17324
rect 11011 17284 11020 17324
rect 11060 17284 12068 17324
rect 12220 17284 14996 17324
rect 4300 17240 4340 17284
rect 1987 17200 1996 17240
rect 2036 17200 2179 17240
rect 2219 17200 2228 17240
rect 3322 17200 3331 17240
rect 3371 17200 4012 17240
rect 4052 17200 4061 17240
rect 4282 17200 4291 17240
rect 4331 17200 4340 17240
rect 4474 17200 4483 17240
rect 4532 17200 4663 17240
rect 4841 17200 4963 17240
rect 5012 17200 5021 17240
rect 6113 17156 6153 17284
rect 6499 17200 6508 17240
rect 6548 17200 7892 17240
rect 8297 17200 8323 17240
rect 8363 17200 8428 17240
rect 8468 17200 8477 17240
rect 8681 17200 8803 17240
rect 8852 17200 8861 17240
rect 3034 17116 3043 17156
rect 3083 17116 3380 17156
rect 3802 17116 3811 17156
rect 3851 17116 4780 17156
rect 4820 17116 4829 17156
rect 5242 17147 5548 17156
rect 3340 17072 3380 17116
rect 5242 17107 5251 17147
rect 5291 17116 5548 17147
rect 5588 17116 5597 17156
rect 6010 17147 6153 17156
rect 5291 17107 5300 17116
rect 5242 17106 5300 17107
rect 6010 17107 6019 17147
rect 6059 17116 6153 17147
rect 6211 17116 6220 17156
rect 6260 17116 6341 17156
rect 6691 17116 6700 17156
rect 6740 17116 7124 17156
rect 7171 17116 7180 17156
rect 7220 17116 7364 17156
rect 6059 17107 6068 17116
rect 6010 17106 6068 17107
rect 6301 17072 6341 17116
rect 7084 17072 7124 17116
rect 2275 17032 2284 17072
rect 2324 17032 2333 17072
rect 3113 17032 3244 17072
rect 3284 17032 3293 17072
rect 3340 17032 3479 17072
rect 3519 17032 3528 17072
rect 3619 17032 3628 17072
rect 3668 17032 3724 17072
rect 3764 17032 3799 17072
rect 4195 17032 4204 17072
rect 4244 17032 4588 17072
rect 4628 17032 4637 17072
rect 4780 17032 4963 17072
rect 5003 17032 5012 17072
rect 5068 17063 5108 17072
rect 2284 16484 2324 17032
rect 3610 16948 3619 16988
rect 3659 16948 4684 16988
rect 4724 16948 4733 16988
rect 4780 16904 4820 17032
rect 5338 17032 5347 17072
rect 5387 17032 5396 17072
rect 5443 17032 5452 17072
rect 5521 17032 5623 17072
rect 5733 17032 5742 17072
rect 5782 17032 5827 17072
rect 5878 17032 5887 17072
rect 5927 17032 5961 17072
rect 6106 17032 6115 17072
rect 6155 17032 6204 17072
rect 6282 17032 6291 17072
rect 6331 17032 6341 17072
rect 5068 16904 5108 17023
rect 5356 16988 5396 17032
rect 5740 16988 5780 17032
rect 5921 16988 5961 17032
rect 5251 16948 5260 16988
rect 5300 16948 5396 16988
rect 5731 16948 5740 16988
rect 5780 16948 5789 16988
rect 5921 16948 5932 16988
rect 5972 16948 5983 16988
rect 6164 16904 6204 17032
rect 6490 17031 6499 17071
rect 6539 17031 6571 17071
rect 6787 17032 6796 17072
rect 6836 17032 6967 17072
rect 7066 17032 7075 17072
rect 7115 17032 7124 17072
rect 7180 17063 7220 17072
rect 6531 16988 6571 17031
rect 6499 16948 6508 16988
rect 6548 16948 6571 16988
rect 7180 16904 7220 17023
rect 7324 17063 7364 17116
rect 7852 17072 7892 17200
rect 8428 17156 8468 17200
rect 8428 17116 8789 17156
rect 8749 17072 8789 17116
rect 8908 17072 8948 17284
rect 12220 17240 12260 17284
rect 16871 17240 16911 17368
rect 18700 17368 19508 17408
rect 19891 17368 19900 17408
rect 20268 17368 20277 17408
rect 22060 17368 22868 17408
rect 22915 17368 22924 17408
rect 22964 17368 26708 17408
rect 27665 17368 27674 17408
rect 28042 17368 28051 17408
rect 18700 17324 18740 17368
rect 22828 17324 22868 17368
rect 16963 17284 16972 17324
rect 17012 17284 18740 17324
rect 20140 17284 22732 17324
rect 22772 17284 22781 17324
rect 22828 17284 23692 17324
rect 23732 17284 23741 17324
rect 23875 17284 23884 17324
rect 23924 17284 28108 17324
rect 28148 17284 28820 17324
rect 20140 17240 20180 17284
rect 9164 17200 9388 17240
rect 9428 17200 10252 17240
rect 10292 17200 10301 17240
rect 10531 17200 10540 17240
rect 10580 17200 12172 17240
rect 12212 17200 12260 17240
rect 12451 17200 12460 17240
rect 12500 17200 12739 17240
rect 12779 17200 13036 17240
rect 13076 17200 13085 17240
rect 13219 17200 13228 17240
rect 13268 17200 13891 17240
rect 13931 17200 13940 17240
rect 15216 17200 15724 17240
rect 15764 17200 15773 17240
rect 15898 17200 15907 17240
rect 15947 17200 15956 17240
rect 16099 17200 16108 17240
rect 16148 17200 16300 17240
rect 16340 17200 16349 17240
rect 16649 17200 16771 17240
rect 16820 17200 16829 17240
rect 16871 17200 17492 17240
rect 17716 17200 17725 17240
rect 17765 17200 18412 17240
rect 18452 17200 18461 17240
rect 18595 17200 18604 17240
rect 18644 17200 18892 17240
rect 18932 17200 18941 17240
rect 19939 17200 19948 17240
rect 19988 17200 20180 17240
rect 20602 17200 20611 17240
rect 20651 17200 20660 17240
rect 20707 17200 20716 17240
rect 20756 17200 21196 17240
rect 21236 17200 21245 17240
rect 21571 17200 21580 17240
rect 21620 17200 21955 17240
rect 21995 17200 22004 17240
rect 22156 17200 24268 17240
rect 24308 17200 24317 17240
rect 25001 17200 25132 17240
rect 25172 17200 25181 17240
rect 26164 17200 26173 17240
rect 26213 17200 26956 17240
rect 26996 17200 27005 17240
rect 27139 17200 27148 17240
rect 27188 17200 27197 17240
rect 27331 17200 27340 17240
rect 27380 17200 27532 17240
rect 27572 17200 27581 17240
rect 8995 17116 9004 17156
rect 9044 17116 9053 17156
rect 7445 17032 7454 17072
rect 7494 17032 7508 17072
rect 7627 17032 7636 17072
rect 7676 17032 7695 17072
rect 7852 17032 7984 17072
rect 8024 17032 8044 17072
rect 8084 17032 8093 17072
rect 8145 17032 8154 17072
rect 8194 17032 8203 17072
rect 8266 17032 8275 17072
rect 8315 17032 8324 17072
rect 7324 17014 7364 17023
rect 7468 16988 7508 17032
rect 7655 16988 7695 17032
rect 8154 16988 8194 17032
rect 8279 16988 8319 17032
rect 8387 17021 8396 17061
rect 8436 17021 8445 17061
rect 8532 17021 8541 17061
rect 8581 17030 8590 17061
rect 8731 17032 8740 17072
rect 8780 17032 8789 17072
rect 8890 17032 8899 17072
rect 8939 17032 8948 17072
rect 9004 17072 9044 17116
rect 9164 17072 9204 17200
rect 9292 17116 9484 17156
rect 9524 17116 9533 17156
rect 9580 17116 10540 17156
rect 10580 17116 10589 17156
rect 11020 17116 11404 17156
rect 11444 17116 11453 17156
rect 12076 17116 13324 17156
rect 13364 17116 13373 17156
rect 13603 17116 13612 17156
rect 13652 17116 13996 17156
rect 14036 17147 14228 17156
rect 14036 17116 14179 17147
rect 9292 17072 9332 17116
rect 9580 17072 9620 17116
rect 11020 17072 11060 17116
rect 12076 17072 12116 17116
rect 14170 17107 14179 17116
rect 14219 17107 14228 17147
rect 14170 17106 14228 17107
rect 9004 17032 9016 17072
rect 9056 17032 9091 17072
rect 9146 17032 9155 17072
rect 9195 17032 9204 17072
rect 9274 17032 9283 17072
rect 9323 17032 9332 17072
rect 9523 17032 9532 17072
rect 9572 17032 9620 17072
rect 9929 17032 10003 17072
rect 10043 17032 10060 17072
rect 10100 17032 10109 17072
rect 10243 17032 10252 17072
rect 10292 17032 10627 17072
rect 10667 17032 10676 17072
rect 11011 17032 11020 17072
rect 11060 17032 11069 17072
rect 11390 17032 11500 17072
rect 11552 17032 11570 17072
rect 11683 17032 11692 17072
rect 11732 17032 11884 17072
rect 11924 17032 11933 17072
rect 12058 17032 12067 17072
rect 12107 17032 12116 17072
rect 12163 17032 12172 17072
rect 12212 17032 12343 17072
rect 12538 17032 12547 17072
rect 12587 17032 12596 17072
rect 12643 17032 12652 17072
rect 12692 17032 12979 17072
rect 13019 17032 13228 17072
rect 13268 17032 13277 17072
rect 13385 17032 13516 17072
rect 13556 17032 13565 17072
rect 13612 17032 13708 17072
rect 13748 17032 13757 17072
rect 13882 17032 13891 17072
rect 13931 17032 13940 17072
rect 8581 17021 8660 17030
rect 7459 16948 7468 16988
rect 7508 16948 7541 16988
rect 7655 16948 7852 16988
rect 7892 16948 7901 16988
rect 8125 16948 8194 16988
rect 8236 16948 8319 16988
rect 7468 16904 7508 16948
rect 8125 16904 8165 16948
rect 4003 16864 4012 16904
rect 4052 16864 4492 16904
rect 4532 16864 4541 16904
rect 4771 16864 4780 16904
rect 4820 16864 4829 16904
rect 5068 16864 6220 16904
rect 6260 16864 6269 16904
rect 7180 16864 7372 16904
rect 7412 16864 7421 16904
rect 7468 16864 8165 16904
rect 8236 16820 8276 16948
rect 8396 16904 8436 17021
rect 8550 16990 8660 17021
rect 8620 16904 8660 16990
rect 8908 16988 8948 17032
rect 9532 16988 9572 17032
rect 9667 16990 9676 17030
rect 9716 16990 9725 17030
rect 8908 16948 9572 16988
rect 8396 16864 8428 16904
rect 8468 16864 8477 16904
rect 8620 16864 8924 16904
rect 2467 16780 2476 16820
rect 2516 16780 2572 16820
rect 2612 16780 2647 16820
rect 5722 16780 5731 16820
rect 5771 16780 5780 16820
rect 6595 16780 6604 16820
rect 6644 16780 7075 16820
rect 7115 16780 7180 16820
rect 7220 16780 7284 16820
rect 7843 16780 7852 16820
rect 7892 16780 8276 16820
rect 5740 16652 5780 16780
rect 3103 16612 3112 16652
rect 3480 16612 3489 16652
rect 3619 16612 3628 16652
rect 3668 16612 5780 16652
rect 6115 16528 6124 16568
rect 6164 16528 8564 16568
rect 8524 16484 8564 16528
rect 8884 16484 8924 16864
rect 9676 16652 9716 16990
rect 12556 16988 12596 17032
rect 13612 16988 13652 17032
rect 13900 16988 13940 17032
rect 13996 17063 14036 17072
rect 14266 17032 14275 17072
rect 14315 17032 14324 17072
rect 14371 17032 14380 17072
rect 14449 17032 14551 17072
rect 15216 17032 15256 17200
rect 15916 17156 15956 17200
rect 17452 17156 17492 17200
rect 20620 17156 20660 17200
rect 22156 17156 22196 17200
rect 15400 17116 15436 17156
rect 15476 17116 15485 17156
rect 15593 17116 15628 17156
rect 15668 17147 15764 17156
rect 15668 17116 15715 17147
rect 15436 17072 15476 17116
rect 15706 17107 15715 17116
rect 15755 17107 15764 17147
rect 15916 17116 16436 17156
rect 16963 17116 16972 17156
rect 17012 17116 17396 17156
rect 17452 17116 17876 17156
rect 15706 17106 15764 17107
rect 16396 17072 16436 17116
rect 17356 17072 17396 17116
rect 17836 17072 17876 17116
rect 15296 17032 15305 17072
rect 15429 17032 15438 17072
rect 15478 17032 15487 17072
rect 15532 17063 15583 17072
rect 9833 16948 9868 16988
rect 9908 16948 9964 16988
rect 10004 16948 10013 16988
rect 10531 16948 10540 16988
rect 10580 16948 10828 16988
rect 10868 16948 11347 16988
rect 11387 16948 11396 16988
rect 12556 16948 13036 16988
rect 13076 16948 13085 16988
rect 13171 16948 13180 16988
rect 13220 16948 13229 16988
rect 13603 16948 13612 16988
rect 13652 16948 13661 16988
rect 13853 16948 13900 16988
rect 13940 16948 13949 16988
rect 9763 16864 9772 16904
rect 9812 16864 9868 16904
rect 9908 16864 9943 16904
rect 12510 16864 12519 16904
rect 12559 16864 12596 16904
rect 10409 16780 10444 16820
rect 10484 16780 10540 16820
rect 10580 16780 10589 16820
rect 11395 16780 11404 16820
rect 11444 16780 12172 16820
rect 12212 16780 12221 16820
rect 9676 16612 10000 16652
rect 10877 16612 10886 16652
rect 11254 16612 11263 16652
rect 9960 16484 10000 16612
rect 12556 16568 12596 16864
rect 13180 16820 13220 16948
rect 13996 16904 14036 17023
rect 14284 16988 14324 17032
rect 15572 17023 15583 17063
rect 15798 17032 15807 17072
rect 15847 17032 15856 17072
rect 15979 17032 15988 17072
rect 16052 17032 16168 17072
rect 16210 17032 16219 17072
rect 16259 17032 16340 17072
rect 16387 17032 16396 17072
rect 16436 17032 16445 17072
rect 16492 17032 16612 17072
rect 16652 17032 16661 17072
rect 16762 17032 16771 17072
rect 16811 17032 16820 17072
rect 16879 17032 16888 17072
rect 16928 17032 16937 17072
rect 17020 17063 17060 17072
rect 15532 17014 15583 17023
rect 14284 16948 14668 16988
rect 14708 16948 14717 16988
rect 15082 16948 15091 16988
rect 15131 16948 15340 16988
rect 15380 16948 15389 16988
rect 15543 16904 15583 17014
rect 15816 16988 15856 17032
rect 16300 16988 16340 17032
rect 16492 16988 16532 17032
rect 16780 16988 16820 17032
rect 15811 16948 15820 16988
rect 15860 16948 15903 16988
rect 16195 16948 16204 16988
rect 16244 16948 16340 16988
rect 16483 16948 16492 16988
rect 16532 16948 16541 16988
rect 16675 16948 16684 16988
rect 16724 16948 16820 16988
rect 13996 16864 14476 16904
rect 14516 16864 16396 16904
rect 16436 16864 16445 16904
rect 13180 16780 14092 16820
rect 14132 16780 14141 16820
rect 16888 16736 16928 17032
rect 17146 17032 17155 17072
rect 17195 17032 17204 17072
rect 17347 17032 17356 17072
rect 17396 17032 17405 17072
rect 17539 17032 17548 17072
rect 17588 17032 17597 17072
rect 17818 17032 17827 17072
rect 17867 17032 17876 17072
rect 17932 17116 18499 17156
rect 18539 17116 18548 17156
rect 18604 17116 19124 17156
rect 19651 17116 19660 17156
rect 19700 17116 19852 17156
rect 19892 17116 19901 17156
rect 20323 17116 20332 17156
rect 20372 17116 20468 17156
rect 20620 17116 21044 17156
rect 21297 17116 21306 17156
rect 21346 17116 22196 17156
rect 22627 17116 22636 17156
rect 22676 17116 23308 17156
rect 23348 17116 23357 17156
rect 17932 17063 17972 17116
rect 18604 17072 18644 17116
rect 19084 17072 19124 17116
rect 20428 17072 20468 17116
rect 21004 17072 21044 17116
rect 23404 17072 23444 17200
rect 27148 17156 27188 17200
rect 23683 17116 23692 17156
rect 23732 17116 23828 17156
rect 23875 17116 23884 17156
rect 23924 17116 24181 17156
rect 23788 17072 23828 17116
rect 24141 17072 24181 17116
rect 24266 17116 24844 17156
rect 24884 17116 24893 17156
rect 25228 17116 26324 17156
rect 26698 17116 26707 17156
rect 26747 17116 27615 17156
rect 27715 17116 27724 17156
rect 27764 17116 27793 17156
rect 24266 17072 24306 17116
rect 25228 17072 25268 17116
rect 26284 17072 26324 17116
rect 27575 17072 27615 17116
rect 27724 17072 27764 17116
rect 28780 17072 28820 17284
rect 29539 17200 29548 17240
rect 29588 17200 29731 17240
rect 29771 17200 29780 17240
rect 29897 17200 30028 17240
rect 30068 17200 30077 17240
rect 29836 17116 31756 17156
rect 31796 17116 31805 17156
rect 29836 17072 29876 17116
rect 17020 16988 17060 17023
rect 17020 16948 17068 16988
rect 17108 16948 17117 16988
rect 17164 16904 17204 17032
rect 17548 16988 17588 17032
rect 18267 17032 18316 17072
rect 18356 17032 18398 17072
rect 18438 17032 18447 17072
rect 18508 17032 18604 17072
rect 18644 17032 18653 17072
rect 18700 17063 18740 17072
rect 17932 17014 17972 17023
rect 17251 16948 17260 16988
rect 17300 16948 17588 16988
rect 17164 16864 17300 16904
rect 18089 16864 18220 16904
rect 18260 16864 18269 16904
rect 12739 16696 12748 16736
rect 12788 16696 16928 16736
rect 13123 16612 13132 16652
rect 13172 16612 13516 16652
rect 13556 16612 13565 16652
rect 13900 16612 16204 16652
rect 16244 16612 16253 16652
rect 13900 16568 13940 16612
rect 10051 16528 10060 16568
rect 10100 16528 10580 16568
rect 11971 16528 11980 16568
rect 12020 16528 13900 16568
rect 13940 16528 13949 16568
rect 1507 16444 1516 16484
rect 1556 16444 2324 16484
rect 3619 16444 3628 16484
rect 3668 16444 4876 16484
rect 4916 16444 4925 16484
rect 5452 16444 5836 16484
rect 5876 16444 5885 16484
rect 6979 16444 6988 16484
rect 7028 16444 8372 16484
rect 8515 16444 8524 16484
rect 8564 16444 8573 16484
rect 8884 16444 8899 16484
rect 8939 16444 8948 16484
rect 9187 16444 9196 16484
rect 9236 16444 9245 16484
rect 9292 16444 9676 16484
rect 9716 16444 9725 16484
rect 9960 16444 10100 16484
rect 1420 16276 2188 16316
rect 2228 16276 2237 16316
rect 1420 16232 1460 16276
rect 2284 16232 2324 16444
rect 3340 16360 5356 16400
rect 5396 16360 5405 16400
rect 3340 16232 3380 16360
rect 5452 16316 5492 16444
rect 8332 16400 8372 16444
rect 9196 16400 9236 16444
rect 9292 16400 9332 16444
rect 10060 16400 10100 16444
rect 5539 16360 5548 16400
rect 5588 16360 5597 16400
rect 5896 16360 6220 16400
rect 6260 16360 6269 16400
rect 6700 16360 8276 16400
rect 8332 16360 8756 16400
rect 4042 16307 5492 16316
rect 4042 16267 4051 16307
rect 4091 16276 5492 16307
rect 4091 16267 4100 16276
rect 4042 16266 4100 16267
rect 5548 16232 5588 16360
rect 5896 16316 5936 16360
rect 6700 16316 6740 16360
rect 5884 16276 5936 16316
rect 5990 16276 6028 16316
rect 6068 16276 6077 16316
rect 6691 16276 6700 16316
rect 6740 16276 6749 16316
rect 7166 16276 7180 16316
rect 7220 16276 7229 16316
rect 7485 16276 7564 16316
rect 7604 16276 8044 16316
rect 8084 16276 8093 16316
rect 5884 16232 5924 16276
rect 5990 16232 6030 16276
rect 7180 16232 7220 16276
rect 7645 16232 7685 16276
rect 8236 16232 8276 16360
rect 8416 16276 8428 16316
rect 8468 16276 8477 16316
rect 8416 16232 8456 16276
rect 8716 16232 8756 16360
rect 8908 16360 9236 16400
rect 9283 16360 9292 16400
rect 9332 16360 9341 16400
rect 9475 16360 9484 16400
rect 9524 16360 10016 16400
rect 10060 16360 10484 16400
rect 8908 16232 8948 16360
rect 9976 16316 10016 16360
rect 10444 16316 10484 16360
rect 10540 16316 10580 16528
rect 17260 16484 17300 16864
rect 18508 16820 18548 17032
rect 17443 16780 17452 16820
rect 17492 16780 18548 16820
rect 18804 17032 18892 17072
rect 18932 17032 18935 17072
rect 18975 17032 18984 17072
rect 19066 17063 19124 17072
rect 18700 16904 18740 17023
rect 19066 17023 19075 17063
rect 19115 17023 19124 17063
rect 19171 17032 19180 17072
rect 19220 17032 19229 17072
rect 19363 17032 19372 17072
rect 19412 17032 19468 17072
rect 19508 17032 19543 17072
rect 19786 17032 19795 17072
rect 19835 17032 19844 17072
rect 20138 17032 20236 17072
rect 20300 17032 20318 17072
rect 20410 17032 20419 17072
rect 20459 17032 20468 17072
rect 20524 17032 20536 17072
rect 20576 17032 20585 17072
rect 20631 17063 20708 17072
rect 19066 17022 19124 17023
rect 19180 16904 19220 17032
rect 19804 16988 19844 17032
rect 19804 16948 20332 16988
rect 20372 16948 20381 16988
rect 20524 16904 20564 17032
rect 18700 16864 19220 16904
rect 20131 16864 20140 16904
rect 20180 16864 20564 16904
rect 20631 17023 20668 17063
rect 20794 17032 20803 17072
rect 20843 17032 20899 17072
rect 20986 17032 20995 17072
rect 21035 17032 21044 17072
rect 21091 17032 21100 17072
rect 21140 17032 21271 17072
rect 21676 17032 21868 17072
rect 21908 17032 21917 17072
rect 22051 17032 22060 17072
rect 22100 17032 22156 17072
rect 22196 17032 22231 17072
rect 22409 17032 22540 17072
rect 22580 17032 22589 17072
rect 22819 17032 22828 17072
rect 22868 17032 22877 17072
rect 23011 17032 23020 17072
rect 23060 17032 23191 17072
rect 23350 17032 23359 17072
rect 23399 17032 23444 17072
rect 23491 17032 23500 17072
rect 23540 17032 23596 17072
rect 23636 17032 23671 17072
rect 23779 17032 23788 17072
rect 23828 17032 23837 17072
rect 24126 17032 24135 17072
rect 24175 17032 24184 17072
rect 24250 17063 24308 17072
rect 20631 17014 20708 17023
rect 20631 16904 20671 17014
rect 20812 16988 20852 17032
rect 21676 16988 21716 17032
rect 22540 16988 22580 17032
rect 20803 16948 20812 16988
rect 20852 16948 20861 16988
rect 20908 16948 21580 16988
rect 21620 16948 21629 16988
rect 21676 16948 21964 16988
rect 22004 16948 22013 16988
rect 22147 16948 22156 16988
rect 22196 16948 22580 16988
rect 22828 16988 22868 17032
rect 24250 17023 24259 17063
rect 24299 17023 24308 17063
rect 24355 17032 24364 17072
rect 24408 17032 24535 17072
rect 24643 17032 24652 17072
rect 24692 17032 24701 17072
rect 24768 17032 24777 17072
rect 24817 17032 24884 17072
rect 24931 17032 24940 17072
rect 24980 17032 25228 17072
rect 25268 17032 25277 17072
rect 25456 17032 25465 17072
rect 25505 17032 25708 17072
rect 25748 17032 25757 17072
rect 25804 17032 25830 17072
rect 25870 17032 25891 17072
rect 25948 17032 25957 17072
rect 25997 17032 26057 17072
rect 26124 17032 26188 17072
rect 26228 17032 26275 17072
rect 26315 17032 26324 17072
rect 26380 17063 26420 17072
rect 24250 17022 24308 17023
rect 22828 16948 22924 16988
rect 22964 16948 22973 16988
rect 23107 16948 23116 16988
rect 23156 16948 23242 16988
rect 23282 16948 23692 16988
rect 23732 16948 23741 16988
rect 20908 16904 20948 16948
rect 20631 16864 20948 16904
rect 21353 16864 21484 16904
rect 21524 16864 21533 16904
rect 18700 16736 18740 16864
rect 19651 16780 19660 16820
rect 19700 16780 21580 16820
rect 21620 16780 21629 16820
rect 21676 16736 21716 16948
rect 24652 16904 24692 17032
rect 24844 16988 24884 17032
rect 25804 16988 25844 17032
rect 26017 16988 26057 17032
rect 26921 17032 27052 17072
rect 27092 17032 27101 17072
rect 27148 17032 27173 17072
rect 27213 17032 27222 17072
rect 27566 17032 27575 17072
rect 27615 17032 27624 17072
rect 27688 17032 27697 17072
rect 27737 17032 27764 17072
rect 27811 17032 27820 17072
rect 27860 17032 27869 17072
rect 28003 17032 28012 17072
rect 28052 17032 28684 17072
rect 28724 17032 28733 17072
rect 28780 17032 28876 17072
rect 28916 17032 28925 17072
rect 29731 17032 29740 17072
rect 29780 17032 29836 17072
rect 29876 17032 29911 17072
rect 30089 17032 30220 17072
rect 30260 17032 30269 17072
rect 24844 16948 25132 16988
rect 25172 16948 25181 16988
rect 25354 16979 25612 16988
rect 25354 16939 25363 16979
rect 25403 16948 25612 16979
rect 25652 16948 25661 16988
rect 25795 16948 25804 16988
rect 25844 16948 25853 16988
rect 26017 16948 26284 16988
rect 26324 16948 26333 16988
rect 25403 16939 25412 16948
rect 25354 16938 25412 16939
rect 22819 16864 22828 16904
rect 22868 16864 23020 16904
rect 23060 16864 23116 16904
rect 23156 16864 23165 16904
rect 23395 16864 23404 16904
rect 23444 16864 24692 16904
rect 24739 16864 24748 16904
rect 24788 16864 24919 16904
rect 26380 16820 26420 17023
rect 27148 16988 27188 17032
rect 27148 16948 27436 16988
rect 27476 16948 27485 16988
rect 27820 16904 27860 17032
rect 28291 16948 28300 16988
rect 28340 16948 30740 16988
rect 26842 16864 26851 16904
rect 26891 16864 26900 16904
rect 27043 16864 27052 16904
rect 27092 16864 27860 16904
rect 27916 16864 28204 16904
rect 28244 16864 28253 16904
rect 29923 16864 29932 16904
rect 29972 16864 30604 16904
rect 30644 16864 30653 16904
rect 23587 16780 23596 16820
rect 23636 16780 23980 16820
rect 24020 16780 24029 16820
rect 25987 16780 25996 16820
rect 26036 16780 26045 16820
rect 26284 16780 26420 16820
rect 26860 16820 26900 16864
rect 27916 16820 27956 16864
rect 30700 16820 30740 16948
rect 30857 16864 30988 16904
rect 31028 16864 31037 16904
rect 26860 16780 27956 16820
rect 28003 16780 28012 16820
rect 28052 16780 28108 16820
rect 28148 16780 28183 16820
rect 30307 16780 30316 16820
rect 30356 16780 30365 16820
rect 30700 16780 30932 16820
rect 18508 16696 18740 16736
rect 20323 16696 20332 16736
rect 20372 16696 21716 16736
rect 15235 16444 15244 16484
rect 15284 16444 15764 16484
rect 17251 16444 17260 16484
rect 17300 16444 17309 16484
rect 17923 16444 17932 16484
rect 17972 16444 18316 16484
rect 18356 16444 18365 16484
rect 15724 16400 15764 16444
rect 18508 16400 18548 16696
rect 18651 16612 18660 16652
rect 19028 16612 19037 16652
rect 19363 16612 19372 16652
rect 19412 16612 22060 16652
rect 22100 16612 22109 16652
rect 20044 16444 20236 16484
rect 20276 16444 21196 16484
rect 21236 16444 21245 16484
rect 23779 16444 23788 16484
rect 23828 16444 24076 16484
rect 24116 16444 24125 16484
rect 25123 16444 25132 16484
rect 25172 16444 25411 16484
rect 25451 16444 25460 16484
rect 15017 16360 15052 16400
rect 15092 16360 15148 16400
rect 15188 16360 15197 16400
rect 15715 16360 15724 16400
rect 15764 16360 15773 16400
rect 16387 16360 16396 16400
rect 16436 16360 18548 16400
rect 18979 16360 18988 16400
rect 19028 16360 19412 16400
rect 9259 16276 9388 16316
rect 9430 16276 9439 16316
rect 9976 16276 10148 16316
rect 10243 16276 10252 16316
rect 10292 16276 10301 16316
rect 10435 16276 10444 16316
rect 10484 16276 10493 16316
rect 10540 16276 10659 16316
rect 10699 16276 10708 16316
rect 11107 16276 11116 16316
rect 11156 16276 11308 16316
rect 11348 16276 11357 16316
rect 11500 16276 11828 16316
rect 12617 16276 12700 16316
rect 12740 16276 12748 16316
rect 12788 16276 12797 16316
rect 13315 16276 13324 16316
rect 13364 16276 13652 16316
rect 14275 16276 14284 16316
rect 14324 16276 14420 16316
rect 14467 16276 14476 16316
rect 14516 16276 15052 16316
rect 15092 16276 15244 16316
rect 15284 16276 15293 16316
rect 15340 16276 15436 16316
rect 15476 16276 15628 16316
rect 15668 16276 15677 16316
rect 15820 16276 16108 16316
rect 16148 16276 16361 16316
rect 16483 16276 16492 16316
rect 16532 16276 16684 16316
rect 16724 16276 16733 16316
rect 16841 16276 16924 16316
rect 16964 16276 16972 16316
rect 17012 16276 17021 16316
rect 17635 16276 17644 16316
rect 17684 16276 17972 16316
rect 19145 16276 19276 16316
rect 19316 16276 19325 16316
rect 1411 16192 1420 16232
rect 1460 16192 1469 16232
rect 1612 16165 1621 16205
rect 1661 16165 1700 16205
rect 1834 16192 1843 16232
rect 1883 16192 1996 16232
rect 2036 16192 2045 16232
rect 2179 16192 2188 16232
rect 2228 16192 2324 16232
rect 2476 16192 2755 16232
rect 2795 16192 2804 16232
rect 2851 16192 2860 16232
rect 2900 16192 3380 16232
rect 3427 16192 3436 16232
rect 3476 16192 3628 16232
rect 3668 16192 3677 16232
rect 3907 16192 3916 16232
rect 3956 16192 3965 16232
rect 4144 16192 4153 16232
rect 4193 16192 4340 16232
rect 4483 16192 4492 16232
rect 4532 16192 4972 16232
rect 5012 16192 5021 16232
rect 5225 16192 5356 16232
rect 5396 16192 5405 16232
rect 5548 16192 5731 16232
rect 5771 16192 5780 16232
rect 5866 16192 5875 16232
rect 5915 16192 5924 16232
rect 5972 16192 5981 16232
rect 6021 16192 6030 16232
rect 6076 16192 6101 16232
rect 6141 16192 6150 16232
rect 6211 16192 6220 16232
rect 6289 16192 6508 16232
rect 6548 16192 6557 16232
rect 6665 16192 6796 16232
rect 6836 16192 6845 16232
rect 6892 16192 6915 16232
rect 6955 16192 6964 16232
rect 7024 16192 7033 16232
rect 7073 16192 7082 16232
rect 7180 16192 7204 16232
rect 7244 16192 7253 16232
rect 7354 16192 7363 16232
rect 7403 16192 7412 16232
rect 7480 16192 7489 16232
rect 7529 16192 7538 16232
rect 7637 16192 7646 16232
rect 7686 16192 7695 16232
rect 7738 16192 7747 16232
rect 7787 16192 7852 16232
rect 7892 16192 7927 16232
rect 7978 16192 7987 16232
rect 8027 16192 8036 16232
rect 8122 16192 8131 16232
rect 8171 16192 8180 16232
rect 8236 16192 8248 16232
rect 8288 16192 8297 16232
rect 8378 16192 8387 16232
rect 8427 16192 8456 16232
rect 8502 16192 8515 16232
rect 8555 16192 8564 16232
rect 8707 16192 8716 16232
rect 8756 16192 8765 16232
rect 8890 16192 8899 16232
rect 8939 16192 8948 16232
rect 9004 16192 9052 16232
rect 9092 16192 9101 16232
rect 9208 16192 9217 16232
rect 9257 16192 9266 16232
rect 9426 16192 9509 16232
rect 9549 16192 9558 16232
rect 1660 16148 1700 16165
rect 1660 16108 1804 16148
rect 1844 16108 1853 16148
rect 2476 16064 2516 16192
rect 3916 16148 3956 16192
rect 4300 16148 4340 16192
rect 6076 16148 6116 16192
rect 3331 16108 3340 16148
rect 3380 16108 3820 16148
rect 3860 16108 3869 16148
rect 3916 16108 4108 16148
rect 4148 16108 4157 16148
rect 4282 16108 4291 16148
rect 4331 16108 4340 16148
rect 4579 16108 4588 16148
rect 4628 16108 5300 16148
rect 5923 16108 5932 16148
rect 5972 16108 6116 16148
rect 5260 16064 5300 16108
rect 6892 16064 6932 16192
rect 7042 16148 7082 16192
rect 7372 16148 7412 16192
rect 7042 16108 7084 16148
rect 7124 16108 7133 16148
rect 7235 16108 7412 16148
rect 7493 16148 7533 16192
rect 7996 16148 8036 16192
rect 7493 16108 7564 16148
rect 7604 16108 7613 16148
rect 7996 16108 8044 16148
rect 8084 16108 8093 16148
rect 2275 16024 2284 16064
rect 2324 16024 2516 16064
rect 3139 16024 3148 16064
rect 3188 16024 3197 16064
rect 3322 16024 3331 16064
rect 3371 16024 4012 16064
rect 4052 16024 4579 16064
rect 4619 16024 4684 16064
rect 4724 16024 4733 16064
rect 5129 16024 5251 16064
rect 5300 16024 5309 16064
rect 6202 16024 6211 16064
rect 6251 16024 6700 16064
rect 6740 16024 6932 16064
rect 67 15772 76 15812
rect 116 15772 500 15812
rect 0 15644 400 15664
rect 460 15644 500 15772
rect 2380 15728 2420 16024
rect 3148 15980 3188 16024
rect 7235 15980 7275 16108
rect 7354 16024 7363 16064
rect 7403 16024 7948 16064
rect 7988 16024 7997 16064
rect 8140 15980 8180 16192
rect 8502 16148 8542 16192
rect 9004 16148 9044 16192
rect 9217 16148 9257 16192
rect 9426 16148 9466 16192
rect 8419 16108 8428 16148
rect 8468 16108 8542 16148
rect 8707 16108 8716 16148
rect 8756 16108 9044 16148
rect 9091 16108 9100 16148
rect 9140 16108 9257 16148
rect 9315 16108 9466 16148
rect 9652 16148 9692 16243
rect 9732 16203 9741 16243
rect 10108 16232 10148 16276
rect 10252 16232 10292 16276
rect 11500 16232 11540 16276
rect 11788 16232 11828 16276
rect 13612 16232 13652 16276
rect 14380 16232 14420 16276
rect 15340 16232 15380 16276
rect 15820 16232 15860 16276
rect 16321 16232 16361 16276
rect 17932 16274 17972 16276
rect 17932 16265 18015 16274
rect 17932 16234 17975 16265
rect 9864 16192 9873 16232
rect 9913 16192 9922 16232
rect 9994 16205 10003 16232
rect 9976 16192 10003 16205
rect 10043 16192 10052 16232
rect 9652 16108 9676 16148
rect 9716 16108 9725 16148
rect 9315 16064 9355 16108
rect 9868 16064 9908 16192
rect 9976 16165 10052 16192
rect 10234 16192 10243 16232
rect 10283 16192 10339 16232
rect 10531 16192 10540 16232
rect 10580 16192 10589 16232
rect 10768 16192 10777 16232
rect 10817 16192 10868 16232
rect 10915 16192 10924 16232
rect 10964 16192 11212 16232
rect 11252 16192 11261 16232
rect 11308 16192 11331 16232
rect 11371 16192 11380 16232
rect 11424 16192 11449 16232
rect 11489 16192 11540 16232
rect 11587 16192 11596 16232
rect 11636 16192 11645 16232
rect 11779 16192 11788 16232
rect 11828 16192 12076 16232
rect 12116 16192 12125 16232
rect 12535 16192 12544 16232
rect 12584 16192 13228 16232
rect 13268 16192 13277 16232
rect 13453 16192 13462 16232
rect 13502 16192 13511 16232
rect 13603 16192 13612 16232
rect 13652 16192 13661 16232
rect 13769 16192 13900 16232
rect 13940 16192 13949 16232
rect 14266 16192 14275 16232
rect 14315 16192 14324 16232
rect 14380 16192 14572 16232
rect 14612 16192 14621 16232
rect 14899 16192 14908 16232
rect 14948 16192 14957 16232
rect 15092 16192 15148 16232
rect 15188 16192 15223 16232
rect 15263 16192 15295 16232
rect 15340 16192 15363 16232
rect 15403 16192 15412 16232
rect 15475 16192 15484 16232
rect 15524 16192 15533 16232
rect 15619 16192 15628 16232
rect 15668 16192 15785 16232
rect 15825 16192 15860 16232
rect 15946 16192 15955 16232
rect 15995 16192 16156 16232
rect 16196 16192 16204 16232
rect 16244 16192 16253 16232
rect 16312 16192 16321 16232
rect 16361 16192 16370 16232
rect 16588 16192 16613 16232
rect 16653 16192 16662 16232
rect 16759 16192 16768 16232
rect 16808 16192 16817 16232
rect 16867 16192 16876 16232
rect 16916 16192 17452 16232
rect 17492 16192 17501 16232
rect 17827 16192 17836 16232
rect 17876 16192 17885 16232
rect 19372 16232 19412 16360
rect 19747 16276 19756 16316
rect 19796 16276 19948 16316
rect 19988 16276 19997 16316
rect 20044 16232 20084 16444
rect 22243 16360 22252 16400
rect 22292 16360 22301 16400
rect 25027 16360 25036 16400
rect 25076 16360 25268 16400
rect 21475 16276 21484 16316
rect 21524 16276 21533 16316
rect 21737 16276 21868 16316
rect 21908 16276 21917 16316
rect 22252 16232 22292 16360
rect 25057 16276 25132 16316
rect 25172 16276 25181 16316
rect 25057 16274 25097 16276
rect 25036 16265 25097 16274
rect 17975 16216 18015 16225
rect 18307 16192 18316 16232
rect 18356 16192 18595 16232
rect 18635 16192 19180 16232
rect 19220 16192 19229 16232
rect 19363 16192 19372 16232
rect 19412 16192 19421 16232
rect 19468 16192 19491 16232
rect 19531 16192 19540 16232
rect 19597 16192 19606 16232
rect 19646 16192 20084 16232
rect 20236 16192 20323 16232
rect 20363 16192 20372 16232
rect 22252 16192 22387 16232
rect 22427 16192 22436 16232
rect 22915 16192 22924 16232
rect 22964 16192 23060 16232
rect 23107 16192 23116 16232
rect 23156 16192 23252 16232
rect 23299 16192 23308 16232
rect 23348 16192 23596 16232
rect 23636 16192 23645 16232
rect 23779 16192 23788 16232
rect 23828 16192 23959 16232
rect 24067 16192 24076 16232
rect 24116 16192 24212 16232
rect 24259 16192 24268 16232
rect 24308 16192 24439 16232
rect 24607 16192 24652 16232
rect 24692 16192 24738 16232
rect 24778 16192 24787 16232
rect 24922 16203 24931 16232
rect 24971 16203 24980 16232
rect 25076 16234 25097 16265
rect 25228 16232 25268 16360
rect 25996 16316 26036 16780
rect 26284 16736 26324 16780
rect 26275 16696 26284 16736
rect 26324 16696 26333 16736
rect 30316 16652 30356 16780
rect 26425 16612 26434 16652
rect 26802 16612 26811 16652
rect 26947 16612 26956 16652
rect 26996 16612 30356 16652
rect 27523 16528 27532 16568
rect 27572 16528 30836 16568
rect 30796 16484 30836 16528
rect 27427 16444 27436 16484
rect 27476 16444 30068 16484
rect 30787 16444 30796 16484
rect 30836 16444 30845 16484
rect 26380 16360 27052 16400
rect 27092 16360 27101 16400
rect 26380 16316 26420 16360
rect 30028 16316 30068 16444
rect 30892 16400 30932 16780
rect 30211 16360 30220 16400
rect 30260 16360 30316 16400
rect 30356 16360 30391 16400
rect 30700 16360 30932 16400
rect 25507 16276 25516 16316
rect 25556 16276 25756 16316
rect 25796 16276 25805 16316
rect 25996 16276 26179 16316
rect 26219 16276 26228 16316
rect 26371 16276 26380 16316
rect 26420 16276 26429 16316
rect 26956 16276 27340 16316
rect 27380 16276 27389 16316
rect 28073 16276 28195 16316
rect 28244 16276 28253 16316
rect 29923 16276 29932 16316
rect 29972 16276 29981 16316
rect 30028 16276 30115 16316
rect 30155 16276 30164 16316
rect 25402 16234 25411 16274
rect 25451 16234 25460 16274
rect 25036 16216 25076 16225
rect 24838 16192 24931 16203
rect 10108 16183 10148 16192
rect 9976 16148 10016 16165
rect 10540 16148 10580 16192
rect 10828 16148 10868 16192
rect 11308 16148 11348 16192
rect 11500 16148 11540 16192
rect 11596 16148 11636 16192
rect 13471 16148 13511 16192
rect 14284 16148 14324 16192
rect 14908 16148 14948 16192
rect 9955 16108 9964 16148
rect 10004 16108 10016 16148
rect 10243 16108 10252 16148
rect 10292 16108 10580 16148
rect 10819 16108 10828 16148
rect 10868 16108 10877 16148
rect 11284 16108 11308 16148
rect 11348 16108 11357 16148
rect 11491 16108 11500 16148
rect 11540 16108 11549 16148
rect 11596 16108 12460 16148
rect 12500 16108 12509 16148
rect 12739 16108 12748 16148
rect 12788 16108 12797 16148
rect 13471 16108 13708 16148
rect 13748 16108 13804 16148
rect 13844 16108 14324 16148
rect 14380 16108 14948 16148
rect 15255 16148 15295 16192
rect 15484 16148 15524 16192
rect 16588 16148 16628 16192
rect 15255 16108 15524 16148
rect 16387 16108 16396 16148
rect 16436 16108 16628 16148
rect 16777 16148 16817 16192
rect 17836 16148 17876 16192
rect 19468 16148 19508 16192
rect 19607 16148 19647 16192
rect 16777 16108 16972 16148
rect 17012 16108 17021 16148
rect 17836 16108 17932 16148
rect 17972 16108 17981 16148
rect 18124 16108 19508 16148
rect 19555 16108 19564 16148
rect 19604 16108 19647 16148
rect 12748 16064 12788 16108
rect 14380 16064 14420 16108
rect 3148 15940 6836 15980
rect 7145 15940 7276 15980
rect 7316 15940 8180 15980
rect 9100 16024 9355 16064
rect 9475 16024 9484 16064
rect 9524 16024 9763 16064
rect 9803 16024 9812 16064
rect 9868 16024 10444 16064
rect 10484 16024 10493 16064
rect 11683 16024 11692 16064
rect 11732 16024 11741 16064
rect 11788 16024 12788 16064
rect 13258 16024 13267 16064
rect 13307 16024 14420 16064
rect 14467 16024 14476 16064
rect 14516 16024 14525 16064
rect 4343 15856 4352 15896
rect 4720 15856 4729 15896
rect 3916 15772 4012 15812
rect 4052 15772 4061 15812
rect 4108 15772 5164 15812
rect 5204 15772 5213 15812
rect 3916 15728 3956 15772
rect 4108 15728 4148 15772
rect 6796 15728 6836 15940
rect 6883 15856 6892 15896
rect 6932 15856 8660 15896
rect 8620 15812 8660 15856
rect 9100 15812 9140 16024
rect 11692 15896 11732 16024
rect 9283 15856 9292 15896
rect 9332 15856 11404 15896
rect 11444 15856 11453 15896
rect 11500 15856 11732 15896
rect 8620 15772 8948 15812
rect 9100 15772 10503 15812
rect 10915 15772 10924 15812
rect 10964 15772 10973 15812
rect 7738 15730 7747 15770
rect 7787 15730 7802 15770
rect 7762 15728 7802 15730
rect 1865 15688 1996 15728
rect 2036 15688 2045 15728
rect 2356 15688 2365 15728
rect 2405 15688 2420 15728
rect 3401 15688 3427 15728
rect 3467 15688 3532 15728
rect 3572 15688 3581 15728
rect 3898 15688 3907 15728
rect 3947 15688 3956 15728
rect 4099 15688 4108 15728
rect 4148 15688 4157 15728
rect 4588 15688 4876 15728
rect 4916 15688 4925 15728
rect 5059 15688 5068 15728
rect 5108 15688 5251 15728
rect 5291 15688 5300 15728
rect 5347 15688 5356 15728
rect 5396 15688 5443 15728
rect 5483 15688 5527 15728
rect 6796 15688 7220 15728
rect 7354 15688 7363 15728
rect 7403 15688 7564 15728
rect 7604 15688 7613 15728
rect 7762 15688 8812 15728
rect 8852 15688 8861 15728
rect 0 15604 500 15644
rect 2476 15604 2860 15644
rect 2900 15604 2909 15644
rect 3610 15604 3619 15644
rect 3659 15604 4340 15644
rect 0 15584 400 15604
rect 2476 15560 2516 15604
rect 4300 15560 4340 15604
rect 4450 15604 4492 15644
rect 4532 15604 4541 15644
rect 4450 15560 4490 15604
rect 4588 15560 4628 15688
rect 4675 15604 4684 15644
rect 4724 15604 4916 15644
rect 4963 15604 4972 15644
rect 5012 15604 5452 15644
rect 5492 15604 5501 15644
rect 5548 15604 6220 15644
rect 6260 15604 6269 15644
rect 6883 15604 6892 15644
rect 6932 15604 7076 15644
rect 4876 15560 4916 15604
rect 5548 15560 5588 15604
rect 7036 15560 7076 15604
rect 7180 15560 7220 15688
rect 7651 15604 7660 15644
rect 7700 15604 7802 15644
rect 7762 15602 7802 15604
rect 7762 15562 7784 15602
rect 7824 15562 7833 15602
rect 8908 15560 8948 15772
rect 9292 15688 10060 15728
rect 10100 15688 10109 15728
rect 9292 15560 9332 15688
rect 10463 15644 10503 15772
rect 10924 15686 10964 15772
rect 11500 15728 11540 15856
rect 11788 15812 11828 16024
rect 13276 15980 13316 16024
rect 12739 15940 12748 15980
rect 12788 15940 13316 15980
rect 14476 15896 14516 16024
rect 14908 15896 14948 16108
rect 16588 16064 16628 16108
rect 18124 16064 18164 16108
rect 16588 16024 17260 16064
rect 17300 16024 17539 16064
rect 17579 16024 17588 16064
rect 18115 16024 18124 16064
rect 18164 16024 18173 16064
rect 18595 16024 18604 16064
rect 18644 16024 18796 16064
rect 18836 16024 18845 16064
rect 20236 15980 20276 16192
rect 23020 16148 23060 16192
rect 23212 16148 23252 16192
rect 24172 16148 24212 16192
rect 24838 16163 24940 16192
rect 24980 16163 24989 16203
rect 25219 16192 25228 16232
rect 25268 16192 25277 16232
rect 25420 16148 25460 16234
rect 26956 16232 26996 16276
rect 30700 16232 30740 16360
rect 31075 16276 31084 16316
rect 31124 16276 31133 16316
rect 31084 16232 31124 16276
rect 25591 16192 25600 16232
rect 25640 16192 25804 16232
rect 25844 16192 25853 16232
rect 26050 16192 26059 16232
rect 26099 16192 26228 16232
rect 26275 16192 26284 16232
rect 26324 16192 26455 16232
rect 26650 16223 26668 16232
rect 26188 16148 26228 16192
rect 26650 16183 26659 16223
rect 26708 16192 26839 16232
rect 26947 16192 26956 16232
rect 26996 16192 27005 16232
rect 27305 16192 27436 16232
rect 27476 16192 27485 16232
rect 27619 16192 27628 16232
rect 27668 16192 27677 16232
rect 29580 16192 29644 16232
rect 29684 16192 29731 16232
rect 29771 16192 29876 16232
rect 30691 16192 30700 16232
rect 30740 16192 30749 16232
rect 30883 16192 30892 16232
rect 30932 16192 30941 16232
rect 31037 16192 31073 16232
rect 31113 16192 31124 16232
rect 31267 16192 31276 16232
rect 31316 16192 31756 16232
rect 31796 16192 31805 16232
rect 26699 16183 26708 16192
rect 26650 16182 26708 16183
rect 27628 16148 27668 16192
rect 22051 16108 22060 16148
rect 22100 16108 22588 16148
rect 22628 16108 22637 16148
rect 23020 16108 23116 16148
rect 23156 16108 23165 16148
rect 23212 16108 23404 16148
rect 23444 16108 23453 16148
rect 24163 16108 24172 16148
rect 24212 16108 24221 16148
rect 25411 16108 25420 16148
rect 25460 16108 25469 16148
rect 26179 16108 26188 16148
rect 26228 16108 26237 16148
rect 26755 16108 26764 16148
rect 26804 16108 29164 16148
rect 29204 16108 29213 16148
rect 22723 16024 22732 16064
rect 22772 16024 23020 16064
rect 23060 16024 23069 16064
rect 23465 16024 23596 16064
rect 23636 16024 23645 16064
rect 25603 16024 25612 16064
rect 25652 16024 27052 16064
rect 27092 16024 27820 16064
rect 27860 16024 28012 16064
rect 28052 16024 28061 16064
rect 29836 15980 29876 16192
rect 30892 16148 30932 16192
rect 30499 16108 30508 16148
rect 30548 16108 30796 16148
rect 30836 16108 30932 16148
rect 31075 16024 31084 16064
rect 31124 16024 31133 16064
rect 15331 15940 15340 15980
rect 15380 15940 20276 15980
rect 27139 15940 27148 15980
rect 27188 15940 29780 15980
rect 29836 15940 30700 15980
rect 30740 15940 30749 15980
rect 29740 15896 29780 15940
rect 31084 15896 31124 16024
rect 11971 15856 11980 15896
rect 12020 15856 12029 15896
rect 12117 15856 12126 15896
rect 12494 15856 12503 15896
rect 14476 15856 14764 15896
rect 14804 15856 14813 15896
rect 14908 15856 15628 15896
rect 15668 15856 15677 15896
rect 17443 15856 17452 15896
rect 17492 15856 17501 15896
rect 17923 15856 17932 15896
rect 17972 15856 18316 15896
rect 18356 15856 18365 15896
rect 19891 15856 19900 15896
rect 20268 15856 20277 15896
rect 27665 15856 27674 15896
rect 28042 15856 28051 15896
rect 29740 15856 31124 15896
rect 11404 15688 11540 15728
rect 11596 15772 11828 15812
rect 11980 15812 12020 15856
rect 11980 15772 12043 15812
rect 10924 15646 10936 15686
rect 10976 15646 10985 15686
rect 11404 15644 11444 15688
rect 11596 15644 11636 15772
rect 11770 15688 11779 15728
rect 11828 15688 11959 15728
rect 12003 15644 12043 15772
rect 12940 15772 14476 15812
rect 14516 15772 14525 15812
rect 15235 15772 15244 15812
rect 15284 15772 16876 15812
rect 16916 15772 16925 15812
rect 12940 15728 12980 15772
rect 12163 15688 12172 15728
rect 12212 15688 12980 15728
rect 9571 15604 9580 15644
rect 9620 15604 9676 15644
rect 9716 15604 9751 15644
rect 9859 15604 9868 15644
rect 9908 15604 10291 15644
rect 10331 15604 10340 15644
rect 10463 15604 10882 15644
rect 10463 15560 10503 15604
rect 10842 15602 10882 15604
rect 11308 15604 11444 15644
rect 11578 15635 11636 15644
rect 10842 15587 10976 15602
rect 10842 15562 11046 15587
rect 10936 15560 11046 15562
rect 11308 15560 11348 15604
rect 11578 15595 11587 15635
rect 11627 15595 11636 15635
rect 11578 15594 11636 15595
rect 11692 15604 12043 15644
rect 12355 15604 12364 15644
rect 12404 15604 12940 15644
rect 12980 15604 12989 15644
rect 11692 15560 11732 15604
rect 12610 15560 12650 15604
rect 1594 15520 1603 15560
rect 1643 15520 1652 15560
rect 1699 15520 1708 15560
rect 1748 15520 1879 15560
rect 2458 15520 2467 15560
rect 2507 15520 2516 15560
rect 2563 15520 2572 15560
rect 2612 15520 2743 15560
rect 2947 15520 2956 15560
rect 2996 15520 3095 15560
rect 3135 15520 3144 15560
rect 3331 15520 3340 15560
rect 3380 15520 3511 15560
rect 3811 15520 3820 15560
rect 3860 15520 4012 15560
rect 4052 15520 4061 15560
rect 4300 15520 4323 15560
rect 4363 15520 4372 15560
rect 4432 15520 4441 15560
rect 4481 15520 4490 15560
rect 4579 15520 4588 15560
rect 4628 15520 4637 15560
rect 4771 15520 4780 15560
rect 4820 15520 4829 15560
rect 4876 15520 5164 15560
rect 5204 15520 5213 15560
rect 5417 15520 5548 15560
rect 5588 15520 5597 15560
rect 6307 15520 6316 15560
rect 6356 15520 6604 15560
rect 6644 15520 6653 15560
rect 7027 15520 7036 15560
rect 7076 15520 7085 15560
rect 7162 15520 7171 15560
rect 7211 15520 7220 15560
rect 7267 15520 7276 15560
rect 7316 15520 7325 15560
rect 8074 15520 8083 15560
rect 8123 15520 8140 15560
rect 8180 15520 8263 15560
rect 8323 15520 8332 15560
rect 8372 15520 8468 15560
rect 8515 15520 8524 15560
rect 8564 15520 8620 15560
rect 8660 15520 8724 15560
rect 8908 15520 9100 15560
rect 9140 15520 9149 15560
rect 9283 15520 9292 15560
rect 9332 15520 9341 15560
rect 9475 15520 9484 15560
rect 9524 15520 9772 15560
rect 9812 15520 9821 15560
rect 9996 15520 10009 15560
rect 10049 15520 10196 15560
rect 10447 15520 10456 15560
rect 10496 15520 10505 15560
rect 10601 15520 10701 15560
rect 10772 15520 10781 15560
rect 10936 15547 11020 15560
rect 11006 15520 11020 15547
rect 11060 15520 11141 15560
rect 11181 15520 11191 15560
rect 11290 15520 11299 15560
rect 11339 15520 11348 15560
rect 11404 15551 11444 15560
rect 1612 15476 1652 15520
rect 2572 15502 2612 15511
rect 4195 15478 4204 15518
rect 4244 15478 4253 15518
rect 1565 15436 1612 15476
rect 1652 15436 1661 15476
rect 3226 15436 3235 15476
rect 3275 15436 3284 15476
rect 3244 15392 3284 15436
rect 4204 15392 4244 15478
rect 4780 15476 4820 15520
rect 6922 15478 6931 15518
rect 6971 15478 6983 15518
rect 4553 15436 4588 15476
rect 4628 15436 4684 15476
rect 4724 15436 4733 15476
rect 4780 15436 5164 15476
rect 5204 15436 5213 15476
rect 6617 15436 6700 15476
rect 6779 15436 6797 15476
rect 3244 15352 4148 15392
rect 4204 15352 4246 15392
rect 6451 15352 6460 15392
rect 6500 15352 6796 15392
rect 6836 15352 6845 15392
rect 2851 15268 2860 15308
rect 2900 15268 2956 15308
rect 2996 15268 3031 15308
rect 0 15224 400 15244
rect 0 15184 3724 15224
rect 3764 15184 3773 15224
rect 0 15164 400 15184
rect 4108 15140 4148 15352
rect 4206 15308 4246 15352
rect 6943 15308 6983 15478
rect 7276 15392 7316 15520
rect 8428 15476 8468 15520
rect 9100 15476 9140 15520
rect 10156 15476 10196 15520
rect 10847 15478 10856 15518
rect 10896 15478 10905 15518
rect 11674 15520 11683 15560
rect 11723 15520 11732 15560
rect 11851 15520 11860 15560
rect 11924 15520 12040 15560
rect 12355 15520 12364 15560
rect 12404 15520 12413 15560
rect 12592 15520 12601 15560
rect 12641 15520 12650 15560
rect 12739 15520 12748 15560
rect 12788 15520 12892 15560
rect 12932 15520 12941 15560
rect 7817 15436 7948 15476
rect 7988 15436 7997 15476
rect 8419 15436 8428 15476
rect 8468 15436 8477 15476
rect 9100 15436 9196 15476
rect 9236 15436 9245 15476
rect 9898 15467 10060 15476
rect 9898 15427 9907 15467
rect 9947 15436 10060 15467
rect 10100 15436 10109 15476
rect 10156 15436 10636 15476
rect 10676 15436 10685 15476
rect 9947 15427 9956 15436
rect 9898 15426 9956 15427
rect 10856 15392 10896 15478
rect 11404 15476 11444 15511
rect 11011 15436 11020 15476
rect 11060 15436 11116 15476
rect 11156 15436 11191 15476
rect 11395 15436 11404 15476
rect 11444 15436 11491 15476
rect 12259 15436 12268 15476
rect 12308 15436 12317 15476
rect 7276 15352 7852 15392
rect 7892 15352 7901 15392
rect 8236 15352 9236 15392
rect 8236 15308 8276 15352
rect 4195 15268 4204 15308
rect 4244 15268 4253 15308
rect 4963 15268 4972 15308
rect 5012 15268 5021 15308
rect 5731 15268 5740 15308
rect 5780 15268 5932 15308
rect 5972 15268 5981 15308
rect 6943 15268 8276 15308
rect 8323 15268 8332 15308
rect 8372 15268 8381 15308
rect 9091 15268 9100 15308
rect 9140 15268 9149 15308
rect 4972 15224 5012 15268
rect 4579 15184 4588 15224
rect 4628 15184 5012 15224
rect 3103 15100 3112 15140
rect 3480 15100 3489 15140
rect 4108 15100 4972 15140
rect 5012 15100 5021 15140
rect 1603 14932 1612 14972
rect 1652 14932 1948 14972
rect 1988 14932 1997 14972
rect 4073 14932 4195 14972
rect 4244 14932 4253 14972
rect 8332 14888 8372 15268
rect 3980 14879 4876 14888
rect 4020 14848 4876 14879
rect 4916 14848 4925 14888
rect 5262 14848 6028 14888
rect 6068 14848 6548 14888
rect 6883 14848 6892 14888
rect 6932 14848 7364 14888
rect 8094 14848 8103 14888
rect 8143 14848 8372 14888
rect 8515 14848 8524 14888
rect 8564 14848 8716 14888
rect 8756 14848 8765 14888
rect 3980 14830 4020 14839
rect 0 14804 400 14824
rect 0 14764 652 14804
rect 692 14764 701 14804
rect 1324 14764 2764 14804
rect 2804 14764 2813 14804
rect 2947 14764 2956 14804
rect 2996 14764 3148 14804
rect 3188 14764 3284 14804
rect 4579 14764 4588 14804
rect 4628 14764 4964 14804
rect 0 14744 400 14764
rect 1324 14720 1364 14764
rect 2092 14720 2132 14764
rect 3244 14720 3284 14764
rect 3340 14720 3380 14729
rect 4924 14720 4964 14764
rect 1193 14680 1324 14720
rect 1364 14680 1373 14720
rect 1481 14680 1516 14720
rect 1556 14680 1612 14720
rect 1652 14680 1661 14720
rect 1961 14680 2092 14720
rect 2132 14680 2141 14720
rect 2275 14680 2284 14720
rect 2324 14680 2333 14720
rect 3235 14680 3244 14720
rect 3284 14680 3293 14720
rect 3380 14680 3436 14720
rect 3476 14680 3511 14720
rect 3619 14680 3628 14720
rect 3668 14680 4003 14720
rect 4043 14680 4052 14720
rect 4553 14680 4588 14720
rect 4628 14680 4684 14720
rect 4724 14680 4733 14720
rect 4924 14680 4963 14720
rect 5003 14680 5012 14720
rect 5059 14691 5068 14731
rect 5108 14691 5120 14731
rect 5262 14720 5302 14848
rect 6113 14764 6124 14804
rect 6164 14764 6173 14804
rect 6269 14764 6316 14804
rect 6356 14764 6365 14804
rect 5832 14722 5932 14762
rect 2284 14636 2324 14680
rect 3340 14671 3380 14680
rect 5080 14636 5120 14691
rect 5242 14711 5302 14720
rect 5242 14671 5251 14711
rect 5291 14680 5302 14711
rect 5377 14680 5386 14720
rect 5426 14680 5435 14720
rect 5513 14680 5524 14720
rect 5564 14680 5644 14720
rect 5684 14680 5693 14720
rect 5923 14691 5932 14722
rect 5972 14691 5981 14762
rect 6113 14720 6153 14764
rect 6316 14720 6356 14764
rect 6508 14731 6548 14848
rect 7324 14804 7364 14848
rect 6595 14764 6604 14804
rect 6644 14764 6788 14804
rect 7075 14764 7084 14804
rect 7124 14764 7180 14804
rect 7220 14764 7255 14804
rect 7306 14795 7364 14804
rect 6070 14680 6079 14720
rect 6119 14680 6153 14720
rect 6198 14680 6207 14720
rect 6247 14680 6256 14720
rect 6298 14680 6307 14720
rect 6347 14680 6356 14720
rect 6475 14691 6484 14731
rect 6524 14691 6548 14731
rect 6748 14720 6788 14764
rect 7306 14755 7315 14795
rect 7355 14755 7364 14795
rect 7306 14754 7364 14755
rect 7426 14764 7468 14804
rect 7508 14764 7517 14804
rect 8131 14764 8140 14804
rect 8180 14764 8189 14804
rect 8279 14764 8660 14804
rect 8803 14764 8812 14804
rect 8852 14764 8983 14804
rect 7426 14720 7466 14764
rect 8140 14720 8180 14764
rect 6748 14680 7180 14720
rect 7220 14680 7229 14720
rect 7408 14680 7417 14720
rect 7457 14680 7466 14720
rect 7543 14680 7552 14720
rect 7592 14680 8044 14720
rect 8084 14680 8093 14720
rect 8136 14680 8145 14720
rect 8185 14680 8227 14720
rect 5291 14671 5300 14680
rect 5242 14670 5300 14671
rect 1699 14596 1708 14636
rect 1748 14596 2324 14636
rect 2907 14596 2956 14636
rect 2996 14596 3038 14636
rect 3078 14596 3087 14636
rect 4445 14596 4492 14636
rect 4532 14596 4541 14636
rect 5068 14596 5120 14636
rect 5382 14636 5422 14680
rect 6216 14636 6256 14680
rect 5382 14596 5492 14636
rect 6216 14596 6508 14636
rect 6548 14596 6557 14636
rect 2284 14552 2324 14596
rect 4492 14552 4532 14596
rect 1961 14512 2092 14552
rect 2132 14512 2141 14552
rect 2284 14512 2900 14552
rect 3130 14512 3139 14552
rect 3179 14512 4204 14552
rect 4244 14512 4253 14552
rect 4474 14512 4483 14552
rect 4523 14512 4532 14552
rect 4579 14512 4588 14552
rect 4628 14512 4637 14552
rect 4771 14512 4780 14552
rect 4820 14512 4972 14552
rect 5012 14512 5021 14552
rect 2860 14468 2900 14512
rect 4588 14468 4628 14512
rect 2860 14428 4628 14468
rect 5068 14468 5108 14596
rect 5155 14512 5164 14552
rect 5204 14512 5335 14552
rect 5068 14428 5356 14468
rect 5396 14428 5405 14468
rect 0 14384 400 14404
rect 5452 14384 5492 14596
rect 8279 14552 8319 14764
rect 8620 14762 8660 14764
rect 8620 14722 8648 14762
rect 8688 14722 8697 14762
rect 9100 14720 9140 15268
rect 9196 15224 9236 15352
rect 10856 15352 11884 15392
rect 11924 15352 11933 15392
rect 10856 15308 10896 15352
rect 12268 15308 12308 15436
rect 10627 15268 10636 15308
rect 10676 15268 10896 15308
rect 11683 15268 11692 15308
rect 11732 15268 12308 15308
rect 12364 15308 12404 15520
rect 13036 15476 13076 15772
rect 15916 15728 15956 15772
rect 17452 15728 17492 15856
rect 20524 15772 21100 15812
rect 21140 15772 21149 15812
rect 25036 15772 28204 15812
rect 28244 15772 28253 15812
rect 20524 15728 20564 15772
rect 25036 15728 25076 15772
rect 13315 15688 13324 15728
rect 13364 15688 13507 15728
rect 13547 15688 13556 15728
rect 13603 15688 13612 15728
rect 13652 15688 14284 15728
rect 14324 15688 14333 15728
rect 14380 15688 15428 15728
rect 15907 15688 15916 15728
rect 15956 15688 15965 15728
rect 16012 15688 16469 15728
rect 16762 15688 16771 15728
rect 16811 15688 17492 15728
rect 18499 15688 18508 15728
rect 18548 15688 18988 15728
rect 19028 15688 19037 15728
rect 20515 15688 20524 15728
rect 20564 15688 20573 15728
rect 20890 15688 20899 15728
rect 20939 15688 20948 15728
rect 14380 15644 14420 15688
rect 15388 15644 15428 15688
rect 16012 15644 16052 15688
rect 13228 15604 13516 15644
rect 13556 15604 13565 15644
rect 13673 15635 13804 15644
rect 13673 15604 13795 15635
rect 13844 15604 13853 15644
rect 14050 15604 14476 15644
rect 14516 15604 14580 15644
rect 14668 15604 14764 15644
rect 14804 15604 14813 15644
rect 14938 15635 15148 15644
rect 13228 15602 13268 15604
rect 13191 15562 13200 15602
rect 13240 15562 13268 15602
rect 13786 15595 13795 15604
rect 13835 15595 13844 15604
rect 13786 15594 13844 15595
rect 14050 15560 14090 15604
rect 14668 15560 14708 15604
rect 14938 15595 14947 15635
rect 14987 15604 15148 15635
rect 15188 15604 15197 15644
rect 15379 15604 15388 15644
rect 15428 15604 16052 15644
rect 16099 15604 16108 15644
rect 16148 15604 16157 15644
rect 14987 15595 14996 15604
rect 14938 15594 14996 15595
rect 15388 15560 15428 15604
rect 16108 15560 16148 15604
rect 16429 15560 16469 15688
rect 20908 15644 20948 15688
rect 16588 15604 17108 15644
rect 17443 15604 17452 15644
rect 17492 15604 17501 15644
rect 19171 15604 19180 15644
rect 19220 15604 19988 15644
rect 20323 15604 20332 15644
rect 20372 15604 20948 15644
rect 21007 15688 22060 15728
rect 22100 15688 22109 15728
rect 24259 15688 24268 15728
rect 24308 15688 25076 15728
rect 25123 15688 25132 15728
rect 25172 15688 25228 15728
rect 25268 15688 25303 15728
rect 27043 15688 27052 15728
rect 27092 15688 27101 15728
rect 27305 15688 27427 15728
rect 27476 15688 27485 15728
rect 16588 15560 16628 15604
rect 13324 15520 13363 15560
rect 13403 15520 13412 15560
rect 13498 15520 13507 15560
rect 13547 15520 13556 15560
rect 13324 15476 13364 15520
rect 12490 15467 12788 15476
rect 12490 15427 12499 15467
rect 12539 15436 12788 15467
rect 13027 15436 13036 15476
rect 13076 15436 13085 15476
rect 13219 15436 13228 15476
rect 13268 15436 13364 15476
rect 12539 15427 12548 15436
rect 12490 15426 12548 15427
rect 12748 15308 12788 15436
rect 13001 15352 13132 15392
rect 13172 15352 13181 15392
rect 12364 15268 12596 15308
rect 12739 15268 12748 15308
rect 12788 15268 13324 15308
rect 13364 15268 13373 15308
rect 9196 15184 12268 15224
rect 12308 15184 12317 15224
rect 10877 15100 10886 15140
rect 11254 15100 11263 15140
rect 9283 15016 9292 15056
rect 9332 15016 10732 15056
rect 10772 15016 10781 15056
rect 12556 14972 12596 15268
rect 12835 15016 12844 15056
rect 12884 15016 12893 15056
rect 10051 14932 10060 14972
rect 10100 14932 10339 14972
rect 10379 14932 10388 14972
rect 11779 14932 11788 14972
rect 11828 14932 11837 14972
rect 12067 14932 12076 14972
rect 12116 14932 12125 14972
rect 12538 14932 12547 14972
rect 12587 14932 12596 14972
rect 12844 14972 12884 15016
rect 13516 14972 13556 15520
rect 13610 15551 13652 15560
rect 13610 15511 13612 15551
rect 13882 15520 13891 15560
rect 13931 15520 13940 15560
rect 14028 15520 14037 15560
rect 14077 15520 14090 15560
rect 14204 15520 14213 15560
rect 14253 15520 14273 15560
rect 14313 15520 14384 15560
rect 14467 15520 14476 15560
rect 14516 15520 14525 15560
rect 14650 15520 14659 15560
rect 14699 15520 14708 15560
rect 14764 15551 14804 15560
rect 13610 15502 13652 15511
rect 13610 15392 13650 15502
rect 13900 15476 13940 15520
rect 14476 15476 14516 15520
rect 15034 15520 15043 15560
rect 15083 15520 15092 15560
rect 15211 15520 15220 15560
rect 15260 15520 15428 15560
rect 15619 15520 15628 15560
rect 15668 15520 15916 15560
rect 15956 15520 15965 15560
rect 16061 15520 16106 15560
rect 16146 15520 16155 15560
rect 16411 15520 16420 15560
rect 16460 15520 16469 15560
rect 16570 15520 16579 15560
rect 16619 15520 16628 15560
rect 16687 15520 16696 15560
rect 16736 15520 16745 15560
rect 16829 15520 16867 15560
rect 16907 15520 16916 15560
rect 14764 15476 14804 15511
rect 13795 15436 13804 15476
rect 13844 15436 13940 15476
rect 14083 15436 14092 15476
rect 14132 15436 14516 15476
rect 14668 15436 14804 15476
rect 15052 15476 15092 15520
rect 15916 15476 15956 15520
rect 16696 15476 16736 15520
rect 16876 15476 16916 15520
rect 16963 15509 16972 15549
rect 17012 15509 17021 15549
rect 15052 15436 15436 15476
rect 15476 15436 15485 15476
rect 15619 15436 15628 15476
rect 15668 15436 15677 15476
rect 15916 15436 16492 15476
rect 16532 15436 16736 15476
rect 16867 15436 16876 15476
rect 16916 15436 16925 15476
rect 14668 15392 14708 15436
rect 15052 15392 15092 15436
rect 15628 15392 15668 15436
rect 16972 15392 17012 15509
rect 13610 15352 14188 15392
rect 14228 15352 14237 15392
rect 14284 15352 14708 15392
rect 14755 15352 14764 15392
rect 14804 15352 15092 15392
rect 15235 15352 15244 15392
rect 15284 15352 15668 15392
rect 16780 15352 17012 15392
rect 14284 15308 14324 15352
rect 14275 15268 14284 15308
rect 14324 15268 14333 15308
rect 14650 15268 14659 15308
rect 14699 15268 14708 15308
rect 14668 15224 14708 15268
rect 13987 15184 13996 15224
rect 14036 15184 14708 15224
rect 16780 15056 16820 15352
rect 17068 15308 17108 15604
rect 17452 15560 17492 15604
rect 19948 15560 19988 15604
rect 21007 15560 21047 15688
rect 27052 15644 27092 15688
rect 21475 15604 21484 15644
rect 21524 15604 22004 15644
rect 22522 15604 22531 15644
rect 22571 15604 22732 15644
rect 22772 15604 22781 15644
rect 24835 15604 24844 15644
rect 24884 15604 26084 15644
rect 21964 15560 22004 15604
rect 26044 15560 26084 15604
rect 26908 15604 26956 15644
rect 26996 15604 27005 15644
rect 27052 15604 27572 15644
rect 26908 15560 26948 15604
rect 27532 15560 27572 15604
rect 28204 15560 28244 15772
rect 29818 15688 29827 15728
rect 29867 15688 29876 15728
rect 29836 15560 29876 15688
rect 29923 15604 29932 15644
rect 29972 15604 30644 15644
rect 30604 15560 30644 15604
rect 17242 15520 17251 15560
rect 17291 15520 17300 15560
rect 17347 15520 17356 15560
rect 17396 15520 17492 15560
rect 17731 15520 17740 15560
rect 17780 15520 17789 15560
rect 18211 15520 18220 15560
rect 18260 15551 18391 15560
rect 18260 15520 18316 15551
rect 17260 15476 17300 15520
rect 17740 15476 17780 15520
rect 18356 15520 18391 15551
rect 18796 15551 19084 15560
rect 18316 15502 18356 15511
rect 18836 15520 19084 15551
rect 19124 15520 19133 15560
rect 19433 15520 19564 15560
rect 19604 15520 19613 15560
rect 19660 15520 19673 15560
rect 19713 15520 19722 15560
rect 19939 15520 19948 15560
rect 19988 15520 19997 15560
rect 20227 15520 20236 15560
rect 20276 15520 20285 15560
rect 20369 15520 20378 15560
rect 20418 15520 20524 15560
rect 20564 15520 20948 15560
rect 20995 15520 21004 15560
rect 21044 15520 21053 15560
rect 21257 15520 21388 15560
rect 21428 15520 21437 15560
rect 21562 15520 21571 15560
rect 21620 15520 21751 15560
rect 21946 15520 21955 15560
rect 21995 15520 22004 15560
rect 22051 15520 22060 15560
rect 22100 15520 22444 15560
rect 22484 15520 22493 15560
rect 22906 15520 22915 15560
rect 22955 15520 25268 15560
rect 18796 15502 18836 15511
rect 17260 15436 17343 15476
rect 17443 15436 17452 15476
rect 17492 15436 17780 15476
rect 17827 15436 17836 15476
rect 17876 15436 17932 15476
rect 17972 15436 18007 15476
rect 17303 15392 17343 15436
rect 17303 15352 18508 15392
rect 18548 15352 18557 15392
rect 16684 15016 16820 15056
rect 16972 15268 17108 15308
rect 19267 15268 19276 15308
rect 19316 15268 19325 15308
rect 16972 15056 17012 15268
rect 18651 15100 18660 15140
rect 19028 15100 19037 15140
rect 16972 15016 17932 15056
rect 17972 15016 17981 15056
rect 16684 14972 16724 15016
rect 19276 14972 19316 15268
rect 19660 14972 19700 15520
rect 20236 15476 20276 15520
rect 20908 15476 20948 15520
rect 20236 15436 20428 15476
rect 20468 15436 20477 15476
rect 20908 15436 21236 15476
rect 24067 15436 24076 15476
rect 24116 15436 24125 15476
rect 21196 15308 21236 15436
rect 21161 15268 21196 15308
rect 21236 15268 21292 15308
rect 21332 15268 21341 15308
rect 22121 15268 22243 15308
rect 22292 15268 22301 15308
rect 24451 15268 24460 15308
rect 24500 15268 24509 15308
rect 24643 15268 24652 15308
rect 24692 15268 24844 15308
rect 24884 15268 24893 15308
rect 24460 15224 24500 15268
rect 25228 15224 25268 15520
rect 25389 15518 25429 15527
rect 25389 15392 25429 15478
rect 25474 15520 25492 15560
rect 25532 15520 25541 15560
rect 25594 15520 25603 15560
rect 25643 15520 25708 15560
rect 25748 15520 25783 15560
rect 26035 15520 26044 15560
rect 26084 15520 26093 15560
rect 26179 15520 26188 15560
rect 26228 15520 26237 15560
rect 26755 15520 26764 15560
rect 26804 15520 26813 15560
rect 26890 15520 26899 15560
rect 26939 15520 26948 15560
rect 27004 15520 27013 15560
rect 27053 15520 27092 15560
rect 27523 15520 27532 15560
rect 27572 15520 27628 15560
rect 27668 15520 27732 15560
rect 27907 15520 27916 15560
rect 27956 15520 28108 15560
rect 28148 15520 28157 15560
rect 28204 15520 28780 15560
rect 28820 15520 28829 15560
rect 28963 15520 28972 15560
rect 29012 15520 29876 15560
rect 29932 15520 30124 15560
rect 30164 15520 30173 15560
rect 30586 15551 30644 15560
rect 25474 15476 25514 15520
rect 26188 15476 26228 15520
rect 25474 15436 25612 15476
rect 25652 15436 26228 15476
rect 26764 15476 26804 15520
rect 26764 15436 26996 15476
rect 26956 15392 26996 15436
rect 25389 15352 25516 15392
rect 25556 15352 25565 15392
rect 25699 15352 25708 15392
rect 25748 15352 25843 15392
rect 25883 15352 25892 15392
rect 26179 15352 26188 15392
rect 26228 15352 26380 15392
rect 26420 15352 26429 15392
rect 26947 15352 26956 15392
rect 26996 15352 27005 15392
rect 25516 15308 25556 15352
rect 27052 15308 27092 15520
rect 29932 15476 29972 15520
rect 30586 15511 30595 15551
rect 30635 15511 30644 15551
rect 30586 15510 30644 15511
rect 28003 15436 28012 15476
rect 28052 15436 29972 15476
rect 30025 15436 30034 15476
rect 30074 15436 30083 15476
rect 30691 15436 30700 15476
rect 30740 15436 30748 15476
rect 30788 15436 31180 15476
rect 31220 15436 31229 15476
rect 30028 15392 30068 15436
rect 27628 15352 30068 15392
rect 30307 15352 30316 15392
rect 30356 15352 31084 15392
rect 31124 15352 31133 15392
rect 25516 15268 27340 15308
rect 27380 15268 27389 15308
rect 19939 15184 19948 15224
rect 19988 15184 24748 15224
rect 24788 15184 24797 15224
rect 25228 15184 26284 15224
rect 26324 15184 26333 15224
rect 26425 15100 26434 15140
rect 26802 15100 26811 15140
rect 21292 15016 23884 15056
rect 23924 15016 23933 15056
rect 25228 15016 27532 15056
rect 27572 15016 27581 15056
rect 12844 14932 13460 14972
rect 13507 14932 13516 14972
rect 13556 14932 13565 14972
rect 13610 14932 16148 14972
rect 16675 14932 16684 14972
rect 16724 14932 16733 14972
rect 16780 14932 19316 14972
rect 19651 14932 19660 14972
rect 19700 14932 19709 14972
rect 19843 14932 19852 14972
rect 19892 14932 21236 14972
rect 11788 14888 11828 14932
rect 10204 14848 11500 14888
rect 11540 14848 11549 14888
rect 11660 14879 11980 14888
rect 9571 14764 9580 14804
rect 9643 14764 9751 14804
rect 10204 14720 10244 14848
rect 11700 14848 11980 14879
rect 12020 14848 12029 14888
rect 11660 14830 11700 14839
rect 12076 14804 12116 14932
rect 13420 14888 13460 14932
rect 13610 14888 13650 14932
rect 16108 14888 16148 14932
rect 16780 14888 16820 14932
rect 21196 14888 21236 14932
rect 12163 14848 12172 14888
rect 12212 14848 12221 14888
rect 13420 14848 13650 14888
rect 14921 14848 15043 14888
rect 15092 14848 15101 14888
rect 15881 14848 16012 14888
rect 16052 14848 16061 14888
rect 16108 14848 16820 14888
rect 17539 14848 17548 14888
rect 17588 14848 18316 14888
rect 18356 14848 18365 14888
rect 20489 14848 20620 14888
rect 20660 14848 20669 14888
rect 21178 14848 21187 14888
rect 21227 14848 21236 14888
rect 12172 14804 12212 14848
rect 14794 14804 14803 14832
rect 10624 14764 10636 14804
rect 10676 14764 10704 14804
rect 12067 14764 12076 14804
rect 12116 14764 12125 14804
rect 12172 14764 12291 14804
rect 12331 14764 12340 14804
rect 14083 14764 14092 14804
rect 14132 14764 14141 14804
rect 14750 14792 14803 14804
rect 14843 14792 14852 14832
rect 14750 14764 14852 14792
rect 14908 14764 15724 14804
rect 15764 14764 15773 14804
rect 16012 14764 16300 14804
rect 16340 14764 16349 14804
rect 18595 14764 18604 14804
rect 18644 14764 18653 14804
rect 18700 14764 20852 14804
rect 20969 14764 21091 14804
rect 21140 14764 21149 14804
rect 10624 14720 10664 14764
rect 12460 14720 12832 14727
rect 8393 14680 8493 14720
rect 8564 14680 8573 14720
rect 8938 14680 8947 14720
rect 8987 14680 9140 14720
rect 9379 14680 9388 14720
rect 9428 14680 9484 14720
rect 9524 14680 9559 14720
rect 9676 14680 9701 14720
rect 9741 14680 9750 14720
rect 9850 14680 9859 14720
rect 9908 14680 10039 14720
rect 10147 14680 10156 14720
rect 10196 14680 10244 14720
rect 10330 14680 10339 14720
rect 10379 14680 10388 14720
rect 10474 14680 10483 14720
rect 10523 14680 10532 14720
rect 10608 14680 10617 14720
rect 10657 14680 10666 14720
rect 10709 14680 10718 14720
rect 10758 14680 10767 14720
rect 10891 14680 10900 14720
rect 10964 14680 11080 14720
rect 11674 14680 11683 14720
rect 11723 14680 11828 14720
rect 11875 14680 11884 14720
rect 11924 14680 12172 14720
rect 12212 14680 12221 14720
rect 12329 14680 12409 14720
rect 12449 14680 12460 14720
rect 12500 14687 12832 14720
rect 12872 14687 12881 14727
rect 12500 14680 12509 14687
rect 12923 14680 12932 14720
rect 12972 14680 12981 14720
rect 13315 14680 13324 14720
rect 13364 14680 13516 14720
rect 13556 14680 13565 14720
rect 13699 14680 13708 14720
rect 13748 14680 13891 14720
rect 13931 14680 13940 14720
rect 13987 14691 13996 14731
rect 14036 14691 14045 14731
rect 14092 14720 14132 14764
rect 8524 14636 8564 14680
rect 9676 14636 9716 14680
rect 10348 14636 10388 14680
rect 8524 14596 8590 14636
rect 9353 14596 9388 14636
rect 9428 14596 9484 14636
rect 9524 14596 9533 14636
rect 9676 14596 9772 14636
rect 9812 14596 9821 14636
rect 10051 14596 10060 14636
rect 10100 14596 10388 14636
rect 10492 14636 10532 14680
rect 10710 14636 10750 14680
rect 11788 14636 11828 14680
rect 10492 14596 10540 14636
rect 10580 14596 10589 14636
rect 10710 14596 10732 14636
rect 10772 14596 10789 14636
rect 11788 14596 12364 14636
rect 12404 14596 12413 14636
rect 8550 14552 8590 14596
rect 6281 14512 6403 14552
rect 6452 14512 6461 14552
rect 7267 14512 7276 14552
rect 7316 14512 7708 14552
rect 7748 14512 7757 14552
rect 8279 14512 8323 14552
rect 8363 14512 8372 14552
rect 8550 14512 9004 14552
rect 9044 14512 9053 14552
rect 8620 14470 8683 14512
rect 8749 14428 10252 14468
rect 10292 14428 10301 14468
rect 10627 14428 10636 14468
rect 10676 14428 12844 14468
rect 12884 14428 12893 14468
rect 8749 14384 8789 14428
rect 0 14344 596 14384
rect 0 14324 400 14344
rect 556 14300 596 14344
rect 2860 14344 3916 14384
rect 3956 14344 3965 14384
rect 4343 14344 4352 14384
rect 4720 14344 4729 14384
rect 5059 14344 5068 14384
rect 5108 14344 6316 14384
rect 6356 14344 6365 14384
rect 6979 14344 6988 14384
rect 7028 14344 8789 14384
rect 9187 14344 9196 14384
rect 9236 14344 11884 14384
rect 11924 14344 11933 14384
rect 12117 14344 12126 14384
rect 12494 14344 12503 14384
rect 2860 14300 2900 14344
rect 556 14260 1132 14300
rect 1172 14260 1181 14300
rect 1223 14260 2900 14300
rect 3628 14260 6068 14300
rect 1223 14216 1263 14260
rect 3628 14216 3668 14260
rect 643 14176 652 14216
rect 692 14176 1263 14216
rect 1507 14176 1516 14216
rect 1595 14176 1687 14216
rect 2083 14176 2092 14216
rect 2132 14176 2956 14216
rect 2996 14176 3005 14216
rect 3619 14176 3628 14216
rect 3668 14176 3677 14216
rect 3994 14176 4003 14216
rect 4043 14176 4052 14216
rect 5434 14176 5443 14216
rect 5492 14176 5623 14216
rect 5705 14176 5827 14216
rect 5876 14176 5885 14216
rect 4012 14132 4052 14176
rect 1036 14092 1324 14132
rect 1364 14092 1373 14132
rect 2188 14092 4052 14132
rect 4300 14092 5068 14132
rect 5108 14092 5117 14132
rect 5242 14123 5548 14132
rect 1036 14048 1076 14092
rect 2188 14048 2228 14092
rect 2668 14048 2708 14092
rect 4300 14048 4340 14092
rect 1027 14008 1036 14048
rect 1076 14008 1085 14048
rect 1210 14008 1219 14048
rect 1259 14008 1708 14048
rect 1760 14008 1769 14048
rect 1882 14008 1891 14048
rect 1931 14008 1940 14048
rect 2179 14008 2188 14048
rect 2228 14008 2237 14048
rect 2554 14008 2563 14048
rect 2603 14008 2612 14048
rect 2659 14008 2668 14048
rect 2708 14008 2717 14048
rect 3017 14008 3148 14048
rect 3188 14008 3197 14048
rect 3305 14008 3436 14048
rect 3476 14008 3485 14048
rect 4291 14008 4300 14048
rect 4340 14008 4349 14048
rect 4841 14008 4963 14048
rect 5012 14008 5021 14048
rect 5068 14039 5108 14092
rect 5242 14083 5251 14123
rect 5291 14092 5548 14123
rect 5588 14092 5597 14132
rect 5291 14083 5300 14092
rect 5242 14082 5300 14083
rect 0 13964 400 13984
rect 1900 13964 1940 14008
rect 2572 13964 2612 14008
rect 3436 13964 3476 14008
rect 5334 14008 5343 14048
rect 5383 14008 5392 14048
rect 5501 14008 5524 14048
rect 5564 14008 5588 14048
rect 5720 14008 5729 14048
rect 5769 14008 5780 14048
rect 5923 14008 5932 14048
rect 5972 14008 5981 14048
rect 6028 14039 6068 14260
rect 6113 14216 6153 14344
rect 7996 14260 10924 14300
rect 10964 14260 10973 14300
rect 11596 14260 12844 14300
rect 12884 14260 12893 14300
rect 6113 14176 6172 14216
rect 6212 14176 6221 14216
rect 7171 14176 7180 14216
rect 7220 14176 7533 14216
rect 7625 14176 7747 14216
rect 7796 14176 7805 14216
rect 7493 14132 7533 14176
rect 6787 14092 6796 14132
rect 6836 14092 7220 14132
rect 7493 14092 7839 14132
rect 7180 14048 7220 14092
rect 7799 14048 7839 14092
rect 7996 14048 8036 14260
rect 11596 14216 11636 14260
rect 12940 14216 12980 14680
rect 13996 14636 14036 14691
rect 14092 14680 14141 14720
rect 14181 14680 14190 14720
rect 14261 14680 14270 14720
rect 14310 14680 14319 14720
rect 14443 14680 14452 14720
rect 14516 14680 14632 14720
rect 14270 14636 14310 14680
rect 13219 14596 13228 14636
rect 13268 14596 14036 14636
rect 14188 14596 14310 14636
rect 14750 14636 14790 14764
rect 14908 14720 14948 14764
rect 16012 14720 16052 14764
rect 18604 14720 18644 14764
rect 18700 14720 18740 14764
rect 20812 14720 20852 14764
rect 21292 14720 21332 15016
rect 25228 14972 25268 15016
rect 27628 14972 27668 15352
rect 28099 15268 28108 15308
rect 28148 15268 28157 15308
rect 29635 15268 29644 15308
rect 29684 15268 29740 15308
rect 29780 15268 29815 15308
rect 23107 14932 23116 14972
rect 23156 14932 23287 14972
rect 23683 14932 23692 14972
rect 23732 14932 24268 14972
rect 24308 14932 24940 14972
rect 24980 14932 24989 14972
rect 25219 14932 25228 14972
rect 25268 14932 25277 14972
rect 25507 14932 25516 14972
rect 25556 14932 26132 14972
rect 27619 14932 27628 14972
rect 27668 14932 27677 14972
rect 21859 14848 21868 14888
rect 21908 14848 21917 14888
rect 22051 14848 22060 14888
rect 22100 14848 24067 14888
rect 24107 14848 24116 14888
rect 24161 14848 24844 14888
rect 24884 14848 24893 14888
rect 25175 14848 25708 14888
rect 25748 14848 25757 14888
rect 25891 14848 25900 14888
rect 25940 14848 25949 14888
rect 21868 14804 21908 14848
rect 24161 14804 24201 14848
rect 21437 14764 21484 14804
rect 21524 14764 21533 14804
rect 21658 14764 21667 14804
rect 21707 14764 21908 14804
rect 22243 14764 22252 14804
rect 22292 14764 22484 14804
rect 21484 14720 21524 14764
rect 22444 14720 22484 14764
rect 23500 14764 24201 14804
rect 24739 14764 24748 14804
rect 24788 14764 24884 14804
rect 24931 14764 24940 14804
rect 24980 14764 25057 14804
rect 25097 14764 25111 14804
rect 23500 14720 23540 14764
rect 24844 14720 24884 14764
rect 25175 14753 25215 14848
rect 25900 14804 25940 14848
rect 25289 14764 25420 14804
rect 25460 14764 25469 14804
rect 25626 14764 25635 14804
rect 25675 14764 25940 14804
rect 14842 14680 14851 14720
rect 14891 14680 14948 14720
rect 15113 14680 15244 14720
rect 15284 14680 15293 14720
rect 15427 14680 15436 14720
rect 15476 14680 15485 14720
rect 16003 14680 16012 14720
rect 16052 14680 16061 14720
rect 16195 14680 16204 14720
rect 16244 14680 16375 14720
rect 16483 14680 16492 14720
rect 16532 14680 16663 14720
rect 16745 14680 16876 14720
rect 16916 14680 16925 14720
rect 17059 14680 17068 14720
rect 17108 14680 17740 14720
rect 17780 14680 17789 14720
rect 18499 14680 18508 14720
rect 18548 14680 18644 14720
rect 18691 14680 18700 14720
rect 18740 14680 18749 14720
rect 18953 14680 18988 14720
rect 19028 14680 19084 14720
rect 19124 14680 19133 14720
rect 15436 14636 15476 14680
rect 14750 14596 15052 14636
rect 15092 14596 15101 14636
rect 15305 14596 15436 14636
rect 15476 14596 16012 14636
rect 16052 14596 16061 14636
rect 13210 14512 13219 14552
rect 13259 14512 13324 14552
rect 13364 14512 13399 14552
rect 13066 14470 13075 14510
rect 13115 14470 13124 14510
rect 13084 14384 13124 14470
rect 14188 14468 14228 14596
rect 14750 14552 14790 14596
rect 16204 14552 16244 14680
rect 19258 14662 19267 14702
rect 19307 14662 19316 14702
rect 19363 14680 19372 14720
rect 19412 14680 19948 14720
rect 19988 14680 19997 14720
rect 20218 14680 20227 14720
rect 20267 14680 20756 14720
rect 20812 14680 21332 14720
rect 21466 14680 21475 14720
rect 21515 14680 21524 14720
rect 21571 14680 21580 14720
rect 21620 14680 21868 14720
rect 21908 14680 21917 14720
rect 22025 14680 22156 14720
rect 22196 14680 22205 14720
rect 22435 14680 22444 14720
rect 22484 14680 22493 14720
rect 23482 14680 23491 14720
rect 23531 14680 23540 14720
rect 23587 14680 23596 14720
rect 23636 14680 23767 14720
rect 24451 14680 24460 14720
rect 24500 14680 24652 14720
rect 24692 14680 24701 14720
rect 24835 14680 24844 14720
rect 24884 14680 24893 14720
rect 25708 14720 25796 14721
rect 26092 14720 26132 14932
rect 26860 14848 27724 14888
rect 27764 14848 27773 14888
rect 26275 14764 26284 14804
rect 26324 14764 26420 14804
rect 26633 14764 26755 14804
rect 26804 14764 26813 14804
rect 26380 14720 26420 14764
rect 26860 14720 26900 14848
rect 26947 14764 26956 14804
rect 26996 14764 27436 14804
rect 27476 14764 27485 14804
rect 27532 14764 27628 14804
rect 27668 14764 27677 14804
rect 27436 14720 27476 14764
rect 25175 14704 25215 14713
rect 25420 14680 25516 14720
rect 25556 14680 25565 14720
rect 25633 14680 25708 14720
rect 25748 14680 25750 14720
rect 25790 14680 25799 14720
rect 25911 14680 25921 14720
rect 25961 14680 25970 14720
rect 26092 14680 26188 14720
rect 26228 14680 26237 14720
rect 26371 14680 26380 14720
rect 26420 14680 26429 14720
rect 26606 14680 26615 14720
rect 26655 14680 26664 14720
rect 26851 14680 26860 14720
rect 26900 14680 26909 14720
rect 27209 14680 27340 14720
rect 27380 14680 27389 14720
rect 27532 14720 27572 14764
rect 28108 14720 28148 15268
rect 29251 15100 29260 15140
rect 29300 15100 30452 15140
rect 29251 14932 29260 14972
rect 29300 14932 30124 14972
rect 30164 14932 30356 14972
rect 28474 14764 28483 14804
rect 28523 14764 28532 14804
rect 30211 14764 30220 14804
rect 30260 14764 30269 14804
rect 27532 14680 27628 14720
rect 27668 14680 27677 14720
rect 27808 14680 27817 14720
rect 27857 14680 28148 14720
rect 14362 14512 14371 14552
rect 14411 14512 14790 14552
rect 15331 14512 15340 14552
rect 15380 14512 15628 14552
rect 15668 14512 15677 14552
rect 16204 14512 16387 14552
rect 16427 14512 16436 14552
rect 16483 14512 16492 14552
rect 16532 14512 16972 14552
rect 17012 14512 17021 14552
rect 17347 14512 17356 14552
rect 17396 14512 18691 14552
rect 18731 14512 18740 14552
rect 19276 14468 19316 14662
rect 20716 14636 20756 14680
rect 25420 14636 25460 14680
rect 19363 14596 19372 14636
rect 19412 14596 19756 14636
rect 19796 14596 19805 14636
rect 20323 14596 20332 14636
rect 20372 14596 20524 14636
rect 20564 14596 20573 14636
rect 20681 14596 20812 14636
rect 20852 14596 22004 14636
rect 23770 14596 23779 14636
rect 23828 14596 23959 14636
rect 25411 14596 25420 14636
rect 25460 14596 25469 14636
rect 20332 14552 20372 14596
rect 19939 14512 19948 14552
rect 19988 14512 20372 14552
rect 20428 14512 21868 14552
rect 21908 14512 21917 14552
rect 20428 14468 20468 14512
rect 14179 14428 14188 14468
rect 14228 14428 14237 14468
rect 17059 14428 17068 14468
rect 17108 14428 20468 14468
rect 21964 14468 22004 14596
rect 25911 14552 25951 14680
rect 26188 14636 26228 14680
rect 26615 14636 26655 14680
rect 27436 14671 27476 14680
rect 26188 14596 26655 14636
rect 26938 14596 26947 14636
rect 26987 14596 27134 14636
rect 27174 14596 27183 14636
rect 28003 14596 28012 14636
rect 28052 14596 28099 14636
rect 28139 14596 28183 14636
rect 23299 14512 23308 14552
rect 23348 14512 23500 14552
rect 23540 14512 23549 14552
rect 25756 14512 25951 14552
rect 26467 14512 26476 14552
rect 26516 14512 27235 14552
rect 27275 14512 27284 14552
rect 25756 14468 25796 14512
rect 28492 14468 28532 14764
rect 30316 14720 30356 14932
rect 30412 14804 30452 15100
rect 30569 14932 30700 14972
rect 30740 14932 30749 14972
rect 30857 14848 30988 14888
rect 31028 14848 31037 14888
rect 30412 14764 30836 14804
rect 30796 14720 30836 14764
rect 29347 14680 29356 14720
rect 29396 14680 30019 14720
rect 30059 14680 30068 14720
rect 30316 14680 30604 14720
rect 30644 14680 30653 14720
rect 30787 14680 30796 14720
rect 30836 14680 30845 14720
rect 29635 14596 29644 14636
rect 29684 14596 30403 14636
rect 30443 14596 30452 14636
rect 21964 14428 24652 14468
rect 24692 14428 25796 14468
rect 25900 14428 28532 14468
rect 25900 14384 25940 14428
rect 13084 14344 13324 14384
rect 13364 14344 13373 14384
rect 19891 14344 19900 14384
rect 20268 14344 20277 14384
rect 22060 14344 25940 14384
rect 27665 14344 27674 14384
rect 28042 14344 28051 14384
rect 28867 14344 28876 14384
rect 28916 14344 29452 14384
rect 29492 14344 29501 14384
rect 13123 14260 13132 14300
rect 13172 14260 13268 14300
rect 13891 14260 13900 14300
rect 13940 14260 16628 14300
rect 18595 14260 18604 14300
rect 18644 14260 20812 14300
rect 20852 14260 20861 14300
rect 13228 14216 13268 14260
rect 16588 14216 16628 14260
rect 9641 14176 9772 14216
rect 9812 14176 9821 14216
rect 10042 14176 10051 14216
rect 10091 14176 10156 14216
rect 10196 14176 11636 14216
rect 12739 14176 12748 14216
rect 12788 14176 12797 14216
rect 12931 14176 12940 14216
rect 12980 14176 12989 14216
rect 13210 14176 13219 14216
rect 13259 14176 13268 14216
rect 13507 14176 13516 14216
rect 13556 14176 13708 14216
rect 13748 14176 13757 14216
rect 14010 14176 15436 14216
rect 15476 14176 15485 14216
rect 15785 14176 15907 14216
rect 15956 14176 15965 14216
rect 16579 14176 16588 14216
rect 16628 14176 16637 14216
rect 17356 14176 18316 14216
rect 18356 14176 18365 14216
rect 19171 14176 19180 14216
rect 19220 14176 20948 14216
rect 21187 14176 21196 14216
rect 21236 14176 21388 14216
rect 21428 14176 21437 14216
rect 9187 14092 9196 14132
rect 9236 14092 9245 14132
rect 10339 14092 10348 14132
rect 10388 14092 10819 14132
rect 10859 14092 10868 14132
rect 10985 14092 11020 14132
rect 11060 14092 11116 14132
rect 11156 14092 11165 14132
rect 9196 14048 9236 14092
rect 11596 14090 11636 14176
rect 12259 14092 12268 14132
rect 12308 14092 12596 14132
rect 11578 14050 11587 14090
rect 11627 14050 11636 14090
rect 12556 14048 12596 14092
rect 12748 14067 12788 14176
rect 14010 14132 14050 14176
rect 12835 14092 12844 14132
rect 12884 14092 12893 14132
rect 13132 14092 13900 14132
rect 13940 14092 13949 14132
rect 14001 14092 14010 14132
rect 14050 14092 14092 14132
rect 14132 14092 14210 14132
rect 14563 14092 14572 14132
rect 14612 14092 14621 14132
rect 14956 14092 15628 14132
rect 15668 14092 15677 14132
rect 15800 14092 15809 14132
rect 15849 14092 16012 14132
rect 16052 14092 16061 14132
rect 5068 13990 5108 13999
rect 5352 13964 5392 14008
rect 5548 13964 5588 14008
rect 0 13924 1036 13964
rect 1076 13924 1085 13964
rect 1900 13924 2612 13964
rect 2860 13924 3476 13964
rect 4079 13924 4204 13964
rect 4250 13924 4259 13964
rect 5347 13924 5356 13964
rect 5396 13924 5439 13964
rect 5539 13924 5548 13964
rect 5588 13924 5597 13964
rect 0 13904 400 13924
rect 1210 13756 1219 13796
rect 1259 13756 1268 13796
rect 0 13544 400 13564
rect 0 13504 652 13544
rect 692 13504 701 13544
rect 0 13484 400 13504
rect 1228 13292 1268 13756
rect 2284 13292 2324 13924
rect 2860 13880 2900 13924
rect 5740 13880 5780 14008
rect 2842 13840 2851 13880
rect 2891 13840 2900 13880
rect 4387 13840 4396 13880
rect 4436 13840 5780 13880
rect 5932 13880 5972 14008
rect 6403 14008 6412 14048
rect 6452 14008 7075 14048
rect 7115 14008 7124 14048
rect 7171 14008 7180 14048
rect 7220 14008 7229 14048
rect 7459 14008 7468 14048
rect 7508 14008 7684 14048
rect 7724 14008 7733 14048
rect 7799 14008 7821 14048
rect 7861 14008 7870 14048
rect 7978 14008 7987 14048
rect 8027 14008 8036 14048
rect 8122 14008 8131 14048
rect 8171 14008 8180 14048
rect 8244 14008 8253 14048
rect 8293 14008 8620 14048
rect 8660 14008 8812 14048
rect 8852 14008 8861 14048
rect 8986 14008 8995 14048
rect 9035 14008 9044 14048
rect 9091 14008 9100 14048
rect 9140 14008 9149 14048
rect 9196 14008 9292 14048
rect 9332 14008 9341 14048
rect 9408 14008 9417 14048
rect 9457 14008 9466 14048
rect 9571 14008 9580 14048
rect 9620 14008 9772 14048
rect 9812 14008 9821 14048
rect 9929 14008 9964 14048
rect 10004 14008 10060 14048
rect 10100 14008 10109 14048
rect 10356 14008 10444 14048
rect 10484 14008 10487 14048
rect 10527 14008 10536 14048
rect 10685 14008 10713 14048
rect 10753 14028 10762 14048
rect 10753 14008 10763 14028
rect 11011 14008 11020 14048
rect 11060 14008 11107 14048
rect 11177 14008 11212 14048
rect 11252 14008 11308 14048
rect 11348 14008 11357 14048
rect 11683 14008 11692 14048
rect 11753 14008 11863 14048
rect 11971 14008 11980 14048
rect 12045 14008 12151 14048
rect 12233 14008 12364 14048
rect 12404 14008 12413 14048
rect 12547 14008 12556 14048
rect 12596 14008 12605 14048
rect 12734 14027 12743 14067
rect 12783 14027 12792 14067
rect 12844 14048 12884 14092
rect 13132 14048 13172 14092
rect 14572 14048 14612 14092
rect 12844 14008 12940 14048
rect 12980 14008 12989 14048
rect 13123 14008 13132 14048
rect 13172 14008 13181 14048
rect 13315 14008 13324 14048
rect 13364 14008 13373 14048
rect 13690 14008 13699 14048
rect 13739 14008 13748 14048
rect 13795 14008 13804 14048
rect 13844 14008 13975 14048
rect 14153 14008 14284 14048
rect 14324 14008 14333 14048
rect 14464 14008 14473 14048
rect 14513 14008 14526 14048
rect 14572 14008 14620 14048
rect 14660 14008 14669 14048
rect 6028 13990 6068 13999
rect 6403 13924 6412 13964
rect 6452 13924 6796 13964
rect 6836 13924 6845 13964
rect 7084 13880 7124 14008
rect 8140 13964 8180 14008
rect 7555 13924 7564 13964
rect 7604 13924 8180 13964
rect 5932 13840 6068 13880
rect 7084 13840 8524 13880
rect 8564 13840 8573 13880
rect 8707 13840 8716 13880
rect 8756 13840 8908 13880
rect 8948 13840 8957 13880
rect 6028 13628 6068 13840
rect 7241 13756 7363 13796
rect 7412 13756 7421 13796
rect 3103 13588 3112 13628
rect 3480 13588 3489 13628
rect 4963 13588 4972 13628
rect 5012 13588 7756 13628
rect 7796 13588 7805 13628
rect 7948 13588 8812 13628
rect 8852 13588 8861 13628
rect 7948 13544 7988 13588
rect 6787 13504 6796 13544
rect 6836 13504 7988 13544
rect 8035 13504 8044 13544
rect 8084 13504 8660 13544
rect 8009 13420 8131 13460
rect 8180 13420 8189 13460
rect 8620 13376 8660 13504
rect 9004 13460 9044 14008
rect 9100 13964 9140 14008
rect 9100 13924 9332 13964
rect 9292 13880 9332 13924
rect 9426 13880 9466 14008
rect 10718 13988 10763 14008
rect 10723 13964 10763 13988
rect 11020 13964 11060 14008
rect 10482 13924 10540 13964
rect 10580 13924 10613 13964
rect 10653 13924 10662 13964
rect 10723 13924 10732 13964
rect 10772 13924 10781 13964
rect 11011 13924 11020 13964
rect 11060 13924 11069 13964
rect 11875 13924 11884 13964
rect 11924 13924 12076 13964
rect 12116 13924 12125 13964
rect 12835 13924 12844 13964
rect 12884 13924 12940 13964
rect 12980 13924 13015 13964
rect 13324 13880 13364 14008
rect 13708 13964 13748 14008
rect 13603 13924 13612 13964
rect 13652 13924 13748 13964
rect 14486 13880 14526 14008
rect 14755 13966 14764 14006
rect 14804 13966 14813 14006
rect 14764 13880 14804 13966
rect 14956 13964 14996 14092
rect 17356 14048 17396 14176
rect 20908 14132 20948 14176
rect 17740 14092 18604 14132
rect 18644 14092 18653 14132
rect 19555 14092 19564 14132
rect 19604 14092 19988 14132
rect 17740 14048 17780 14092
rect 19948 14048 19988 14092
rect 20236 14092 20852 14132
rect 20908 14092 21379 14132
rect 21419 14092 21428 14132
rect 20236 14048 20276 14092
rect 20812 14048 20852 14092
rect 15043 14008 15052 14048
rect 15117 14008 15223 14048
rect 15388 14008 15436 14048
rect 15476 14023 15485 14048
rect 15476 14008 15560 14023
rect 15616 14008 15625 14048
rect 15665 14008 15724 14048
rect 15764 14008 15805 14048
rect 15881 14008 15916 14048
rect 15956 14008 16012 14048
rect 16052 14008 16061 14048
rect 16204 14045 16492 14048
rect 15388 13983 15560 14008
rect 16105 14005 16114 14045
rect 16154 14008 16492 14045
rect 16532 14008 16541 14048
rect 16745 14008 16771 14048
rect 16811 14008 16876 14048
rect 16916 14008 16925 14048
rect 17260 14039 17396 14048
rect 16154 14005 16244 14008
rect 17300 14008 17396 14039
rect 17443 14008 17452 14048
rect 17492 14008 17740 14048
rect 17780 14008 17789 14048
rect 18124 14008 18220 14048
rect 18260 14008 18269 14048
rect 18329 14008 18338 14048
rect 18378 14008 18508 14048
rect 18548 14008 18557 14048
rect 18682 14008 18691 14048
rect 18740 14008 18871 14048
rect 19843 14008 19852 14048
rect 19892 14008 19901 14048
rect 19948 14008 19961 14048
rect 20001 14008 20010 14048
rect 20105 14008 20236 14048
rect 20276 14008 20285 14048
rect 20393 14008 20524 14048
rect 20564 14008 20573 14048
rect 20812 14008 21484 14048
rect 21524 14008 21571 14048
rect 21611 14008 21620 14048
rect 22060 14039 22100 14344
rect 22540 14260 23060 14300
rect 23107 14260 23116 14300
rect 23156 14260 29780 14300
rect 22540 14048 22580 14260
rect 23020 14216 23060 14260
rect 29740 14216 29780 14260
rect 23020 14176 23692 14216
rect 23732 14176 23741 14216
rect 23875 14176 23884 14216
rect 23924 14176 25708 14216
rect 25748 14176 25757 14216
rect 29513 14176 29644 14216
rect 29684 14176 29693 14216
rect 29740 14176 30844 14216
rect 30884 14176 30893 14216
rect 26188 14092 29212 14132
rect 29252 14092 29356 14132
rect 29396 14092 29412 14132
rect 29731 14092 29740 14132
rect 29780 14092 29789 14132
rect 30115 14092 30124 14132
rect 30164 14092 30257 14132
rect 26188 14048 26228 14092
rect 29739 14048 29779 14092
rect 30217 14048 30257 14092
rect 17260 13990 17300 13999
rect 15520 13964 15560 13983
rect 14947 13924 14956 13964
rect 14996 13924 15005 13964
rect 15520 13924 15668 13964
rect 17731 13924 17740 13964
rect 17780 13924 17836 13964
rect 17876 13924 17911 13964
rect 15628 13880 15668 13924
rect 18124 13880 18164 14008
rect 19852 13964 19892 14008
rect 22409 14008 22540 14048
rect 22580 14008 22589 14048
rect 22889 14008 23020 14048
rect 23060 14008 23069 14048
rect 22060 13990 22100 13999
rect 23116 13989 23133 14029
rect 23173 13989 23182 14029
rect 23395 14008 23404 14048
rect 23444 14008 23453 14048
rect 23587 14008 23596 14048
rect 23636 14008 23788 14048
rect 23828 14008 24268 14048
rect 24308 14008 24317 14048
rect 26170 14008 26179 14048
rect 26219 14008 26228 14048
rect 26668 14008 27043 14048
rect 27083 14008 27092 14048
rect 27139 14008 27148 14048
rect 27188 14008 27319 14048
rect 27427 14008 27436 14048
rect 27476 14008 27619 14048
rect 27659 14008 27668 14048
rect 27907 14008 27916 14048
rect 27956 14008 28195 14048
rect 28235 14008 28244 14048
rect 28291 14008 28300 14048
rect 28340 14008 28876 14048
rect 28916 14008 28925 14048
rect 29023 14008 29032 14048
rect 29072 14008 29108 14048
rect 29155 14008 29164 14048
rect 29204 14008 29548 14048
rect 29588 14008 29597 14048
rect 29693 14008 29739 14048
rect 29779 14008 29788 14048
rect 30112 14008 30121 14048
rect 30161 14008 30257 14048
rect 18307 13924 18316 13964
rect 18356 13924 19756 13964
rect 19796 13924 19805 13964
rect 19852 13924 20620 13964
rect 20660 13924 20669 13964
rect 22505 13924 22636 13964
rect 22676 13924 22685 13964
rect 9283 13840 9292 13880
rect 9332 13840 9341 13880
rect 9426 13840 10252 13880
rect 10292 13840 10301 13880
rect 11657 13840 11788 13880
rect 11828 13840 11837 13880
rect 12355 13840 12364 13880
rect 12404 13840 12844 13880
rect 12884 13840 12893 13880
rect 13324 13840 13516 13880
rect 13556 13840 14420 13880
rect 14467 13840 14476 13880
rect 14516 13840 14526 13880
rect 14659 13840 14668 13880
rect 14708 13840 14804 13880
rect 14851 13840 14860 13880
rect 14900 13840 15532 13880
rect 15572 13840 15581 13880
rect 15628 13840 16396 13880
rect 16436 13840 16445 13880
rect 16963 13840 16972 13880
rect 17012 13840 17548 13880
rect 17588 13840 18164 13880
rect 19084 13840 21580 13880
rect 21620 13840 22156 13880
rect 22196 13840 22205 13880
rect 14380 13796 14420 13840
rect 19084 13796 19124 13840
rect 9379 13756 9388 13796
rect 9428 13756 10868 13796
rect 10915 13756 10924 13796
rect 10964 13756 14284 13796
rect 14324 13756 14333 13796
rect 14380 13756 15148 13796
rect 15188 13756 15197 13796
rect 15427 13756 15436 13796
rect 15476 13756 17740 13796
rect 17780 13756 17789 13796
rect 18953 13756 19084 13796
rect 19124 13756 19133 13796
rect 19555 13756 19564 13796
rect 19604 13756 19613 13796
rect 19747 13756 19756 13796
rect 19796 13756 22636 13796
rect 22676 13756 22685 13796
rect 10828 13712 10868 13756
rect 19564 13712 19604 13756
rect 23116 13712 23156 13989
rect 23404 13964 23444 14008
rect 23404 13924 24364 13964
rect 24404 13924 24413 13964
rect 24521 13924 24643 13964
rect 24692 13924 24701 13964
rect 26179 13924 26188 13964
rect 26228 13924 26237 13964
rect 26476 13924 26563 13964
rect 26603 13924 26612 13964
rect 26476 13796 26516 13924
rect 26668 13880 26708 14008
rect 29068 13964 29108 14008
rect 29884 13966 29932 14006
rect 29972 13966 29981 14006
rect 29884 13964 29924 13966
rect 28867 13924 28876 13964
rect 28916 13924 29108 13964
rect 29452 13924 29924 13964
rect 30953 13924 31084 13964
rect 31124 13924 31133 13964
rect 26668 13840 27916 13880
rect 27956 13840 27965 13880
rect 29452 13796 29492 13924
rect 24259 13756 24268 13796
rect 24308 13756 24652 13796
rect 24692 13756 25612 13796
rect 25652 13756 25661 13796
rect 25804 13756 26516 13796
rect 27322 13756 27331 13796
rect 27371 13756 29492 13796
rect 29548 13840 30316 13880
rect 30356 13840 30365 13880
rect 9763 13672 9772 13712
rect 9812 13672 10060 13712
rect 10100 13672 10109 13712
rect 10828 13672 11348 13712
rect 11395 13672 11404 13712
rect 11444 13672 19604 13712
rect 22147 13672 22156 13712
rect 22196 13672 23156 13712
rect 11308 13628 11348 13672
rect 10877 13588 10886 13628
rect 11254 13588 11263 13628
rect 11308 13588 16492 13628
rect 16532 13588 16541 13628
rect 18651 13588 18660 13628
rect 19028 13588 19037 13628
rect 19948 13588 23884 13628
rect 23924 13588 23933 13628
rect 9091 13504 9100 13544
rect 9140 13504 10484 13544
rect 16099 13504 16108 13544
rect 16148 13504 16163 13544
rect 10444 13460 10484 13504
rect 9004 13420 9571 13460
rect 9611 13420 9620 13460
rect 9955 13420 9964 13460
rect 10004 13420 10339 13460
rect 10379 13420 10388 13460
rect 10444 13420 12020 13460
rect 12739 13420 12748 13460
rect 12788 13420 13516 13460
rect 13556 13420 13565 13460
rect 14249 13420 14275 13460
rect 14315 13420 14380 13460
rect 14420 13420 14429 13460
rect 15113 13420 15244 13460
rect 15284 13420 15293 13460
rect 16003 13420 16012 13460
rect 16052 13420 16075 13460
rect 11980 13376 12020 13420
rect 6412 13336 6892 13376
rect 6932 13336 6941 13376
rect 7660 13336 8564 13376
rect 8620 13336 11875 13376
rect 11915 13336 11924 13376
rect 11980 13336 13748 13376
rect 14563 13336 14572 13376
rect 14612 13336 14804 13376
rect 15811 13336 15820 13376
rect 15860 13336 15869 13376
rect 1228 13252 2083 13292
rect 2123 13252 2132 13292
rect 2275 13252 2284 13292
rect 2324 13252 2333 13292
rect 4300 13252 5164 13292
rect 5204 13252 5213 13292
rect 5609 13252 5740 13292
rect 5780 13252 5789 13292
rect 5897 13283 6028 13292
rect 5897 13252 5971 13283
rect 4300 13208 4340 13252
rect 5962 13243 5971 13252
rect 6011 13252 6028 13283
rect 6068 13252 6077 13292
rect 6211 13252 6220 13292
rect 6260 13252 6302 13292
rect 6011 13243 6020 13252
rect 5962 13242 6020 13243
rect 1549 13168 1558 13208
rect 1598 13168 1612 13208
rect 1652 13168 1738 13208
rect 1934 13168 1943 13208
rect 1983 13168 1992 13208
rect 2083 13168 2092 13208
rect 2132 13168 2188 13208
rect 2228 13168 2263 13208
rect 2380 13168 2572 13208
rect 2612 13168 2621 13208
rect 2755 13168 2764 13208
rect 2804 13168 3043 13208
rect 3083 13168 3092 13208
rect 3139 13168 3148 13208
rect 3188 13168 3197 13208
rect 4169 13168 4300 13208
rect 4340 13168 4349 13208
rect 4426 13168 4435 13208
rect 4475 13168 4532 13208
rect 0 13124 400 13144
rect 1943 13124 1983 13168
rect 2380 13124 2420 13168
rect 0 13084 940 13124
rect 980 13084 989 13124
rect 1372 13084 1983 13124
rect 2179 13084 2188 13124
rect 2228 13084 2420 13124
rect 0 13064 400 13084
rect 1372 13040 1412 13084
rect 3148 13040 3188 13168
rect 1315 13000 1324 13040
rect 1403 13000 1495 13040
rect 2563 13000 2572 13040
rect 2612 13000 3188 13040
rect 3305 13000 3436 13040
rect 3476 13000 3485 13040
rect 4320 13000 4396 13040
rect 4436 13000 4445 13040
rect 4396 12956 4436 13000
rect 4204 12916 4436 12956
rect 4492 12956 4532 13168
rect 4588 13168 4804 13208
rect 4844 13168 4853 13208
rect 4968 13168 4977 13208
rect 5017 13168 5026 13208
rect 5080 13168 5089 13208
rect 5129 13168 5138 13208
rect 5242 13179 5251 13219
rect 5291 13179 5300 13219
rect 6220 13208 6260 13252
rect 6412 13208 6452 13336
rect 6665 13252 6787 13292
rect 6836 13252 6845 13292
rect 6979 13252 6988 13292
rect 7028 13252 7159 13292
rect 7468 13208 7508 13217
rect 7660 13208 7700 13336
rect 8524 13292 8564 13336
rect 13708 13292 13748 13336
rect 14764 13292 14804 13336
rect 8524 13252 8899 13292
rect 8939 13252 8948 13292
rect 9065 13252 9100 13292
rect 9140 13252 9196 13292
rect 9236 13252 9245 13292
rect 11417 13252 11500 13292
rect 11540 13283 11588 13292
rect 8285 13210 8332 13250
rect 8372 13241 8456 13250
rect 8372 13210 8416 13241
rect 4588 13040 4628 13168
rect 4972 13124 5012 13168
rect 4930 13084 4972 13124
rect 5012 13084 5021 13124
rect 5080 13040 5120 13168
rect 5260 13124 5300 13179
rect 5364 13168 5373 13208
rect 5413 13168 5422 13208
rect 5705 13168 5836 13208
rect 5876 13168 5885 13208
rect 6067 13168 6076 13208
rect 6116 13168 6125 13208
rect 6206 13168 6215 13208
rect 6255 13168 6264 13208
rect 6394 13168 6403 13208
rect 6443 13168 6452 13208
rect 6595 13168 6604 13208
rect 6644 13168 6647 13208
rect 6687 13168 6775 13208
rect 6883 13168 6892 13208
rect 6932 13168 7316 13208
rect 7363 13168 7372 13208
rect 7412 13168 7468 13208
rect 7508 13168 7651 13208
rect 7691 13168 7700 13208
rect 7747 13168 7756 13208
rect 7796 13168 7852 13208
rect 7892 13168 7927 13208
rect 8524 13208 8564 13252
rect 9868 13208 9908 13217
rect 10339 13210 10348 13250
rect 10388 13241 10664 13250
rect 11530 13243 11539 13252
rect 11579 13243 11588 13283
rect 12643 13252 12652 13292
rect 12692 13252 12980 13292
rect 13699 13252 13708 13292
rect 13748 13252 13757 13292
rect 14755 13252 14764 13292
rect 14804 13252 14813 13292
rect 14860 13252 15148 13292
rect 15188 13252 15197 13292
rect 15244 13252 15436 13292
rect 15476 13252 15485 13292
rect 11530 13242 11588 13243
rect 10388 13210 10624 13241
rect 8416 13192 8456 13201
rect 8506 13168 8515 13208
rect 8555 13168 8564 13208
rect 8707 13168 8716 13208
rect 8756 13168 8759 13208
rect 8799 13168 8887 13208
rect 8995 13168 9004 13208
rect 9044 13168 9053 13208
rect 9737 13168 9772 13208
rect 9812 13168 9868 13208
rect 12940 13208 12980 13252
rect 14572 13208 14612 13217
rect 14860 13208 14900 13252
rect 15244 13208 15284 13252
rect 10624 13192 10664 13201
rect 10714 13168 10723 13208
rect 10763 13168 10828 13208
rect 10868 13168 10903 13208
rect 11273 13168 11404 13208
rect 11444 13168 11453 13208
rect 11632 13168 11641 13208
rect 11681 13168 12212 13208
rect 12259 13168 12268 13208
rect 12308 13168 12556 13208
rect 12596 13168 12605 13208
rect 12922 13168 12931 13208
rect 12971 13168 12980 13208
rect 13027 13168 13036 13208
rect 13076 13168 13228 13208
rect 13268 13168 13795 13208
rect 13835 13168 13844 13208
rect 14083 13168 14092 13208
rect 14132 13168 14270 13208
rect 14310 13168 14319 13208
rect 14441 13168 14572 13208
rect 14612 13168 14621 13208
rect 14851 13168 14860 13208
rect 14900 13168 14909 13208
rect 14970 13168 14979 13208
rect 15019 13168 15028 13208
rect 15088 13168 15097 13208
rect 15137 13168 15188 13208
rect 15235 13168 15244 13208
rect 15284 13168 15293 13208
rect 15360 13168 15369 13208
rect 15409 13168 15418 13208
rect 15523 13168 15532 13208
rect 15572 13168 15628 13208
rect 15668 13168 15703 13208
rect 5382 13124 5422 13168
rect 5251 13084 5260 13124
rect 5300 13084 5336 13124
rect 5382 13084 5684 13124
rect 4579 13000 4588 13040
rect 4628 13000 4637 13040
rect 4745 13000 4867 13040
rect 4916 13000 4925 13040
rect 5080 13000 5452 13040
rect 5492 13000 5501 13040
rect 5644 12956 5684 13084
rect 6076 13040 6116 13168
rect 7276 13124 7316 13168
rect 7468 13159 7508 13168
rect 9004 13124 9044 13168
rect 9868 13159 9908 13168
rect 12172 13124 12212 13168
rect 7157 13084 7166 13124
rect 7206 13084 7215 13124
rect 7258 13084 7267 13124
rect 7307 13084 7316 13124
rect 7564 13084 7756 13124
rect 7796 13084 7805 13124
rect 7913 13084 7962 13124
rect 8002 13084 8044 13124
rect 8084 13084 8093 13124
rect 8524 13084 9044 13124
rect 9435 13084 9484 13124
rect 9524 13084 9566 13124
rect 9606 13084 9615 13124
rect 9955 13084 9964 13124
rect 10004 13084 11308 13124
rect 11348 13084 11357 13124
rect 11849 13084 11971 13124
rect 12020 13084 12029 13124
rect 12172 13084 12748 13124
rect 12788 13084 12797 13124
rect 6019 13000 6028 13040
rect 6068 13000 6116 13040
rect 6185 13000 6316 13040
rect 6356 13000 6365 13040
rect 7166 12956 7206 13084
rect 7564 13040 7604 13084
rect 8524 13040 8564 13084
rect 12940 13040 12980 13168
rect 14572 13159 14612 13168
rect 14275 13084 14284 13124
rect 14324 13084 14476 13124
rect 14516 13084 14525 13124
rect 7363 13000 7372 13040
rect 7412 13000 7604 13040
rect 7843 13000 7852 13040
rect 7892 13000 8564 13040
rect 8649 13000 8658 13040
rect 8698 13000 8812 13040
rect 8852 13000 9100 13040
rect 9140 13000 9149 13040
rect 9763 13000 9772 13040
rect 9812 13000 9868 13040
rect 9908 13000 9943 13040
rect 10435 13000 10444 13040
rect 10484 13000 10843 13040
rect 10883 13000 10892 13040
rect 11779 13000 11788 13040
rect 11828 13000 12364 13040
rect 12404 13000 12692 13040
rect 12940 13000 13411 13040
rect 13451 13000 13460 13040
rect 13603 13000 13612 13040
rect 13652 13000 14420 13040
rect 12652 12956 12692 13000
rect 14380 12956 14420 13000
rect 14979 12956 15019 13168
rect 15148 13124 15188 13168
rect 15378 13124 15418 13168
rect 15820 13124 15860 13336
rect 16035 13292 16075 13420
rect 16123 13376 16163 13504
rect 16285 13504 17644 13544
rect 17684 13504 19180 13544
rect 19220 13504 19229 13544
rect 16123 13336 16196 13376
rect 16026 13252 16035 13292
rect 16075 13252 16084 13292
rect 16156 13250 16196 13336
rect 16147 13210 16156 13250
rect 16196 13210 16205 13250
rect 16285 13229 16325 13504
rect 16972 13420 19084 13460
rect 19124 13420 19133 13460
rect 19555 13420 19564 13460
rect 19604 13420 19852 13460
rect 19892 13420 19901 13460
rect 16378 13252 16387 13292
rect 16436 13252 16567 13292
rect 16276 13208 16325 13229
rect 16972 13208 17012 13420
rect 19948 13376 19988 13588
rect 25804 13460 25844 13756
rect 26425 13588 26434 13628
rect 26802 13588 26811 13628
rect 20969 13420 21100 13460
rect 21140 13420 21149 13460
rect 21283 13420 21292 13460
rect 21332 13420 23060 13460
rect 23369 13420 23491 13460
rect 23540 13420 23549 13460
rect 24355 13420 24364 13460
rect 24404 13420 24460 13460
rect 24500 13420 24535 13460
rect 25795 13420 25804 13460
rect 25844 13420 25853 13460
rect 27689 13420 27820 13460
rect 27860 13420 27869 13460
rect 17932 13336 18316 13376
rect 18356 13336 19508 13376
rect 17932 13292 17972 13336
rect 17923 13252 17932 13292
rect 17972 13252 17981 13292
rect 18499 13252 18508 13292
rect 18548 13252 18557 13292
rect 17452 13208 17492 13217
rect 18513 13208 18553 13252
rect 19468 13208 19508 13336
rect 15907 13168 15916 13208
rect 15956 13168 15965 13208
rect 16258 13168 16267 13208
rect 16307 13189 16325 13208
rect 16307 13168 16316 13189
rect 16483 13168 16492 13208
rect 16532 13168 16780 13208
rect 16820 13168 16829 13208
rect 16954 13168 16963 13208
rect 17003 13168 17012 13208
rect 17321 13168 17452 13208
rect 17492 13168 17501 13208
rect 17635 13168 17644 13208
rect 17684 13168 18028 13208
rect 18068 13168 18077 13208
rect 18281 13168 18316 13208
rect 18356 13168 18412 13208
rect 18452 13168 18461 13208
rect 18504 13168 18513 13208
rect 18553 13168 18595 13208
rect 19075 13168 19084 13208
rect 19124 13168 19180 13208
rect 19220 13168 19255 13208
rect 19450 13168 19459 13208
rect 19499 13168 19508 13208
rect 19564 13336 19988 13376
rect 21475 13336 21484 13376
rect 21524 13336 21533 13376
rect 21676 13336 22540 13376
rect 22580 13336 22589 13376
rect 15916 13124 15956 13168
rect 17452 13159 17492 13168
rect 18028 13124 18068 13168
rect 19564 13124 19604 13336
rect 21484 13292 21524 13336
rect 20428 13252 21524 13292
rect 20428 13208 20468 13252
rect 21100 13208 21140 13252
rect 21676 13208 21716 13336
rect 21868 13252 22636 13292
rect 22676 13252 22685 13292
rect 20419 13168 20428 13208
rect 20468 13168 20477 13208
rect 20524 13199 20620 13208
rect 20564 13168 20620 13199
rect 20660 13168 20695 13208
rect 20803 13168 20812 13208
rect 20852 13168 20861 13208
rect 21091 13168 21100 13208
rect 21140 13168 21149 13208
rect 21283 13168 21292 13208
rect 21332 13168 21341 13208
rect 21676 13168 21772 13208
rect 21812 13168 21821 13208
rect 21868 13199 21908 13252
rect 23020 13208 23060 13420
rect 23945 13336 24076 13376
rect 24116 13336 24125 13376
rect 24259 13336 24268 13376
rect 24308 13336 25364 13376
rect 25324 13208 25364 13336
rect 25938 13252 26092 13292
rect 26132 13252 26141 13292
rect 26275 13252 26284 13292
rect 26324 13252 26419 13292
rect 26459 13252 26468 13292
rect 26899 13252 26908 13292
rect 26948 13252 27148 13292
rect 27188 13252 27197 13292
rect 29548 13272 29588 13840
rect 29923 13756 29932 13796
rect 29972 13756 29981 13796
rect 29932 13292 29972 13756
rect 30595 13336 30604 13376
rect 30644 13336 30796 13376
rect 30836 13336 30845 13376
rect 29722 13252 29731 13292
rect 29771 13252 29972 13292
rect 30604 13252 31276 13292
rect 31316 13252 31325 13292
rect 25938 13208 25978 13252
rect 30604 13208 30644 13252
rect 20524 13150 20564 13159
rect 20812 13124 20852 13168
rect 21292 13124 21332 13168
rect 22025 13168 22156 13208
rect 22196 13168 22205 13208
rect 22313 13168 22444 13208
rect 22484 13168 22493 13208
rect 23020 13168 23452 13208
rect 23492 13168 23501 13208
rect 23587 13168 23596 13208
rect 23636 13168 23645 13208
rect 23875 13168 23884 13208
rect 23924 13168 25132 13208
rect 25172 13168 25181 13208
rect 25306 13168 25315 13208
rect 25355 13168 25364 13208
rect 25795 13168 25804 13208
rect 25844 13168 25853 13208
rect 25920 13168 25929 13208
rect 25969 13168 25978 13208
rect 26083 13168 26092 13208
rect 26132 13168 26141 13208
rect 26462 13168 26572 13208
rect 26624 13168 26642 13208
rect 26743 13168 26752 13208
rect 26792 13168 26801 13208
rect 29225 13168 29347 13208
rect 29396 13168 29405 13208
rect 29644 13168 29875 13208
rect 29915 13168 29924 13208
rect 30403 13168 30412 13208
rect 30452 13168 30461 13208
rect 30595 13168 30604 13208
rect 30644 13168 30653 13208
rect 31049 13168 31180 13208
rect 31220 13168 31229 13208
rect 21868 13150 21908 13159
rect 23596 13124 23636 13168
rect 15148 13084 15244 13124
rect 15284 13084 15293 13124
rect 15378 13084 15532 13124
rect 15572 13084 15581 13124
rect 15811 13084 15820 13124
rect 15860 13084 15869 13124
rect 15916 13084 16579 13124
rect 16619 13084 16628 13124
rect 18028 13084 19564 13124
rect 19604 13084 19613 13124
rect 20812 13084 21332 13124
rect 22819 13084 22828 13124
rect 22868 13084 23636 13124
rect 24172 13084 25623 13124
rect 25663 13084 25672 13124
rect 20812 13040 20852 13084
rect 16483 13000 16492 13040
rect 16532 13000 16780 13040
rect 16820 13000 16829 13040
rect 17356 13000 20092 13040
rect 20132 13000 20141 13040
rect 20227 13000 20236 13040
rect 20276 13000 20852 13040
rect 23107 13000 23116 13040
rect 23156 13000 23287 13040
rect 17356 12956 17396 13000
rect 24172 12956 24212 13084
rect 25804 13040 25844 13168
rect 26092 13124 26132 13168
rect 25891 13084 25900 13124
rect 25940 13084 26132 13124
rect 24835 13000 24844 13040
rect 24884 13000 25228 13040
rect 25268 13000 25411 13040
rect 25451 13000 25460 13040
rect 25507 13000 25516 13040
rect 25556 13000 25844 13040
rect 26761 13040 26801 13168
rect 29644 13124 29684 13168
rect 30412 13124 30452 13168
rect 27418 13084 27427 13124
rect 27467 13084 29684 13124
rect 29731 13084 29740 13124
rect 29780 13084 30452 13124
rect 26761 13000 26956 13040
rect 26996 13000 30076 13040
rect 30116 13000 30125 13040
rect 30220 13000 30595 13040
rect 30635 13000 30644 13040
rect 30220 12956 30260 13000
rect 4492 12916 4820 12956
rect 5644 12916 6892 12956
rect 6932 12916 8620 12956
rect 8660 12916 9388 12956
rect 9428 12916 12596 12956
rect 12652 12916 12844 12956
rect 12884 12916 13996 12956
rect 14036 12916 14045 12956
rect 14371 12916 14380 12956
rect 14420 12916 14496 12956
rect 14979 12916 15947 12956
rect 16195 12916 16204 12956
rect 16244 12916 17396 12956
rect 17635 12916 17644 12956
rect 17684 12916 20428 12956
rect 20468 12916 20477 12956
rect 23299 12916 23308 12956
rect 23348 12916 24212 12956
rect 28579 12916 28588 12956
rect 28628 12916 30260 12956
rect 2380 12748 2900 12788
rect 0 12704 400 12724
rect 2380 12704 2420 12748
rect 2860 12704 2900 12748
rect 4204 12704 4244 12916
rect 4343 12832 4352 12872
rect 4720 12832 4729 12872
rect 4780 12788 4820 12916
rect 12556 12872 12596 12916
rect 4588 12748 4820 12788
rect 5740 12832 11404 12872
rect 11444 12832 11453 12872
rect 12117 12832 12126 12872
rect 12494 12832 12503 12872
rect 12556 12832 12652 12872
rect 12692 12832 12701 12872
rect 4588 12704 4628 12748
rect 0 12664 1036 12704
rect 1076 12664 1085 12704
rect 1219 12664 1228 12704
rect 1268 12664 1277 12704
rect 1987 12664 1996 12704
rect 2036 12664 2045 12704
rect 2371 12664 2380 12704
rect 2420 12664 2429 12704
rect 2860 12664 4148 12704
rect 4204 12664 4291 12704
rect 4331 12664 4340 12704
rect 4570 12664 4579 12704
rect 4619 12664 4628 12704
rect 0 12644 400 12664
rect 1228 12620 1268 12664
rect 1228 12580 1748 12620
rect 1708 12536 1748 12580
rect 1996 12536 2036 12664
rect 2481 12580 2490 12620
rect 2530 12580 2947 12620
rect 2987 12580 2996 12620
rect 4108 12536 4148 12664
rect 5740 12620 5780 12832
rect 5827 12748 5836 12788
rect 5876 12748 6356 12788
rect 6316 12704 6356 12748
rect 6604 12748 10292 12788
rect 5897 12664 5932 12704
rect 5972 12664 6028 12704
rect 6068 12664 6077 12704
rect 6307 12664 6316 12704
rect 6356 12664 6365 12704
rect 4204 12580 5780 12620
rect 6028 12580 6316 12620
rect 6356 12580 6365 12620
rect 4204 12536 4244 12580
rect 6028 12536 6068 12580
rect 6604 12536 6644 12748
rect 7555 12664 7564 12704
rect 7604 12664 7613 12704
rect 7747 12664 7756 12704
rect 7796 12664 9009 12704
rect 9449 12664 9571 12704
rect 9620 12664 9629 12704
rect 9676 12664 9964 12704
rect 10004 12664 10013 12704
rect 7564 12536 7604 12664
rect 8969 12620 9009 12664
rect 9676 12620 9716 12664
rect 8332 12580 8812 12620
rect 8852 12580 8861 12620
rect 8969 12580 9716 12620
rect 9850 12611 10156 12620
rect 8332 12536 8372 12580
rect 8969 12536 9009 12580
rect 9850 12571 9859 12611
rect 9899 12580 10156 12611
rect 10196 12580 10205 12620
rect 9899 12571 9908 12580
rect 9850 12570 9908 12571
rect 931 12496 940 12536
rect 980 12496 989 12536
rect 1066 12496 1075 12536
rect 1115 12496 1324 12536
rect 1364 12496 1373 12536
rect 1594 12496 1603 12536
rect 1643 12496 1652 12536
rect 1699 12496 1708 12536
rect 1748 12496 1879 12536
rect 1996 12496 2179 12536
rect 2219 12496 2228 12536
rect 2275 12496 2284 12536
rect 2324 12496 2615 12536
rect 2655 12496 2664 12536
rect 2851 12496 2860 12536
rect 2900 12496 2909 12536
rect 3828 12496 3916 12536
rect 3956 12496 3959 12536
rect 3999 12496 4008 12536
rect 4090 12496 4099 12536
rect 4139 12496 4148 12536
rect 4195 12496 4204 12536
rect 4244 12496 4253 12536
rect 4771 12496 4780 12536
rect 4820 12496 4829 12536
rect 4937 12496 5068 12536
rect 5108 12496 5117 12536
rect 5251 12496 5260 12536
rect 5300 12496 5309 12536
rect 5443 12496 5452 12536
rect 5492 12496 5501 12536
rect 5705 12496 5836 12536
rect 5876 12496 5885 12536
rect 6010 12496 6019 12536
rect 6059 12496 6068 12536
rect 6222 12496 6231 12536
rect 6271 12496 6341 12536
rect 6394 12496 6403 12536
rect 6443 12496 6644 12536
rect 6691 12496 6700 12536
rect 6740 12496 7084 12536
rect 7124 12496 7133 12536
rect 7337 12496 7468 12536
rect 7508 12496 7517 12536
rect 7564 12496 8194 12536
rect 8314 12496 8323 12536
rect 8363 12496 8372 12536
rect 8611 12496 8620 12536
rect 8660 12496 8668 12536
rect 8708 12496 8791 12536
rect 8960 12496 8969 12536
rect 9009 12496 9018 12536
rect 9065 12496 9139 12536
rect 9179 12496 9196 12536
rect 9236 12496 9245 12536
rect 9379 12496 9388 12536
rect 9428 12496 9571 12536
rect 9611 12496 9620 12536
rect 9676 12527 9716 12536
rect 940 12452 980 12496
rect 1612 12452 1652 12496
rect 2188 12452 2228 12496
rect 940 12412 1516 12452
rect 1556 12412 1565 12452
rect 1612 12412 2092 12452
rect 2132 12412 2141 12452
rect 2188 12412 2755 12452
rect 2795 12412 2804 12452
rect 2860 12200 2900 12496
rect 4780 12452 4820 12496
rect 5260 12452 5300 12496
rect 4745 12412 4876 12452
rect 4916 12412 5300 12452
rect 5452 12452 5492 12496
rect 6301 12452 6341 12496
rect 8154 12452 8194 12496
rect 9942 12496 9951 12536
rect 9991 12496 10004 12536
rect 9676 12452 9716 12487
rect 9964 12452 10004 12496
rect 10123 12485 10132 12525
rect 10172 12485 10196 12525
rect 5452 12412 5780 12452
rect 6301 12412 6892 12452
rect 6932 12412 6941 12452
rect 7913 12412 7939 12452
rect 7979 12412 8044 12452
rect 8084 12412 8093 12452
rect 8154 12412 8515 12452
rect 8555 12412 8620 12452
rect 8660 12412 8724 12452
rect 8803 12412 8812 12452
rect 8852 12412 8983 12452
rect 9667 12412 9676 12452
rect 9716 12412 9763 12452
rect 9955 12412 9964 12452
rect 10004 12412 10047 12452
rect 5452 12368 5492 12412
rect 5740 12368 5780 12412
rect 10156 12368 10196 12485
rect 5059 12328 5068 12368
rect 5108 12328 5492 12368
rect 5731 12328 5740 12368
rect 5780 12328 5789 12368
rect 6595 12328 6604 12368
rect 6644 12328 8035 12368
rect 8075 12328 8084 12368
rect 8777 12328 8908 12368
rect 8948 12328 8957 12368
rect 10060 12328 10196 12368
rect 10252 12368 10292 12748
rect 12796 12748 14092 12788
rect 14132 12748 14141 12788
rect 12796 12704 12836 12748
rect 15907 12704 15947 12916
rect 19891 12832 19900 12872
rect 20268 12832 20277 12872
rect 21187 12832 21196 12872
rect 21236 12832 24076 12872
rect 24116 12832 24125 12872
rect 27665 12832 27674 12872
rect 28042 12832 28051 12872
rect 18892 12748 23060 12788
rect 28387 12748 28396 12788
rect 28436 12748 30316 12788
rect 30356 12748 30365 12788
rect 10723 12664 10732 12704
rect 10772 12664 11011 12704
rect 11051 12664 11060 12704
rect 11491 12664 11500 12704
rect 11540 12664 11692 12704
rect 11732 12664 11741 12704
rect 12787 12664 12796 12704
rect 12836 12664 12845 12704
rect 13315 12664 13324 12704
rect 13364 12664 13708 12704
rect 13748 12664 13757 12704
rect 14563 12664 14572 12704
rect 14612 12664 15052 12704
rect 15092 12664 15739 12704
rect 15779 12664 15788 12704
rect 15907 12664 16012 12704
rect 16052 12664 16061 12704
rect 16771 12664 16780 12704
rect 16820 12664 17020 12704
rect 17060 12664 17069 12704
rect 18403 12664 18412 12704
rect 18452 12664 18691 12704
rect 18731 12664 18740 12704
rect 10348 12580 11788 12620
rect 11828 12580 11837 12620
rect 11884 12580 12268 12620
rect 12308 12580 12317 12620
rect 12643 12580 12652 12620
rect 12692 12580 12712 12620
rect 14668 12580 15532 12620
rect 15572 12580 15581 12620
rect 16483 12580 16492 12620
rect 16532 12580 16723 12620
rect 16763 12580 16772 12620
rect 17068 12580 17452 12620
rect 17492 12580 18028 12620
rect 18068 12580 18077 12620
rect 18412 12580 18796 12620
rect 18836 12580 18845 12620
rect 10348 12536 10388 12580
rect 11884 12536 11924 12580
rect 12652 12536 12692 12580
rect 14668 12536 14708 12580
rect 17068 12536 17108 12580
rect 10339 12496 10348 12536
rect 10388 12496 10397 12536
rect 10444 12496 10463 12536
rect 10503 12496 10512 12536
rect 10627 12496 10636 12536
rect 10676 12496 10924 12536
rect 10964 12496 10973 12536
rect 11033 12496 11116 12536
rect 11156 12496 11164 12536
rect 11204 12496 11213 12536
rect 11299 12496 11308 12536
rect 11348 12496 11357 12536
rect 11587 12496 11596 12536
rect 11636 12496 11645 12536
rect 11824 12496 11833 12536
rect 11873 12496 11924 12536
rect 11971 12496 11980 12536
rect 12020 12496 12116 12536
rect 12163 12496 12172 12536
rect 12212 12496 12343 12536
rect 12607 12496 12616 12536
rect 12656 12496 12692 12536
rect 12924 12496 12940 12536
rect 12980 12496 13084 12536
rect 13124 12496 13133 12536
rect 13385 12496 13420 12536
rect 13460 12496 13516 12536
rect 13556 12496 13565 12536
rect 13673 12496 13804 12536
rect 13844 12496 13853 12536
rect 13987 12496 13996 12536
rect 14036 12496 14041 12536
rect 14081 12496 14476 12536
rect 14516 12496 14525 12536
rect 14650 12496 14659 12536
rect 14699 12496 14708 12536
rect 14755 12496 14764 12536
rect 14804 12496 15052 12536
rect 15092 12496 15101 12536
rect 15389 12496 15436 12536
rect 15476 12527 15560 12536
rect 15476 12496 15520 12527
rect 10252 12328 10348 12368
rect 10388 12328 10397 12368
rect 10060 12284 10100 12328
rect 4963 12244 4972 12284
rect 5012 12244 5260 12284
rect 5300 12244 5309 12284
rect 9955 12244 9964 12284
rect 10004 12244 10100 12284
rect 2860 12160 8332 12200
rect 8372 12160 9868 12200
rect 9908 12160 9917 12200
rect 10444 12116 10484 12496
rect 11308 12368 11348 12496
rect 11596 12452 11636 12496
rect 11395 12412 11404 12452
rect 11444 12412 11636 12452
rect 11722 12443 11780 12452
rect 11722 12403 11731 12443
rect 11771 12403 11780 12443
rect 11722 12402 11780 12403
rect 11740 12368 11780 12402
rect 11308 12328 11500 12368
rect 11540 12328 11549 12368
rect 11740 12328 11980 12368
rect 12020 12328 12029 12368
rect 12076 12284 12116 12496
rect 15811 12496 15820 12536
rect 15860 12496 15916 12536
rect 15956 12496 15991 12536
rect 16099 12496 16108 12536
rect 16148 12496 16204 12536
rect 16244 12496 16279 12536
rect 16909 12496 16918 12536
rect 16958 12496 17108 12536
rect 17155 12496 17164 12536
rect 17204 12496 17335 12536
rect 17453 12496 17879 12536
rect 17919 12496 17928 12536
rect 18115 12496 18124 12536
rect 18164 12496 18173 12536
rect 18220 12496 18316 12536
rect 18356 12496 18365 12536
rect 15520 12478 15560 12487
rect 15610 12454 15619 12494
rect 15659 12454 15668 12494
rect 13315 12412 13324 12452
rect 13364 12412 13923 12452
rect 13963 12412 13972 12452
rect 14371 12412 14380 12452
rect 14420 12412 15480 12452
rect 15440 12368 15480 12412
rect 15628 12368 15668 12454
rect 15916 12452 15956 12496
rect 17453 12452 17493 12496
rect 15916 12412 16396 12452
rect 16436 12412 16445 12452
rect 16963 12412 16972 12452
rect 17012 12412 17493 12452
rect 17635 12412 17644 12452
rect 17684 12412 18019 12452
rect 18059 12412 18068 12452
rect 18124 12368 18164 12496
rect 18220 12452 18260 12496
rect 18412 12452 18452 12580
rect 18499 12496 18508 12536
rect 18548 12496 18590 12536
rect 18630 12496 18679 12536
rect 18892 12527 18932 12748
rect 20227 12664 20236 12704
rect 20276 12664 22444 12704
rect 22484 12664 22493 12704
rect 23020 12620 23060 12748
rect 29251 12664 29260 12704
rect 29300 12664 29740 12704
rect 29780 12664 29789 12704
rect 22156 12580 22924 12620
rect 22964 12580 22973 12620
rect 23020 12580 24116 12620
rect 22156 12536 22196 12580
rect 19651 12496 19660 12536
rect 19700 12496 21676 12536
rect 21716 12496 21725 12536
rect 22138 12496 22147 12536
rect 22187 12496 22196 12536
rect 23053 12496 23062 12536
rect 23102 12496 23116 12536
rect 23156 12496 23242 12536
rect 18892 12478 18932 12487
rect 18211 12412 18220 12452
rect 18260 12412 18269 12452
rect 18403 12412 18412 12452
rect 18452 12412 18461 12452
rect 19459 12412 19468 12452
rect 19508 12412 19570 12452
rect 19610 12412 19639 12452
rect 20515 12412 20524 12452
rect 20564 12412 20611 12452
rect 20651 12412 20695 12452
rect 15113 12328 15235 12368
rect 15284 12328 15293 12368
rect 15440 12328 16876 12368
rect 16916 12328 16925 12368
rect 17347 12328 17356 12368
rect 17396 12328 18164 12368
rect 20076 12328 20140 12368
rect 20180 12328 20236 12368
rect 20276 12328 20285 12368
rect 11299 12244 11308 12284
rect 11348 12244 13219 12284
rect 13259 12244 15820 12284
rect 15860 12244 15869 12284
rect 19459 12244 19468 12284
rect 19508 12244 19517 12284
rect 20419 12244 20428 12284
rect 20468 12244 21100 12284
rect 21140 12244 21149 12284
rect 19468 12200 19508 12244
rect 11491 12160 11500 12200
rect 11540 12160 19508 12200
rect 3103 12076 3112 12116
rect 3480 12076 3489 12116
rect 5731 12076 5740 12116
rect 5780 12076 6124 12116
rect 6164 12076 6173 12116
rect 9091 12076 9100 12116
rect 9140 12076 10484 12116
rect 10877 12076 10886 12116
rect 11254 12076 11263 12116
rect 13027 12076 13036 12116
rect 13076 12076 17068 12116
rect 17108 12076 18412 12116
rect 18452 12076 18461 12116
rect 18651 12076 18660 12116
rect 19028 12076 19037 12116
rect 19171 12076 19180 12116
rect 19220 12076 21580 12116
rect 21620 12076 21629 12116
rect 18412 12032 18452 12076
rect 9955 11992 9964 12032
rect 10004 11992 10100 12032
rect 10060 11948 10100 11992
rect 12940 11992 13228 12032
rect 13268 11992 13277 12032
rect 13507 11992 13516 12032
rect 13556 11992 15572 12032
rect 12940 11948 12980 11992
rect 1411 11908 1420 11948
rect 1460 11908 1940 11948
rect 2083 11908 2092 11948
rect 2132 11908 2284 11948
rect 2324 11908 2333 11948
rect 2860 11908 3916 11948
rect 3956 11908 3965 11948
rect 4745 11908 4780 11948
rect 4820 11908 4876 11948
rect 4916 11908 4925 11948
rect 5609 11908 5644 11948
rect 5684 11908 5740 11948
rect 5780 11908 5789 11948
rect 6595 11908 6604 11948
rect 6644 11908 6796 11948
rect 6836 11908 6845 11948
rect 7166 11908 7180 11948
rect 7220 11908 7988 11948
rect 9353 11908 9475 11948
rect 9524 11908 9533 11948
rect 10051 11908 10060 11948
rect 10100 11908 10109 11948
rect 11587 11908 11596 11948
rect 11636 11908 11779 11948
rect 11819 11908 11828 11948
rect 12922 11908 12931 11948
rect 12971 11908 12980 11948
rect 1036 11824 1420 11864
rect 1460 11824 1469 11864
rect 1036 11696 1076 11824
rect 1900 11696 1940 11908
rect 2860 11864 2900 11908
rect 7166 11864 7206 11908
rect 1996 11824 2900 11864
rect 3331 11824 3340 11864
rect 3380 11824 3389 11864
rect 6115 11824 6124 11864
rect 6164 11824 7206 11864
rect 7258 11824 7267 11864
rect 7307 11824 7316 11864
rect 1996 11780 2036 11824
rect 3340 11780 3380 11824
rect 7276 11780 7316 11824
rect 1987 11740 1996 11780
rect 2036 11740 2045 11780
rect 3340 11740 4532 11780
rect 4492 11738 4532 11740
rect 5164 11740 5836 11780
rect 5876 11740 5885 11780
rect 6988 11740 7084 11780
rect 7124 11740 7133 11780
rect 7241 11740 7372 11780
rect 7412 11740 7762 11780
rect 7802 11740 7811 11780
rect 4492 11729 4536 11738
rect 4492 11698 4496 11729
rect 748 11656 940 11696
rect 980 11656 989 11696
rect 1036 11656 1123 11696
rect 1163 11656 1172 11696
rect 1314 11656 1323 11696
rect 1363 11656 1411 11696
rect 1469 11656 1515 11696
rect 1555 11656 1564 11696
rect 1651 11656 1660 11696
rect 1700 11656 1709 11696
rect 1786 11656 1795 11696
rect 1835 11656 1844 11696
rect 1891 11656 1900 11696
rect 1940 11656 1949 11696
rect 2057 11656 2188 11696
rect 2228 11656 2237 11696
rect 2371 11656 2380 11696
rect 2420 11656 2668 11696
rect 2708 11656 2717 11696
rect 3139 11656 3148 11696
rect 3188 11656 3197 11696
rect 3401 11656 3532 11696
rect 3572 11656 3581 11696
rect 3881 11656 3916 11696
rect 3956 11656 4012 11696
rect 4052 11656 4061 11696
rect 4378 11656 4387 11696
rect 4427 11656 4436 11696
rect 5164 11696 5204 11740
rect 6988 11696 7028 11740
rect 7948 11696 7988 11908
rect 12940 11864 12980 11908
rect 8667 11824 10348 11864
rect 10388 11824 10397 11864
rect 10492 11824 11884 11864
rect 11924 11824 11933 11864
rect 12508 11824 12980 11864
rect 13132 11908 13708 11948
rect 13748 11908 13757 11948
rect 14851 11908 14860 11948
rect 14900 11908 15340 11948
rect 15380 11908 15389 11948
rect 8667 11738 8707 11824
rect 9484 11740 9868 11780
rect 9908 11740 9917 11780
rect 8650 11698 8659 11738
rect 8699 11698 8708 11738
rect 9484 11696 9524 11740
rect 4496 11680 4536 11689
rect 4867 11656 4876 11696
rect 4916 11656 4972 11696
rect 5012 11656 5047 11696
rect 5155 11656 5164 11696
rect 5204 11656 5213 11696
rect 5338 11656 5347 11696
rect 5387 11656 5740 11696
rect 5780 11656 5789 11696
rect 5897 11656 5932 11696
rect 5972 11656 6028 11696
rect 6068 11656 6077 11696
rect 6185 11656 6307 11696
rect 6356 11656 6365 11696
rect 6970 11656 6979 11696
rect 7019 11656 7028 11696
rect 7075 11656 7084 11696
rect 7124 11656 7796 11696
rect 7843 11656 7852 11696
rect 7892 11656 7988 11696
rect 8777 11656 8800 11696
rect 8840 11656 8908 11696
rect 8948 11656 8957 11696
rect 9283 11656 9292 11696
rect 9332 11656 9341 11696
rect 9466 11656 9475 11696
rect 9515 11656 9524 11696
rect 9850 11656 9859 11696
rect 9899 11656 9908 11696
rect 9955 11656 9964 11717
rect 10004 11696 10013 11717
rect 10492 11696 10532 11824
rect 12508 11780 12548 11824
rect 13132 11780 13172 11908
rect 13507 11824 13516 11864
rect 13556 11824 14380 11864
rect 14420 11824 14429 11864
rect 14476 11824 15146 11864
rect 10579 11740 10588 11780
rect 10628 11740 11788 11780
rect 11828 11740 11837 11780
rect 12490 11771 12548 11780
rect 12490 11731 12499 11771
rect 12539 11731 12548 11771
rect 12937 11740 12946 11780
rect 12986 11740 13172 11780
rect 13219 11740 13228 11780
rect 13268 11740 13603 11780
rect 13643 11740 13652 11780
rect 12490 11730 12548 11731
rect 12076 11696 12116 11705
rect 14476 11696 14516 11824
rect 15106 11780 15146 11824
rect 14851 11740 14860 11780
rect 14900 11740 14996 11780
rect 14572 11696 14612 11705
rect 14956 11696 14996 11740
rect 15106 11740 15244 11780
rect 15284 11740 15293 11780
rect 15427 11740 15436 11780
rect 15476 11740 15485 11780
rect 15106 11696 15146 11740
rect 15436 11696 15476 11740
rect 10004 11656 10114 11696
rect 10243 11656 10252 11696
rect 10292 11656 10301 11696
rect 10423 11656 10432 11696
rect 10472 11656 10532 11696
rect 11011 11656 11020 11696
rect 11060 11656 11069 11696
rect 11177 11656 11308 11696
rect 11348 11656 11357 11696
rect 12233 11656 12364 11696
rect 12404 11656 12413 11696
rect 12592 11656 12601 11696
rect 12641 11656 12652 11696
rect 12692 11656 12781 11696
rect 13027 11656 13036 11696
rect 13076 11656 13316 11696
rect 13385 11656 13483 11696
rect 13556 11656 13565 11696
rect 13699 11656 13708 11696
rect 13748 11656 14420 11696
rect 14467 11656 14476 11696
rect 14516 11656 14525 11696
rect 14822 11656 14831 11696
rect 14871 11656 14900 11696
rect 14952 11656 14961 11696
rect 15001 11656 15010 11696
rect 15082 11656 15091 11696
rect 15131 11656 15146 11696
rect 15226 11656 15235 11696
rect 15275 11656 15305 11696
rect 15348 11656 15357 11696
rect 15397 11656 15476 11696
rect 15532 11696 15572 11992
rect 15820 11992 16108 12032
rect 16148 11992 16157 12032
rect 16867 11992 16876 12032
rect 16916 11992 18356 12032
rect 18412 11992 19028 12032
rect 19555 11992 19564 12032
rect 19604 11992 21044 12032
rect 15820 11696 15860 11992
rect 16090 11908 16099 11948
rect 16139 11908 16588 11948
rect 16628 11908 16637 11948
rect 17155 11908 17164 11948
rect 17204 11908 17356 11948
rect 17396 11908 17405 11948
rect 18089 11908 18115 11948
rect 18155 11908 18220 11948
rect 18260 11908 18269 11948
rect 18316 11864 18356 11992
rect 18499 11908 18508 11948
rect 18548 11908 18595 11948
rect 18635 11908 18679 11948
rect 15916 11824 17588 11864
rect 18316 11824 18548 11864
rect 15916 11780 15956 11824
rect 15907 11740 15916 11780
rect 15956 11740 15965 11780
rect 16072 11740 16108 11780
rect 16148 11740 16159 11780
rect 16119 11696 16159 11740
rect 16328 11696 16368 11824
rect 16867 11740 16876 11780
rect 16916 11740 17012 11780
rect 16972 11696 17012 11740
rect 15532 11656 15575 11696
rect 15615 11656 15624 11696
rect 15706 11656 15715 11696
rect 15755 11656 15764 11696
rect 15811 11656 15820 11696
rect 15860 11656 15991 11696
rect 16101 11656 16110 11696
rect 16150 11656 16159 11696
rect 16204 11656 16217 11696
rect 16257 11656 16266 11696
rect 16328 11656 16357 11696
rect 16397 11656 16406 11696
rect 16474 11656 16483 11696
rect 16523 11656 16579 11696
rect 16651 11656 16660 11696
rect 16700 11656 16820 11696
rect 16954 11656 16963 11696
rect 17003 11656 17012 11696
rect 17059 11677 17068 11717
rect 17108 11677 17239 11717
rect 17548 11696 17588 11824
rect 18414 11696 18454 11705
rect 18508 11696 18548 11824
rect 18988 11780 19028 11992
rect 19075 11908 19084 11948
rect 19124 11908 20428 11948
rect 20468 11908 20477 11948
rect 20899 11908 20908 11948
rect 20948 11908 20957 11948
rect 20908 11864 20948 11908
rect 20236 11824 20716 11864
rect 20756 11824 20948 11864
rect 18988 11740 19219 11780
rect 19259 11740 19268 11780
rect 19747 11740 19756 11780
rect 19796 11740 19987 11780
rect 20027 11740 20036 11780
rect 20236 11738 20276 11824
rect 20521 11740 20530 11780
rect 20570 11740 20908 11780
rect 20948 11740 20957 11780
rect 18892 11696 18932 11705
rect 20170 11698 20179 11738
rect 20219 11698 20276 11738
rect 21004 11696 21044 11992
rect 21545 11908 21676 11948
rect 21716 11908 21725 11948
rect 21964 11864 22004 12432
rect 22522 12412 22531 12452
rect 22571 12412 22580 12452
rect 22627 12412 22636 12452
rect 22676 12412 22828 12452
rect 22907 12412 22916 12452
rect 23753 12412 23875 12452
rect 23924 12412 23933 12452
rect 22540 11948 22580 12412
rect 23491 12244 23500 12284
rect 23540 12244 23549 12284
rect 23500 12032 23540 12244
rect 24076 12116 24116 12580
rect 25420 12580 26284 12620
rect 26324 12580 26804 12620
rect 28387 12580 28396 12620
rect 28436 12580 28588 12620
rect 28628 12580 28637 12620
rect 29539 12580 29548 12620
rect 29588 12580 30124 12620
rect 30164 12580 30173 12620
rect 25420 12536 25460 12580
rect 26764 12536 26804 12580
rect 25402 12496 25411 12536
rect 25451 12496 25460 12536
rect 25699 12496 25708 12536
rect 25748 12496 25996 12536
rect 26036 12496 26045 12536
rect 26092 12496 26188 12536
rect 26228 12496 26237 12536
rect 26746 12496 26755 12536
rect 26795 12496 26804 12536
rect 27235 12496 27244 12536
rect 27284 12496 29644 12536
rect 29684 12496 29693 12536
rect 29740 12496 29817 12536
rect 29857 12496 29866 12536
rect 30019 12496 30028 12536
rect 30068 12496 30077 12536
rect 30124 12496 30220 12536
rect 30260 12496 31660 12536
rect 31700 12496 31709 12536
rect 26092 12452 26132 12496
rect 29548 12452 29588 12496
rect 29740 12452 29780 12496
rect 25623 12200 25663 12452
rect 25786 12412 25795 12452
rect 25835 12412 25844 12452
rect 25891 12412 25900 12452
rect 25940 12412 26132 12452
rect 26179 12412 26188 12452
rect 26228 12412 26380 12452
rect 26420 12412 26429 12452
rect 25804 12368 25844 12412
rect 28012 12368 28052 12432
rect 28169 12412 28300 12452
rect 28340 12412 28349 12452
rect 28675 12412 28684 12452
rect 28724 12412 29396 12452
rect 29539 12412 29548 12452
rect 29588 12412 29597 12452
rect 29731 12412 29740 12452
rect 29780 12412 29789 12452
rect 29356 12368 29396 12412
rect 30028 12368 30068 12496
rect 30124 12452 30164 12496
rect 30115 12412 30124 12452
rect 30164 12412 30173 12452
rect 30508 12412 31372 12452
rect 31412 12412 31421 12452
rect 30508 12368 30548 12412
rect 25804 12328 25996 12368
rect 26036 12328 26045 12368
rect 28012 12328 28876 12368
rect 28916 12328 28925 12368
rect 29251 12328 29260 12368
rect 29300 12328 29309 12368
rect 29356 12328 30068 12368
rect 30499 12328 30508 12368
rect 30548 12328 30557 12368
rect 30691 12328 30700 12368
rect 30740 12328 30892 12368
rect 30932 12328 30941 12368
rect 28553 12244 28588 12284
rect 28628 12244 28684 12284
rect 28724 12244 28733 12284
rect 29260 12200 29300 12328
rect 25623 12160 29300 12200
rect 29356 12160 30508 12200
rect 30548 12160 30557 12200
rect 24076 12076 25460 12116
rect 26425 12076 26434 12116
rect 26802 12076 26811 12116
rect 26947 12076 26956 12116
rect 26996 12076 28876 12116
rect 28916 12076 28925 12116
rect 23500 11992 25268 12032
rect 22540 11908 23491 11948
rect 23531 11908 23540 11948
rect 23945 11908 24076 11948
rect 24116 11908 24125 11948
rect 21955 11824 21964 11864
rect 22004 11824 22013 11864
rect 22828 11824 24172 11864
rect 24212 11824 24221 11864
rect 24316 11855 24460 11864
rect 21091 11740 21100 11780
rect 21140 11740 21244 11780
rect 21284 11740 21293 11780
rect 22828 11696 22868 11824
rect 24356 11824 24460 11855
rect 24500 11824 24509 11864
rect 24316 11806 24356 11815
rect 24407 11740 25132 11780
rect 25172 11740 25181 11780
rect 24407 11696 24447 11740
rect 25228 11696 25268 11992
rect 25420 11948 25460 12076
rect 29356 12032 29396 12160
rect 28588 11992 29396 12032
rect 28588 11948 28628 11992
rect 25420 11908 27148 11948
rect 27188 11908 27197 11948
rect 28579 11908 28588 11948
rect 28628 11908 28637 11948
rect 29059 11908 29068 11948
rect 29108 11908 29155 11948
rect 29195 11908 29239 11948
rect 29923 11908 29932 11948
rect 29972 11908 30316 11948
rect 30356 11908 30365 11948
rect 30569 11908 30700 11948
rect 30740 11908 30749 11948
rect 26572 11824 27532 11864
rect 27572 11824 28148 11864
rect 29251 11824 29260 11864
rect 29300 11824 29356 11864
rect 29396 11824 29431 11864
rect 29539 11824 29548 11864
rect 29588 11824 29597 11864
rect 30307 11824 30316 11864
rect 30356 11824 30548 11864
rect 30857 11824 30892 11864
rect 30932 11824 30988 11864
rect 31028 11824 31037 11864
rect 25507 11740 25516 11780
rect 25556 11740 25603 11780
rect 25643 11740 25687 11780
rect 26572 11696 26612 11824
rect 26659 11740 26668 11780
rect 26708 11740 27250 11780
rect 27290 11740 27299 11780
rect 28108 11696 28148 11824
rect 29548 11780 29588 11824
rect 28195 11740 28204 11780
rect 28244 11740 29012 11780
rect 29059 11740 29068 11780
rect 29108 11740 29396 11780
rect 29443 11740 29452 11780
rect 29492 11740 29501 11780
rect 29548 11740 29780 11780
rect 28972 11696 29012 11740
rect 29356 11696 29396 11740
rect 29452 11696 29492 11740
rect 29740 11696 29780 11740
rect 30220 11740 30412 11780
rect 30452 11740 30461 11780
rect 30220 11696 30260 11740
rect 30508 11696 30548 11824
rect 17539 11656 17548 11696
rect 17588 11656 17597 11696
rect 17722 11656 17731 11696
rect 17780 11656 17911 11696
rect 18283 11656 18412 11696
rect 18454 11656 18461 11696
rect 18508 11656 18796 11696
rect 18836 11656 18845 11696
rect 19171 11656 19180 11696
rect 19220 11656 19384 11696
rect 19424 11656 19433 11696
rect 20611 11656 20620 11696
rect 20660 11656 20791 11696
rect 21004 11656 21043 11696
rect 21083 11656 21092 11696
rect 21763 11656 21772 11696
rect 21812 11656 22636 11696
rect 22676 11656 22685 11696
rect 22819 11656 22828 11696
rect 22868 11656 22877 11696
rect 22985 11656 23116 11696
rect 23156 11656 23165 11696
rect 23299 11656 23308 11696
rect 23348 11656 23357 11696
rect 23482 11656 23491 11696
rect 23540 11656 23671 11696
rect 24250 11656 24259 11696
rect 24299 11656 24447 11696
rect 24643 11656 24652 11696
rect 24692 11656 25132 11696
rect 25172 11656 25181 11696
rect 25228 11656 25996 11696
rect 26036 11656 26045 11696
rect 26345 11656 26476 11696
rect 26516 11656 26525 11696
rect 26572 11656 26860 11696
rect 26900 11656 26909 11696
rect 27331 11656 27340 11696
rect 27380 11656 27511 11696
rect 27833 11656 27916 11696
rect 27956 11656 27964 11696
rect 28004 11656 28013 11696
rect 28099 11656 28108 11696
rect 28148 11656 28157 11696
rect 28387 11656 28396 11696
rect 28436 11656 28588 11696
rect 28628 11656 28637 11696
rect 28771 11656 28780 11696
rect 28820 11656 28829 11696
rect 28963 11656 28972 11696
rect 29012 11656 29021 11696
rect 29068 11656 29141 11696
rect 29181 11656 29190 11696
rect 29347 11656 29356 11696
rect 29396 11656 29405 11696
rect 29452 11656 29548 11696
rect 29588 11656 29597 11696
rect 29731 11656 29740 11696
rect 29780 11656 29789 11696
rect 29923 11656 29932 11696
rect 29972 11656 29981 11696
rect 30211 11656 30220 11696
rect 30260 11656 30269 11696
rect 30403 11656 30412 11696
rect 30452 11656 30604 11696
rect 30644 11656 30708 11696
rect 30787 11656 30796 11696
rect 30836 11656 31756 11696
rect 31796 11656 31805 11696
rect 748 11276 788 11656
rect 1324 11612 1364 11656
rect 1516 11612 1556 11656
rect 1660 11612 1700 11656
rect 1804 11612 1844 11656
rect 3148 11612 3188 11656
rect 3916 11612 3956 11656
rect 1315 11572 1324 11612
rect 1364 11572 1373 11612
rect 1507 11572 1516 11612
rect 1556 11572 1565 11612
rect 1660 11572 1708 11612
rect 1748 11572 1757 11612
rect 1804 11572 2284 11612
rect 2324 11572 2333 11612
rect 2755 11572 2764 11612
rect 2804 11572 2813 11612
rect 3148 11572 3956 11612
rect 4396 11612 4436 11656
rect 7756 11612 7796 11656
rect 9292 11612 9332 11656
rect 9868 11612 9908 11656
rect 10252 11612 10292 11656
rect 11020 11612 11060 11656
rect 12076 11612 12116 11656
rect 4396 11572 4892 11612
rect 4937 11572 5068 11612
rect 5108 11572 5117 11612
rect 5417 11572 5452 11612
rect 5492 11572 5548 11612
rect 5588 11572 5597 11612
rect 5649 11572 5658 11612
rect 5698 11572 5932 11612
rect 5972 11572 5981 11612
rect 6403 11572 6412 11612
rect 6452 11572 6548 11612
rect 6609 11572 6618 11612
rect 6658 11572 7660 11612
rect 7700 11572 7709 11612
rect 7756 11572 8716 11612
rect 8756 11572 9196 11612
rect 9236 11572 9245 11612
rect 9292 11572 9812 11612
rect 9868 11572 10292 11612
rect 10339 11572 10348 11612
rect 10388 11572 10636 11612
rect 10676 11572 11060 11612
rect 11768 11572 11777 11612
rect 11817 11572 11884 11612
rect 11924 11572 11948 11612
rect 12067 11572 12076 11612
rect 12116 11572 12163 11612
rect 2764 11528 2804 11572
rect 4852 11528 4892 11572
rect 6508 11528 6548 11572
rect 9772 11528 9812 11572
rect 905 11488 1036 11528
rect 1076 11488 1085 11528
rect 1219 11488 1228 11528
rect 1268 11488 2563 11528
rect 2603 11488 2804 11528
rect 2851 11488 2860 11528
rect 2900 11488 2909 11528
rect 3034 11488 3043 11528
rect 3083 11488 3532 11528
rect 3572 11488 3581 11528
rect 4003 11488 4012 11528
rect 4052 11488 4204 11528
rect 4244 11519 4375 11528
rect 4244 11488 4291 11519
rect 2860 11444 2900 11488
rect 2860 11404 2956 11444
rect 2996 11404 3005 11444
rect 3052 11360 3092 11488
rect 4282 11479 4291 11488
rect 4331 11488 4375 11519
rect 4852 11488 4876 11528
rect 4916 11488 4925 11528
rect 5818 11488 5827 11528
rect 5867 11488 6220 11528
rect 6260 11488 6269 11528
rect 6508 11488 7555 11528
rect 7595 11488 7948 11528
rect 7988 11488 7997 11528
rect 8131 11488 8140 11528
rect 8180 11488 8467 11528
rect 8507 11488 8516 11528
rect 8947 11488 8956 11528
rect 8996 11488 9100 11528
rect 9140 11488 9149 11528
rect 9772 11488 10156 11528
rect 10196 11488 10732 11528
rect 10772 11488 10924 11528
rect 10964 11488 10973 11528
rect 11369 11488 11500 11528
rect 11540 11488 11549 11528
rect 11971 11488 11980 11528
rect 12020 11488 12268 11528
rect 12308 11488 12317 11528
rect 4331 11479 4340 11488
rect 4282 11478 4340 11479
rect 12268 11444 12308 11488
rect 12268 11404 13036 11444
rect 13076 11404 13085 11444
rect 13276 11360 13316 11656
rect 14380 11612 14420 11656
rect 13411 11572 13420 11612
rect 13460 11572 13795 11612
rect 13835 11572 13844 11612
rect 14083 11572 14092 11612
rect 14132 11572 14271 11612
rect 14311 11572 14320 11612
rect 14362 11572 14371 11612
rect 14411 11572 14420 11612
rect 14572 11612 14612 11656
rect 14860 11612 14900 11656
rect 15265 11612 15305 11656
rect 15724 11612 15764 11656
rect 16204 11612 16244 11656
rect 16492 11612 16532 11656
rect 14572 11572 14804 11612
rect 14860 11572 15148 11612
rect 15188 11572 15197 11612
rect 15265 11572 15436 11612
rect 15476 11572 15485 11612
rect 15724 11572 16012 11612
rect 16052 11572 16061 11612
rect 16179 11572 16204 11612
rect 16244 11572 16253 11612
rect 16483 11572 16492 11612
rect 16532 11572 16541 11612
rect 14092 11528 14132 11572
rect 13507 11488 13516 11528
rect 13556 11488 14132 11528
rect 14764 11528 14804 11572
rect 16780 11528 16820 11656
rect 18414 11647 18454 11656
rect 18892 11612 18932 11656
rect 23308 11612 23348 11656
rect 17635 11572 17644 11612
rect 17684 11572 18110 11612
rect 18150 11572 18159 11612
rect 18499 11572 18508 11612
rect 18548 11572 18590 11612
rect 18630 11572 18679 11612
rect 18892 11572 22492 11612
rect 22532 11572 22541 11612
rect 23273 11572 23404 11612
rect 23444 11572 25900 11612
rect 25940 11572 25949 11612
rect 28780 11528 28820 11656
rect 29068 11612 29108 11656
rect 29932 11612 29972 11656
rect 28867 11572 28876 11612
rect 28916 11572 29836 11612
rect 29876 11572 29885 11612
rect 29932 11572 31468 11612
rect 31508 11572 31517 11612
rect 14764 11488 16588 11528
rect 16628 11488 16637 11528
rect 16771 11488 16780 11528
rect 16820 11519 16951 11528
rect 16820 11488 16867 11519
rect 16858 11479 16867 11488
rect 16907 11488 16951 11519
rect 18307 11488 18316 11528
rect 18356 11488 18700 11528
rect 18740 11488 18749 11528
rect 24931 11488 24940 11528
rect 24980 11488 24989 11528
rect 26249 11488 26371 11528
rect 26420 11488 26429 11528
rect 27427 11488 27436 11528
rect 27476 11488 27811 11528
rect 27851 11488 27860 11528
rect 28780 11488 29932 11528
rect 29972 11488 29981 11528
rect 16907 11479 16916 11488
rect 16858 11478 16916 11479
rect 24940 11444 24980 11488
rect 16972 11404 21716 11444
rect 24259 11404 24268 11444
rect 24308 11404 24980 11444
rect 25027 11404 25036 11444
rect 25076 11404 28916 11444
rect 16972 11360 17012 11404
rect 21676 11360 21716 11404
rect 1699 11320 1708 11360
rect 1748 11320 3092 11360
rect 4343 11320 4352 11360
rect 4720 11320 4729 11360
rect 6403 11320 6412 11360
rect 6452 11320 10100 11360
rect 12117 11320 12126 11360
rect 12494 11320 12503 11360
rect 12931 11320 12940 11360
rect 12980 11320 17012 11360
rect 19891 11320 19900 11360
rect 20268 11320 20277 11360
rect 21667 11320 21676 11360
rect 21716 11320 25516 11360
rect 25556 11320 25565 11360
rect 27665 11320 27674 11360
rect 28042 11320 28051 11360
rect 10060 11276 10100 11320
rect 588 11236 652 11276
rect 692 11236 2188 11276
rect 2228 11236 3764 11276
rect 3724 11234 3764 11236
rect 5164 11236 9606 11276
rect 9955 11236 9964 11276
rect 10004 11236 10013 11276
rect 10060 11236 19372 11276
rect 19412 11236 19421 11276
rect 22924 11236 25036 11276
rect 25076 11236 25085 11276
rect 3724 11194 3811 11234
rect 3851 11194 3860 11234
rect 5164 11192 5204 11236
rect 9566 11192 9606 11236
rect 9964 11192 10004 11236
rect 22924 11192 22964 11236
rect 1795 11152 1804 11192
rect 1844 11152 2284 11192
rect 2324 11152 2333 11192
rect 2755 11152 2764 11192
rect 2804 11152 2813 11192
rect 5146 11152 5155 11192
rect 5195 11152 5204 11192
rect 5801 11152 5923 11192
rect 5972 11152 5981 11192
rect 6604 11152 7028 11192
rect 7529 11152 7660 11192
rect 7700 11152 7709 11192
rect 8419 11152 8428 11192
rect 8468 11152 8812 11192
rect 8852 11152 8861 11192
rect 9466 11152 9475 11192
rect 9515 11152 9524 11192
rect 9566 11152 10051 11192
rect 10091 11152 10100 11192
rect 10243 11152 10252 11192
rect 10292 11152 10732 11192
rect 10772 11152 10781 11192
rect 10915 11152 10924 11192
rect 10964 11152 11308 11192
rect 11348 11152 11357 11192
rect 11753 11152 11884 11192
rect 11924 11152 11933 11192
rect 13193 11152 13324 11192
rect 13364 11152 13373 11192
rect 13594 11152 13603 11192
rect 13643 11152 13804 11192
rect 13844 11152 13853 11192
rect 14467 11152 14476 11192
rect 14516 11152 14860 11192
rect 14900 11152 14909 11192
rect 15139 11152 15148 11192
rect 15188 11152 15820 11192
rect 15860 11152 15869 11192
rect 16003 11152 16012 11192
rect 16052 11152 17740 11192
rect 17780 11152 17789 11192
rect 18281 11152 18403 11192
rect 18452 11152 18461 11192
rect 18691 11152 18700 11192
rect 18740 11152 18796 11192
rect 18836 11152 18871 11192
rect 20611 11152 20620 11192
rect 20660 11152 21091 11192
rect 21131 11152 21140 11192
rect 22570 11152 22579 11192
rect 22619 11152 22964 11192
rect 23395 11152 23404 11192
rect 23444 11152 24364 11192
rect 24404 11152 24413 11192
rect 24460 11152 25411 11192
rect 25451 11152 25460 11192
rect 26537 11152 26668 11192
rect 26708 11152 26717 11192
rect 27130 11152 27139 11192
rect 27179 11152 27340 11192
rect 27380 11152 27389 11192
rect 2764 11108 2804 11152
rect 931 11068 940 11108
rect 980 11068 1556 11108
rect 2764 11068 2900 11108
rect 2947 11068 2956 11108
rect 2996 11068 3284 11108
rect 1516 11024 1556 11068
rect 2860 11024 2900 11068
rect 3244 11024 3284 11068
rect 4977 11068 5164 11108
rect 5204 11068 5213 11108
rect 4977 11024 5017 11068
rect 6604 11024 6644 11152
rect 6988 11108 7028 11152
rect 9484 11108 9524 11152
rect 6691 11068 6700 11108
rect 6740 11068 6836 11108
rect 6988 11068 8044 11108
rect 8084 11068 8093 11108
rect 9484 11068 9868 11108
rect 9908 11068 9917 11108
rect 9964 11068 10156 11108
rect 10196 11068 10580 11108
rect 11472 11068 11500 11108
rect 11540 11068 11828 11108
rect 6796 11024 6836 11068
rect 7756 11024 7796 11068
rect 9964 11024 10004 11068
rect 10540 11024 10580 11068
rect 11548 11024 11588 11068
rect 11788 11024 11828 11068
rect 12840 11068 13612 11108
rect 13652 11068 13661 11108
rect 13891 11068 13900 11108
rect 13940 11068 13949 11108
rect 14266 11068 14275 11108
rect 14315 11068 15340 11108
rect 15380 11068 15389 11108
rect 15619 11068 15628 11108
rect 15668 11068 15956 11108
rect 835 10984 844 11024
rect 884 10984 893 11024
rect 1027 10984 1036 11024
rect 1076 10984 1228 11024
rect 1268 10984 1277 11024
rect 1402 10984 1411 11024
rect 1451 10984 1460 11024
rect 1507 10984 1516 11024
rect 1556 10984 1844 11024
rect 2467 10984 2476 11024
rect 2516 10984 2525 11024
rect 2602 10984 2611 11024
rect 2651 10984 2668 11024
rect 2708 10984 2791 11024
rect 2860 10984 3139 11024
rect 3179 10984 3188 11024
rect 3235 10984 3244 11024
rect 3284 10984 3841 11024
rect 3881 10984 3890 11024
rect 4073 10984 4147 11024
rect 4187 10984 4204 11024
rect 4244 10984 4253 11024
rect 4834 10984 4843 11024
rect 4883 10984 5017 11024
rect 5059 10984 5068 11024
rect 5108 10984 5239 11024
rect 5539 10984 5548 11024
rect 5588 10984 5591 11024
rect 5631 10984 5719 11024
rect 5827 10984 5836 11024
rect 5876 10984 6644 11024
rect 6691 10984 6700 11024
rect 6740 10984 6749 11024
rect 6796 10984 6883 11024
rect 6923 10984 6932 11024
rect 6988 10984 7036 11024
rect 7076 10984 7085 11024
rect 7171 10984 7180 11024
rect 7241 10984 7351 11024
rect 7459 10984 7468 11024
rect 7533 10984 7639 11024
rect 7747 10984 7756 11024
rect 7796 10984 7805 11024
rect 7939 10984 7948 11024
rect 8013 10984 8119 11024
rect 8393 10984 8524 11024
rect 8564 10984 8573 11024
rect 8752 10984 8761 11024
rect 8801 10984 8908 11024
rect 8948 10984 8957 11024
rect 9571 10984 9580 11024
rect 9620 10984 9751 11024
rect 9946 10984 9955 11024
rect 9995 10984 10004 11024
rect 10257 10984 10266 11024
rect 10306 10984 10444 11024
rect 10484 10984 10493 11024
rect 10540 10984 10583 11024
rect 10623 10984 10632 11024
rect 11203 10984 11212 11024
rect 11252 10984 11404 11024
rect 11444 10984 11453 11024
rect 11530 11015 11588 11024
rect 844 10940 884 10984
rect 844 10900 940 10940
rect 980 10900 989 10940
rect 1420 10436 1460 10984
rect 931 10396 940 10436
rect 980 10396 989 10436
rect 1420 10396 1660 10436
rect 1700 10396 1709 10436
rect 940 10352 980 10396
rect 652 10312 980 10352
rect 652 10184 692 10312
rect 1804 10268 1844 10984
rect 2476 10940 2516 10984
rect 3148 10940 3188 10984
rect 6700 10940 6740 10984
rect 6988 10940 7028 10984
rect 10444 10940 10484 10984
rect 11530 10975 11539 11015
rect 11579 10975 11588 11015
rect 11632 10984 11641 11024
rect 11681 10984 11732 11024
rect 11779 10984 11788 11024
rect 11828 10984 11837 11024
rect 11971 10984 11980 11024
rect 12020 10984 12151 11024
rect 12202 10984 12211 11024
rect 12251 10984 12748 11024
rect 12788 10984 12797 11024
rect 11530 10974 11588 10975
rect 2476 10900 2572 10940
rect 2612 10900 2621 10940
rect 3148 10900 4012 10940
rect 4052 10900 4061 10940
rect 4841 10900 4963 10940
rect 5012 10900 5021 10940
rect 5609 10900 5731 10940
rect 5780 10900 6028 10940
rect 6068 10900 6077 10940
rect 6700 10900 6988 10940
rect 7028 10900 7037 10940
rect 7241 10900 7372 10940
rect 7412 10900 7421 10940
rect 7651 10900 7660 10940
rect 7700 10900 7875 10940
rect 7915 10900 7924 10940
rect 8512 10900 8620 10940
rect 8683 10900 8692 10940
rect 9772 10900 10484 10940
rect 11692 10940 11732 10984
rect 11692 10900 12652 10940
rect 12692 10900 12701 10940
rect 9772 10856 9812 10900
rect 12840 10856 12880 11068
rect 13036 11024 13076 11068
rect 13900 11024 13940 11068
rect 14476 11024 14516 11068
rect 14860 11024 14900 11068
rect 15916 11024 15956 11068
rect 16780 11024 16820 11152
rect 17548 11068 17836 11108
rect 17876 11068 17885 11108
rect 18019 11068 18028 11108
rect 18068 11068 18508 11108
rect 18548 11068 19028 11108
rect 21571 11068 21580 11108
rect 21620 11068 22868 11108
rect 12922 10984 12931 11024
rect 12971 10984 12980 11024
rect 13027 10984 13036 11024
rect 13076 10984 13085 11024
rect 13385 10984 13505 11024
rect 13556 10984 13565 11024
rect 13699 10984 13708 11024
rect 13748 10984 13757 11024
rect 13804 11015 13851 11024
rect 3907 10816 3916 10856
rect 3956 10816 5068 10856
rect 5108 10816 5117 10856
rect 7267 10816 7276 10856
rect 7316 10816 8428 10856
rect 8468 10816 8477 10856
rect 9763 10816 9772 10856
rect 9812 10816 9821 10856
rect 10252 10816 12880 10856
rect 12940 10856 12980 10984
rect 13708 10940 13748 10984
rect 13844 10975 13851 11015
rect 13900 10984 13943 11024
rect 13983 10984 13992 11024
rect 14057 10984 14188 11024
rect 14228 10984 14237 11024
rect 14467 10984 14476 11024
rect 14516 10984 14525 11024
rect 14659 10984 14668 11024
rect 14708 10984 14717 11024
rect 14851 10984 14860 11024
rect 14900 10984 14909 11024
rect 14956 10984 15043 11024
rect 15083 10984 15235 11024
rect 15275 10984 15284 11024
rect 15412 10984 15532 11024
rect 15583 10984 15592 11024
rect 15715 10984 15724 11024
rect 15764 10984 15773 11024
rect 15907 10984 15916 11024
rect 15956 10984 15965 11024
rect 16762 10984 16771 11024
rect 16811 10984 16820 11024
rect 16867 10984 16876 11024
rect 16916 10984 17047 11024
rect 17321 10984 17452 11024
rect 17492 10984 17501 11024
rect 13804 10966 13851 10975
rect 13027 10900 13036 10940
rect 13076 10900 13748 10940
rect 13811 10940 13851 10966
rect 14668 10940 14708 10984
rect 14956 10940 14996 10984
rect 15724 10940 15764 10984
rect 13811 10900 13900 10940
rect 13940 10900 13949 10940
rect 14074 10900 14083 10940
rect 14123 10900 14132 10940
rect 14668 10900 14996 10940
rect 15052 10900 15764 10940
rect 15916 10940 15956 10984
rect 15916 10900 16972 10940
rect 17012 10900 17021 10940
rect 14092 10856 14132 10900
rect 12940 10816 14132 10856
rect 10252 10772 10292 10816
rect 3418 10732 3427 10772
rect 3467 10732 3532 10772
rect 3572 10732 3607 10772
rect 6874 10732 6883 10772
rect 6923 10732 7180 10772
rect 7220 10732 7229 10772
rect 10243 10732 10252 10772
rect 10292 10732 10301 10772
rect 12307 10732 12316 10772
rect 12356 10732 12556 10772
rect 12596 10732 12605 10772
rect 5548 10648 7564 10688
rect 7604 10648 7613 10688
rect 7660 10648 12748 10688
rect 12788 10648 12797 10688
rect 3103 10564 3112 10604
rect 3480 10564 3489 10604
rect 5548 10520 5588 10648
rect 7660 10604 7700 10648
rect 5635 10564 5644 10604
rect 5684 10564 7700 10604
rect 9571 10564 9580 10604
rect 9620 10564 9908 10604
rect 10877 10564 10886 10604
rect 11254 10564 11263 10604
rect 3820 10480 5588 10520
rect 8515 10480 8524 10520
rect 8564 10480 9524 10520
rect 3331 10396 3340 10436
rect 3380 10396 3389 10436
rect 3340 10352 3380 10396
rect 2266 10312 2275 10352
rect 2315 10312 2900 10352
rect 3340 10312 3764 10352
rect 2860 10268 2900 10312
rect 931 10228 940 10268
rect 980 10228 1708 10268
rect 1748 10228 1757 10268
rect 1804 10228 2420 10268
rect 2467 10228 2476 10268
rect 2516 10228 2659 10268
rect 2699 10228 2708 10268
rect 2860 10228 3619 10268
rect 3659 10228 3668 10268
rect 1036 10184 1076 10228
rect 2380 10184 2420 10228
rect 2860 10184 2900 10228
rect 3724 10184 3764 10312
rect 3820 10268 3860 10480
rect 9484 10436 9524 10480
rect 5242 10396 5251 10436
rect 5291 10396 5548 10436
rect 5588 10396 5597 10436
rect 6281 10396 6316 10436
rect 6356 10396 6412 10436
rect 6452 10396 7660 10436
rect 7700 10396 7709 10436
rect 8899 10396 8908 10436
rect 8948 10396 9052 10436
rect 9092 10396 9101 10436
rect 9475 10396 9484 10436
rect 9524 10396 9533 10436
rect 4012 10312 6220 10352
rect 6260 10312 6269 10352
rect 6892 10312 9428 10352
rect 3811 10228 3820 10268
rect 3860 10228 3869 10268
rect 4012 10184 4052 10312
rect 6892 10268 6932 10312
rect 4099 10228 4108 10268
rect 4148 10228 5876 10268
rect 5836 10184 5876 10228
rect 6076 10228 6932 10268
rect 7049 10228 7171 10268
rect 7220 10228 7229 10268
rect 8899 10228 8908 10268
rect 8948 10228 9332 10268
rect 643 10144 652 10184
rect 692 10144 701 10184
rect 835 10144 844 10184
rect 884 10144 893 10184
rect 1027 10144 1036 10184
rect 1076 10144 1085 10184
rect 1289 10144 1420 10184
rect 1460 10144 1469 10184
rect 1795 10144 1804 10184
rect 1844 10144 1987 10184
rect 2027 10144 2036 10184
rect 2083 10144 2092 10184
rect 2132 10144 2263 10184
rect 2380 10144 2524 10184
rect 2564 10144 2573 10184
rect 2668 10144 2764 10184
rect 2804 10144 2813 10184
rect 2860 10144 3043 10184
rect 3083 10144 3092 10184
rect 3139 10144 3148 10184
rect 3188 10144 3499 10184
rect 3572 10144 3581 10184
rect 3715 10144 3724 10184
rect 3764 10144 3773 10184
rect 4003 10144 4012 10184
rect 4052 10144 4061 10184
rect 4387 10144 4396 10184
rect 4436 10144 4445 10184
rect 4492 10144 4963 10184
rect 5003 10144 5012 10184
rect 5059 10144 5068 10184
rect 5108 10144 5239 10184
rect 5513 10144 5548 10184
rect 5588 10144 5644 10184
rect 5684 10144 5693 10184
rect 5827 10144 5836 10184
rect 5876 10144 5885 10184
rect 844 10100 884 10144
rect 643 10060 652 10100
rect 692 10060 884 10100
rect 1027 10060 1036 10100
rect 1076 10060 2476 10100
rect 2516 10060 2525 10100
rect 826 9976 835 10016
rect 875 9976 2092 10016
rect 2132 9976 2141 10016
rect 2668 9848 2708 10144
rect 2842 10060 2851 10100
rect 2900 10060 3031 10100
rect 3305 10060 3354 10100
rect 3394 10060 3436 10100
rect 3476 10060 3485 10100
rect 3043 9892 3052 9932
rect 3092 9892 3820 9932
rect 3860 9892 3869 9932
rect 4012 9848 4052 10144
rect 4396 9932 4436 10144
rect 4492 10016 4532 10144
rect 4972 10100 5012 10144
rect 4972 10060 5260 10100
rect 5300 10060 5309 10100
rect 6076 10016 6116 10228
rect 9292 10184 9332 10228
rect 9388 10184 9428 10312
rect 9868 10326 9908 10564
rect 13324 10436 13364 10816
rect 10025 10396 10147 10436
rect 10196 10396 10205 10436
rect 10252 10396 11404 10436
rect 11444 10396 11453 10436
rect 13306 10396 13315 10436
rect 13355 10396 13364 10436
rect 14860 10436 14900 10900
rect 15052 10856 15092 10900
rect 15034 10816 15043 10856
rect 15083 10816 15092 10856
rect 15532 10816 17108 10856
rect 15532 10772 15572 10816
rect 15523 10732 15532 10772
rect 15572 10732 15581 10772
rect 16963 10732 16972 10772
rect 17012 10732 17021 10772
rect 14860 10396 14908 10436
rect 14948 10396 14957 10436
rect 16627 10396 16636 10436
rect 16676 10396 16780 10436
rect 16820 10396 16829 10436
rect 9868 10286 9916 10326
rect 9956 10286 9965 10326
rect 10252 10184 10292 10396
rect 11497 10228 11506 10268
rect 11546 10228 11980 10268
rect 12059 10228 12068 10268
rect 12364 10228 12652 10268
rect 12692 10228 12940 10268
rect 12980 10228 12989 10268
rect 12364 10184 12404 10228
rect 16972 10184 17012 10732
rect 17068 10184 17108 10816
rect 17548 10436 17588 11068
rect 18988 11024 19028 11068
rect 22828 11024 22868 11068
rect 22924 11024 22964 11152
rect 23011 11068 23020 11108
rect 23060 11068 23356 11108
rect 23396 11068 23405 11108
rect 23884 11068 24259 11108
rect 24299 11068 24308 11108
rect 23884 11024 23924 11068
rect 24460 11024 24500 11152
rect 25420 11108 25460 11152
rect 24547 11068 24556 11108
rect 24596 11068 24605 11108
rect 24742 11068 25132 11108
rect 25172 11068 25224 11108
rect 25420 11068 25940 11108
rect 24556 11024 24596 11068
rect 24742 11024 24782 11068
rect 25132 11024 25172 11068
rect 25900 11024 25940 11068
rect 26284 11068 26380 11108
rect 26420 11068 26429 11108
rect 26284 11024 26324 11068
rect 17722 10984 17731 11024
rect 17771 10984 17780 11024
rect 17827 10984 17836 11024
rect 17876 10984 18302 11024
rect 18342 10984 18351 11024
rect 18604 11015 18644 11024
rect 17740 10940 17780 10984
rect 18970 10984 18979 11024
rect 19019 10984 19028 11024
rect 19555 10984 19564 11024
rect 19604 10984 19948 11024
rect 19988 10984 19997 11024
rect 20585 10984 20716 11024
rect 20756 10984 20765 11024
rect 21065 10984 21196 11024
rect 21236 10984 21245 11024
rect 21571 10984 21580 11024
rect 21620 10984 22060 11024
rect 22100 10984 22109 11024
rect 22330 11015 22388 11024
rect 17740 10900 18220 10940
rect 18260 10900 18269 10940
rect 18604 10856 18644 10975
rect 21580 10940 21620 10984
rect 22330 10975 22339 11015
rect 22379 10975 22388 11015
rect 22435 10984 22444 11024
rect 22484 10984 22540 11024
rect 22580 10984 22624 11024
rect 22819 10984 22828 11024
rect 22868 10984 22877 11024
rect 22924 10984 22947 11024
rect 22987 10984 22996 11024
rect 23059 10984 23068 11024
rect 23108 10984 23117 11024
rect 23194 11015 23212 11024
rect 22330 10974 22388 10975
rect 19459 10900 19468 10940
rect 19508 10900 21620 10940
rect 22348 10940 22388 10974
rect 23068 10940 23108 10984
rect 23194 10975 23203 11015
rect 23252 10984 23383 11024
rect 23587 10984 23596 11024
rect 23636 10984 23639 11024
rect 23679 10984 23767 11024
rect 23875 10984 23884 11024
rect 23924 10984 23933 11024
rect 24152 10984 24161 11024
rect 24201 10984 24282 11024
rect 24329 10984 24460 11024
rect 24500 10984 24509 11024
rect 24556 10984 24638 11024
rect 24678 10984 24687 11024
rect 24739 10984 24748 11024
rect 24788 10984 24797 11024
rect 23243 10975 23252 10984
rect 23194 10974 23252 10975
rect 22348 10900 22732 10940
rect 22772 10900 22781 10940
rect 23020 10900 23108 10940
rect 23770 10900 23779 10940
rect 23819 10900 23828 10940
rect 23971 10900 23980 10940
rect 24020 10900 24151 10940
rect 17993 10816 18124 10856
rect 18164 10816 18173 10856
rect 18604 10816 19024 10856
rect 19064 10816 19084 10856
rect 19124 10816 19133 10856
rect 20131 10816 20140 10856
rect 20180 10816 22051 10856
rect 22091 10816 22100 10856
rect 23020 10772 23060 10900
rect 19276 10732 19555 10772
rect 19595 10732 19604 10772
rect 20314 10732 20323 10772
rect 20363 10732 20372 10772
rect 22531 10732 22540 10772
rect 22580 10732 23060 10772
rect 19276 10688 19316 10732
rect 20332 10688 20372 10732
rect 18403 10648 18412 10688
rect 18452 10648 19124 10688
rect 19171 10648 19180 10688
rect 19220 10648 19316 10688
rect 19363 10648 19372 10688
rect 19412 10648 20372 10688
rect 19084 10604 19124 10648
rect 18651 10564 18660 10604
rect 19028 10564 19037 10604
rect 19084 10564 21580 10604
rect 21620 10564 21629 10604
rect 17731 10480 17740 10520
rect 17780 10480 20468 10520
rect 20428 10436 20468 10480
rect 20812 10480 23692 10520
rect 23732 10480 23741 10520
rect 17242 10396 17251 10436
rect 17291 10396 17588 10436
rect 17644 10396 20372 10436
rect 20428 10396 20668 10436
rect 20708 10396 20717 10436
rect 17644 10268 17684 10396
rect 20332 10352 20372 10396
rect 20812 10352 20852 10480
rect 23788 10436 23828 10900
rect 24242 10856 24282 10984
rect 24945 10982 24985 10991
rect 25090 10984 25099 11024
rect 25139 10984 25172 11024
rect 25315 10984 25324 11024
rect 25364 10984 25429 11024
rect 25481 10984 25612 11024
rect 25652 10984 25661 11024
rect 25891 10984 25900 11024
rect 25940 10984 25949 11024
rect 26266 10984 26275 11024
rect 26315 10984 26324 11024
rect 26371 10984 26380 11024
rect 26420 10984 26429 11024
rect 27427 10984 27436 11024
rect 27476 10984 27820 11024
rect 27860 10984 27869 11024
rect 28457 10984 28588 11024
rect 28628 10984 28637 11024
rect 24460 10966 24500 10975
rect 24941 10942 24945 10982
rect 24941 10933 24985 10942
rect 24233 10816 24364 10856
rect 24404 10816 24844 10856
rect 24884 10816 24893 10856
rect 24941 10772 24981 10933
rect 25210 10900 25219 10940
rect 25259 10900 25268 10940
rect 25228 10856 25268 10900
rect 25123 10816 25132 10856
rect 25172 10816 25268 10856
rect 25389 10856 25429 10984
rect 26380 10940 26420 10984
rect 26275 10900 26284 10940
rect 26324 10900 26420 10940
rect 27305 10900 27346 10940
rect 27386 10900 27436 10940
rect 27476 10900 27485 10940
rect 28876 10856 28916 11404
rect 30115 11320 30124 11360
rect 30164 11320 30260 11360
rect 28963 11236 28972 11276
rect 29012 11236 29684 11276
rect 29644 11192 29684 11236
rect 29321 11152 29356 11192
rect 29396 11152 29452 11192
rect 29492 11152 29501 11192
rect 29635 11152 29644 11192
rect 29684 11152 29693 11192
rect 29827 11152 29836 11192
rect 29876 11152 29885 11192
rect 29993 11152 30124 11192
rect 30164 11152 30173 11192
rect 29539 11068 29548 11108
rect 29588 11068 29597 11108
rect 29548 11024 29588 11068
rect 29836 11051 29876 11152
rect 29829 11043 29876 11051
rect 29129 10984 29260 11024
rect 29300 10984 29309 11024
rect 29434 10984 29443 11024
rect 29483 10984 29588 11024
rect 29635 10984 29644 11024
rect 29684 10984 29693 11024
rect 29820 11003 29829 11043
rect 29869 11003 29878 11043
rect 30220 11024 30260 11320
rect 30211 10984 30220 11024
rect 30260 10984 30269 11024
rect 29644 10940 29684 10984
rect 29932 10942 30028 10982
rect 30068 10942 30077 10982
rect 29932 10940 29972 10942
rect 29635 10900 29644 10940
rect 29684 10900 29731 10940
rect 29827 10900 29836 10940
rect 29876 10900 29972 10940
rect 25389 10816 26860 10856
rect 26900 10816 26909 10856
rect 28867 10816 28876 10856
rect 28916 10816 28925 10856
rect 30281 10816 30412 10856
rect 30452 10816 30461 10856
rect 30665 10816 30796 10856
rect 30836 10816 30845 10856
rect 25389 10772 25429 10816
rect 24941 10732 25429 10772
rect 25603 10732 25612 10772
rect 25652 10732 25661 10772
rect 26083 10732 26092 10772
rect 26132 10732 28195 10772
rect 28235 10732 28244 10772
rect 21571 10396 21580 10436
rect 21620 10396 22051 10436
rect 22091 10396 22100 10436
rect 23788 10396 23980 10436
rect 24020 10396 24029 10436
rect 24905 10396 25036 10436
rect 25076 10396 25085 10436
rect 19354 10312 19363 10352
rect 19403 10312 20236 10352
rect 20276 10312 20285 10352
rect 20332 10312 20852 10352
rect 20995 10312 21004 10352
rect 21044 10312 22732 10352
rect 22772 10312 22781 10352
rect 22828 10312 23155 10352
rect 23195 10312 23204 10352
rect 17155 10228 17164 10268
rect 17204 10228 17213 10268
rect 17417 10228 17548 10268
rect 17588 10228 17597 10268
rect 17644 10228 17763 10268
rect 17803 10228 17812 10268
rect 18019 10228 18028 10268
rect 18068 10228 18220 10268
rect 18260 10228 18269 10268
rect 19180 10228 19468 10268
rect 19508 10228 19517 10268
rect 19651 10228 19660 10268
rect 19700 10228 20010 10268
rect 21187 10228 21196 10268
rect 21236 10228 21245 10268
rect 22531 10228 22540 10268
rect 22580 10228 22732 10268
rect 22772 10228 22781 10268
rect 17164 10184 17204 10228
rect 19180 10184 19220 10228
rect 19970 10226 20010 10228
rect 19970 10186 19996 10226
rect 20036 10186 20045 10226
rect 21196 10184 21236 10228
rect 22828 10184 22868 10312
rect 25612 10268 25652 10732
rect 26425 10564 26434 10604
rect 26802 10564 26811 10604
rect 27689 10396 27811 10436
rect 27860 10396 27869 10436
rect 27523 10312 27532 10352
rect 27572 10312 28244 10352
rect 28361 10312 28492 10352
rect 28532 10312 28541 10352
rect 30281 10312 30412 10352
rect 30452 10312 30461 10352
rect 30665 10312 30796 10352
rect 30836 10312 30845 10352
rect 22954 10259 23644 10268
rect 22954 10219 22963 10259
rect 23003 10228 23644 10259
rect 23684 10228 23693 10268
rect 25129 10228 25138 10268
rect 25178 10228 25652 10268
rect 25842 10228 25900 10268
rect 25940 10228 26002 10268
rect 26042 10228 26764 10268
rect 26804 10228 26813 10268
rect 26860 10228 27052 10268
rect 27092 10228 27101 10268
rect 27148 10228 28052 10268
rect 23003 10219 23012 10228
rect 22954 10218 23012 10219
rect 24141 10184 24181 10193
rect 26860 10184 26900 10228
rect 27148 10184 27188 10228
rect 28012 10184 28052 10228
rect 28108 10184 28148 10193
rect 6316 10144 6460 10184
rect 6500 10144 6509 10184
rect 6595 10144 6604 10184
rect 6644 10144 7031 10184
rect 7071 10144 7080 10184
rect 7267 10144 7276 10184
rect 7316 10144 7447 10184
rect 7817 10144 7948 10184
rect 7988 10144 8140 10184
rect 8180 10144 8189 10184
rect 8297 10144 8428 10184
rect 8468 10144 8477 10184
rect 8681 10144 8812 10184
rect 8852 10144 8861 10184
rect 8995 10144 9004 10184
rect 9044 10144 9187 10184
rect 9227 10144 9236 10184
rect 9283 10144 9292 10184
rect 9332 10144 9341 10184
rect 9388 10144 9495 10184
rect 9535 10144 9716 10184
rect 9859 10144 9868 10184
rect 9908 10144 9955 10184
rect 9995 10144 10292 10184
rect 10615 10144 10624 10184
rect 10664 10144 11308 10184
rect 11348 10144 11357 10184
rect 11587 10144 11596 10184
rect 11636 10144 11884 10184
rect 11924 10144 11933 10184
rect 12355 10144 12364 10184
rect 12404 10144 12413 10184
rect 12617 10144 12652 10184
rect 12692 10144 12748 10184
rect 12788 10144 12797 10184
rect 13018 10144 13027 10184
rect 13067 10144 13076 10184
rect 13123 10144 13132 10184
rect 13172 10144 13420 10184
rect 13460 10144 13556 10184
rect 13687 10144 13696 10184
rect 13748 10144 13876 10184
rect 14345 10144 14476 10184
rect 14516 10144 14525 10184
rect 14755 10144 14764 10184
rect 14804 10144 14813 10184
rect 15017 10144 15148 10184
rect 15188 10144 15197 10184
rect 15523 10144 15532 10184
rect 15572 10144 15628 10184
rect 15668 10144 15703 10184
rect 15881 10144 16012 10184
rect 16052 10144 16061 10184
rect 16387 10144 16396 10184
rect 16436 10144 16445 10184
rect 16954 10144 16963 10184
rect 17003 10144 17012 10184
rect 17059 10144 17068 10184
rect 17108 10144 17117 10184
rect 17164 10144 17644 10184
rect 17684 10144 17693 10184
rect 17827 10144 17836 10184
rect 17901 10144 18007 10184
rect 18115 10144 18124 10184
rect 18164 10144 18173 10184
rect 18220 10144 18243 10184
rect 18283 10144 18292 10184
rect 18352 10144 18361 10184
rect 18401 10144 18508 10184
rect 18548 10144 18557 10184
rect 19171 10144 19180 10184
rect 19220 10144 19229 10184
rect 19354 10144 19363 10184
rect 19412 10144 19543 10184
rect 19625 10144 19756 10184
rect 19796 10144 19805 10184
rect 19852 10144 19875 10184
rect 19915 10144 19924 10184
rect 20995 10144 21004 10184
rect 21044 10144 21236 10184
rect 21283 10144 21292 10184
rect 21332 10144 21463 10184
rect 21545 10144 21580 10184
rect 21620 10144 21676 10184
rect 21716 10144 21725 10184
rect 21772 10144 22444 10184
rect 22484 10144 22493 10184
rect 22819 10144 22828 10184
rect 22868 10144 22877 10184
rect 23056 10144 23065 10184
rect 23105 10144 23116 10184
rect 23156 10144 23245 10184
rect 23308 10144 23356 10184
rect 23396 10144 23405 10184
rect 23491 10144 23500 10184
rect 23540 10144 23671 10184
rect 23779 10144 23788 10184
rect 23828 10144 23959 10184
rect 24010 10144 24076 10184
rect 24116 10144 24141 10184
rect 24235 10144 24244 10184
rect 24284 10144 24293 10184
rect 24355 10144 24364 10184
rect 24408 10144 24535 10184
rect 25219 10144 25228 10184
rect 25268 10144 25844 10184
rect 26083 10144 26092 10184
rect 26132 10144 26141 10184
rect 26851 10144 26860 10184
rect 26900 10144 26909 10184
rect 27139 10144 27148 10184
rect 27188 10144 27197 10184
rect 27322 10144 27331 10184
rect 27371 10144 27380 10184
rect 6316 10100 6356 10144
rect 6163 10060 6172 10100
rect 6212 10060 6356 10100
rect 8428 10100 8468 10144
rect 8428 10060 9388 10100
rect 9428 10060 9437 10100
rect 9676 10016 9716 10144
rect 13036 10100 13076 10144
rect 13516 10100 13556 10144
rect 14764 10100 14804 10144
rect 12960 10060 13036 10100
rect 13076 10060 13085 10100
rect 13516 10060 14324 10100
rect 14764 10060 15820 10100
rect 15860 10060 15869 10100
rect 14284 10016 14324 10060
rect 4483 9976 4492 10016
rect 4532 9976 4541 10016
rect 4963 9976 4972 10016
rect 5012 9976 6116 10016
rect 7354 9976 7363 10016
rect 7403 9976 7660 10016
rect 7700 9976 7709 10016
rect 7834 9976 7843 10016
rect 7883 9976 7892 10016
rect 8009 9976 8140 10016
rect 8180 9976 8189 10016
rect 9676 9976 10156 10016
rect 10196 9976 10780 10016
rect 10820 9976 10828 10016
rect 10868 9976 10980 10016
rect 13843 9976 13852 10016
rect 13892 9976 13996 10016
rect 14036 9976 14045 10016
rect 14266 9976 14275 10016
rect 14315 9976 14324 10016
rect 7852 9932 7892 9976
rect 16396 9932 16436 10144
rect 18124 10100 18164 10144
rect 18077 10060 18124 10100
rect 18164 10060 18173 10100
rect 18220 10016 18260 10144
rect 19852 10100 19892 10144
rect 21772 10100 21812 10144
rect 18307 10060 18316 10100
rect 18356 10060 19660 10100
rect 19700 10060 19709 10100
rect 19852 10060 20620 10100
rect 20660 10060 20669 10100
rect 21436 10060 21812 10100
rect 22234 10060 22243 10100
rect 22283 10060 22484 10100
rect 21436 10016 21476 10060
rect 22444 10016 22484 10060
rect 23308 10016 23348 10144
rect 24141 10135 24181 10144
rect 24242 10016 24282 10144
rect 25804 10016 25844 10144
rect 26092 10100 26132 10144
rect 27340 10100 27380 10144
rect 26092 10060 27380 10100
rect 27436 10144 27628 10184
rect 27668 10144 27677 10184
rect 28003 10144 28012 10184
rect 28052 10144 28061 10184
rect 28204 10184 28244 10312
rect 28204 10144 29356 10184
rect 29396 10144 29405 10184
rect 26668 10016 26708 10060
rect 27436 10016 27476 10144
rect 28108 10100 28148 10144
rect 27523 10060 27532 10100
rect 27572 10060 27806 10100
rect 27846 10060 27855 10100
rect 27916 10060 28148 10100
rect 17827 9976 17836 10016
rect 17876 9976 18260 10016
rect 18796 9976 21476 10016
rect 21545 9976 21676 10016
rect 21716 9976 22348 10016
rect 22388 9976 22397 10016
rect 22444 9976 22636 10016
rect 22676 9976 23348 10016
rect 23779 9976 23788 10016
rect 23828 9976 24282 10016
rect 25786 9976 25795 10016
rect 25835 9976 25844 10016
rect 26650 9976 26659 10016
rect 26699 9976 26708 10016
rect 26755 9976 26764 10016
rect 26804 9976 27476 10016
rect 4396 9892 4876 9932
rect 4916 9892 5492 9932
rect 7171 9892 7180 9932
rect 7220 9892 8524 9932
rect 8564 9892 8573 9932
rect 16265 9892 16396 9932
rect 16436 9892 17548 9932
rect 17588 9892 18412 9932
rect 18452 9892 18461 9932
rect 5452 9848 5492 9892
rect 940 9808 2708 9848
rect 2764 9808 4052 9848
rect 4343 9808 4352 9848
rect 4720 9808 4729 9848
rect 5443 9808 5452 9848
rect 5492 9808 5501 9848
rect 12117 9808 12126 9848
rect 12494 9808 12503 9848
rect 940 9680 980 9808
rect 2764 9764 2804 9808
rect 18796 9764 18836 9976
rect 27916 9932 27956 10060
rect 28003 9976 28012 10016
rect 28052 9976 28108 10016
rect 28148 9976 28183 10016
rect 28553 9976 28684 10016
rect 28724 9976 28733 10016
rect 26947 9892 26956 9932
rect 26996 9892 27956 9932
rect 19891 9808 19900 9848
rect 20268 9808 20277 9848
rect 27665 9808 27674 9848
rect 28042 9808 28051 9848
rect 1507 9724 1516 9764
rect 1556 9724 2476 9764
rect 2516 9724 2804 9764
rect 2860 9724 4108 9764
rect 4148 9724 4157 9764
rect 8803 9724 8812 9764
rect 8852 9724 9236 9764
rect 2860 9680 2900 9724
rect 9196 9680 9236 9724
rect 9772 9724 11252 9764
rect 9772 9680 9812 9724
rect 931 9640 940 9680
rect 980 9640 989 9680
rect 1673 9640 1804 9680
rect 1844 9640 1853 9680
rect 2284 9640 2900 9680
rect 3139 9640 3148 9680
rect 3188 9640 4204 9680
rect 4244 9640 4253 9680
rect 4762 9640 4771 9680
rect 4811 9640 5164 9680
rect 5204 9640 5213 9680
rect 6970 9640 6979 9680
rect 7019 9640 7276 9680
rect 7316 9640 7325 9680
rect 7651 9640 7660 9680
rect 7700 9640 8276 9680
rect 8489 9640 8524 9680
rect 8564 9640 8620 9680
rect 8660 9640 9004 9680
rect 9044 9640 9053 9680
rect 9187 9640 9196 9680
rect 9236 9640 9245 9680
rect 9754 9640 9763 9680
rect 9803 9640 9812 9680
rect 10313 9640 10444 9680
rect 10484 9640 10493 9680
rect 10906 9640 10915 9680
rect 10955 9640 10964 9680
rect 2284 9512 2324 9640
rect 2371 9556 2380 9596
rect 2420 9556 3284 9596
rect 3811 9556 3820 9596
rect 3860 9556 3869 9596
rect 4018 9556 4108 9596
rect 4148 9556 4157 9596
rect 4218 9556 6260 9596
rect 6307 9556 6316 9596
rect 6356 9556 6604 9596
rect 6644 9556 6653 9596
rect 7171 9556 7180 9596
rect 7220 9556 7316 9596
rect 3244 9539 3284 9556
rect 3244 9512 3369 9539
rect 3820 9512 3860 9556
rect 4018 9512 4058 9556
rect 4218 9512 4258 9556
rect 6220 9512 6260 9556
rect 7276 9512 7316 9556
rect 7468 9556 7948 9596
rect 7988 9556 7997 9596
rect 7468 9512 7508 9556
rect 8236 9512 8276 9640
rect 9196 9596 9236 9640
rect 10924 9596 10964 9640
rect 9196 9556 9620 9596
rect 9580 9512 9620 9556
rect 10636 9556 10964 9596
rect 10636 9512 10676 9556
rect 11212 9512 11252 9724
rect 13996 9724 14804 9764
rect 15907 9724 15916 9764
rect 15956 9724 18836 9764
rect 13996 9680 14036 9724
rect 12259 9640 12268 9680
rect 12308 9640 12692 9680
rect 13577 9640 13699 9680
rect 13748 9640 13757 9680
rect 13987 9640 13996 9680
rect 14036 9640 14045 9680
rect 14467 9640 14476 9680
rect 14516 9640 14668 9680
rect 14708 9640 14717 9680
rect 11971 9556 11980 9596
rect 12020 9556 12116 9596
rect 12355 9556 12364 9596
rect 12404 9556 12413 9596
rect 12076 9512 12116 9556
rect 12364 9512 12404 9556
rect 12652 9512 12692 9640
rect 13315 9556 13324 9596
rect 13364 9556 14188 9596
rect 14228 9556 14237 9596
rect 14668 9512 14708 9640
rect 14764 9596 14804 9724
rect 15017 9640 15148 9680
rect 15188 9640 15197 9680
rect 15619 9640 15628 9680
rect 15668 9640 15811 9680
rect 15851 9640 15860 9680
rect 17513 9640 17644 9680
rect 17684 9640 17693 9680
rect 17818 9640 17827 9680
rect 17867 9640 17876 9680
rect 18682 9640 18691 9680
rect 18731 9640 18740 9680
rect 17836 9596 17876 9640
rect 18700 9596 18740 9640
rect 14764 9556 15255 9596
rect 15295 9556 15304 9596
rect 15401 9556 15532 9596
rect 15572 9556 15581 9596
rect 17260 9556 17876 9596
rect 18028 9556 18740 9596
rect 17260 9512 17300 9556
rect 18028 9512 18068 9556
rect 18796 9512 18836 9724
rect 20236 9724 23116 9764
rect 23156 9724 23636 9764
rect 23683 9724 23692 9764
rect 23732 9724 24500 9764
rect 20236 9680 20276 9724
rect 23596 9680 23636 9724
rect 24460 9680 24500 9724
rect 20218 9640 20227 9680
rect 20267 9640 20276 9680
rect 20777 9640 20899 9680
rect 20948 9640 20957 9680
rect 21658 9640 21667 9680
rect 21707 9640 21716 9680
rect 23011 9640 23020 9680
rect 23060 9640 23069 9680
rect 23273 9640 23404 9680
rect 23444 9640 23453 9680
rect 23587 9640 23596 9680
rect 23636 9640 24020 9680
rect 24259 9640 24268 9680
rect 24308 9640 24317 9680
rect 24442 9640 24451 9680
rect 24491 9640 24500 9680
rect 25721 9640 25804 9680
rect 25883 9640 25901 9680
rect 25987 9640 25996 9680
rect 26036 9640 26516 9680
rect 27401 9640 27436 9680
rect 27476 9640 27532 9680
rect 27572 9640 27581 9680
rect 21676 9596 21716 9640
rect 23020 9596 23060 9640
rect 18892 9556 19372 9596
rect 19412 9556 19700 9596
rect 643 9472 652 9512
rect 692 9472 940 9512
rect 980 9472 989 9512
rect 1123 9472 1132 9512
rect 1172 9472 1181 9512
rect 1315 9472 1324 9512
rect 1364 9472 1516 9512
rect 1556 9472 1565 9512
rect 1699 9472 1708 9512
rect 1748 9472 2284 9512
rect 2324 9472 2333 9512
rect 2471 9472 2480 9512
rect 2520 9472 2563 9512
rect 2659 9472 2668 9512
rect 2708 9472 2839 9512
rect 2947 9472 2956 9512
rect 2996 9472 3005 9512
rect 3052 9472 3095 9512
rect 3135 9472 3144 9512
rect 3244 9499 3340 9512
rect 3329 9472 3340 9499
rect 3380 9472 3389 9512
rect 3497 9472 3532 9512
rect 3572 9472 3628 9512
rect 3668 9472 3677 9512
rect 3744 9472 3753 9512
rect 3793 9472 3860 9512
rect 3907 9472 3916 9512
rect 3956 9472 3965 9512
rect 4018 9472 4108 9512
rect 4148 9472 4157 9512
rect 4218 9472 4300 9512
rect 4340 9472 4349 9512
rect 4675 9472 4684 9512
rect 4724 9472 4855 9512
rect 5059 9472 5068 9512
rect 5108 9472 5111 9512
rect 5151 9472 5239 9512
rect 5347 9472 5356 9512
rect 5396 9472 5644 9512
rect 5684 9472 5693 9512
rect 5801 9472 5827 9512
rect 5867 9472 5932 9512
rect 5972 9472 5981 9512
rect 6089 9472 6220 9512
rect 6260 9472 6269 9512
rect 6403 9472 6412 9512
rect 6452 9472 6583 9512
rect 6691 9472 6700 9512
rect 6740 9472 6796 9512
rect 6836 9472 6871 9512
rect 6979 9472 6988 9512
rect 7028 9472 7159 9512
rect 7210 9472 7219 9512
rect 7259 9472 7316 9512
rect 7363 9472 7372 9512
rect 7412 9472 7468 9512
rect 7508 9472 7572 9512
rect 7651 9472 7660 9512
rect 7700 9472 8131 9512
rect 8171 9472 8180 9512
rect 8227 9472 8236 9512
rect 8276 9472 8407 9512
rect 8515 9472 8524 9512
rect 8564 9472 8716 9512
rect 8756 9472 8765 9512
rect 8969 9472 9100 9512
rect 9140 9472 9149 9512
rect 9300 9472 9388 9512
rect 9428 9472 9431 9512
rect 9471 9472 9480 9512
rect 9562 9472 9571 9512
rect 9611 9472 9620 9512
rect 9667 9472 9676 9512
rect 9716 9472 9725 9512
rect 10217 9472 10294 9512
rect 10334 9472 10348 9512
rect 10388 9472 10397 9512
rect 10531 9472 10540 9512
rect 10580 9472 10589 9512
rect 10636 9472 10659 9512
rect 10699 9472 10708 9512
rect 10768 9472 10777 9512
rect 10817 9472 10868 9512
rect 11177 9472 11212 9512
rect 11252 9472 11308 9512
rect 11348 9472 11357 9512
rect 11849 9472 11884 9512
rect 11924 9472 11980 9512
rect 12020 9472 12029 9512
rect 12076 9472 12119 9512
rect 12159 9472 12168 9512
rect 12364 9472 12407 9512
rect 12447 9472 12456 9512
rect 12643 9472 12652 9512
rect 12692 9472 12701 9512
rect 12748 9472 13036 9512
rect 13076 9472 13228 9512
rect 13268 9472 13277 9512
rect 13411 9472 13420 9512
rect 13460 9472 13591 9512
rect 13769 9472 13804 9512
rect 13844 9472 13900 9512
rect 13940 9472 13949 9512
rect 14179 9472 14188 9512
rect 14228 9472 14237 9512
rect 14441 9472 14572 9512
rect 14612 9472 14621 9512
rect 14668 9472 14947 9512
rect 14987 9472 14996 9512
rect 15043 9472 15052 9512
rect 15092 9472 15101 9512
rect 15427 9472 15436 9512
rect 15476 9472 15485 9512
rect 15619 9472 15628 9512
rect 15668 9472 15799 9512
rect 16099 9472 16108 9512
rect 16148 9472 16396 9512
rect 16436 9472 16445 9512
rect 17242 9472 17251 9512
rect 17291 9472 17300 9512
rect 17347 9472 17356 9512
rect 17396 9472 17405 9512
rect 18004 9472 18013 9512
rect 18053 9472 18068 9512
rect 18115 9472 18124 9512
rect 18164 9472 18295 9512
rect 18787 9472 18796 9512
rect 18836 9472 18845 9512
rect 1132 9428 1172 9472
rect 1708 9428 1748 9472
rect 2480 9428 2520 9472
rect 2956 9428 2996 9472
rect 1132 9388 1324 9428
rect 1364 9388 1748 9428
rect 2467 9388 2476 9428
rect 2516 9388 2525 9428
rect 2909 9388 2956 9428
rect 2996 9388 3005 9428
rect 3052 9344 3092 9472
rect 3916 9428 3956 9472
rect 4435 9430 4444 9470
rect 4484 9430 4493 9470
rect 3139 9388 3148 9428
rect 3188 9388 3221 9428
rect 3261 9388 3319 9428
rect 3427 9388 3436 9428
rect 3476 9388 3485 9428
rect 3916 9388 4244 9428
rect 2083 9304 2092 9344
rect 2132 9304 3092 9344
rect 2537 9220 2668 9260
rect 2708 9220 2717 9260
rect 3436 9176 3476 9388
rect 4204 9260 4244 9388
rect 4439 9344 4479 9430
rect 4570 9388 4579 9428
rect 4619 9388 4628 9428
rect 5129 9388 5251 9428
rect 5300 9388 5309 9428
rect 5443 9388 5452 9428
rect 5492 9388 7468 9428
rect 7508 9388 7517 9428
rect 4588 9344 4628 9388
rect 9676 9344 9716 9472
rect 9763 9388 9772 9428
rect 9812 9388 10099 9428
rect 10139 9388 10157 9428
rect 4291 9304 4300 9344
rect 4340 9304 4479 9344
rect 4579 9304 4588 9344
rect 4628 9304 4675 9344
rect 5443 9304 5452 9344
rect 5492 9304 5872 9344
rect 5912 9304 9100 9344
rect 9140 9304 9149 9344
rect 9379 9304 9388 9344
rect 9428 9304 9716 9344
rect 10540 9344 10580 9472
rect 10828 9428 10868 9472
rect 12748 9428 12788 9472
rect 14188 9428 14228 9472
rect 10723 9388 10732 9428
rect 10772 9388 10868 9428
rect 11113 9388 11122 9428
rect 11162 9388 12364 9428
rect 12404 9388 12413 9428
rect 12460 9388 12533 9428
rect 12573 9388 12582 9428
rect 12739 9388 12748 9428
rect 12788 9388 12797 9428
rect 13699 9388 13708 9428
rect 13748 9388 14228 9428
rect 10540 9304 11348 9344
rect 3619 9220 3628 9260
rect 3668 9220 3724 9260
rect 3764 9220 3799 9260
rect 4204 9220 6700 9260
rect 6740 9220 6749 9260
rect 11011 9220 11020 9260
rect 11060 9220 11069 9260
rect 11020 9176 11060 9220
rect 3436 9136 6124 9176
rect 6164 9136 6173 9176
rect 10732 9136 11060 9176
rect 3103 9052 3112 9092
rect 3480 9052 3489 9092
rect 7660 8968 9580 9008
rect 9620 8968 9629 9008
rect 0 8924 400 8944
rect 7660 8924 7700 8968
rect 0 8884 556 8924
rect 596 8884 605 8924
rect 1027 8884 1036 8924
rect 1076 8884 2572 8924
rect 2612 8884 2621 8924
rect 3322 8884 3331 8924
rect 3371 8884 4684 8924
rect 4724 8884 4733 8924
rect 5827 8884 5836 8924
rect 5876 8884 6364 8924
rect 6404 8884 6413 8924
rect 7651 8884 7660 8924
rect 7700 8884 7709 8924
rect 8419 8884 8428 8924
rect 8468 8884 10636 8924
rect 10676 8884 10685 8924
rect 0 8864 400 8884
rect 643 8800 652 8840
rect 692 8800 940 8840
rect 980 8800 989 8840
rect 2956 8800 3724 8840
rect 3764 8800 3773 8840
rect 5356 8800 6988 8840
rect 7028 8800 7037 8840
rect 9091 8800 9100 8840
rect 9140 8831 9284 8840
rect 9140 8800 9244 8831
rect 2956 8756 2996 8800
rect 1987 8716 1996 8756
rect 2036 8716 2045 8756
rect 2938 8716 2947 8756
rect 2987 8716 2996 8756
rect 3628 8716 4588 8756
rect 4628 8716 4637 8756
rect 4777 8716 4786 8756
rect 4826 8716 5260 8756
rect 5300 8716 5309 8756
rect 3628 8672 3668 8716
rect 5356 8672 5396 8800
rect 9244 8782 9284 8791
rect 6028 8716 6604 8756
rect 6644 8716 6653 8756
rect 9667 8716 9676 8756
rect 9716 8716 9964 8756
rect 10004 8716 10013 8756
rect 6028 8672 6068 8716
rect 2554 8632 2563 8672
rect 2603 8632 2708 8672
rect 2668 8588 2708 8632
rect 2860 8632 3052 8672
rect 3092 8632 3101 8672
rect 3209 8632 3329 8672
rect 3380 8632 3389 8672
rect 3497 8632 3628 8672
rect 3668 8632 3677 8672
rect 3785 8632 3820 8672
rect 3860 8632 3916 8672
rect 3956 8632 3965 8672
rect 4195 8632 4204 8672
rect 4244 8632 4628 8672
rect 4867 8632 4876 8672
rect 4916 8632 5396 8672
rect 5443 8632 5452 8672
rect 5492 8632 5623 8672
rect 5674 8632 5683 8672
rect 5723 8632 5780 8672
rect 6019 8632 6028 8672
rect 6068 8632 6077 8672
rect 6124 8632 6604 8672
rect 6644 8632 6932 8672
rect 6979 8632 6988 8672
rect 7028 8632 7180 8672
rect 7220 8632 7267 8672
rect 7307 8632 7316 8672
rect 7363 8639 7372 8679
rect 7416 8639 7543 8679
rect 10732 8672 10772 9136
rect 10877 9052 10886 9092
rect 11254 9052 11263 9092
rect 11308 8924 11348 9304
rect 12460 9176 12500 9388
rect 15052 9344 15092 9472
rect 15436 9428 15476 9472
rect 15139 9388 15148 9428
rect 15188 9388 15476 9428
rect 16009 9388 16018 9428
rect 16058 9388 16108 9428
rect 16148 9388 16189 9428
rect 16771 9388 16780 9428
rect 16820 9388 17260 9428
rect 17300 9388 17309 9428
rect 16780 9344 16820 9388
rect 13891 9304 13900 9344
rect 13940 9304 14572 9344
rect 14612 9304 14621 9344
rect 15052 9304 15820 9344
rect 15860 9304 16820 9344
rect 17356 9260 17396 9472
rect 18892 9428 18932 9556
rect 19660 9512 19700 9556
rect 21100 9556 21716 9596
rect 22589 9556 22636 9596
rect 22676 9556 22685 9596
rect 23020 9556 23788 9596
rect 23828 9556 23924 9596
rect 21100 9512 21140 9556
rect 22636 9512 22676 9556
rect 23884 9512 23924 9556
rect 23980 9512 24020 9640
rect 24268 9512 24308 9640
rect 24931 9556 24940 9596
rect 24980 9556 25214 9596
rect 25254 9556 25263 9596
rect 25306 9556 25315 9596
rect 25355 9556 25900 9596
rect 25940 9556 25949 9596
rect 26153 9556 26284 9596
rect 26324 9556 26333 9596
rect 26476 9512 26516 9640
rect 26947 9556 26956 9596
rect 26996 9556 27340 9596
rect 27380 9556 27389 9596
rect 19171 9472 19180 9512
rect 19220 9472 19372 9512
rect 19412 9472 19468 9512
rect 19508 9472 19517 9512
rect 19651 9472 19660 9512
rect 19700 9472 19709 9512
rect 19843 9472 19852 9512
rect 19892 9472 20515 9512
rect 20555 9472 20564 9512
rect 21076 9472 21085 9512
rect 21125 9472 21140 9512
rect 21187 9472 21196 9512
rect 21236 9472 21367 9512
rect 21955 9472 21964 9512
rect 22004 9472 22135 9512
rect 22618 9472 22627 9512
rect 22667 9472 22676 9512
rect 22723 9472 22732 9512
rect 22772 9472 23012 9512
rect 23081 9472 23203 9512
rect 23252 9472 23261 9512
rect 23369 9472 23500 9512
rect 23540 9472 23549 9512
rect 23866 9472 23875 9512
rect 23915 9472 23924 9512
rect 23971 9472 23980 9512
rect 24020 9472 24029 9512
rect 24268 9472 24604 9512
rect 24644 9472 24653 9512
rect 24739 9472 24748 9512
rect 24788 9472 24797 9512
rect 25289 9472 25420 9512
rect 25460 9472 25469 9512
rect 25516 9503 25708 9512
rect 22972 9428 23012 9472
rect 23500 9428 23540 9472
rect 17443 9388 17452 9428
rect 17492 9388 18932 9428
rect 20122 9388 20131 9428
rect 20171 9388 20332 9428
rect 20372 9388 20381 9428
rect 20620 9388 20707 9428
rect 20747 9388 20756 9428
rect 21859 9388 21868 9428
rect 21914 9388 22039 9428
rect 22889 9388 23020 9428
rect 23060 9388 23540 9428
rect 20620 9260 20660 9388
rect 17251 9220 17260 9260
rect 17300 9220 17396 9260
rect 19459 9220 19468 9260
rect 19508 9220 19996 9260
rect 20036 9220 20660 9260
rect 12460 9136 21676 9176
rect 21716 9136 21725 9176
rect 18651 9052 18660 9092
rect 19028 9052 19037 9092
rect 11875 8968 11884 9008
rect 11924 8968 13132 9008
rect 13172 8968 19180 9008
rect 19220 8968 19229 9008
rect 20620 8968 21868 9008
rect 21908 8968 21917 9008
rect 11107 8884 11116 8924
rect 11156 8884 11348 8924
rect 13507 8884 13516 8924
rect 13556 8884 13565 8924
rect 15340 8884 15916 8924
rect 15956 8884 15965 8924
rect 16483 8884 16492 8924
rect 16532 8884 17108 8924
rect 17242 8884 17251 8924
rect 17300 8884 17431 8924
rect 19747 8884 19756 8924
rect 19796 8884 20035 8924
rect 20075 8884 20084 8924
rect 13516 8840 13556 8884
rect 10819 8800 10828 8840
rect 10868 8831 12260 8840
rect 10868 8800 12220 8831
rect 12442 8800 12451 8840
rect 12491 8800 13036 8840
rect 13076 8800 13085 8840
rect 13132 8800 13556 8840
rect 14179 8800 14188 8840
rect 14228 8800 14237 8840
rect 12220 8782 12260 8791
rect 13132 8756 13172 8800
rect 14188 8756 14228 8800
rect 15340 8756 15380 8884
rect 17068 8840 17108 8884
rect 16858 8800 16867 8840
rect 16907 8800 16916 8840
rect 17068 8800 17300 8840
rect 19651 8800 19660 8840
rect 19700 8800 19747 8840
rect 19787 8800 19831 8840
rect 16876 8756 16916 8800
rect 11299 8716 11308 8756
rect 11348 8716 12020 8756
rect 12355 8716 12364 8756
rect 12404 8716 12652 8756
rect 12692 8716 13172 8756
rect 13219 8716 13228 8756
rect 13268 8716 14228 8756
rect 15005 8716 15052 8756
rect 15092 8716 15101 8756
rect 15148 8716 15380 8756
rect 15427 8716 15436 8756
rect 15476 8716 15532 8756
rect 15572 8716 15607 8756
rect 15811 8716 15820 8756
rect 15860 8716 16532 8756
rect 16771 8716 16780 8756
rect 16820 8716 16829 8756
rect 16876 8716 17108 8756
rect 7651 8632 7660 8672
rect 7700 8632 8131 8672
rect 8171 8632 8180 8672
rect 8227 8632 8236 8672
rect 8276 8632 8407 8672
rect 9274 8632 9283 8672
rect 9323 8632 9484 8672
rect 9524 8632 9533 8672
rect 9629 8632 9643 8672
rect 9683 8632 9692 8672
rect 9754 8632 9763 8672
rect 9803 8632 9812 8672
rect 9859 8632 9868 8672
rect 9908 8632 10039 8672
rect 10313 8632 10336 8672
rect 10376 8632 10444 8672
rect 10484 8632 10493 8672
rect 10732 8632 10819 8672
rect 10859 8632 10868 8672
rect 10924 8632 11788 8672
rect 11828 8632 11924 8672
rect 2860 8588 2900 8632
rect 3628 8623 3668 8632
rect 2668 8548 2900 8588
rect 0 8504 400 8524
rect 4588 8504 4628 8632
rect 5740 8588 5780 8632
rect 5059 8548 5068 8588
rect 5108 8548 5780 8588
rect 0 8464 460 8504
rect 500 8464 509 8504
rect 3523 8464 3532 8504
rect 3572 8464 4300 8504
rect 4340 8464 4349 8504
rect 4570 8464 4579 8504
rect 4619 8464 4876 8504
rect 4916 8464 4925 8504
rect 5177 8464 5260 8504
rect 5300 8464 5308 8504
rect 5348 8464 5357 8504
rect 0 8444 400 8464
rect 4343 8296 4352 8336
rect 4720 8296 4729 8336
rect 5740 8252 5780 8548
rect 6124 8504 6164 8632
rect 6892 8588 6932 8632
rect 9652 8588 9692 8632
rect 6892 8548 7220 8588
rect 8131 8548 8140 8588
rect 8180 8548 8439 8588
rect 8479 8548 8488 8588
rect 9353 8548 9388 8588
rect 9428 8548 9484 8588
rect 9524 8548 9533 8588
rect 9652 8548 9676 8588
rect 9716 8548 9725 8588
rect 7180 8504 7220 8548
rect 9772 8504 9812 8632
rect 10924 8588 10964 8632
rect 6115 8464 6124 8504
rect 6164 8464 6173 8504
rect 7162 8495 7220 8504
rect 7162 8455 7171 8495
rect 7211 8455 7220 8495
rect 9187 8464 9196 8504
rect 9236 8464 9812 8504
rect 10156 8548 10492 8588
rect 10532 8548 10964 8588
rect 11081 8548 11130 8588
rect 11170 8548 11212 8588
rect 11252 8548 11261 8588
rect 7162 8454 7220 8455
rect 3340 8212 3532 8252
rect 3572 8212 3581 8252
rect 5740 8212 6356 8252
rect 7459 8212 7468 8252
rect 7508 8212 8180 8252
rect 9859 8212 9868 8252
rect 9908 8212 10004 8252
rect 3340 8168 3380 8212
rect 6316 8168 6356 8212
rect 643 8128 652 8168
rect 692 8128 1468 8168
rect 1508 8128 3043 8168
rect 3083 8128 3092 8168
rect 3331 8128 3340 8168
rect 3380 8128 3389 8168
rect 3619 8128 3628 8168
rect 3668 8128 3811 8168
rect 3851 8128 3860 8168
rect 3907 8128 3916 8168
rect 3956 8128 4972 8168
rect 5012 8128 5021 8168
rect 5635 8128 5644 8168
rect 5684 8128 5827 8168
rect 5867 8128 5876 8168
rect 6298 8128 6307 8168
rect 6347 8128 6356 8168
rect 6595 8128 6604 8168
rect 6644 8128 7372 8168
rect 7412 8128 7421 8168
rect 7651 8128 7660 8168
rect 7700 8128 7709 8168
rect 0 8084 400 8104
rect 0 8044 844 8084
rect 884 8044 893 8084
rect 0 8024 400 8044
rect 2668 8000 2708 8128
rect 2755 8044 2764 8084
rect 2804 8044 3820 8084
rect 3860 8044 3869 8084
rect 4876 8044 7412 8084
rect 4876 8000 4916 8044
rect 7372 8000 7412 8044
rect 7660 8000 7700 8128
rect 8140 8000 8180 8212
rect 9964 8168 10004 8212
rect 8969 8128 9091 8168
rect 9140 8128 9149 8168
rect 9667 8128 9676 8168
rect 9716 8128 9859 8168
rect 9899 8128 9908 8168
rect 9955 8128 9964 8168
rect 10004 8128 10013 8168
rect 10156 8084 10196 8548
rect 10723 8464 10732 8504
rect 10772 8464 10915 8504
rect 10955 8464 10964 8504
rect 11561 8464 11683 8504
rect 11732 8464 11741 8504
rect 10732 8168 10772 8464
rect 11884 8420 11924 8632
rect 11980 8588 12020 8716
rect 15052 8672 15092 8716
rect 15148 8672 15188 8716
rect 16492 8672 16532 8716
rect 16780 8672 16820 8716
rect 17068 8672 17108 8716
rect 17260 8672 17300 8800
rect 19459 8716 19468 8756
rect 19508 8716 19555 8756
rect 19468 8672 19508 8716
rect 19756 8672 19796 8800
rect 20332 8672 20372 8681
rect 20620 8672 20660 8968
rect 20899 8884 20908 8924
rect 20948 8884 21772 8924
rect 21812 8884 21821 8924
rect 21955 8884 21964 8924
rect 22004 8884 22868 8924
rect 23011 8884 23020 8924
rect 23060 8884 23191 8924
rect 22828 8840 22868 8884
rect 22819 8800 22828 8840
rect 22868 8800 23404 8840
rect 23444 8800 24652 8840
rect 24692 8800 24701 8840
rect 22723 8716 22732 8756
rect 22772 8716 22781 8756
rect 24748 8672 24788 9472
rect 25556 9472 25708 9503
rect 25748 9472 25757 9512
rect 25886 9472 25996 9512
rect 26048 9472 26057 9512
rect 26135 9472 26171 9512
rect 26211 9472 26220 9512
rect 26374 9472 26383 9512
rect 26423 9472 26516 9512
rect 26563 9472 26572 9512
rect 26612 9472 26633 9512
rect 26746 9472 26755 9512
rect 26795 9472 26804 9512
rect 26921 9472 27052 9512
rect 27092 9472 27101 9512
rect 27280 9472 27289 9512
rect 27329 9472 27532 9512
rect 27572 9472 28684 9512
rect 28724 9472 28733 9512
rect 29225 9472 29347 9512
rect 29396 9472 29405 9512
rect 25516 9454 25556 9463
rect 26135 9344 26175 9472
rect 25315 9304 25324 9344
rect 25364 9304 26175 9344
rect 26593 9260 26633 9472
rect 26764 9428 26804 9472
rect 26764 9388 26956 9428
rect 26996 9388 27005 9428
rect 27052 9419 27244 9428
rect 27052 9388 27187 9419
rect 27052 9344 27092 9388
rect 27178 9379 27187 9388
rect 27227 9388 27244 9419
rect 27284 9388 27293 9428
rect 28483 9388 28492 9428
rect 28532 9388 28541 9428
rect 29722 9388 29731 9428
rect 29771 9388 29780 9428
rect 27227 9379 27236 9388
rect 27178 9378 27236 9379
rect 26746 9304 26755 9344
rect 26795 9304 27092 9344
rect 26593 9220 26860 9260
rect 26900 9220 26909 9260
rect 26425 9052 26434 9092
rect 26802 9052 26811 9092
rect 29740 8924 29780 9388
rect 28195 8884 28204 8924
rect 28244 8884 29780 8924
rect 25708 8800 28396 8840
rect 28436 8800 28445 8840
rect 25129 8716 25138 8756
rect 25178 8716 25612 8756
rect 25652 8716 25661 8756
rect 25708 8672 25748 8800
rect 25865 8716 25948 8756
rect 25988 8716 25996 8756
rect 26036 8716 27188 8756
rect 27148 8672 27188 8716
rect 27244 8672 27284 8681
rect 12137 8632 12259 8672
rect 12308 8632 12317 8672
rect 12364 8632 12835 8672
rect 12875 8632 12884 8672
rect 12940 8632 13564 8672
rect 13604 8632 13652 8672
rect 13699 8632 13708 8672
rect 13748 8632 13879 8672
rect 13996 8632 14188 8672
rect 14228 8632 14237 8672
rect 14371 8632 14380 8672
rect 14420 8632 14764 8672
rect 14804 8632 14813 8672
rect 15034 8632 15043 8672
rect 15083 8632 15092 8672
rect 15139 8632 15148 8672
rect 15188 8632 15197 8672
rect 15244 8632 15628 8672
rect 15668 8632 15677 8672
rect 15724 8632 15747 8672
rect 15787 8632 15796 8672
rect 15856 8632 15865 8672
rect 15905 8632 15956 8672
rect 16186 8632 16195 8672
rect 16235 8632 16291 8672
rect 16483 8632 16492 8672
rect 16532 8632 16541 8672
rect 16675 8632 16684 8672
rect 16724 8632 16733 8672
rect 16780 8632 16867 8672
rect 16907 8632 16916 8672
rect 17059 8632 17068 8672
rect 17108 8632 17117 8672
rect 17242 8632 17251 8672
rect 17291 8632 17300 8672
rect 17801 8632 17878 8672
rect 17918 8632 17932 8672
rect 17972 8632 17981 8672
rect 18499 8632 18508 8672
rect 18548 8632 18557 8672
rect 18641 8632 18650 8672
rect 18690 8632 19180 8672
rect 19220 8632 19229 8672
rect 19450 8632 19459 8672
rect 19499 8632 19508 8672
rect 19555 8632 19564 8672
rect 19604 8632 19613 8672
rect 19756 8632 20236 8672
rect 20276 8632 20285 8672
rect 20602 8632 20611 8672
rect 20651 8632 20660 8672
rect 21466 8632 21475 8672
rect 21515 8632 21676 8672
rect 21716 8632 22924 8672
rect 22964 8632 22973 8672
rect 24163 8632 24172 8672
rect 24212 8632 24221 8672
rect 24425 8632 24556 8672
rect 24596 8632 24605 8672
rect 24652 8632 24788 8672
rect 24835 8632 24844 8672
rect 24884 8632 25228 8672
rect 25268 8632 25420 8672
rect 25460 8632 25469 8672
rect 25708 8632 25804 8672
rect 25844 8632 25853 8672
rect 26755 8632 26764 8672
rect 26804 8632 27092 8672
rect 27139 8632 27148 8672
rect 27188 8632 27197 8672
rect 27401 8632 27436 8672
rect 27476 8632 27532 8672
rect 27572 8632 27581 8672
rect 28099 8632 28108 8672
rect 28148 8632 29068 8672
rect 29108 8632 29117 8672
rect 12364 8588 12404 8632
rect 11980 8548 12404 8588
rect 11971 8464 11980 8504
rect 12020 8464 12844 8504
rect 12884 8464 12893 8504
rect 12940 8420 12980 8632
rect 13612 8588 13652 8632
rect 13996 8588 14036 8632
rect 15244 8588 15284 8632
rect 15724 8588 15764 8632
rect 15916 8588 15956 8632
rect 16204 8588 16244 8632
rect 16684 8588 16724 8632
rect 18508 8588 18548 8632
rect 13123 8548 13132 8588
rect 13172 8548 13181 8588
rect 13612 8548 14036 8588
rect 15235 8548 15244 8588
rect 15284 8548 15293 8588
rect 15340 8548 15351 8588
rect 15391 8548 15400 8588
rect 15628 8548 15764 8588
rect 15907 8548 15916 8588
rect 15956 8548 15965 8588
rect 16195 8548 16204 8588
rect 16244 8548 16253 8588
rect 16608 8548 16684 8588
rect 16724 8548 17683 8588
rect 17723 8548 18220 8588
rect 18260 8548 18548 8588
rect 19564 8588 19604 8632
rect 20332 8588 20372 8632
rect 19564 8548 19756 8588
rect 19796 8548 19805 8588
rect 19939 8548 19948 8588
rect 19988 8548 20030 8588
rect 20070 8548 20119 8588
rect 20332 8548 20620 8588
rect 20660 8548 20669 8588
rect 20788 8548 20908 8588
rect 20959 8548 20968 8588
rect 21082 8548 21091 8588
rect 21140 8548 21271 8588
rect 11884 8380 12980 8420
rect 13132 8336 13172 8548
rect 15340 8504 15380 8548
rect 13987 8464 13996 8504
rect 14036 8464 15436 8504
rect 15476 8464 15540 8504
rect 15628 8420 15668 8548
rect 18665 8464 18796 8504
rect 18836 8464 18845 8504
rect 20698 8464 20707 8504
rect 20747 8464 22156 8504
rect 22196 8464 22205 8504
rect 15043 8380 15052 8420
rect 15092 8380 15668 8420
rect 24172 8420 24212 8632
rect 24652 8504 24692 8632
rect 27052 8588 27092 8632
rect 27244 8588 27284 8632
rect 26811 8548 26860 8588
rect 26900 8548 26942 8588
rect 26982 8548 26991 8588
rect 27034 8548 27043 8588
rect 27083 8548 27092 8588
rect 27139 8548 27148 8588
rect 27188 8548 27284 8588
rect 24643 8464 24652 8504
rect 24692 8464 24701 8504
rect 24922 8464 24931 8504
rect 24971 8464 24980 8504
rect 26083 8464 26092 8504
rect 26132 8464 26263 8504
rect 24940 8420 24980 8464
rect 24172 8380 24652 8420
rect 24692 8380 24980 8420
rect 12117 8296 12126 8336
rect 12494 8296 12503 8336
rect 13132 8296 19372 8336
rect 19412 8296 19421 8336
rect 19891 8296 19900 8336
rect 20268 8296 20277 8336
rect 27665 8296 27674 8336
rect 28042 8296 28051 8336
rect 14668 8212 16436 8252
rect 17539 8212 17548 8252
rect 17588 8212 18356 8252
rect 24835 8212 24844 8252
rect 24884 8212 25268 8252
rect 10723 8128 10732 8168
rect 10772 8128 10781 8168
rect 11273 8128 11404 8168
rect 11444 8128 11453 8168
rect 12643 8128 12652 8168
rect 12692 8128 13132 8168
rect 13172 8128 13181 8168
rect 8227 8044 8236 8084
rect 8276 8044 10196 8084
rect 11587 8044 11596 8084
rect 11636 8044 11980 8084
rect 12020 8044 12029 8084
rect 12175 8044 12184 8084
rect 12224 8044 12268 8084
rect 12308 8044 12355 8084
rect 13018 8044 13027 8084
rect 13067 8044 13324 8084
rect 13364 8044 13556 8084
rect 8620 8000 8660 8044
rect 9292 8000 9332 8044
rect 11692 8000 11732 8044
rect 13516 8000 13556 8044
rect 14270 8044 14516 8084
rect 14270 8000 14310 8044
rect 14476 8000 14516 8044
rect 14668 8000 14708 8212
rect 15811 8128 15820 8168
rect 15860 8128 15916 8168
rect 15956 8128 15991 8168
rect 16073 8128 16195 8168
rect 16244 8128 16253 8168
rect 16204 8084 16244 8128
rect 14755 8044 14764 8084
rect 14804 8044 15188 8084
rect 15148 8000 15188 8044
rect 15724 8044 16244 8084
rect 16396 8084 16436 8212
rect 17530 8128 17539 8168
rect 17579 8128 18028 8168
rect 18068 8128 18077 8168
rect 18202 8128 18211 8168
rect 18251 8128 18260 8168
rect 18220 8084 18260 8128
rect 16396 8044 16780 8084
rect 16820 8044 16829 8084
rect 17452 8044 18260 8084
rect 15724 8000 15764 8044
rect 16396 8000 16436 8044
rect 17452 8000 17492 8044
rect 18316 8000 18356 8212
rect 19747 8128 19756 8168
rect 19796 8128 20131 8168
rect 20171 8128 20180 8168
rect 20297 8128 20332 8168
rect 20372 8128 20428 8168
rect 20468 8128 20477 8168
rect 20969 8128 21100 8168
rect 21140 8128 21149 8168
rect 18787 8044 18796 8084
rect 18836 8044 20084 8084
rect 20044 8000 20084 8044
rect 20140 8044 20564 8084
rect 22025 8044 22147 8084
rect 22196 8044 22205 8084
rect 23945 8044 23980 8084
rect 24020 8075 24116 8084
rect 24020 8044 24067 8075
rect 259 7935 268 7975
rect 308 7935 317 7975
rect 931 7960 940 8000
rect 980 7991 1364 8000
rect 980 7960 1315 7991
rect 1306 7951 1315 7960
rect 1355 7951 1364 7991
rect 2659 7960 2668 8000
rect 2708 7960 2717 8000
rect 2842 7960 2851 8000
rect 2891 7960 2956 8000
rect 2996 7960 3148 8000
rect 3188 7960 3197 8000
rect 3907 7960 3916 8000
rect 3956 7960 4108 8000
rect 4148 7960 4157 8000
rect 4836 7960 4845 8000
rect 4885 7960 4916 8000
rect 4963 7960 4972 8000
rect 5033 7960 5143 8000
rect 5251 7960 5260 8000
rect 5325 7960 5431 8000
rect 5923 7960 5932 8000
rect 5972 7960 5981 8000
rect 6403 7960 6412 8000
rect 6452 7960 6604 8000
rect 6644 7960 6653 8000
rect 7116 7960 7180 8000
rect 7220 7960 7267 8000
rect 7307 7960 7316 8000
rect 7363 7960 7372 8000
rect 7412 7960 7543 8000
rect 7660 7960 8035 8000
rect 8075 7960 8084 8000
rect 8131 7960 8140 8000
rect 8180 7960 8428 8000
rect 8468 7960 8477 8000
rect 8611 7960 8620 8000
rect 8660 7960 8669 8000
rect 8803 7960 8812 8000
rect 8852 7960 8983 8000
rect 9283 7960 9292 8000
rect 9332 7960 9341 8000
rect 9449 7960 9580 8000
rect 9620 7960 9629 8000
rect 9754 7960 9763 8000
rect 9803 7960 9812 8000
rect 10065 7960 10074 8000
rect 10114 7960 10123 8000
rect 10243 7960 10252 8000
rect 10292 7960 10423 8000
rect 10505 7960 10636 8000
rect 10676 7960 10685 8000
rect 11369 7960 11404 8000
rect 11444 7960 11500 8000
rect 11540 7960 11549 8000
rect 11692 7960 11717 8000
rect 11757 7960 11766 8000
rect 11866 7960 11875 8000
rect 11915 7960 11924 8000
rect 12067 7960 12076 8000
rect 12116 7960 12695 8000
rect 12735 7960 12744 8000
rect 12876 7960 12931 8000
rect 12971 7960 13036 8000
rect 13076 7960 13111 8000
rect 13219 7960 13228 8000
rect 13268 7960 13276 8000
rect 13316 7960 13399 8000
rect 13516 7960 13577 8000
rect 13617 7960 13626 8000
rect 13699 7960 13708 8000
rect 13771 7960 14310 8000
rect 14467 7960 14476 8000
rect 14516 7960 14525 8000
rect 14602 7960 14611 8000
rect 14651 7960 14956 8000
rect 14996 7960 15005 8000
rect 15139 7960 15148 8000
rect 15188 7960 15319 8000
rect 15370 7960 15379 8000
rect 15419 7960 15428 8000
rect 15715 7960 15724 8000
rect 15764 7960 15773 8000
rect 16387 7960 16396 8000
rect 16436 7960 16445 8000
rect 16553 7960 16684 8000
rect 16724 7960 16733 8000
rect 17155 7960 17164 8000
rect 17204 7960 17207 8000
rect 17247 7960 17335 8000
rect 17443 7960 17452 8000
rect 17492 7960 17501 8000
rect 17635 7960 17644 8000
rect 17684 7960 17740 8000
rect 17780 7960 17815 8000
rect 18019 7960 18028 8000
rect 18068 7960 18220 8000
rect 18260 7960 18269 8000
rect 18316 7960 18364 8000
rect 18404 7960 18413 8000
rect 18499 7960 18508 8000
rect 18548 7960 18557 8000
rect 19258 7960 19267 8000
rect 19307 7960 19316 8000
rect 19363 7960 19372 8000
rect 19412 7960 19799 8000
rect 19839 7960 19848 8000
rect 20035 7960 20044 8000
rect 20084 7960 20093 8000
rect 1306 7950 1364 7951
rect 268 7832 308 7935
rect 5932 7916 5972 7960
rect 2851 7876 2860 7916
rect 2900 7876 4018 7916
rect 4058 7876 4067 7916
rect 4867 7876 4876 7916
rect 4916 7876 5164 7916
rect 5204 7876 5213 7916
rect 5932 7876 7220 7916
rect 7180 7832 7220 7876
rect 7276 7832 7316 7960
rect 8044 7916 8084 7960
rect 9772 7916 9812 7960
rect 8044 7876 8332 7916
rect 8372 7876 8381 7916
rect 9187 7876 9196 7916
rect 9236 7876 9812 7916
rect 10074 7916 10114 7960
rect 11884 7916 11924 7960
rect 15378 7916 15418 7960
rect 18220 7916 18260 7960
rect 18508 7916 18548 7960
rect 10074 7876 10156 7916
rect 10196 7876 11212 7916
rect 11252 7876 11261 7916
rect 11610 7876 11619 7916
rect 11659 7876 11788 7916
rect 11828 7876 11924 7916
rect 12713 7876 12835 7916
rect 12884 7876 12893 7916
rect 13289 7876 13420 7916
rect 13460 7876 13469 7916
rect 13516 7876 15820 7916
rect 15860 7876 15869 7916
rect 17338 7876 17347 7916
rect 17387 7876 17396 7916
rect 18220 7876 18548 7916
rect 19276 7916 19316 7960
rect 19276 7876 19939 7916
rect 19979 7876 19988 7916
rect 13516 7832 13556 7876
rect 17356 7832 17396 7876
rect 268 7792 500 7832
rect 1865 7792 1996 7832
rect 2036 7792 2045 7832
rect 5059 7792 5068 7832
rect 5108 7792 7124 7832
rect 7171 7792 7180 7832
rect 7220 7792 7229 7832
rect 7276 7792 8140 7832
rect 8180 7792 8189 7832
rect 9571 7792 9580 7832
rect 9620 7792 11500 7832
rect 11540 7792 11549 7832
rect 13507 7792 13516 7832
rect 13556 7792 13565 7832
rect 17356 7792 17740 7832
rect 17780 7792 17789 7832
rect 0 7664 400 7684
rect 460 7664 500 7792
rect 7084 7748 7124 7792
rect 5923 7708 5932 7748
rect 5972 7708 6124 7748
rect 6164 7708 6892 7748
rect 6932 7708 6941 7748
rect 7084 7708 8044 7748
rect 8084 7708 8093 7748
rect 8314 7708 8323 7748
rect 8363 7708 8372 7748
rect 8489 7708 8620 7748
rect 8660 7708 8669 7748
rect 9475 7708 9484 7748
rect 9524 7708 10060 7748
rect 10100 7708 10109 7748
rect 12163 7708 12172 7748
rect 12212 7708 12221 7748
rect 14537 7708 14659 7748
rect 14708 7708 14717 7748
rect 14825 7708 14956 7748
rect 14996 7708 15005 7748
rect 0 7624 500 7664
rect 8332 7664 8372 7708
rect 12172 7664 12212 7708
rect 8332 7624 9676 7664
rect 9716 7624 9725 7664
rect 11395 7624 11404 7664
rect 11444 7624 12212 7664
rect 0 7604 400 7624
rect 3103 7540 3112 7580
rect 3480 7540 3489 7580
rect 10877 7540 10886 7580
rect 11254 7540 11263 7580
rect 18651 7540 18660 7580
rect 19028 7540 19037 7580
rect 9379 7456 9388 7496
rect 9428 7456 9475 7496
rect 9388 7412 9428 7456
rect 19372 7412 19412 7876
rect 20140 7832 20180 8044
rect 20524 8000 20564 8044
rect 24058 8035 24067 8044
rect 24107 8035 24116 8075
rect 24163 8044 24172 8084
rect 24212 8044 24260 8084
rect 24355 8044 24364 8084
rect 24404 8044 24596 8084
rect 24643 8044 24652 8084
rect 24692 8044 24730 8084
rect 24058 8034 24116 8035
rect 24220 8000 24260 8044
rect 24556 8000 24596 8044
rect 24690 8002 24730 8044
rect 24940 8044 25132 8084
rect 25172 8044 25181 8084
rect 24940 8010 24980 8044
rect 24652 8000 24730 8002
rect 24844 8000 24980 8010
rect 25228 8008 25268 8212
rect 27977 8128 28108 8168
rect 28148 8128 28157 8168
rect 25786 8044 25795 8084
rect 25835 8044 26092 8084
rect 26132 8044 26141 8084
rect 25214 8000 25268 8008
rect 20297 7960 20428 8000
rect 20468 7960 20477 8000
rect 20524 7960 20659 8000
rect 20699 7960 21388 8000
rect 21428 7960 21437 8000
rect 21641 7960 21772 8000
rect 21812 7960 21821 8000
rect 22697 7960 22828 8000
rect 22868 7960 22877 8000
rect 23177 7960 23308 8000
rect 23348 7960 23357 8000
rect 23657 7960 23779 8000
rect 23828 7960 23837 8000
rect 23884 7991 23924 8000
rect 24162 7960 24171 8000
rect 24211 7960 24260 8000
rect 23884 7916 23924 7951
rect 24331 7949 24340 7989
rect 24380 7949 24404 7989
rect 24533 7960 24542 8000
rect 24582 7960 24596 8000
rect 24643 7960 24652 8000
rect 24692 7962 24730 8000
rect 24692 7960 24701 7962
rect 24835 7960 24844 8000
rect 24884 7970 24980 8000
rect 24884 7960 24893 7970
rect 25022 7960 25031 8000
rect 25071 7960 25080 8000
rect 25207 7960 25216 8000
rect 25256 7968 25268 8000
rect 25256 7960 25265 7968
rect 25315 7960 25324 8000
rect 25364 7960 25420 8000
rect 25460 7960 25495 8000
rect 25603 7960 25612 8000
rect 25652 7960 25661 8000
rect 26170 7960 26179 8000
rect 26228 7960 26359 8000
rect 20554 7907 20812 7916
rect 20554 7867 20563 7907
rect 20603 7876 20812 7907
rect 20852 7876 20861 7916
rect 23209 7876 23218 7916
rect 23258 7876 23348 7916
rect 23683 7876 23692 7916
rect 23732 7876 23924 7916
rect 24364 7916 24404 7949
rect 25036 7916 25076 7960
rect 24364 7876 24844 7916
rect 24884 7876 24893 7916
rect 25027 7876 25036 7916
rect 25076 7876 25118 7916
rect 20603 7867 20612 7876
rect 20554 7866 20612 7867
rect 19546 7792 19555 7832
rect 19595 7792 20180 7832
rect 20611 7708 20620 7748
rect 20660 7708 23116 7748
rect 23156 7708 23165 7748
rect 20419 7456 20428 7496
rect 20468 7456 21236 7496
rect 21196 7412 21236 7456
rect 163 7372 172 7412
rect 212 7372 500 7412
rect 5897 7372 6028 7412
rect 6068 7372 6077 7412
rect 6124 7372 7180 7412
rect 7220 7372 7229 7412
rect 8026 7372 8035 7412
rect 8075 7372 9196 7412
rect 9236 7372 9245 7412
rect 9379 7372 9388 7412
rect 9428 7372 9437 7412
rect 10121 7372 10252 7412
rect 10292 7372 10301 7412
rect 14467 7372 14476 7412
rect 14516 7372 17164 7412
rect 17204 7372 17213 7412
rect 18970 7372 18979 7412
rect 19019 7372 19276 7412
rect 19316 7372 19325 7412
rect 19372 7372 19660 7412
rect 19700 7372 19709 7412
rect 20681 7372 20812 7412
rect 20852 7372 20861 7412
rect 21178 7372 21187 7412
rect 21227 7372 21236 7412
rect 23308 7412 23348 7876
rect 24364 7832 24404 7876
rect 25612 7832 25652 7960
rect 23395 7792 23404 7832
rect 23444 7792 24404 7832
rect 24547 7792 24556 7832
rect 24596 7792 24940 7832
rect 24980 7792 24989 7832
rect 25210 7792 25219 7832
rect 25259 7792 25652 7832
rect 27436 7832 27476 7896
rect 27436 7792 28300 7832
rect 28340 7792 28349 7832
rect 23770 7708 23779 7748
rect 23819 7708 24364 7748
rect 24404 7708 24413 7748
rect 24547 7708 24556 7748
rect 24596 7708 25420 7748
rect 25460 7708 25469 7748
rect 26755 7708 26764 7748
rect 26804 7708 27724 7748
rect 27764 7708 27773 7748
rect 26425 7540 26434 7580
rect 26802 7540 26811 7580
rect 23308 7372 23356 7412
rect 23396 7372 23405 7412
rect 0 7244 400 7264
rect 460 7244 500 7372
rect 6124 7328 6164 7372
rect 2860 7288 3628 7328
rect 3668 7288 3677 7328
rect 4073 7288 4204 7328
rect 4244 7288 4253 7328
rect 4300 7319 6164 7328
rect 4300 7288 4652 7319
rect 2860 7244 2900 7288
rect 0 7204 500 7244
rect 2122 7204 2131 7244
rect 2171 7204 2476 7244
rect 2516 7204 2525 7244
rect 2764 7204 2900 7244
rect 3340 7204 3916 7244
rect 3956 7204 3965 7244
rect 0 7184 400 7204
rect 2764 7160 2804 7204
rect 3244 7160 3284 7169
rect 2317 7120 2326 7160
rect 2366 7120 2516 7160
rect 2563 7120 2572 7160
rect 2612 7120 2804 7160
rect 2851 7120 2860 7160
rect 2900 7120 3244 7160
rect 2476 6992 2516 7120
rect 3244 7111 3284 7120
rect 2860 7036 2942 7076
rect 2982 7036 2991 7076
rect 2860 6992 2900 7036
rect 3340 6992 3380 7204
rect 4300 7160 4340 7288
rect 4692 7288 6164 7319
rect 7171 7288 7180 7328
rect 7220 7288 9388 7328
rect 9428 7288 9437 7328
rect 12883 7288 12892 7328
rect 12932 7288 12980 7328
rect 18490 7288 18499 7328
rect 18539 7288 18548 7328
rect 20899 7288 20908 7328
rect 20948 7288 21716 7328
rect 22339 7288 22348 7328
rect 22388 7319 22519 7328
rect 22420 7288 22519 7319
rect 22723 7288 22732 7328
rect 22772 7288 23500 7328
rect 23540 7288 23549 7328
rect 4652 7270 4692 7279
rect 12940 7244 12980 7288
rect 18508 7244 18548 7288
rect 21676 7244 21716 7288
rect 22380 7270 22420 7279
rect 4813 7204 5644 7244
rect 5684 7204 5693 7244
rect 5980 7204 6452 7244
rect 8035 7204 8044 7244
rect 8084 7204 9484 7244
rect 9524 7204 9533 7244
rect 9763 7204 9772 7244
rect 9812 7204 10354 7244
rect 10394 7204 10403 7244
rect 11020 7204 11636 7244
rect 12940 7204 13420 7244
rect 13460 7204 13469 7244
rect 15724 7204 16012 7244
rect 16052 7204 16061 7244
rect 16169 7204 16204 7244
rect 16244 7204 16300 7244
rect 16340 7204 16349 7244
rect 16675 7204 16684 7244
rect 16724 7204 17588 7244
rect 18508 7204 18836 7244
rect 19651 7204 19660 7244
rect 19700 7204 20852 7244
rect 21667 7204 21676 7244
rect 21716 7204 21725 7244
rect 22243 7204 22252 7244
rect 22292 7204 22301 7244
rect 22732 7204 23596 7244
rect 23636 7204 23645 7244
rect 25132 7204 25516 7244
rect 25556 7204 25565 7244
rect 26467 7204 26476 7244
rect 26516 7204 26860 7244
rect 26900 7204 26909 7244
rect 27331 7204 27340 7244
rect 27380 7204 27389 7244
rect 4813 7160 4853 7204
rect 3427 7120 3436 7160
rect 3476 7120 3485 7160
rect 3619 7120 3628 7160
rect 3668 7120 3820 7160
rect 3860 7120 4012 7160
rect 4052 7120 4340 7160
rect 4666 7120 4675 7160
rect 4715 7120 4853 7160
rect 5059 7120 5068 7160
rect 5108 7120 5239 7160
rect 3436 7076 3476 7120
rect 5980 7076 6020 7204
rect 6412 7160 6452 7204
rect 6883 7162 6892 7202
rect 6932 7162 7063 7202
rect 6100 7120 6109 7160
rect 6149 7120 6164 7160
rect 6214 7120 6223 7160
rect 6263 7120 6356 7160
rect 6412 7120 6787 7160
rect 6827 7120 6836 7160
rect 9292 7160 9332 7204
rect 9772 7160 9812 7204
rect 11020 7160 11060 7204
rect 11596 7160 11636 7204
rect 13228 7160 13268 7204
rect 15724 7160 15764 7204
rect 16012 7160 16052 7204
rect 17548 7160 17588 7204
rect 18796 7160 18836 7204
rect 20812 7160 20852 7204
rect 21484 7160 21524 7169
rect 22252 7160 22292 7204
rect 22732 7160 22772 7204
rect 25132 7202 25172 7204
rect 25066 7162 25075 7202
rect 25115 7162 25172 7202
rect 27340 7160 27380 7204
rect 6892 7144 6932 7153
rect 7564 7120 7747 7160
rect 7787 7120 7796 7160
rect 7843 7120 7852 7160
rect 7892 7120 7901 7160
rect 8201 7120 8323 7160
rect 8372 7120 8381 7160
rect 8611 7120 8620 7160
rect 8671 7120 8791 7160
rect 9065 7120 9100 7160
rect 9140 7120 9187 7160
rect 9227 7120 9245 7160
rect 9289 7120 9298 7160
rect 9338 7120 9347 7160
rect 9763 7120 9772 7160
rect 9812 7120 9888 7160
rect 9955 7120 9964 7160
rect 10004 7120 10444 7160
rect 10484 7120 11060 7160
rect 11107 7120 11116 7160
rect 11156 7120 11287 7160
rect 11491 7120 11500 7160
rect 11540 7120 11549 7160
rect 11596 7120 11692 7160
rect 11732 7120 12268 7160
rect 12308 7120 12317 7160
rect 12521 7120 12652 7160
rect 12692 7120 12701 7160
rect 13210 7120 13219 7160
rect 13259 7120 13268 7160
rect 13315 7120 13324 7160
rect 13364 7120 13495 7160
rect 14170 7120 14179 7160
rect 14219 7120 14668 7160
rect 14708 7120 14851 7160
rect 14891 7120 14900 7160
rect 14947 7120 14956 7160
rect 14996 7120 15092 7160
rect 6124 7076 6164 7120
rect 3436 7036 4108 7076
rect 4148 7036 4157 7076
rect 4867 7036 4876 7076
rect 4916 7036 6020 7076
rect 6115 7036 6124 7076
rect 6164 7036 6196 7076
rect 2441 6952 2467 6992
rect 2507 6952 2572 6992
rect 2612 6952 2621 6992
rect 2755 6952 2764 6992
rect 2804 6952 2900 6992
rect 3034 6952 3043 6992
rect 3083 6952 3092 6992
rect 3139 6952 3148 6992
rect 3188 6952 3380 6992
rect 3785 6952 3916 6992
rect 3956 6952 3965 6992
rect 5731 6952 5740 6992
rect 5780 6952 5789 6992
rect 3052 6908 3092 6952
rect 3052 6868 3340 6908
rect 3380 6868 3389 6908
rect 0 6824 400 6844
rect 0 6784 748 6824
rect 788 6784 797 6824
rect 4343 6784 4352 6824
rect 4720 6784 4729 6824
rect 0 6764 400 6784
rect 2764 6616 3052 6656
rect 3092 6616 3101 6656
rect 4937 6616 5068 6656
rect 5108 6616 5117 6656
rect 2764 6572 2804 6616
rect 5740 6572 5780 6952
rect 2746 6532 2755 6572
rect 2795 6532 2804 6572
rect 2947 6532 2956 6572
rect 2996 6532 3188 6572
rect 3148 6488 3188 6532
rect 5644 6532 5780 6572
rect 5980 6572 6020 7036
rect 6316 6992 6356 7120
rect 6220 6952 6356 6992
rect 6403 6952 6412 6992
rect 6452 6983 6740 6992
rect 6452 6952 6691 6983
rect 6220 6656 6260 6952
rect 6682 6943 6691 6952
rect 6731 6943 6740 6983
rect 6682 6942 6740 6943
rect 6211 6616 6220 6656
rect 6260 6616 6269 6656
rect 5980 6532 6068 6572
rect 6979 6532 6988 6572
rect 7028 6532 7418 6572
rect 5644 6488 5684 6532
rect 6028 6488 6068 6532
rect 7378 6490 7418 6532
rect 2371 6448 2380 6488
rect 2420 6448 2429 6488
rect 2563 6448 2572 6488
rect 2637 6448 2743 6488
rect 3130 6448 3139 6488
rect 3179 6448 4780 6488
rect 4820 6448 5452 6488
rect 5492 6448 5501 6488
rect 5581 6448 5590 6488
rect 5630 6448 5684 6488
rect 5801 6448 5932 6488
rect 5972 6448 5981 6488
rect 6028 6448 6071 6488
rect 6111 6448 6120 6488
rect 6281 6448 6412 6488
rect 6452 6448 6461 6488
rect 6508 6448 6527 6488
rect 6567 6448 6576 6488
rect 6691 6448 6700 6488
rect 6740 6448 6871 6488
rect 7145 6448 7267 6488
rect 7316 6448 7325 6488
rect 7369 6450 7378 6490
rect 7418 6450 7427 6490
rect 0 6404 400 6424
rect 0 6364 1132 6404
rect 1172 6364 1181 6404
rect 2153 6364 2284 6404
rect 2324 6364 2333 6404
rect 0 6344 400 6364
rect 2380 6152 2420 6448
rect 6508 6404 6548 6448
rect 2506 6395 2668 6404
rect 2506 6355 2515 6395
rect 2555 6364 2668 6395
rect 2708 6364 2717 6404
rect 4195 6364 4204 6404
rect 4244 6364 4253 6404
rect 5386 6364 5395 6404
rect 5435 6364 5548 6404
rect 5588 6364 5597 6404
rect 5731 6364 5740 6404
rect 5780 6364 6548 6404
rect 2555 6355 2564 6364
rect 2506 6354 2564 6355
rect 7564 6320 7604 7120
rect 7852 6656 7892 7120
rect 11116 7076 11156 7120
rect 8515 7036 8524 7076
rect 8564 7036 11156 7076
rect 8297 6952 8419 6992
rect 8468 6952 8477 6992
rect 9946 6952 9955 6992
rect 9995 6952 10004 6992
rect 10138 6952 10147 6992
rect 10187 6952 10444 6992
rect 10484 6952 10493 6992
rect 9676 6700 9868 6740
rect 9908 6700 9917 6740
rect 9676 6656 9716 6700
rect 7651 6616 7660 6656
rect 7700 6616 7892 6656
rect 8803 6616 8812 6656
rect 8852 6616 9484 6656
rect 9524 6616 9533 6656
rect 9667 6616 9676 6656
rect 9716 6616 9725 6656
rect 9850 6616 9859 6656
rect 9899 6616 9908 6656
rect 7852 6488 7892 6616
rect 9868 6572 9908 6616
rect 8122 6532 8131 6572
rect 8171 6532 9292 6572
rect 9332 6532 9341 6572
rect 9431 6532 9908 6572
rect 9964 6572 10004 6952
rect 11500 6740 11540 7120
rect 12940 7036 14284 7076
rect 14324 7036 14333 7076
rect 14481 7036 14490 7076
rect 14530 7036 14956 7076
rect 14996 7036 15005 7076
rect 11587 6952 11596 6992
rect 11636 6952 11767 6992
rect 12117 6784 12126 6824
rect 12494 6784 12503 6824
rect 11500 6700 11828 6740
rect 11788 6656 11828 6700
rect 12940 6656 12980 7036
rect 13603 6952 13612 6992
rect 13652 6952 13661 6992
rect 13612 6656 13652 6952
rect 14284 6908 14324 7036
rect 15052 6908 15092 7120
rect 15244 7120 15628 7160
rect 15668 7120 15677 7160
rect 15244 6992 15284 7120
rect 15724 7111 15764 7120
rect 15820 7120 15863 7160
rect 15903 7120 15912 7160
rect 15994 7120 16003 7160
rect 16043 7120 16052 7160
rect 16099 7120 16108 7160
rect 16148 7120 16157 7160
rect 16265 7120 16396 7160
rect 16436 7120 16445 7160
rect 16579 7120 16588 7160
rect 16628 7120 17068 7160
rect 17108 7120 17117 7160
rect 17434 7120 17443 7160
rect 17483 7120 17493 7160
rect 17539 7120 17548 7160
rect 17588 7120 17597 7160
rect 17836 7120 18211 7160
rect 18251 7120 18260 7160
rect 18307 7120 18316 7160
rect 18356 7120 18365 7160
rect 18796 7120 18940 7160
rect 18980 7120 18989 7160
rect 19075 7120 19084 7160
rect 19124 7120 19220 7160
rect 19267 7120 19276 7160
rect 19316 7120 19708 7160
rect 19748 7120 19757 7160
rect 19843 7120 19852 7160
rect 19892 7120 19901 7160
rect 19948 7120 20524 7160
rect 20564 7120 20611 7160
rect 20651 7120 20660 7160
rect 20707 7120 20716 7160
rect 20756 7120 20765 7160
rect 20812 7120 21182 7160
rect 21222 7120 21231 7160
rect 21641 7120 21772 7160
rect 21812 7120 21821 7160
rect 21868 7120 21891 7160
rect 21931 7120 21955 7160
rect 22000 7120 22009 7160
rect 22049 7120 22156 7160
rect 22196 7120 22205 7160
rect 22252 7120 22339 7160
rect 22379 7120 22388 7160
rect 22723 7120 22732 7160
rect 22772 7120 22781 7160
rect 23011 7120 23020 7160
rect 23060 7120 23156 7160
rect 23203 7120 23212 7160
rect 23252 7120 24064 7160
rect 24104 7120 24268 7160
rect 24308 7120 24317 7160
rect 25219 7120 25228 7160
rect 25268 7120 25277 7160
rect 25411 7120 25420 7160
rect 25460 7120 25591 7160
rect 25987 7120 25996 7160
rect 26036 7120 26135 7160
rect 26175 7120 26184 7160
rect 26266 7120 26275 7160
rect 26315 7120 26324 7160
rect 26371 7120 26380 7160
rect 26420 7120 26551 7160
rect 27113 7120 27235 7160
rect 27284 7120 27293 7160
rect 27340 7120 27543 7160
rect 27583 7120 27592 7160
rect 15416 7036 15425 7076
rect 15476 7036 15596 7076
rect 15820 6992 15860 7120
rect 16108 7076 16148 7120
rect 15235 6952 15244 6992
rect 15284 6952 15293 6992
rect 15514 6952 15523 6992
rect 15563 6952 15572 6992
rect 15619 6952 15628 6992
rect 15668 6952 15860 6992
rect 16035 7036 16148 7076
rect 17453 7076 17493 7120
rect 17453 7036 17548 7076
rect 17588 7036 17597 7076
rect 14284 6868 15092 6908
rect 15532 6908 15572 6952
rect 16035 6908 16075 7036
rect 17836 6992 17876 7120
rect 18316 7076 18356 7120
rect 18220 7036 18356 7076
rect 16387 6952 16396 6992
rect 16436 6952 16972 6992
rect 17012 6952 17021 6992
rect 17827 6952 17836 6992
rect 17876 6952 17885 6992
rect 18220 6908 18260 7036
rect 15532 6868 16075 6908
rect 17155 6868 17164 6908
rect 17204 6868 18260 6908
rect 14563 6700 14572 6740
rect 14612 6700 18356 6740
rect 11779 6616 11788 6656
rect 11828 6616 11837 6656
rect 12250 6616 12259 6656
rect 12299 6616 12980 6656
rect 13315 6616 13324 6656
rect 13364 6616 13373 6656
rect 13612 6616 13699 6656
rect 13739 6616 13748 6656
rect 11788 6572 11828 6616
rect 13324 6572 13364 6616
rect 9964 6532 10772 6572
rect 11788 6532 12308 6572
rect 13324 6532 13652 6572
rect 13865 6532 13914 6572
rect 13954 6532 13996 6572
rect 14036 6532 14045 6572
rect 14371 6532 14380 6572
rect 14420 6532 15244 6572
rect 15284 6532 15293 6572
rect 9431 6488 9471 6532
rect 10732 6488 10772 6532
rect 7810 6448 7819 6488
rect 7859 6448 7892 6488
rect 8035 6448 8044 6488
rect 8084 6448 8215 6488
rect 8323 6448 8332 6488
rect 8372 6448 8524 6488
rect 8564 6448 8573 6488
rect 8707 6448 8716 6488
rect 8756 6448 8852 6488
rect 9379 6448 9388 6488
rect 9428 6448 9471 6488
rect 9514 6448 9523 6488
rect 9563 6448 9676 6488
rect 9716 6448 9725 6488
rect 9881 6448 9964 6488
rect 10004 6448 10012 6488
rect 10052 6448 10061 6488
rect 10147 6448 10156 6488
rect 10196 6448 10205 6488
rect 10435 6448 10444 6488
rect 10484 6448 10583 6488
rect 10623 6448 10632 6488
rect 10732 6448 10828 6488
rect 10868 6448 10877 6488
rect 11386 6448 11395 6488
rect 11435 6448 11444 6488
rect 11491 6448 11500 6488
rect 11540 6448 11596 6488
rect 11636 6448 11671 6488
rect 11796 6448 11884 6488
rect 11924 6448 11927 6488
rect 11967 6448 11976 6488
rect 12041 6448 12172 6488
rect 12212 6448 12221 6488
rect 7930 6364 7939 6404
rect 7979 6364 7988 6404
rect 7948 6320 7988 6364
rect 4588 6280 7988 6320
rect 8812 6320 8852 6448
rect 10156 6404 10196 6448
rect 11404 6404 11444 6448
rect 12268 6404 12308 6532
rect 13612 6488 13652 6532
rect 15340 6488 15380 6700
rect 18316 6656 18356 6700
rect 19180 6656 19220 7120
rect 19852 7076 19892 7120
rect 19555 7036 19564 7076
rect 19604 7036 19892 7076
rect 19948 6992 19988 7120
rect 15977 6616 16108 6656
rect 16148 6616 16157 6656
rect 16771 6616 16780 6656
rect 16820 6616 16876 6656
rect 16916 6616 16951 6656
rect 18316 6616 18988 6656
rect 19028 6616 19037 6656
rect 19162 6616 19171 6656
rect 19211 6616 19220 6656
rect 19756 6952 19988 6992
rect 15724 6532 15820 6572
rect 15860 6532 15869 6572
rect 15916 6532 16396 6572
rect 16436 6532 16445 6572
rect 16492 6532 17972 6572
rect 15724 6488 15764 6532
rect 15916 6488 15956 6532
rect 16492 6488 16532 6532
rect 17932 6488 17972 6532
rect 18316 6488 18356 6616
rect 19756 6572 19796 6952
rect 20716 6908 20756 7120
rect 21257 7036 21388 7076
rect 21428 7036 21437 7076
rect 21484 6992 21524 7120
rect 21868 7076 21908 7120
rect 23116 7076 23156 7120
rect 25228 7076 25268 7120
rect 26284 7076 26324 7120
rect 21859 7036 21868 7076
rect 21908 7036 21917 7076
rect 22339 7036 22348 7076
rect 22388 7036 23020 7076
rect 23060 7036 23069 7076
rect 23116 7036 23404 7076
rect 23444 7036 24220 7076
rect 24260 7036 24269 7076
rect 24364 7036 25268 7076
rect 25315 7036 25324 7076
rect 25364 7036 27148 7076
rect 27188 7036 27197 7076
rect 27305 7036 27436 7076
rect 27476 7036 27485 7076
rect 20995 6952 21004 6992
rect 21044 6952 21524 6992
rect 22025 6952 22156 6992
rect 22196 6952 23980 6992
rect 24020 6952 24029 6992
rect 20716 6868 21772 6908
rect 21812 6868 21821 6908
rect 19891 6784 19900 6824
rect 20268 6784 20277 6824
rect 20140 6700 21004 6740
rect 21044 6700 21053 6740
rect 19930 6616 19939 6656
rect 19979 6616 19988 6656
rect 18412 6532 19796 6572
rect 12713 6448 12844 6488
rect 12884 6448 12893 6488
rect 13001 6448 13036 6488
rect 13076 6448 13132 6488
rect 13172 6448 13181 6488
rect 13594 6448 13603 6488
rect 13643 6448 13652 6488
rect 13699 6448 13708 6488
rect 13748 6448 14039 6488
rect 14079 6448 14088 6488
rect 14275 6448 14284 6488
rect 14324 6448 14333 6488
rect 14467 6448 14476 6488
rect 14516 6448 15038 6488
rect 15078 6448 15087 6488
rect 15340 6479 15436 6488
rect 9475 6364 9484 6404
rect 9524 6364 10196 6404
rect 10627 6364 10636 6404
rect 10676 6364 10723 6404
rect 10763 6364 10807 6404
rect 10915 6364 10924 6404
rect 10964 6364 10973 6404
rect 11404 6364 11540 6404
rect 12058 6364 12067 6404
rect 12107 6364 12308 6404
rect 13612 6404 13652 6448
rect 13612 6364 14179 6404
rect 14219 6364 14228 6404
rect 8812 6280 9772 6320
rect 9812 6280 9821 6320
rect 4588 6236 4628 6280
rect 8812 6236 8852 6280
rect 10924 6236 10964 6364
rect 11500 6236 11540 6364
rect 14284 6320 14324 6448
rect 15380 6448 15436 6479
rect 15476 6448 15540 6488
rect 15706 6448 15715 6488
rect 15755 6448 15764 6488
rect 15811 6448 15820 6488
rect 15860 6448 15956 6488
rect 16291 6448 16300 6488
rect 16340 6448 16492 6488
rect 16532 6448 16541 6488
rect 16675 6448 16684 6488
rect 16724 6448 16733 6488
rect 16963 6448 16972 6488
rect 17012 6448 17164 6488
rect 17204 6448 17213 6488
rect 17392 6448 17401 6488
rect 17441 6448 17548 6488
rect 17588 6448 17597 6488
rect 17923 6448 17932 6488
rect 17972 6448 17981 6488
rect 18307 6448 18316 6488
rect 18356 6448 18365 6488
rect 15340 6430 15380 6439
rect 15820 6404 15860 6448
rect 14371 6364 14380 6404
rect 14420 6364 14429 6404
rect 15523 6364 15532 6404
rect 15572 6364 15860 6404
rect 16684 6404 16724 6448
rect 16684 6364 17068 6404
rect 17108 6364 17117 6404
rect 17164 6364 17283 6404
rect 17323 6364 17332 6404
rect 13900 6280 14324 6320
rect 13900 6236 13940 6280
rect 14380 6236 14420 6364
rect 17164 6320 17204 6364
rect 15994 6280 16003 6320
rect 16043 6280 17204 6320
rect 3331 6196 3340 6236
rect 3380 6196 4628 6236
rect 4675 6196 4684 6236
rect 4724 6196 5836 6236
rect 5876 6196 5885 6236
rect 6281 6196 6412 6236
rect 6452 6196 6461 6236
rect 6595 6196 6604 6236
rect 6644 6196 7276 6236
rect 7316 6196 8852 6236
rect 9379 6196 9388 6236
rect 9428 6196 9964 6236
rect 10004 6196 10013 6236
rect 10924 6196 11444 6236
rect 11500 6196 11884 6236
rect 11924 6196 12652 6236
rect 12692 6196 12701 6236
rect 12940 6196 13844 6236
rect 13891 6196 13900 6236
rect 13940 6196 13949 6236
rect 14083 6196 14092 6236
rect 14132 6196 14420 6236
rect 15034 6196 15043 6236
rect 15083 6196 16300 6236
rect 16340 6196 16349 6236
rect 2380 6112 7948 6152
rect 7988 6112 7997 6152
rect 8044 6112 10060 6152
rect 10100 6112 10109 6152
rect 8044 6068 8084 6112
rect 11404 6068 11444 6196
rect 12940 6068 12980 6196
rect 3103 6028 3112 6068
rect 3480 6028 3489 6068
rect 6691 6028 6700 6068
rect 6740 6028 8084 6068
rect 9283 6028 9292 6068
rect 9332 6028 10388 6068
rect 10877 6028 10886 6068
rect 11254 6028 11263 6068
rect 11404 6028 12980 6068
rect 13804 6068 13844 6196
rect 15811 6112 15820 6152
rect 15860 6112 17068 6152
rect 17108 6112 17117 6152
rect 18412 6068 18452 6532
rect 19948 6488 19988 6616
rect 20140 6488 20180 6700
rect 24364 6656 24404 7036
rect 24451 6952 24460 6992
rect 24500 6952 24883 6992
rect 24923 6952 25228 6992
rect 25268 6952 25277 6992
rect 27322 6952 27331 6992
rect 27371 6952 27532 6992
rect 27572 6952 27581 6992
rect 27665 6784 27674 6824
rect 28042 6784 28051 6824
rect 20986 6616 20995 6656
rect 21035 6616 21196 6656
rect 21236 6616 21245 6656
rect 21641 6616 21763 6656
rect 21812 6616 21821 6656
rect 22121 6616 22243 6656
rect 22292 6616 22301 6656
rect 23299 6616 23308 6656
rect 23348 6616 23875 6656
rect 23915 6616 23924 6656
rect 23971 6616 23980 6656
rect 24020 6616 24151 6656
rect 24355 6616 24364 6656
rect 24404 6616 24413 6656
rect 20707 6532 20716 6572
rect 20756 6532 21236 6572
rect 21196 6488 21236 6532
rect 21388 6532 21868 6572
rect 21908 6532 21917 6572
rect 21964 6532 22156 6572
rect 22196 6532 22205 6572
rect 23395 6532 23404 6572
rect 23444 6532 24208 6572
rect 21388 6488 21428 6532
rect 19459 6448 19468 6488
rect 19508 6448 19988 6488
rect 20116 6448 20125 6488
rect 20165 6448 20180 6488
rect 20227 6448 20236 6488
rect 20276 6448 20407 6488
rect 20532 6448 20620 6488
rect 20660 6448 20663 6488
rect 20703 6448 20712 6488
rect 20899 6448 20908 6488
rect 20948 6448 21079 6488
rect 21187 6448 21196 6488
rect 21236 6448 21245 6488
rect 21370 6448 21379 6488
rect 21419 6448 21428 6488
rect 21475 6448 21484 6488
rect 21524 6448 21533 6488
rect 21915 6448 21924 6488
rect 21964 6448 22004 6532
rect 24168 6488 24208 6532
rect 22051 6448 22060 6488
rect 22100 6448 22109 6488
rect 22217 6448 22348 6488
rect 22388 6448 22397 6488
rect 23465 6448 23596 6488
rect 23636 6448 23645 6488
rect 23768 6448 23777 6488
rect 23817 6448 23828 6488
rect 23945 6448 24076 6488
rect 24116 6448 24125 6488
rect 24168 6448 24263 6488
rect 24303 6448 24312 6488
rect 24442 6448 24451 6488
rect 24500 6448 24631 6488
rect 19267 6364 19276 6404
rect 19316 6364 19378 6404
rect 19418 6364 20803 6404
rect 20843 6364 20852 6404
rect 21161 6280 21292 6320
rect 21332 6280 21341 6320
rect 13804 6028 18452 6068
rect 18513 6196 18556 6236
rect 18596 6196 18605 6236
rect 0 5984 400 6004
rect 0 5944 460 5984
rect 500 5944 509 5984
rect 0 5924 400 5944
rect 5609 5860 5740 5900
rect 5780 5860 5789 5900
rect 9667 5860 9676 5900
rect 9716 5860 9908 5900
rect 2668 5776 2900 5816
rect 4867 5776 4876 5816
rect 4916 5776 5204 5816
rect 6499 5776 6508 5816
rect 6548 5776 8180 5816
rect 8873 5776 9004 5816
rect 9044 5776 9053 5816
rect 2668 5732 2708 5776
rect 2572 5692 2708 5732
rect 2860 5732 2900 5776
rect 5164 5732 5204 5776
rect 6508 5732 6548 5776
rect 8140 5732 8180 5776
rect 9868 5732 9908 5860
rect 10348 5816 10388 6028
rect 10435 5860 10444 5900
rect 10484 5860 14228 5900
rect 14345 5860 14380 5900
rect 14420 5860 14476 5900
rect 14516 5860 14525 5900
rect 14921 5860 15043 5900
rect 15092 5860 15101 5900
rect 14188 5816 14228 5860
rect 18513 5816 18553 6196
rect 21484 6152 21524 6448
rect 22060 6404 22100 6448
rect 23788 6404 23828 6448
rect 24076 6430 24116 6439
rect 22060 6364 22580 6404
rect 23779 6364 23788 6404
rect 23828 6364 23864 6404
rect 22540 6320 22580 6364
rect 23788 6320 23828 6364
rect 22531 6280 22540 6320
rect 22580 6280 23828 6320
rect 22793 6196 22924 6236
rect 22964 6196 22973 6236
rect 24442 6196 24451 6236
rect 24491 6196 24500 6236
rect 24460 6152 24500 6196
rect 21484 6112 24500 6152
rect 18651 6028 18660 6068
rect 19028 6028 19037 6068
rect 19555 6028 19564 6068
rect 19604 6028 22252 6068
rect 22292 6028 22301 6068
rect 26425 6028 26434 6068
rect 26802 6028 26811 6068
rect 21085 5944 21388 5984
rect 21428 5944 23636 5984
rect 20489 5860 20611 5900
rect 20660 5860 20669 5900
rect 20777 5860 20908 5900
rect 20948 5860 20957 5900
rect 21085 5816 21125 5944
rect 23596 5900 23636 5944
rect 22051 5860 22060 5900
rect 22100 5860 22348 5900
rect 22388 5860 23212 5900
rect 23252 5860 23261 5900
rect 23465 5860 23596 5900
rect 23636 5860 23645 5900
rect 10348 5776 12940 5816
rect 12980 5776 12989 5816
rect 13411 5776 13420 5816
rect 13460 5776 13469 5816
rect 14188 5776 18452 5816
rect 18513 5776 18740 5816
rect 20227 5776 20236 5816
rect 20276 5776 21125 5816
rect 23020 5776 23788 5816
rect 23828 5776 23837 5816
rect 13420 5732 13460 5776
rect 2860 5692 3668 5732
rect 2275 5608 2284 5648
rect 2324 5608 2462 5648
rect 2502 5608 2511 5648
rect 2572 5564 2612 5692
rect 2764 5648 2804 5657
rect 3628 5648 3668 5692
rect 4108 5692 5108 5732
rect 5164 5692 6548 5732
rect 6691 5692 6700 5732
rect 6740 5692 8044 5732
rect 8084 5692 8093 5732
rect 8140 5692 8660 5732
rect 9868 5692 10659 5732
rect 10699 5692 11156 5732
rect 13420 5692 14132 5732
rect 2659 5608 2668 5648
rect 2708 5608 2764 5648
rect 2804 5608 2839 5648
rect 2938 5608 2947 5648
rect 2996 5608 3127 5648
rect 3619 5608 3628 5648
rect 3668 5608 3677 5648
rect 3785 5608 3907 5648
rect 3956 5608 3965 5648
rect 2764 5599 2804 5608
rect 3916 5564 3956 5608
rect 4108 5564 4148 5692
rect 5068 5648 5108 5692
rect 8620 5648 8660 5692
rect 11116 5648 11156 5692
rect 4195 5608 4204 5648
rect 4244 5608 4563 5648
rect 4603 5608 4623 5648
rect 4674 5608 4683 5648
rect 4723 5608 4780 5648
rect 4820 5608 4863 5648
rect 5059 5608 5068 5648
rect 5108 5608 5117 5648
rect 6106 5608 6115 5648
rect 6155 5608 6164 5648
rect 6211 5608 6220 5648
rect 6260 5608 6391 5648
rect 6473 5608 6604 5648
rect 6644 5608 6653 5648
rect 6787 5608 6796 5648
rect 6836 5608 6988 5648
rect 7028 5608 7123 5648
rect 7163 5608 7188 5648
rect 7309 5608 7318 5648
rect 7358 5608 7459 5648
rect 7499 5608 7508 5648
rect 8131 5608 8140 5648
rect 8180 5608 8189 5648
rect 8611 5608 8620 5648
rect 8660 5608 8669 5648
rect 9257 5608 9379 5648
rect 9428 5608 9437 5648
rect 9763 5608 9772 5648
rect 9812 5608 10060 5648
rect 10100 5608 10109 5648
rect 10531 5608 10540 5648
rect 10580 5608 10589 5648
rect 10768 5608 10777 5648
rect 10817 5608 10964 5648
rect 11098 5608 11107 5648
rect 11147 5608 11156 5648
rect 11203 5608 11212 5648
rect 11252 5608 11444 5648
rect 11491 5608 11500 5648
rect 11540 5608 11644 5648
rect 11684 5608 11693 5648
rect 11753 5608 11834 5648
rect 11874 5608 11884 5648
rect 11924 5608 11933 5648
rect 12137 5608 12172 5648
rect 12212 5608 12268 5648
rect 12308 5608 12317 5648
rect 12425 5608 12556 5648
rect 12596 5608 12605 5648
rect 12835 5608 12844 5648
rect 12884 5608 13027 5648
rect 13067 5608 13076 5648
rect 13135 5615 13144 5655
rect 13184 5615 13268 5655
rect 14092 5648 14132 5692
rect 14380 5692 14900 5732
rect 15235 5692 15244 5732
rect 15284 5692 15860 5732
rect 16291 5692 16300 5732
rect 16340 5692 17780 5732
rect 14380 5648 14420 5692
rect 14860 5648 14900 5692
rect 15820 5648 15860 5692
rect 17740 5648 17780 5692
rect 18412 5648 18452 5776
rect 18700 5648 18740 5776
rect 18883 5692 18892 5732
rect 18932 5692 19564 5732
rect 19604 5692 19613 5732
rect 19564 5648 19604 5692
rect 20428 5648 20468 5776
rect 20620 5692 20812 5732
rect 20852 5692 20861 5732
rect 20620 5648 20660 5692
rect 20908 5648 20948 5776
rect 23020 5732 23060 5776
rect 21161 5692 21292 5732
rect 21332 5692 21341 5732
rect 22944 5692 23060 5732
rect 4583 5564 4623 5608
rect 6124 5564 6164 5608
rect 2554 5524 2563 5564
rect 2603 5524 2612 5564
rect 3523 5524 3532 5564
rect 3572 5524 3956 5564
rect 4099 5524 4108 5564
rect 4148 5524 4157 5564
rect 4209 5524 4218 5564
rect 4258 5524 4532 5564
rect 4583 5524 5588 5564
rect 6077 5524 6124 5564
rect 6164 5524 6173 5564
rect 6394 5524 6403 5564
rect 6443 5524 7564 5564
rect 7604 5524 7613 5564
rect 4492 5480 4532 5524
rect 5548 5480 5588 5524
rect 2508 5440 2572 5480
rect 2612 5440 2668 5480
rect 2708 5440 4003 5480
rect 4043 5440 4204 5480
rect 4244 5440 4253 5480
rect 4492 5440 4588 5480
rect 4628 5440 4637 5480
rect 5539 5440 5548 5480
rect 5588 5440 6124 5480
rect 6164 5440 6173 5480
rect 4588 5396 4628 5440
rect 4588 5356 6988 5396
rect 7028 5356 7037 5396
rect 4343 5272 4352 5312
rect 4720 5272 4729 5312
rect 6115 5272 6124 5312
rect 6164 5272 7180 5312
rect 7220 5272 7229 5312
rect 8140 5144 8180 5608
rect 8524 5524 8948 5564
rect 9353 5524 9484 5564
rect 9524 5524 9533 5564
rect 9681 5524 9690 5564
rect 9730 5524 9859 5564
rect 9899 5524 9908 5564
rect 10313 5524 10444 5564
rect 10484 5524 10493 5564
rect 8524 5480 8564 5524
rect 8908 5480 8948 5524
rect 10540 5480 10580 5608
rect 10924 5564 10964 5608
rect 11404 5564 11444 5608
rect 12172 5564 12212 5608
rect 12844 5564 12884 5608
rect 10924 5524 11444 5564
rect 11971 5524 11980 5564
rect 12020 5524 12212 5564
rect 12652 5524 12884 5564
rect 8393 5440 8515 5480
rect 8564 5440 8573 5480
rect 8803 5440 8812 5480
rect 8852 5440 8861 5480
rect 8908 5440 10147 5480
rect 10187 5440 10196 5480
rect 10540 5440 11308 5480
rect 11348 5440 11357 5480
rect 5068 5104 6412 5144
rect 6452 5104 6461 5144
rect 7363 5104 7372 5144
rect 7412 5104 8180 5144
rect 5068 5060 5108 5104
rect 5050 5020 5059 5060
rect 5099 5020 5108 5060
rect 5321 5020 5452 5060
rect 5492 5020 8468 5060
rect 5452 4976 5492 5020
rect 8428 4976 8468 5020
rect 5434 4936 5443 4976
rect 5483 4936 5492 4976
rect 5635 4936 5644 4976
rect 5684 4936 7316 4976
rect 6211 4852 6220 4892
rect 6260 4852 6269 4892
rect 7276 4724 7316 4936
rect 7372 4967 7604 4976
rect 7372 4936 7555 4967
rect 7372 4808 7412 4936
rect 7546 4927 7555 4936
rect 7595 4927 7604 4967
rect 8410 4936 8419 4976
rect 8459 4936 8468 4976
rect 8812 4976 8852 5440
rect 11404 5144 11444 5524
rect 12652 5480 12692 5524
rect 11491 5440 11500 5480
rect 11540 5440 11788 5480
rect 11828 5440 11837 5480
rect 11971 5440 11980 5480
rect 12020 5440 12172 5480
rect 12212 5440 12221 5480
rect 12643 5440 12652 5480
rect 12692 5440 12701 5480
rect 12809 5471 12940 5480
rect 12809 5440 12931 5471
rect 12980 5440 12989 5480
rect 12922 5431 12931 5440
rect 12971 5431 12980 5440
rect 12922 5430 12980 5431
rect 12117 5272 12126 5312
rect 12494 5272 12503 5312
rect 13228 5144 13268 5615
rect 13673 5608 13804 5648
rect 13844 5608 13853 5648
rect 14074 5608 14083 5648
rect 14123 5608 14132 5648
rect 14371 5608 14380 5648
rect 14420 5608 14429 5648
rect 14746 5608 14755 5648
rect 14795 5608 14804 5648
rect 14851 5608 14860 5648
rect 14900 5608 14909 5648
rect 15353 5608 15436 5648
rect 15476 5608 15484 5648
rect 15524 5608 15533 5648
rect 15619 5608 15628 5648
rect 15668 5608 15764 5648
rect 15820 5608 16204 5648
rect 16244 5608 16253 5648
rect 16300 5608 16323 5648
rect 16363 5608 16372 5648
rect 16432 5608 16441 5648
rect 16481 5608 16492 5648
rect 16532 5608 16684 5648
rect 16724 5608 16733 5648
rect 16937 5608 17068 5648
rect 17108 5608 17117 5648
rect 17164 5608 17635 5648
rect 17675 5608 17684 5648
rect 17731 5608 17740 5648
rect 17780 5608 17789 5648
rect 18281 5608 18412 5648
rect 18452 5608 18461 5648
rect 18569 5608 18700 5648
rect 18740 5608 18796 5648
rect 18836 5608 18845 5648
rect 19075 5608 19084 5648
rect 19124 5608 19180 5648
rect 19220 5608 19255 5648
rect 19555 5608 19564 5648
rect 19604 5608 19613 5648
rect 20419 5608 20428 5648
rect 20468 5608 20477 5648
rect 20602 5608 20611 5648
rect 20651 5608 20660 5648
rect 20803 5608 20812 5648
rect 20852 5608 20948 5648
rect 20995 5608 21004 5648
rect 21044 5608 21175 5648
rect 21658 5608 21667 5648
rect 21716 5608 21847 5648
rect 14092 5564 14132 5608
rect 14764 5564 14804 5608
rect 14092 5524 14804 5564
rect 14860 5564 14900 5608
rect 15724 5564 15764 5608
rect 16300 5564 16340 5608
rect 14860 5524 15380 5564
rect 15523 5524 15532 5564
rect 15572 5524 15764 5564
rect 15811 5524 15820 5564
rect 15860 5524 16340 5564
rect 15340 5480 15380 5524
rect 17164 5480 17204 5608
rect 17260 5524 20908 5564
rect 20948 5524 20957 5564
rect 13603 5440 13612 5480
rect 13652 5440 13661 5480
rect 13882 5440 13891 5480
rect 13931 5440 14380 5480
rect 14420 5440 14429 5480
rect 15322 5440 15331 5480
rect 15371 5440 15380 5480
rect 16099 5440 16108 5480
rect 16148 5440 16204 5480
rect 16244 5440 16279 5480
rect 17155 5440 17164 5480
rect 17204 5440 17213 5480
rect 13612 5396 13652 5440
rect 17260 5396 17300 5524
rect 17993 5440 18028 5480
rect 18068 5440 18124 5480
rect 18164 5440 18173 5480
rect 18298 5440 18307 5480
rect 18347 5440 18356 5480
rect 18979 5440 18988 5480
rect 19028 5440 19037 5480
rect 19084 5440 19267 5480
rect 19307 5440 19316 5480
rect 20227 5440 20236 5480
rect 20276 5440 20285 5480
rect 13612 5356 17300 5396
rect 13612 5144 13652 5356
rect 18316 5312 18356 5440
rect 16003 5272 16012 5312
rect 16052 5272 18356 5312
rect 18412 5188 18892 5228
rect 18932 5188 18941 5228
rect 18412 5144 18452 5188
rect 10339 5104 10348 5144
rect 10388 5104 11252 5144
rect 11386 5104 11395 5144
rect 11435 5104 11444 5144
rect 11971 5104 11980 5144
rect 12020 5104 12259 5144
rect 12299 5104 12308 5144
rect 12547 5104 12556 5144
rect 12596 5104 13268 5144
rect 13324 5104 13652 5144
rect 15401 5104 15532 5144
rect 15572 5104 15581 5144
rect 18403 5104 18412 5144
rect 18452 5104 18461 5144
rect 18569 5104 18691 5144
rect 18740 5104 18749 5144
rect 11212 4976 11252 5104
rect 12643 5020 12652 5060
rect 12692 5020 12701 5060
rect 12826 5020 12835 5060
rect 12875 5020 13219 5060
rect 13259 5020 13268 5060
rect 12652 4976 12692 5020
rect 12931 4976 12980 4978
rect 13324 4976 13364 5104
rect 18988 5060 19028 5440
rect 13612 5020 15340 5060
rect 15380 5020 16532 5060
rect 16675 5020 16684 5060
rect 16724 5020 18836 5060
rect 18897 5020 18906 5060
rect 18946 5020 19028 5060
rect 13612 4976 13652 5020
rect 16492 4976 16532 5020
rect 18796 4976 18836 5020
rect 19084 4976 19124 5440
rect 20236 5396 20276 5440
rect 20236 5356 20372 5396
rect 19891 5272 19900 5312
rect 20268 5272 20277 5312
rect 20332 4976 20372 5356
rect 21436 5272 23404 5312
rect 23444 5272 23453 5312
rect 27665 5272 27674 5312
rect 28042 5272 28051 5312
rect 21436 5144 21476 5272
rect 21955 5188 21964 5228
rect 22004 5188 22013 5228
rect 21964 5144 22004 5188
rect 21427 5104 21436 5144
rect 21476 5104 21485 5144
rect 21737 5104 21868 5144
rect 21908 5104 21917 5144
rect 21964 5104 22252 5144
rect 22292 5104 22301 5144
rect 20995 5020 21004 5060
rect 21044 5020 21716 5060
rect 21969 5020 21978 5060
rect 22018 5020 22924 5060
rect 22964 5020 22973 5060
rect 21676 4976 21716 5020
rect 8812 4936 10892 4976
rect 11203 4936 11212 4976
rect 11252 4936 11261 4976
rect 11561 4936 11692 4976
rect 11732 4936 11741 4976
rect 12355 4936 12364 4976
rect 12404 4936 12556 4976
rect 12596 4936 12605 4976
rect 12652 4936 12738 4976
rect 12778 4936 12787 4976
rect 12922 4936 12931 4976
rect 12971 4936 12980 4976
rect 13027 4936 13036 4976
rect 13076 4936 13364 4976
rect 13594 4936 13603 4976
rect 13643 4936 13652 4976
rect 16474 4936 16483 4976
rect 16523 4936 16532 4976
rect 18403 4936 18412 4976
rect 18452 4936 18595 4976
rect 18635 4936 18644 4976
rect 18796 4936 19124 4976
rect 7546 4926 7604 4927
rect 7660 4852 7708 4892
rect 7748 4852 7757 4892
rect 7913 4852 8044 4892
rect 8084 4852 8093 4892
rect 8995 4852 9004 4892
rect 9044 4852 9053 4892
rect 7363 4768 7372 4808
rect 7412 4768 7421 4808
rect 7660 4724 7700 4852
rect 10051 4768 10060 4808
rect 10100 4768 10540 4808
rect 10580 4768 10589 4808
rect 6979 4684 6988 4724
rect 7028 4684 7037 4724
rect 7276 4684 7700 4724
rect 9571 4684 9580 4724
rect 9620 4684 9964 4724
rect 10004 4684 10013 4724
rect 10217 4684 10348 4724
rect 10388 4684 10397 4724
rect 6988 4640 7028 4684
rect 10852 4640 10892 4936
rect 12364 4892 12404 4936
rect 11593 4852 11602 4892
rect 11642 4852 11884 4892
rect 11924 4852 12404 4892
rect 12931 4808 12971 4936
rect 14371 4852 14380 4892
rect 14420 4852 14429 4892
rect 15017 4852 15148 4892
rect 15188 4852 15197 4892
rect 15977 4852 16108 4892
rect 16148 4852 16157 4892
rect 17155 4852 17164 4892
rect 17204 4852 17213 4892
rect 17923 4852 17932 4892
rect 17972 4852 18028 4892
rect 18068 4852 18103 4892
rect 19084 4808 19124 4936
rect 20122 4967 20372 4976
rect 20122 4927 20131 4967
rect 20171 4936 20372 4967
rect 20777 4936 20908 4976
rect 20948 4936 20957 4976
rect 21004 4936 21104 4976
rect 21144 4936 21153 4976
rect 21257 4936 21292 4976
rect 21332 4936 21388 4976
rect 21428 4936 21437 4976
rect 21658 4936 21667 4976
rect 21707 4936 21716 4976
rect 21763 4936 21772 4976
rect 21812 4936 21943 4976
rect 22147 4936 22156 4976
rect 22196 4936 22205 4976
rect 22339 4936 22348 4976
rect 22388 4936 22519 4976
rect 20171 4927 20180 4936
rect 20122 4926 20180 4927
rect 21004 4892 21044 4936
rect 20236 4852 20284 4892
rect 20324 4852 21044 4892
rect 22156 4892 22196 4936
rect 22156 4852 24460 4892
rect 24500 4852 24509 4892
rect 20236 4808 20276 4852
rect 12931 4768 13228 4808
rect 13268 4768 13277 4808
rect 19084 4768 20276 4808
rect 20908 4808 20948 4852
rect 20908 4768 21772 4808
rect 21812 4768 21821 4808
rect 22156 4724 22196 4852
rect 18883 4684 18892 4724
rect 18932 4684 19276 4724
rect 19316 4684 19325 4724
rect 20995 4684 21004 4724
rect 21044 4684 22196 4724
rect 6988 4600 8716 4640
rect 8756 4600 8765 4640
rect 10852 4600 13804 4640
rect 13844 4600 13853 4640
rect 17059 4600 17068 4640
rect 17108 4600 20812 4640
rect 20852 4600 20861 4640
rect 3103 4516 3112 4556
rect 3480 4516 3489 4556
rect 10877 4516 10886 4556
rect 11254 4516 11263 4556
rect 18651 4516 18660 4556
rect 19028 4516 19037 4556
rect 26425 4516 26434 4556
rect 26802 4516 26811 4556
rect 7939 4432 7948 4472
rect 7988 4432 15244 4472
rect 15284 4432 15293 4472
rect 7843 4348 7852 4388
rect 7892 4348 8044 4388
rect 8084 4348 8093 4388
rect 13097 4348 13228 4388
rect 13268 4348 13277 4388
rect 14284 4348 15148 4388
rect 15188 4348 15197 4388
rect 15977 4348 16108 4388
rect 16148 4348 16157 4388
rect 14284 4304 14324 4348
rect 6089 4264 6220 4304
rect 6260 4264 6269 4304
rect 7171 4264 7180 4304
rect 7220 4264 8476 4304
rect 8516 4264 8525 4304
rect 11491 4264 11500 4304
rect 11540 4264 11788 4304
rect 11828 4264 11837 4304
rect 13577 4264 13708 4304
rect 13748 4264 13757 4304
rect 13891 4264 13900 4304
rect 13940 4264 14324 4304
rect 14371 4264 14380 4304
rect 14420 4264 14476 4304
rect 14516 4264 14551 4304
rect 17033 4264 17164 4304
rect 17204 4264 17213 4304
rect 7564 4180 8259 4220
rect 8299 4180 8308 4220
rect 8515 4180 8524 4220
rect 8564 4180 9811 4220
rect 9851 4180 9860 4220
rect 10579 4180 10588 4220
rect 10628 4180 11980 4220
rect 12020 4180 12029 4220
rect 13228 4180 13804 4220
rect 13844 4180 14132 4220
rect 14275 4180 14284 4220
rect 14324 4180 15187 4220
rect 15227 4180 15236 4220
rect 7564 4136 7604 4180
rect 8524 4136 8564 4180
rect 13228 4136 13268 4180
rect 14092 4136 14132 4180
rect 14284 4136 14324 4180
rect 7433 4096 7555 4136
rect 7604 4096 7613 4136
rect 7939 4096 7948 4136
rect 7988 4096 8140 4136
rect 8180 4096 8189 4136
rect 8332 4096 8377 4136
rect 8417 4096 8564 4136
rect 8611 4096 8620 4136
rect 8660 4096 8716 4136
rect 8756 4096 8791 4136
rect 9929 4096 10006 4136
rect 10046 4096 10060 4136
rect 10100 4096 10109 4136
rect 10339 4096 10348 4136
rect 10427 4096 10519 4136
rect 11561 4096 11692 4136
rect 11732 4096 11741 4136
rect 11875 4096 11884 4136
rect 11924 4096 12055 4136
rect 13219 4096 13228 4136
rect 13268 4096 13277 4136
rect 13411 4096 13420 4136
rect 13460 4096 13469 4136
rect 13769 4096 13804 4136
rect 13844 4096 13900 4136
rect 13940 4096 13949 4136
rect 14083 4096 14092 4136
rect 14132 4096 14141 4136
rect 14188 4096 14324 4136
rect 15373 4096 15382 4136
rect 15422 4096 15532 4136
rect 15572 4096 15581 4136
rect 15689 4096 15811 4136
rect 15860 4096 15869 4136
rect 16073 4096 16122 4136
rect 16162 4096 16204 4136
rect 16244 4096 16253 4136
rect 7857 4012 7866 4052
rect 7906 4012 8044 4052
rect 8084 4012 8093 4052
rect 8332 3968 8372 4096
rect 11692 4052 11732 4096
rect 13420 4052 13460 4096
rect 14188 4052 14228 4096
rect 15820 4052 15860 4096
rect 11692 4012 14228 4052
rect 14284 4012 15860 4052
rect 15907 4012 15916 4052
rect 15956 4012 16684 4052
rect 16724 4012 16733 4052
rect 14284 3968 14324 4012
rect 7642 3928 7651 3968
rect 7691 3928 8372 3968
rect 13699 3928 13708 3968
rect 13748 3928 13987 3968
rect 14027 3928 14036 3968
rect 14275 3928 14284 3968
rect 14324 3928 14333 3968
rect 4343 3760 4352 3800
rect 4720 3760 4729 3800
rect 12117 3760 12126 3800
rect 12494 3760 12503 3800
rect 19891 3760 19900 3800
rect 20268 3760 20277 3800
rect 27665 3760 27674 3800
rect 28042 3760 28051 3800
rect 3103 3004 3112 3044
rect 3480 3004 3489 3044
rect 10877 3004 10886 3044
rect 11254 3004 11263 3044
rect 18651 3004 18660 3044
rect 19028 3004 19037 3044
rect 26425 3004 26434 3044
rect 26802 3004 26811 3044
rect 4343 2248 4352 2288
rect 4720 2248 4729 2288
rect 12117 2248 12126 2288
rect 12494 2248 12503 2288
rect 19891 2248 19900 2288
rect 20268 2248 20277 2288
rect 27665 2248 27674 2288
rect 28042 2248 28051 2288
rect 3103 1492 3112 1532
rect 3480 1492 3489 1532
rect 10877 1492 10886 1532
rect 11254 1492 11263 1532
rect 18651 1492 18660 1532
rect 19028 1492 19037 1532
rect 26425 1492 26434 1532
rect 26802 1492 26811 1532
rect 4343 736 4352 776
rect 4720 736 4729 776
rect 12117 736 12126 776
rect 12494 736 12503 776
rect 19891 736 19900 776
rect 20268 736 20277 776
rect 27665 736 27674 776
rect 28042 736 28051 776
<< via2 >>
rect 16396 28624 16436 28664
rect 9100 28540 9140 28580
rect 29260 28540 29300 28580
rect 30028 28540 30068 28580
rect 2956 28456 2996 28496
rect 9196 28456 9236 28496
rect 13900 28456 13940 28496
rect 25516 28456 25556 28496
rect 1804 28372 1844 28412
rect 7084 28372 7124 28412
rect 6796 28204 6836 28244
rect 2764 28120 2804 28160
rect 3532 28120 3572 28160
rect 8236 28120 8276 28160
rect 27724 28120 27764 28160
rect 30988 28120 31028 28160
rect 1900 28036 1940 28076
rect 5932 28036 5972 28076
rect 2188 27952 2228 27992
rect 2956 27952 2996 27992
rect 4352 27952 4720 27992
rect 12126 27952 12494 27992
rect 14092 27952 14132 27992
rect 19900 27952 20268 27992
rect 25228 27952 25268 27992
rect 27674 27952 28042 27992
rect 5452 27868 5492 27908
rect 10636 27868 10676 27908
rect 26956 27868 26996 27908
rect 6988 27784 7028 27824
rect 25420 27784 25460 27824
rect 1900 27700 1940 27740
rect 2476 27700 2516 27740
rect 6700 27700 6740 27740
rect 9292 27700 9332 27740
rect 10060 27700 10100 27740
rect 12940 27700 12980 27740
rect 17068 27700 17108 27740
rect 29260 27700 29300 27740
rect 1804 27616 1844 27656
rect 2668 27616 2708 27656
rect 3148 27616 3179 27656
rect 3179 27616 3188 27656
rect 4396 27616 4436 27656
rect 5740 27616 5780 27656
rect 7372 27616 7412 27656
rect 11308 27616 11348 27656
rect 12172 27616 12212 27656
rect 2188 27532 2228 27572
rect 2956 27532 2996 27572
rect 6508 27532 6548 27572
rect 7468 27532 7508 27572
rect 9580 27532 9620 27572
rect 10540 27532 10580 27572
rect 14188 27532 14228 27572
rect 15340 27616 15380 27656
rect 15628 27616 15668 27656
rect 19180 27616 19220 27656
rect 22348 27616 22379 27656
rect 22379 27616 22388 27656
rect 26860 27616 26900 27656
rect 29356 27616 29396 27656
rect 30124 27616 30164 27656
rect 30412 27616 30452 27656
rect 15052 27532 15092 27572
rect 15724 27532 15764 27572
rect 21100 27532 21140 27572
rect 21964 27532 22004 27572
rect 22540 27532 22580 27572
rect 24940 27532 24980 27572
rect 26956 27532 26996 27572
rect 27340 27532 27380 27572
rect 30604 27532 30644 27572
rect 30892 27532 30932 27572
rect 2092 27448 2132 27488
rect 2380 27448 2411 27488
rect 2411 27448 2420 27488
rect 2764 27448 2804 27488
rect 3532 27448 3572 27488
rect 14860 27448 14900 27488
rect 19084 27448 19124 27488
rect 8620 27364 8660 27404
rect 10732 27364 10772 27404
rect 15820 27364 15860 27404
rect 16108 27364 16148 27404
rect 17548 27364 17579 27404
rect 17579 27364 17588 27404
rect 20428 27364 20468 27404
rect 21196 27364 21236 27404
rect 23404 27364 23444 27404
rect 25900 27364 25940 27404
rect 27916 27364 27956 27404
rect 29164 27364 29204 27404
rect 29644 27364 29684 27404
rect 3916 27280 3956 27320
rect 8524 27280 8564 27320
rect 10348 27280 10388 27320
rect 12076 27280 12116 27320
rect 14764 27280 14804 27320
rect 14956 27280 14996 27320
rect 23308 27280 23348 27320
rect 3112 27196 3480 27236
rect 10886 27196 11254 27236
rect 18660 27196 19028 27236
rect 26434 27196 26802 27236
rect 10444 27112 10484 27152
rect 13516 27112 13556 27152
rect 21004 27112 21044 27152
rect 2092 27028 2132 27068
rect 6700 27028 6731 27068
rect 6731 27028 6740 27068
rect 9580 27028 9620 27068
rect 11212 27028 11252 27068
rect 12076 27028 12116 27068
rect 13420 27028 13460 27068
rect 19180 27028 19220 27068
rect 19372 27028 19412 27068
rect 21964 27028 22004 27068
rect 26860 27028 26900 27068
rect 30124 27028 30164 27068
rect 2860 26944 2900 26984
rect 6508 26944 6548 26984
rect 8524 26944 8564 26984
rect 3244 26860 3275 26900
rect 3275 26860 3284 26900
rect 3532 26860 3572 26900
rect 7948 26860 7988 26900
rect 2668 26776 2699 26816
rect 2699 26776 2708 26816
rect 2860 26776 2900 26816
rect 4588 26776 4628 26816
rect 5068 26776 5108 26816
rect 5548 26776 5588 26816
rect 5932 26776 5972 26816
rect 6508 26776 6548 26816
rect 6892 26797 6932 26837
rect 7180 26776 7220 26816
rect 8620 26776 8660 26816
rect 11692 26944 11732 26984
rect 13324 26944 13364 26984
rect 15724 26944 15764 26984
rect 10924 26860 10964 26900
rect 12172 26860 12212 26900
rect 18316 26860 18356 26900
rect 18508 26860 18548 26900
rect 19372 26860 19412 26900
rect 23404 26860 23444 26900
rect 30124 26860 30164 26900
rect 5260 26692 5300 26732
rect 5644 26692 5684 26732
rect 7084 26692 7124 26732
rect 8140 26692 8180 26732
rect 8332 26692 8372 26732
rect 10444 26776 10484 26816
rect 12556 26776 12596 26816
rect 13324 26776 13345 26816
rect 13345 26776 13364 26816
rect 13804 26776 13844 26816
rect 17068 26776 17099 26816
rect 17099 26776 17108 26816
rect 1516 26608 1556 26648
rect 1900 26608 1940 26648
rect 3340 26608 3380 26648
rect 4684 26608 4724 26648
rect 5452 26608 5483 26648
rect 5483 26608 5492 26648
rect 19660 26776 19700 26816
rect 20332 26776 20372 26816
rect 21196 26776 21236 26816
rect 21484 26776 21524 26816
rect 23116 26776 23156 26816
rect 24076 26776 24116 26816
rect 25900 26776 25940 26816
rect 27052 26776 27092 26816
rect 27916 26776 27956 26816
rect 29356 26776 29396 26816
rect 7564 26608 7604 26648
rect 10732 26692 10772 26732
rect 12652 26692 12692 26732
rect 13516 26692 13556 26732
rect 13996 26692 14036 26732
rect 15052 26692 15083 26732
rect 15083 26692 15092 26732
rect 17548 26692 17588 26732
rect 17740 26692 17780 26732
rect 9580 26608 9620 26648
rect 10156 26608 10196 26648
rect 10348 26608 10379 26648
rect 10379 26608 10388 26648
rect 11116 26608 11156 26648
rect 11596 26608 11636 26648
rect 8428 26524 8468 26564
rect 11788 26524 11828 26564
rect 2092 26440 2132 26480
rect 4352 26440 4720 26480
rect 7756 26440 7796 26480
rect 7948 26440 7988 26480
rect 10444 26440 10484 26480
rect 5164 26356 5204 26396
rect 5356 26356 5396 26396
rect 11884 26356 11924 26396
rect 12460 26608 12500 26648
rect 12940 26608 12980 26648
rect 13708 26608 13748 26648
rect 13900 26608 13940 26648
rect 18412 26608 18452 26648
rect 18892 26608 18932 26648
rect 20140 26608 20180 26648
rect 20428 26608 20459 26648
rect 20459 26608 20468 26648
rect 12844 26524 12884 26564
rect 17356 26524 17396 26564
rect 18508 26524 18548 26564
rect 12126 26440 12494 26480
rect 18988 26440 19028 26480
rect 12652 26356 12692 26396
rect 24748 26692 24788 26732
rect 26284 26692 26324 26732
rect 30700 26692 30740 26732
rect 23596 26608 23636 26648
rect 24556 26608 24596 26648
rect 25804 26608 25844 26648
rect 28300 26608 28340 26648
rect 29164 26608 29204 26648
rect 30028 26608 30068 26648
rect 19900 26440 20268 26480
rect 5068 26272 5108 26312
rect 8140 26272 8180 26312
rect 11116 26272 11156 26312
rect 14668 26272 14708 26312
rect 16300 26272 16340 26312
rect 2476 26188 2516 26228
rect 2956 26188 2996 26228
rect 5548 26188 5588 26228
rect 6508 26188 6539 26228
rect 6539 26188 6548 26228
rect 9580 26188 9620 26228
rect 19084 26272 19124 26312
rect 12844 26188 12884 26228
rect 13324 26188 13364 26228
rect 13516 26188 13556 26228
rect 13900 26188 13931 26228
rect 13931 26188 13940 26228
rect 16972 26188 17012 26228
rect 18412 26188 18452 26228
rect 18892 26188 18932 26228
rect 31084 26608 31124 26648
rect 28204 26524 28244 26564
rect 27674 26440 28042 26480
rect 23884 26356 23924 26396
rect 22636 26272 22676 26312
rect 25516 26272 25547 26312
rect 25547 26272 25556 26312
rect 25228 26188 25268 26228
rect 25420 26188 25460 26228
rect 30124 26356 30164 26396
rect 25996 26272 26036 26312
rect 27820 26272 27860 26312
rect 26188 26188 26228 26228
rect 2860 26135 2900 26144
rect 2860 26104 2891 26135
rect 2891 26104 2900 26135
rect 3340 26104 3380 26144
rect 4012 26104 4052 26144
rect 4780 26104 4820 26144
rect 5164 26104 5204 26144
rect 6892 26104 6923 26144
rect 6923 26104 6932 26144
rect 9388 26104 9419 26144
rect 9419 26104 9428 26144
rect 12460 26104 12500 26144
rect 2188 26020 2228 26060
rect 2476 26020 2516 26060
rect 5356 26020 5396 26060
rect 5740 26020 5780 26060
rect 1132 25936 1172 25976
rect 1516 25936 1556 25976
rect 1900 25936 1940 25976
rect 5260 25936 5300 25976
rect 13420 26104 13449 26144
rect 13449 26104 13460 26144
rect 13804 26104 13844 26144
rect 15340 26104 15380 26144
rect 19084 26104 19124 26144
rect 20812 26104 20852 26144
rect 22348 26104 22388 26144
rect 24364 26104 24404 26144
rect 25036 26135 25076 26144
rect 6796 26020 6836 26060
rect 8236 26020 8276 26060
rect 11404 26020 11444 26060
rect 11788 25936 11828 25976
rect 14860 26020 14900 26060
rect 18220 26020 18260 26060
rect 18508 26020 18548 26060
rect 25036 26104 25067 26135
rect 25067 26104 25076 26135
rect 25708 26104 25748 26144
rect 26764 26104 26804 26144
rect 27340 26104 27380 26144
rect 30604 26272 30644 26312
rect 28780 26188 28820 26228
rect 29356 26188 29396 26228
rect 19756 26020 19796 26060
rect 20140 26020 20180 26060
rect 24844 26020 24884 26060
rect 25900 26020 25940 26060
rect 26380 26020 26420 26060
rect 28972 26020 29012 26060
rect 29164 26020 29204 26060
rect 13804 25936 13844 25976
rect 17548 25936 17588 25976
rect 18412 25936 18452 25976
rect 19468 25936 19508 25976
rect 21388 25936 21428 25976
rect 24076 25936 24116 25976
rect 26956 25936 26996 25976
rect 28108 25936 28148 25976
rect 3052 25852 3092 25892
rect 5452 25852 5492 25892
rect 5932 25852 5972 25892
rect 8332 25852 8372 25892
rect 8620 25852 8660 25892
rect 12652 25852 12692 25892
rect 22828 25852 22868 25892
rect 23788 25852 23828 25892
rect 30892 25852 30932 25892
rect 2860 25768 2900 25808
rect 6892 25768 6932 25808
rect 15244 25768 15284 25808
rect 17644 25768 17684 25808
rect 844 25348 884 25388
rect 1228 25348 1268 25388
rect 3112 25684 3480 25724
rect 3724 25684 3764 25724
rect 7564 25684 7604 25724
rect 9004 25684 9044 25724
rect 10886 25684 11254 25724
rect 18660 25684 19028 25724
rect 21292 25684 21332 25724
rect 26092 25684 26132 25724
rect 26434 25684 26802 25724
rect 7468 25600 7508 25640
rect 16876 25600 16916 25640
rect 18124 25600 18164 25640
rect 21772 25600 21812 25640
rect 23884 25600 23924 25640
rect 8140 25516 8180 25556
rect 11692 25516 11732 25556
rect 1612 25432 1652 25472
rect 5452 25432 5492 25472
rect 10060 25432 10100 25472
rect 10636 25432 10676 25472
rect 11788 25432 11828 25472
rect 16108 25516 16148 25556
rect 21580 25516 21620 25556
rect 23980 25516 24020 25556
rect 14188 25432 14228 25472
rect 19084 25432 19124 25472
rect 25228 25432 25268 25472
rect 2572 25348 2612 25388
rect 3244 25348 3284 25388
rect 5260 25348 5300 25388
rect 5644 25348 5684 25388
rect 6988 25348 7028 25388
rect 7180 25348 7220 25388
rect 9100 25348 9140 25388
rect 10732 25348 10772 25388
rect 12556 25348 12596 25388
rect 13324 25348 13364 25388
rect 13804 25348 13844 25388
rect 14668 25348 14708 25388
rect 16108 25348 16148 25388
rect 17548 25348 17588 25388
rect 2380 25264 2420 25304
rect 2956 25264 2996 25304
rect 5740 25264 5780 25304
rect 5932 25295 5972 25304
rect 5932 25264 5972 25295
rect 6508 25264 6548 25304
rect 6892 25264 6932 25304
rect 8332 25264 8344 25304
rect 8344 25264 8372 25304
rect 9292 25264 9332 25304
rect 10444 25264 10484 25304
rect 10828 25264 10867 25304
rect 10867 25264 10868 25304
rect 11404 25264 11444 25304
rect 11692 25264 11732 25304
rect 25708 25463 25748 25472
rect 25708 25432 25716 25463
rect 25716 25432 25748 25463
rect 26956 25432 26996 25472
rect 21772 25348 21812 25388
rect 23692 25348 23732 25388
rect 26284 25348 26324 25388
rect 26860 25348 26900 25388
rect 13228 25264 13256 25304
rect 13256 25264 13268 25304
rect 14860 25264 14879 25304
rect 14879 25264 14900 25304
rect 15148 25264 15188 25304
rect 16204 25264 16244 25304
rect 17068 25264 17108 25304
rect 18988 25264 19028 25304
rect 21484 25264 21524 25304
rect 21676 25264 21716 25304
rect 22348 25264 22388 25304
rect 25420 25264 25445 25304
rect 25445 25264 25460 25304
rect 1324 25180 1364 25220
rect 1612 25180 1652 25220
rect 652 25096 692 25136
rect 1996 25096 2027 25136
rect 2027 25096 2036 25136
rect 3148 25096 3188 25136
rect 5452 25180 5492 25220
rect 8524 25180 8564 25220
rect 5356 25096 5396 25136
rect 11020 25096 11060 25136
rect 2284 25012 2324 25052
rect 11404 25012 11444 25052
rect 12172 25180 12212 25220
rect 12460 25180 12491 25220
rect 12491 25180 12500 25220
rect 12748 25180 12788 25220
rect 13036 25180 13076 25220
rect 17260 25180 17300 25220
rect 18508 25180 18548 25220
rect 20620 25180 20660 25220
rect 21868 25180 21908 25220
rect 22924 25180 22964 25220
rect 12844 25096 12884 25136
rect 14380 25096 14420 25136
rect 15340 25096 15380 25136
rect 19660 25096 19700 25136
rect 20716 25096 20756 25136
rect 22732 25096 22772 25136
rect 11596 25012 11636 25052
rect 4352 24928 4720 24968
rect 8812 24928 8852 24968
rect 12126 24928 12494 24968
rect 10444 24844 10484 24884
rect 10636 24844 10676 24884
rect 11020 24844 11060 24884
rect 1708 24760 1748 24800
rect 11308 24760 11348 24800
rect 13900 24760 13940 24800
rect 4588 24676 4628 24716
rect 7468 24676 7508 24716
rect 15244 25012 15284 25052
rect 23788 25012 23828 25052
rect 19372 24928 19412 24968
rect 19900 24928 20268 24968
rect 17548 24844 17588 24884
rect 20620 24844 20660 24884
rect 16204 24760 16244 24800
rect 19852 24760 19883 24800
rect 19883 24760 19892 24800
rect 20524 24760 20555 24800
rect 20555 24760 20564 24800
rect 21676 24760 21716 24800
rect 21868 24760 21908 24800
rect 23116 24760 23147 24800
rect 23147 24760 23156 24800
rect 23788 24760 23828 24800
rect 9388 24676 9428 24716
rect 9772 24676 9812 24716
rect 13324 24676 13364 24716
rect 13516 24707 13556 24716
rect 13516 24676 13547 24707
rect 13547 24676 13556 24707
rect 13996 24676 14036 24716
rect 14764 24676 14804 24716
rect 17068 24676 17108 24716
rect 25420 25096 25460 25136
rect 25708 25096 25748 25136
rect 25996 25012 26036 25052
rect 27052 25348 27092 25388
rect 27628 25348 27668 25388
rect 27244 25264 27284 25304
rect 28876 25264 28916 25304
rect 29932 25264 29972 25304
rect 26380 25180 26420 25220
rect 26668 25180 26708 25220
rect 27052 25180 27092 25220
rect 28108 25180 28148 25220
rect 28588 25180 28628 25220
rect 26476 25096 26516 25136
rect 27340 25096 27380 25136
rect 29836 25096 29876 25136
rect 18988 24676 19028 24716
rect 2284 24592 2315 24632
rect 2315 24592 2324 24632
rect 2764 24592 2804 24632
rect 4108 24592 4148 24632
rect 5740 24592 5780 24632
rect 8524 24592 8564 24632
rect 9292 24592 9332 24632
rect 9484 24592 9509 24632
rect 9509 24592 9524 24632
rect 14188 24623 14228 24632
rect 14188 24592 14219 24623
rect 14219 24592 14228 24623
rect 14956 24592 14957 24632
rect 14957 24592 14996 24632
rect 15820 24592 15860 24632
rect 21580 24676 21620 24716
rect 23308 24676 23348 24716
rect 26764 24928 26804 24968
rect 28300 25012 28340 25052
rect 30028 25012 30068 25052
rect 27674 24928 28042 24968
rect 28108 24928 28148 24968
rect 30412 24928 30452 24968
rect 31468 24928 31508 24968
rect 24652 24844 24692 24884
rect 25324 24760 25364 24800
rect 28684 24844 28724 24884
rect 30796 24844 30836 24884
rect 24268 24676 24308 24716
rect 24844 24676 24884 24716
rect 25516 24676 25556 24716
rect 26092 24760 26132 24800
rect 26668 24760 26708 24800
rect 28012 24760 28052 24800
rect 28492 24760 28532 24800
rect 28876 24760 28916 24800
rect 30028 24760 30068 24800
rect 18508 24623 18548 24632
rect 1036 24508 1076 24548
rect 8716 24508 8756 24548
rect 9004 24508 9044 24548
rect 10060 24508 10100 24548
rect 13132 24508 13172 24548
rect 13612 24508 13652 24548
rect 14476 24508 14516 24548
rect 17740 24508 17780 24548
rect 18508 24592 18539 24623
rect 18539 24592 18548 24623
rect 19468 24592 19493 24632
rect 19493 24592 19508 24632
rect 20428 24592 20468 24632
rect 21292 24592 21304 24632
rect 21304 24592 21332 24632
rect 18604 24508 18644 24548
rect 19756 24508 19796 24548
rect 21004 24508 21044 24548
rect 21964 24508 22004 24548
rect 23116 24592 23156 24632
rect 23884 24592 23896 24632
rect 23896 24592 23924 24632
rect 24460 24592 24500 24632
rect 26188 24676 26228 24716
rect 26956 24676 26996 24716
rect 27532 24676 27572 24716
rect 28300 24676 28340 24716
rect 29836 24676 29876 24716
rect 25708 24592 25748 24632
rect 26380 24592 26409 24632
rect 26409 24592 26420 24632
rect 27820 24592 27860 24632
rect 29356 24592 29387 24632
rect 29387 24592 29396 24632
rect 22732 24508 22772 24548
rect 23020 24508 23060 24548
rect 23980 24508 24020 24548
rect 24172 24508 24212 24548
rect 24844 24508 24884 24548
rect 26860 24508 26900 24548
rect 27052 24508 27092 24548
rect 27340 24508 27380 24548
rect 28684 24508 28724 24548
rect 28972 24508 29012 24548
rect 29740 24508 29780 24548
rect 11788 24424 11828 24464
rect 12556 24424 12596 24464
rect 13516 24424 13556 24464
rect 15148 24424 15188 24464
rect 18220 24424 18260 24464
rect 20236 24424 20276 24464
rect 21292 24424 21332 24464
rect 21676 24424 21716 24464
rect 22828 24424 22868 24464
rect 23308 24424 23348 24464
rect 26092 24424 26132 24464
rect 26764 24424 26804 24464
rect 28396 24424 28436 24464
rect 364 24340 404 24380
rect 4972 24340 5012 24380
rect 7660 24340 7700 24380
rect 8428 24340 8468 24380
rect 10444 24340 10484 24380
rect 12172 24340 12212 24380
rect 13996 24340 14036 24380
rect 21484 24340 21524 24380
rect 21772 24340 21812 24380
rect 22444 24340 22484 24380
rect 25996 24340 26036 24380
rect 28972 24340 29012 24380
rect 10540 24256 10580 24296
rect 19468 24256 19508 24296
rect 23116 24256 23156 24296
rect 27628 24256 27668 24296
rect 3112 24172 3480 24212
rect 6028 24172 6068 24212
rect 10886 24172 11254 24212
rect 13324 24172 13364 24212
rect 14188 24172 14228 24212
rect 15724 24172 15764 24212
rect 16204 24172 16244 24212
rect 18660 24172 19028 24212
rect 19180 24172 19220 24212
rect 25036 24172 25076 24212
rect 26434 24172 26802 24212
rect 1228 24088 1268 24128
rect 5548 24088 5588 24128
rect 5740 24088 5780 24128
rect 21868 24088 21908 24128
rect 28588 24088 28628 24128
rect 2380 24004 2420 24044
rect 4588 24004 4628 24044
rect 8620 24004 8660 24044
rect 9964 24004 10004 24044
rect 13228 24004 13268 24044
rect 14668 24004 14708 24044
rect 16396 24004 16436 24044
rect 23308 24004 23348 24044
rect 24460 24004 24500 24044
rect 10540 23920 10580 23960
rect 12748 23920 12788 23960
rect 13420 23920 13460 23960
rect 1516 23836 1556 23876
rect 3244 23836 3284 23876
rect 2284 23752 2324 23792
rect 3820 23752 3860 23792
rect 7372 23836 7412 23876
rect 9100 23836 9140 23876
rect 10156 23836 10196 23876
rect 10444 23836 10484 23876
rect 13132 23836 13172 23876
rect 17260 23920 17300 23960
rect 19948 23920 19988 23960
rect 22156 23920 22196 23960
rect 24364 23920 24404 23960
rect 14188 23836 14228 23876
rect 16012 23836 16052 23876
rect 16684 23836 16724 23876
rect 20236 23836 20276 23876
rect 21484 23836 21524 23876
rect 23212 23836 23252 23876
rect 23500 23836 23540 23876
rect 23980 23836 24020 23876
rect 24172 23836 24212 23876
rect 4972 23783 5012 23792
rect 4972 23752 5012 23783
rect 5260 23752 5300 23792
rect 5740 23752 5780 23792
rect 6028 23752 6068 23792
rect 7660 23752 7700 23792
rect 8620 23752 8660 23792
rect 9292 23752 9332 23792
rect 9676 23752 9716 23792
rect 11308 23752 11348 23792
rect 12172 23752 12212 23792
rect 12556 23752 12596 23792
rect 15340 23752 15371 23792
rect 15371 23752 15380 23792
rect 17260 23752 17300 23792
rect 17740 23752 17780 23792
rect 19180 23752 19220 23792
rect 19660 23752 19700 23792
rect 19852 23752 19892 23792
rect 20524 23752 20564 23792
rect 21676 23752 21716 23792
rect 21964 23752 22004 23792
rect 22828 23752 22857 23792
rect 22857 23752 22868 23792
rect 23308 23752 23348 23792
rect 1612 23668 1652 23708
rect 1996 23668 2036 23708
rect 5932 23668 5972 23708
rect 7180 23668 7220 23708
rect 7852 23668 7892 23708
rect 8044 23668 8084 23708
rect 1420 23332 1460 23372
rect 6700 23584 6740 23624
rect 7276 23584 7316 23624
rect 8236 23584 8276 23624
rect 6124 23500 6164 23540
rect 9196 23668 9236 23708
rect 7564 23500 7604 23540
rect 8812 23500 8852 23540
rect 10060 23668 10100 23708
rect 4352 23416 4720 23456
rect 9484 23416 9524 23456
rect 5740 23332 5780 23372
rect 10636 23668 10676 23708
rect 11020 23668 11060 23708
rect 13324 23668 13364 23708
rect 14668 23668 14708 23708
rect 20908 23668 20948 23708
rect 22156 23668 22196 23708
rect 22444 23668 22484 23708
rect 23212 23668 23251 23708
rect 23251 23668 23252 23708
rect 25420 24004 25460 24044
rect 27340 24004 27380 24044
rect 25324 23920 25364 23960
rect 25516 23920 25556 23960
rect 24748 23836 24788 23876
rect 25228 23836 25268 23876
rect 26764 23836 26804 23876
rect 28972 23836 29012 23876
rect 30220 23836 30260 23876
rect 23980 23668 24020 23708
rect 25324 23752 25364 23792
rect 26476 23752 26507 23792
rect 26507 23752 26516 23792
rect 26668 23752 26708 23792
rect 27052 23752 27092 23792
rect 28204 23752 28244 23792
rect 28876 23752 28916 23792
rect 29068 23752 29108 23792
rect 29260 23752 29300 23792
rect 25420 23668 25460 23708
rect 27340 23668 27380 23708
rect 27628 23668 27668 23708
rect 29548 23668 29588 23708
rect 11596 23584 11636 23624
rect 13708 23584 13748 23624
rect 17644 23584 17684 23624
rect 18220 23584 18260 23624
rect 19948 23584 19988 23624
rect 20428 23584 20468 23624
rect 20620 23584 20651 23624
rect 20651 23584 20660 23624
rect 22924 23584 22964 23624
rect 23500 23584 23540 23624
rect 24364 23584 24404 23624
rect 25516 23584 25556 23624
rect 25804 23584 25844 23624
rect 26284 23584 26324 23624
rect 26668 23584 26708 23624
rect 27436 23584 27476 23624
rect 27724 23584 27764 23624
rect 29932 23584 29972 23624
rect 31180 23584 31220 23624
rect 11692 23500 11732 23540
rect 12844 23500 12884 23540
rect 24460 23500 24500 23540
rect 10444 23416 10484 23456
rect 11500 23416 11540 23456
rect 12126 23416 12494 23456
rect 19468 23416 19508 23456
rect 19900 23416 20268 23456
rect 24748 23416 24788 23456
rect 10636 23332 10676 23372
rect 2380 23248 2420 23288
rect 3820 23248 3860 23288
rect 4492 23248 4532 23288
rect 5548 23248 5588 23288
rect 7468 23248 7508 23288
rect 8140 23248 8180 23288
rect 940 23164 980 23204
rect 2668 23164 2708 23204
rect 3244 23164 3284 23204
rect 5068 23164 5108 23204
rect 5644 23164 5684 23204
rect 7564 23164 7604 23204
rect 9004 23164 9044 23204
rect 9676 23164 9716 23204
rect 10252 23164 10292 23204
rect 1612 23080 1643 23120
rect 1643 23080 1652 23120
rect 2092 23080 2121 23120
rect 2121 23080 2132 23120
rect 2284 23080 2324 23120
rect 1036 22912 1067 22952
rect 1067 22912 1076 22952
rect 11116 23248 11156 23288
rect 11788 23248 11828 23288
rect 13132 23248 13172 23288
rect 10732 23164 10772 23204
rect 11404 23164 11444 23204
rect 11884 23164 11924 23204
rect 27674 23416 28042 23456
rect 14380 23248 14420 23288
rect 15244 23332 15284 23372
rect 15724 23332 15764 23372
rect 20524 23332 20564 23372
rect 23308 23332 23348 23372
rect 24364 23332 24404 23372
rect 29932 23332 29972 23372
rect 31180 23332 31220 23372
rect 13516 23164 13556 23204
rect 13804 23164 13844 23204
rect 13996 23164 14036 23204
rect 14668 23164 14708 23204
rect 4108 23080 4148 23120
rect 4396 23080 4436 23120
rect 1900 22996 1940 23036
rect 2188 22996 2228 23036
rect 4204 22996 4244 23036
rect 5164 23080 5204 23120
rect 5452 23080 5492 23120
rect 5740 23080 5780 23120
rect 7468 23080 7508 23120
rect 8236 23080 8276 23120
rect 8908 23080 8948 23120
rect 12844 23080 12884 23120
rect 14188 23080 14228 23120
rect 17836 23248 17876 23288
rect 18220 23248 18251 23288
rect 18251 23248 18260 23288
rect 18508 23248 18548 23288
rect 19180 23248 19220 23288
rect 20236 23248 20276 23288
rect 21292 23248 21332 23288
rect 21772 23248 21812 23288
rect 16204 23164 16244 23204
rect 16684 23164 16715 23204
rect 16715 23164 16724 23204
rect 17260 23164 17300 23204
rect 19660 23164 19700 23204
rect 20428 23164 20468 23204
rect 22156 23164 22196 23204
rect 22348 23164 22388 23204
rect 23212 23164 23252 23204
rect 25036 23164 25076 23204
rect 26188 23164 26228 23204
rect 26956 23164 26996 23204
rect 27148 23164 27188 23204
rect 5260 22996 5283 23036
rect 5283 22996 5300 23036
rect 5836 22996 5876 23036
rect 10252 22996 10292 23036
rect 3436 22912 3476 22952
rect 8524 22912 8555 22952
rect 8555 22912 8564 22952
rect 8812 22912 8852 22952
rect 10540 22996 10580 23036
rect 10828 22996 10868 23036
rect 11308 22996 11348 23036
rect 10636 22912 10676 22952
rect 11788 22996 11828 23036
rect 1708 22828 1748 22868
rect 2956 22828 2996 22868
rect 7948 22828 7988 22868
rect 8716 22828 8756 22868
rect 8908 22828 8948 22868
rect 10060 22828 10100 22868
rect 10828 22828 10868 22868
rect 17452 23080 17492 23120
rect 17740 23080 17780 23120
rect 18028 23080 18068 23120
rect 19564 23080 19604 23120
rect 19756 23080 19796 23120
rect 21292 23080 21332 23120
rect 12076 22996 12116 23036
rect 12268 22996 12308 23036
rect 13612 22996 13652 23036
rect 14380 22996 14403 23036
rect 14403 22996 14420 23036
rect 13996 22912 14027 22952
rect 14027 22912 14036 22952
rect 15436 22996 15476 23036
rect 18220 22996 18260 23036
rect 12364 22828 12404 22868
rect 13036 22828 13076 22868
rect 13324 22828 13364 22868
rect 14092 22828 14132 22868
rect 21484 23080 21515 23120
rect 21515 23080 21524 23120
rect 22060 23080 22100 23120
rect 25132 23080 25172 23120
rect 25324 23080 25364 23120
rect 25516 23080 25547 23120
rect 25547 23080 25556 23120
rect 21772 22996 21812 23036
rect 22156 22996 22196 23036
rect 16012 22912 16052 22952
rect 18316 22912 18356 22952
rect 19276 22912 19316 22952
rect 20908 22912 20948 22952
rect 18220 22828 18260 22868
rect 20716 22828 20756 22868
rect 2572 22744 2612 22784
rect 7756 22744 7796 22784
rect 10444 22744 10484 22784
rect 11788 22744 11828 22784
rect 12172 22744 12212 22784
rect 22540 22744 22580 22784
rect 1036 22660 1076 22700
rect 2764 22660 2804 22700
rect 3112 22660 3480 22700
rect 7852 22660 7892 22700
rect 10886 22660 11254 22700
rect 8428 22576 8468 22616
rect 460 22492 500 22532
rect 6124 22492 6164 22532
rect 6316 22492 6356 22532
rect 7180 22492 7220 22532
rect 7948 22492 7988 22532
rect 8524 22492 8564 22532
rect 9676 22492 9716 22532
rect 10636 22492 10676 22532
rect 11308 22492 11348 22532
rect 11692 22492 11732 22532
rect 2092 22408 2132 22448
rect 4300 22408 4340 22448
rect 4780 22408 4820 22448
rect 5452 22408 5492 22448
rect 556 22324 596 22364
rect 1228 22324 1268 22364
rect 2188 22324 2228 22364
rect 3532 22324 3572 22364
rect 3916 22324 3956 22364
rect 4396 22324 4436 22364
rect 5068 22324 5108 22364
rect 5548 22324 5588 22364
rect 5836 22324 5876 22364
rect 6796 22324 6836 22364
rect 1708 22240 1748 22280
rect 2092 22240 2132 22280
rect 268 22156 308 22196
rect 1420 22156 1460 22196
rect 1324 22072 1364 22112
rect 2284 22072 2324 22112
rect 3436 22240 3476 22280
rect 3724 22240 3764 22280
rect 4972 22240 5012 22280
rect 5452 22240 5492 22280
rect 5740 22240 5780 22280
rect 2668 22156 2708 22196
rect 3340 22156 3380 22196
rect 4204 22156 4244 22196
rect 4876 22156 4916 22196
rect 3148 22072 3179 22112
rect 3179 22072 3188 22112
rect 460 21988 500 22028
rect 1036 21988 1076 22028
rect 1612 21988 1652 22028
rect 7852 22408 7892 22448
rect 8428 22408 8468 22448
rect 10252 22408 10292 22448
rect 7564 22324 7604 22364
rect 24652 22996 24692 23036
rect 28588 23164 28628 23204
rect 26092 23080 26108 23120
rect 26108 23080 26132 23120
rect 26380 23080 26420 23120
rect 27436 23080 27476 23120
rect 27244 22996 27284 23036
rect 27628 22996 27668 23036
rect 27820 22996 27859 23036
rect 27859 22996 27860 23036
rect 28204 22996 28244 23036
rect 29164 23080 29204 23120
rect 29548 23080 29588 23120
rect 30316 23080 30356 23120
rect 31084 23080 31124 23120
rect 25516 22912 25556 22952
rect 26284 22912 26324 22952
rect 27148 22912 27188 22952
rect 27916 22828 27956 22868
rect 31276 22828 31316 22868
rect 27628 22744 27668 22784
rect 18660 22660 19028 22700
rect 19276 22660 19316 22700
rect 26434 22660 26802 22700
rect 14764 22576 14804 22616
rect 16876 22576 16916 22616
rect 22060 22576 22100 22616
rect 23020 22576 23060 22616
rect 26860 22576 26900 22616
rect 30124 22576 30164 22616
rect 17452 22492 17492 22532
rect 21772 22492 21812 22532
rect 22156 22492 22196 22532
rect 23692 22492 23732 22532
rect 24268 22492 24308 22532
rect 25708 22492 25748 22532
rect 26284 22492 26324 22532
rect 27724 22492 27764 22532
rect 10444 22408 10484 22448
rect 7660 22240 7700 22280
rect 8524 22240 8564 22280
rect 9964 22240 10004 22280
rect 10636 22240 10676 22280
rect 12268 22408 12308 22448
rect 18124 22408 18164 22448
rect 19372 22408 19412 22448
rect 22636 22408 22676 22448
rect 26668 22408 26708 22448
rect 29164 22408 29204 22448
rect 11500 22324 11540 22364
rect 14284 22324 14324 22364
rect 18604 22324 18644 22364
rect 18988 22324 19028 22364
rect 19756 22324 19787 22364
rect 19787 22324 19796 22364
rect 21676 22324 21716 22364
rect 11596 22240 11636 22280
rect 11980 22240 12020 22280
rect 12940 22240 12980 22280
rect 13708 22240 13748 22280
rect 14092 22240 14132 22280
rect 15148 22240 15188 22280
rect 15532 22240 15572 22280
rect 15916 22240 15956 22280
rect 17068 22240 17108 22280
rect 18028 22240 18068 22280
rect 18508 22240 18548 22280
rect 20908 22240 20948 22280
rect 22060 22240 22100 22280
rect 22732 22324 22763 22364
rect 22763 22324 22772 22364
rect 23116 22324 23156 22364
rect 23404 22324 23444 22364
rect 25804 22324 25844 22364
rect 26092 22324 26132 22364
rect 22828 22240 22868 22280
rect 23308 22240 23348 22280
rect 23788 22240 23828 22280
rect 6124 22156 6164 22196
rect 6412 22156 6452 22196
rect 6604 22156 6644 22196
rect 7468 22156 7508 22196
rect 9676 22156 9716 22196
rect 10156 22156 10196 22196
rect 10444 22156 10484 22196
rect 13804 22156 13844 22196
rect 16108 22156 16148 22196
rect 18316 22156 18356 22196
rect 19180 22156 19220 22196
rect 21196 22156 21236 22196
rect 22252 22156 22292 22196
rect 5740 22072 5780 22112
rect 8044 22072 8075 22112
rect 8075 22072 8084 22112
rect 8236 22072 8276 22112
rect 10060 22072 10100 22112
rect 10252 22072 10292 22112
rect 12748 22072 12779 22112
rect 12779 22072 12788 22112
rect 13708 22072 13748 22112
rect 18220 22072 18260 22112
rect 18988 22072 19028 22112
rect 20332 22072 20372 22112
rect 20812 22072 20852 22112
rect 22540 22072 22580 22112
rect 7084 21988 7124 22028
rect 10348 21988 10388 22028
rect 28588 22324 28628 22364
rect 30412 22324 30452 22364
rect 31276 22324 31307 22364
rect 31307 22324 31316 22364
rect 23212 22156 23252 22196
rect 25036 22240 25076 22280
rect 25420 22240 25427 22280
rect 25427 22240 25460 22280
rect 25708 22240 25748 22280
rect 27724 22240 27764 22280
rect 27916 22240 27956 22280
rect 28204 22240 28244 22280
rect 28684 22240 28696 22280
rect 28696 22240 28724 22280
rect 29452 22240 29492 22280
rect 24364 22156 24404 22196
rect 24460 22072 24500 22112
rect 21484 21988 21524 22028
rect 25132 22156 25172 22196
rect 25516 22156 25556 22196
rect 25804 22156 25844 22196
rect 23788 21988 23828 22028
rect 26092 22072 26132 22112
rect 26380 22156 26420 22196
rect 26668 22156 26708 22196
rect 26860 22156 26900 22196
rect 29356 22156 29396 22196
rect 26284 22072 26324 22112
rect 27436 22072 27476 22112
rect 29260 21988 29300 22028
rect 4352 21904 4720 21944
rect 7564 21904 7604 21944
rect 8812 21904 8852 21944
rect 12126 21904 12494 21944
rect 19900 21904 20268 21944
rect 24364 21904 24404 21944
rect 25132 21904 25172 21944
rect 26860 21904 26900 21944
rect 27674 21904 28042 21944
rect 3148 21820 3188 21860
rect 3340 21820 3380 21860
rect 1612 21736 1652 21776
rect 1996 21736 2036 21776
rect 3532 21736 3572 21776
rect 4972 21736 5012 21776
rect 2188 21652 2228 21692
rect 3436 21652 3476 21692
rect 4492 21652 4532 21692
rect 6604 21820 6644 21860
rect 9868 21820 9908 21860
rect 13612 21820 13652 21860
rect 17260 21820 17300 21860
rect 22060 21820 22100 21860
rect 23308 21820 23348 21860
rect 25708 21820 25748 21860
rect 27148 21820 27188 21860
rect 6028 21736 6068 21776
rect 6316 21736 6356 21776
rect 7660 21736 7700 21776
rect 9580 21736 9620 21776
rect 1516 21568 1556 21575
rect 1516 21535 1556 21568
rect 1804 21568 1843 21608
rect 1843 21568 1844 21608
rect 3052 21568 3092 21608
rect 460 21484 500 21524
rect 1324 21484 1364 21524
rect 1420 21400 1460 21440
rect 1612 21400 1652 21440
rect 3532 21568 3572 21608
rect 3916 21568 3956 21608
rect 4876 21568 4916 21608
rect 5452 21568 5492 21608
rect 3244 21484 3284 21524
rect 4108 21484 4148 21524
rect 4780 21484 4820 21524
rect 4972 21484 5012 21524
rect 5548 21484 5588 21524
rect 10444 21736 10475 21776
rect 10475 21736 10484 21776
rect 10924 21736 10964 21776
rect 12940 21736 12980 21776
rect 13708 21736 13748 21776
rect 15148 21736 15188 21776
rect 18028 21736 18068 21776
rect 18604 21736 18644 21776
rect 20908 21736 20948 21776
rect 7468 21652 7508 21692
rect 8236 21652 8276 21692
rect 10156 21652 10196 21692
rect 11788 21652 11828 21692
rect 11980 21652 12020 21692
rect 15532 21652 15572 21692
rect 16012 21652 16052 21692
rect 19276 21652 19316 21692
rect 6316 21568 6356 21608
rect 6604 21568 6629 21608
rect 6629 21568 6644 21608
rect 6988 21568 7028 21608
rect 8428 21568 8468 21608
rect 10732 21568 10772 21608
rect 11045 21568 11085 21608
rect 11596 21599 11636 21608
rect 11596 21568 11627 21599
rect 11627 21568 11636 21599
rect 11884 21568 11924 21608
rect 12652 21568 12683 21608
rect 12683 21568 12692 21608
rect 13516 21568 13556 21608
rect 14188 21568 14228 21608
rect 14476 21568 14507 21608
rect 14507 21568 14516 21608
rect 15052 21568 15092 21608
rect 6796 21484 6836 21524
rect 5740 21400 5780 21440
rect 6988 21400 7028 21440
rect 7564 21484 7604 21524
rect 8044 21484 8084 21524
rect 9388 21484 9428 21524
rect 7276 21400 7316 21440
rect 8236 21400 8276 21440
rect 4780 21232 4820 21272
rect 8428 21232 8468 21272
rect 2956 21148 2996 21188
rect 3112 21148 3480 21188
rect 7948 21148 7988 21188
rect 21772 21652 21812 21692
rect 22732 21736 22772 21776
rect 23692 21736 23732 21776
rect 24556 21736 24596 21776
rect 25420 21736 25460 21776
rect 26668 21736 26708 21776
rect 26860 21736 26900 21776
rect 28108 21736 28148 21776
rect 29452 21736 29492 21776
rect 22540 21652 22580 21692
rect 24652 21652 24692 21692
rect 25132 21652 25172 21692
rect 25612 21652 25652 21692
rect 26572 21652 26612 21692
rect 27436 21652 27476 21692
rect 27916 21652 27956 21692
rect 28972 21652 29003 21692
rect 29003 21652 29012 21692
rect 16108 21568 16148 21608
rect 16876 21568 16888 21608
rect 16888 21568 16916 21608
rect 17644 21568 17684 21608
rect 18508 21568 18548 21608
rect 18988 21568 19028 21608
rect 19180 21568 19220 21608
rect 20332 21568 20372 21608
rect 20716 21568 20756 21608
rect 22252 21568 22283 21608
rect 22283 21568 22292 21608
rect 22828 21568 22868 21608
rect 24460 21568 24500 21608
rect 24844 21568 24884 21608
rect 25420 21568 25460 21608
rect 13612 21484 13652 21524
rect 16684 21484 16724 21524
rect 10252 21400 10292 21440
rect 10060 21316 10100 21356
rect 11404 21400 11444 21440
rect 11596 21400 11636 21440
rect 13900 21400 13940 21440
rect 14092 21400 14132 21440
rect 15436 21400 15476 21440
rect 13228 21316 13268 21356
rect 9964 21232 10004 21272
rect 10540 21232 10580 21272
rect 14380 21232 14420 21272
rect 18220 21484 18251 21524
rect 18251 21484 18260 21524
rect 19468 21484 19508 21524
rect 17164 21316 17204 21356
rect 18508 21316 18548 21356
rect 20044 21400 20084 21440
rect 20908 21400 20948 21440
rect 21676 21484 21716 21524
rect 22060 21484 22100 21524
rect 22924 21484 22964 21524
rect 24172 21484 24212 21524
rect 26092 21568 26132 21608
rect 24364 21484 24404 21524
rect 25132 21484 25172 21524
rect 27244 21568 27284 21608
rect 27628 21568 27668 21608
rect 28204 21568 28244 21608
rect 28684 21568 28724 21608
rect 29356 21568 29387 21608
rect 29387 21568 29396 21608
rect 30412 21484 30452 21524
rect 21868 21400 21908 21440
rect 23308 21400 23348 21440
rect 27532 21400 27572 21440
rect 21484 21316 21524 21356
rect 23116 21316 23156 21356
rect 24460 21316 24500 21356
rect 25324 21316 25364 21356
rect 26668 21316 26708 21356
rect 27628 21316 27668 21356
rect 29548 21316 29588 21356
rect 30988 21316 31028 21356
rect 22828 21232 22868 21272
rect 24844 21232 24884 21272
rect 9676 21148 9716 21188
rect 10886 21148 11254 21188
rect 15628 21148 15668 21188
rect 18660 21148 19028 21188
rect 21004 21148 21044 21188
rect 26434 21148 26802 21188
rect 460 20980 500 21020
rect 5068 21064 5108 21104
rect 9100 21064 9140 21104
rect 11596 21064 11636 21104
rect 14860 21064 14900 21104
rect 28684 21064 28724 21104
rect 30316 21064 30356 21104
rect 1228 20980 1268 21020
rect 1420 20980 1460 21020
rect 1420 20812 1460 20852
rect 3244 20896 3284 20936
rect 5548 20980 5588 21020
rect 5068 20896 5108 20936
rect 5740 20896 5780 20936
rect 1900 20812 1940 20852
rect 4396 20812 4436 20852
rect 5164 20812 5204 20852
rect 5548 20812 5588 20852
rect 5836 20812 5876 20852
rect 7372 20980 7412 21020
rect 7948 20980 7988 21020
rect 9196 20980 9236 21020
rect 9388 20980 9428 21020
rect 9676 20980 9716 21020
rect 11884 20980 11924 21020
rect 13900 20980 13940 21020
rect 15436 20980 15476 21020
rect 16972 20980 17012 21020
rect 18892 20980 18932 21020
rect 20428 20980 20468 21020
rect 21292 20980 21332 21020
rect 24556 20980 24596 21020
rect 25804 20980 25844 21020
rect 26860 20980 26900 21020
rect 7276 20896 7316 20936
rect 7564 20896 7604 20936
rect 8236 20896 8276 20936
rect 6220 20812 6260 20852
rect 7468 20812 7508 20852
rect 7660 20812 7700 20852
rect 8620 20812 8660 20852
rect 9580 20812 9620 20852
rect 2188 20728 2228 20768
rect 2572 20728 2574 20768
rect 2574 20728 2612 20768
rect 3532 20728 3572 20768
rect 4012 20728 4052 20768
rect 4588 20728 4628 20768
rect 4972 20728 5003 20768
rect 5003 20728 5012 20768
rect 6796 20728 6836 20768
rect 7276 20728 7316 20768
rect 8236 20728 8276 20768
rect 8524 20728 8564 20768
rect 460 20644 500 20684
rect 2380 20644 2420 20684
rect 2860 20644 2900 20684
rect 5260 20644 5300 20684
rect 6508 20644 6548 20684
rect 7852 20644 7892 20684
rect 1612 20560 1652 20600
rect 1996 20560 2036 20600
rect 2188 20560 2228 20600
rect 2764 20560 2804 20600
rect 3052 20560 3092 20600
rect 3340 20560 3371 20600
rect 3371 20560 3380 20600
rect 3916 20560 3956 20600
rect 4396 20560 4436 20600
rect 5740 20560 5780 20600
rect 6220 20560 6260 20600
rect 6604 20560 6644 20600
rect 8236 20560 8276 20600
rect 9004 20728 9044 20768
rect 9388 20728 9428 20768
rect 15916 20896 15956 20936
rect 14092 20812 14132 20852
rect 14860 20812 14900 20852
rect 11788 20728 11828 20768
rect 12556 20728 12596 20768
rect 12844 20728 12884 20768
rect 13132 20728 13172 20768
rect 13900 20728 13940 20768
rect 19468 20896 19508 20936
rect 21868 20896 21908 20936
rect 27724 20980 27755 21020
rect 27755 20980 27764 21020
rect 28204 20980 28244 21020
rect 25708 20896 25748 20936
rect 17068 20812 17108 20852
rect 17260 20812 17300 20852
rect 18412 20812 18452 20852
rect 18700 20812 18740 20852
rect 19084 20812 19124 20852
rect 19756 20812 19796 20852
rect 21580 20812 21620 20852
rect 21964 20812 22004 20852
rect 24172 20812 24212 20852
rect 25324 20812 25355 20852
rect 25355 20812 25364 20852
rect 25612 20812 25652 20852
rect 28300 20812 28340 20852
rect 29356 20812 29396 20852
rect 14572 20728 14612 20768
rect 15628 20728 15668 20768
rect 16396 20728 16436 20768
rect 17164 20728 17204 20768
rect 18220 20728 18251 20768
rect 18251 20728 18260 20768
rect 18508 20728 18522 20768
rect 18522 20728 18548 20768
rect 20620 20728 20660 20768
rect 20812 20728 20852 20768
rect 22156 20728 22196 20768
rect 23116 20728 23147 20768
rect 23147 20728 23156 20768
rect 26380 20728 26420 20768
rect 26860 20728 26900 20768
rect 11884 20644 11924 20684
rect 12940 20644 12980 20684
rect 13612 20644 13652 20684
rect 14668 20644 14708 20684
rect 15916 20644 15956 20684
rect 16972 20644 17012 20684
rect 17740 20644 17780 20684
rect 9388 20560 9428 20600
rect 11404 20560 11444 20600
rect 15148 20560 15179 20600
rect 15179 20560 15188 20600
rect 15628 20560 15668 20600
rect 16012 20560 16052 20600
rect 18028 20560 18059 20600
rect 18059 20560 18068 20600
rect 18316 20560 18347 20600
rect 18347 20560 18356 20600
rect 19084 20560 19124 20600
rect 940 20476 980 20516
rect 7948 20476 7988 20516
rect 9196 20476 9236 20516
rect 10252 20476 10292 20516
rect 19372 20644 19412 20684
rect 19756 20644 19796 20684
rect 19468 20560 19508 20600
rect 20044 20560 20084 20600
rect 21004 20644 21044 20684
rect 24172 20644 24212 20684
rect 25132 20644 25172 20684
rect 26572 20644 26612 20684
rect 27244 20644 27284 20684
rect 23596 20560 23636 20600
rect 25324 20560 25364 20600
rect 25612 20560 25652 20600
rect 26860 20560 26900 20600
rect 16876 20476 16916 20516
rect 18412 20476 18452 20516
rect 23404 20476 23444 20516
rect 25708 20476 25748 20516
rect 27916 20728 27956 20768
rect 28972 20728 29012 20768
rect 30508 20728 30548 20768
rect 30796 20728 30836 20768
rect 28204 20644 28244 20684
rect 28492 20644 28532 20684
rect 31660 20644 31700 20684
rect 28684 20560 28724 20600
rect 27244 20476 27284 20516
rect 4352 20392 4720 20432
rect 8428 20392 8468 20432
rect 11884 20392 11924 20432
rect 12126 20392 12494 20432
rect 14476 20392 14516 20432
rect 18700 20392 18740 20432
rect 1804 20308 1844 20348
rect 3052 20308 3092 20348
rect 6028 20308 6068 20348
rect 9676 20308 9716 20348
rect 11404 20308 11444 20348
rect 2572 20224 2612 20264
rect 3244 20224 3275 20264
rect 3275 20224 3284 20264
rect 5164 20224 5204 20264
rect 5356 20224 5396 20264
rect 5836 20224 5876 20264
rect 6604 20224 6644 20264
rect 6796 20224 6836 20264
rect 11788 20224 11828 20264
rect 12556 20224 12596 20264
rect 12844 20224 12884 20264
rect 13132 20224 13172 20264
rect 17644 20308 17684 20348
rect 19900 20392 20268 20432
rect 27674 20392 28042 20432
rect 29932 20392 29972 20432
rect 23500 20308 23540 20348
rect 26668 20308 26708 20348
rect 27148 20308 27188 20348
rect 14188 20224 14219 20264
rect 14219 20224 14228 20264
rect 14668 20224 14708 20264
rect 15148 20224 15188 20264
rect 15916 20224 15956 20264
rect 16588 20224 16619 20264
rect 16619 20224 16628 20264
rect 18892 20224 18932 20264
rect 24172 20224 24212 20264
rect 6700 20140 6740 20180
rect 7276 20140 7316 20180
rect 8620 20140 8660 20180
rect 9772 20140 9812 20180
rect 1900 20056 1940 20096
rect 2284 20056 2324 20096
rect 3052 20056 3092 20096
rect 3340 20056 3380 20096
rect 3820 20056 3860 20096
rect 4684 20056 4724 20096
rect 460 19804 500 19844
rect 844 19804 884 19844
rect 5164 20056 5193 20096
rect 5193 20056 5204 20096
rect 5836 20056 5876 20096
rect 6124 20056 6153 20096
rect 6153 20056 6164 20096
rect 6892 20056 6931 20096
rect 6931 20056 6932 20096
rect 7372 20056 7412 20096
rect 8140 20087 8180 20096
rect 8140 20056 8171 20087
rect 8171 20056 8180 20087
rect 8716 20056 8756 20096
rect 9388 20056 9428 20096
rect 4300 19972 4340 20012
rect 5260 19972 5300 20012
rect 6028 19972 6068 20012
rect 6604 19888 6644 19928
rect 8140 19888 8180 19928
rect 13804 20140 13835 20180
rect 13835 20140 13844 20180
rect 16684 20140 16724 20180
rect 17164 20140 17204 20180
rect 19372 20140 19412 20180
rect 20812 20140 20852 20180
rect 24748 20140 24788 20180
rect 26572 20224 26612 20264
rect 28012 20224 28052 20264
rect 28972 20224 29012 20264
rect 26668 20140 26708 20180
rect 28108 20140 28148 20180
rect 29548 20140 29588 20180
rect 29932 20140 29972 20180
rect 12844 20056 12884 20096
rect 13900 20056 13940 20096
rect 14284 20056 14324 20096
rect 15532 20056 15572 20071
rect 15532 20031 15572 20056
rect 12748 19972 12788 20012
rect 14380 19972 14420 20012
rect 14668 19972 14708 20012
rect 15244 19972 15284 20012
rect 13324 19888 13364 19928
rect 13516 19888 13556 19928
rect 16204 19972 16244 20012
rect 16780 19972 16820 20012
rect 17260 19972 17300 20012
rect 17452 19972 17492 20012
rect 16492 19888 16532 19928
rect 17164 19888 17204 19928
rect 2572 19804 2612 19844
rect 4396 19804 4436 19844
rect 5068 19804 5108 19844
rect 7468 19804 7508 19844
rect 7852 19804 7892 19844
rect 13036 19804 13076 19844
rect 13900 19804 13940 19844
rect 14860 19804 14900 19844
rect 15916 19804 15956 19844
rect 17644 19804 17684 19844
rect 19564 20056 19568 20096
rect 19568 20056 19604 20096
rect 22156 20056 22196 20096
rect 23596 20056 23636 20096
rect 24652 20056 24692 20096
rect 25132 20056 25163 20096
rect 25163 20056 25172 20096
rect 18508 19972 18548 20012
rect 19084 19972 19124 20012
rect 19372 19972 19412 20012
rect 21868 19972 21908 20012
rect 19180 19888 19220 19928
rect 19660 19888 19700 19928
rect 18604 19804 18644 19844
rect 2956 19720 2996 19760
rect 6220 19720 6260 19760
rect 11692 19720 11732 19760
rect 14380 19720 14420 19760
rect 17260 19720 17300 19760
rect 18508 19720 18548 19760
rect 20812 19720 20852 19760
rect 3112 19636 3480 19676
rect 10156 19636 10196 19676
rect 10886 19636 11254 19676
rect 11500 19636 11540 19676
rect 4396 19468 4427 19508
rect 4427 19468 4436 19508
rect 6604 19468 6644 19508
rect 652 19384 692 19424
rect 3628 19384 3668 19424
rect 5836 19384 5876 19424
rect 940 19300 980 19340
rect 2188 19300 2228 19340
rect 3724 19300 3764 19340
rect 4588 19300 4628 19340
rect 5260 19300 5300 19340
rect 7180 19552 7220 19592
rect 10732 19468 10772 19508
rect 13420 19468 13460 19508
rect 14572 19468 14612 19508
rect 15148 19468 15188 19508
rect 6220 19300 6260 19340
rect 12652 19384 12692 19424
rect 12940 19384 12980 19424
rect 7660 19300 7700 19340
rect 9196 19300 9236 19340
rect 10636 19300 10676 19340
rect 12748 19300 12788 19340
rect 13228 19300 13268 19340
rect 14668 19300 14708 19340
rect 15148 19300 15188 19340
rect 15916 19300 15939 19340
rect 15939 19300 15956 19340
rect 2380 19216 2420 19256
rect 2764 19216 2804 19256
rect 3052 19216 3092 19256
rect 3532 19216 3572 19256
rect 3820 19216 3860 19256
rect 4300 19216 4340 19256
rect 5068 19216 5108 19256
rect 6124 19216 6164 19256
rect 6604 19216 6644 19256
rect 6892 19216 6921 19256
rect 6921 19216 6932 19256
rect 7756 19216 7796 19256
rect 9004 19216 9044 19256
rect 18660 19636 19028 19676
rect 19564 19468 19604 19508
rect 22828 19804 22868 19844
rect 23020 19720 23060 19760
rect 22636 19552 22676 19592
rect 23308 19552 23348 19592
rect 25324 20056 25364 20096
rect 25516 20056 25556 20096
rect 26572 20056 26612 20096
rect 26860 20056 26900 20096
rect 27532 20056 27572 20096
rect 29452 20056 29492 20096
rect 24748 19972 24788 20012
rect 25804 19972 25844 20012
rect 26956 19972 26996 20012
rect 27244 19972 27284 20012
rect 28108 19972 28148 20012
rect 31372 19972 31412 20012
rect 25132 19888 25172 19928
rect 26380 19888 26420 19928
rect 27148 19888 27188 19928
rect 22348 19384 22388 19424
rect 27628 19804 27668 19844
rect 29644 19804 29684 19844
rect 26860 19720 26900 19760
rect 26434 19636 26802 19676
rect 27148 19384 27188 19424
rect 27724 19552 27764 19592
rect 30316 19552 30356 19592
rect 28204 19468 28244 19508
rect 28492 19468 28532 19508
rect 30508 19468 30548 19508
rect 17452 19300 17492 19340
rect 20140 19300 20180 19340
rect 20716 19300 20756 19340
rect 23116 19300 23156 19340
rect 24556 19300 24596 19340
rect 26572 19300 26612 19340
rect 9772 19216 9812 19256
rect 10156 19216 10196 19256
rect 11308 19216 11348 19256
rect 11788 19216 11828 19256
rect 12556 19216 12596 19256
rect 652 19048 692 19088
rect 3628 19132 3668 19172
rect 4012 19132 4052 19172
rect 2572 19048 2612 19088
rect 3148 19048 3188 19088
rect 3436 18880 3476 18920
rect 5164 19132 5204 19172
rect 5548 19132 5588 19172
rect 6028 19132 6068 19172
rect 6316 19132 6356 19172
rect 6508 19132 6548 19172
rect 7276 19132 7316 19172
rect 8908 19132 8948 19172
rect 13900 19216 13912 19256
rect 13912 19216 13940 19256
rect 14092 19216 14123 19256
rect 14123 19216 14132 19256
rect 14476 19216 14516 19256
rect 14764 19216 14804 19256
rect 15436 19216 15476 19256
rect 16204 19216 16244 19256
rect 16972 19216 16984 19256
rect 16984 19216 17012 19256
rect 17836 19216 17876 19256
rect 28876 19384 28916 19424
rect 27820 19300 27860 19340
rect 28204 19300 28244 19340
rect 30604 19300 30644 19340
rect 18604 19216 18644 19256
rect 19276 19216 19316 19256
rect 19570 19216 19607 19256
rect 19607 19216 19610 19256
rect 21292 19216 21332 19256
rect 21772 19216 21812 19256
rect 22156 19216 22187 19256
rect 22187 19216 22196 19256
rect 22636 19216 22667 19256
rect 22667 19216 22676 19256
rect 22924 19216 22964 19256
rect 23404 19216 23444 19256
rect 23980 19216 23985 19256
rect 23985 19216 24020 19256
rect 24364 19216 24404 19256
rect 24844 19216 24875 19256
rect 24875 19216 24884 19256
rect 25612 19216 25652 19256
rect 26380 19216 26420 19256
rect 27148 19216 27188 19256
rect 28396 19216 28436 19256
rect 29452 19216 29492 19256
rect 9388 19132 9428 19172
rect 10732 19132 10772 19172
rect 13708 19132 13748 19172
rect 14860 19132 14900 19172
rect 4300 19048 4340 19088
rect 6988 19048 7028 19088
rect 8716 19048 8756 19088
rect 9964 19048 10004 19088
rect 11980 19048 12020 19088
rect 13900 19048 13940 19088
rect 6412 18964 6452 19004
rect 15244 19132 15284 19172
rect 16492 19132 16532 19172
rect 19660 19132 19700 19172
rect 20332 19132 20372 19172
rect 20716 19132 20756 19172
rect 22252 19132 22292 19172
rect 4352 18880 4720 18920
rect 9196 18964 9236 19004
rect 10156 18964 10196 19004
rect 13516 18964 13556 19004
rect 14476 18964 14516 19004
rect 8524 18796 8564 18836
rect 8908 18880 8948 18920
rect 12126 18880 12494 18920
rect 13900 18880 13940 18920
rect 15148 18880 15188 18920
rect 9388 18796 9428 18836
rect 16012 19048 16052 19088
rect 17164 19048 17204 19088
rect 15244 18796 15284 18836
rect 16204 18796 16244 18836
rect 3628 18712 3668 18752
rect 5068 18712 5108 18752
rect 5260 18712 5300 18752
rect 6604 18712 6644 18752
rect 6892 18712 6923 18752
rect 6923 18712 6932 18752
rect 7756 18712 7796 18752
rect 11308 18712 11348 18752
rect 11884 18712 11924 18752
rect 12556 18712 12596 18752
rect 13708 18712 13748 18752
rect 14188 18712 14228 18752
rect 8620 18628 8660 18668
rect 8908 18628 8948 18668
rect 9676 18628 9716 18668
rect 10348 18628 10388 18668
rect 10540 18628 10580 18668
rect 3148 18544 3188 18584
rect 4108 18544 4148 18584
rect 4684 18544 4724 18584
rect 4972 18544 5012 18584
rect 5452 18544 5492 18584
rect 6124 18544 6148 18584
rect 6148 18544 6164 18584
rect 6700 18544 6731 18584
rect 6731 18544 6740 18584
rect 7180 18544 7220 18584
rect 7756 18544 7796 18584
rect 8236 18544 8276 18584
rect 9100 18544 9140 18584
rect 10156 18544 10196 18584
rect 1996 18460 2036 18500
rect 3724 18460 3764 18500
rect 4876 18460 4916 18500
rect 5068 18460 5108 18500
rect 6220 18460 6260 18500
rect 6412 18460 6452 18500
rect 7564 18460 7604 18500
rect 14284 18628 14324 18668
rect 18028 19048 18068 19088
rect 20044 19048 20084 19088
rect 14764 18712 14804 18752
rect 15436 18712 15476 18752
rect 16972 18712 17012 18752
rect 18604 18712 18644 18752
rect 19276 18712 19316 18752
rect 15052 18628 15092 18668
rect 16204 18628 16244 18668
rect 16876 18628 16916 18668
rect 11404 18544 11444 18584
rect 12460 18544 12500 18584
rect 12844 18544 12884 18584
rect 13708 18544 13748 18584
rect 14572 18544 14612 18584
rect 15244 18544 15284 18584
rect 16588 18544 16628 18584
rect 17068 18544 17108 18584
rect 8428 18460 8459 18500
rect 8459 18460 8468 18500
rect 9580 18460 9620 18500
rect 8716 18376 8756 18416
rect 11308 18460 11348 18500
rect 12172 18460 12212 18500
rect 2284 18292 2324 18332
rect 6892 18292 6932 18332
rect 7756 18292 7796 18332
rect 8524 18292 8564 18332
rect 9004 18292 9044 18332
rect 13900 18460 13940 18500
rect 14284 18460 14324 18500
rect 12652 18376 12692 18416
rect 13996 18376 14036 18416
rect 14380 18376 14420 18416
rect 14668 18376 14708 18416
rect 10636 18292 10676 18332
rect 6604 18208 6644 18248
rect 9196 18208 9236 18248
rect 1996 17872 2036 17912
rect 2380 17788 2420 17828
rect 3112 18124 3480 18164
rect 10886 18124 11254 18164
rect 11500 18124 11540 18164
rect 12460 18124 12500 18164
rect 6220 18040 6260 18080
rect 3724 17956 3764 17996
rect 7180 17956 7220 17996
rect 2668 17788 2708 17828
rect 3820 17872 3860 17912
rect 4204 17872 4244 17912
rect 4972 17872 5012 17912
rect 5932 17872 5972 17912
rect 6220 17872 6260 17912
rect 2956 17788 2996 17828
rect 5356 17788 5396 17828
rect 9100 18040 9140 18080
rect 11404 18040 11444 18080
rect 12364 18040 12404 18080
rect 6604 17788 6644 17828
rect 2572 17704 2612 17744
rect 3148 17704 3188 17744
rect 4204 17704 4244 17744
rect 4396 17704 4436 17744
rect 4780 17704 4820 17744
rect 5740 17704 5764 17744
rect 5764 17704 5780 17744
rect 7468 17788 7508 17828
rect 8716 17872 8756 17912
rect 9772 17956 9812 17996
rect 11020 17956 11060 17996
rect 11212 17956 11252 17996
rect 9676 17872 9716 17912
rect 11500 17872 11540 17912
rect 8044 17788 8084 17828
rect 8620 17788 8660 17828
rect 10540 17788 10580 17828
rect 10732 17788 10772 17828
rect 15148 18460 15188 18500
rect 15244 18376 15284 18416
rect 15628 18376 15668 18416
rect 14764 18292 14804 18332
rect 19900 18880 20268 18920
rect 23212 18880 23252 18920
rect 23404 18880 23444 18920
rect 21292 18796 21332 18836
rect 24844 19048 24884 19088
rect 25804 19048 25844 19088
rect 26284 19079 26324 19088
rect 26284 19048 26323 19079
rect 26323 19048 26324 19079
rect 27628 19048 27668 19088
rect 31084 19048 31124 19088
rect 26092 18964 26132 19004
rect 30508 18964 30548 19004
rect 25612 18880 25652 18920
rect 27674 18880 28042 18920
rect 28876 18880 28916 18920
rect 29452 18796 29492 18836
rect 29932 18796 29972 18836
rect 20332 18712 20372 18752
rect 23020 18712 23060 18752
rect 23980 18712 24020 18752
rect 24940 18712 24980 18752
rect 25420 18712 25460 18752
rect 27436 18712 27476 18752
rect 20524 18628 20564 18668
rect 22348 18628 22388 18668
rect 23212 18628 23252 18668
rect 23788 18628 23828 18668
rect 24076 18628 24116 18668
rect 25804 18628 25844 18668
rect 26284 18628 26324 18668
rect 26476 18628 26516 18668
rect 29644 18628 29684 18668
rect 30028 18628 30068 18668
rect 16204 18460 16244 18500
rect 17836 18544 17876 18584
rect 18604 18544 18644 18584
rect 19276 18544 19316 18584
rect 16588 18376 16628 18416
rect 17260 18376 17300 18416
rect 18988 18460 19028 18500
rect 16492 18292 16532 18332
rect 17452 18292 17492 18332
rect 12172 17956 12212 17996
rect 12556 17956 12596 17996
rect 14284 17956 14324 17996
rect 14668 17956 14708 17996
rect 13132 17872 13172 17912
rect 13228 17788 13268 17828
rect 13900 17872 13940 17912
rect 14380 17872 14420 17912
rect 13996 17788 14036 17828
rect 14572 17788 14612 17828
rect 20428 18544 20444 18584
rect 20444 18544 20468 18584
rect 20812 18544 20852 18584
rect 21292 18544 21332 18584
rect 21676 18544 21716 18584
rect 19660 18460 19700 18500
rect 20332 18460 20372 18500
rect 21196 18460 21236 18500
rect 21868 18460 21908 18500
rect 18316 18376 18356 18416
rect 21388 18376 21428 18416
rect 18412 18292 18452 18332
rect 23596 18575 23636 18584
rect 23596 18544 23636 18575
rect 23980 18544 24020 18584
rect 24364 18544 24404 18584
rect 26380 18544 26420 18584
rect 26764 18544 26804 18584
rect 22444 18460 22484 18500
rect 23500 18460 23540 18500
rect 24844 18460 24884 18500
rect 24556 18376 24596 18416
rect 25612 18460 25652 18500
rect 26092 18460 26123 18500
rect 26123 18460 26132 18500
rect 27340 18460 27380 18500
rect 30316 18712 30356 18752
rect 30700 18628 30740 18668
rect 29548 18544 29588 18584
rect 30316 18460 30356 18500
rect 26956 18376 26996 18416
rect 27724 18376 27764 18416
rect 29836 18376 29876 18416
rect 22252 18292 22292 18332
rect 22636 18292 22676 18332
rect 24268 18292 24308 18332
rect 15436 18208 15476 18248
rect 17260 18208 17300 18248
rect 21964 18208 22004 18248
rect 23020 18208 23060 18248
rect 23212 18208 23252 18248
rect 24364 18208 24404 18248
rect 18660 18124 19028 18164
rect 19276 18124 19316 18164
rect 17836 18040 17876 18080
rect 20236 18040 20276 18080
rect 20620 18040 20660 18080
rect 20812 18040 20852 18080
rect 21580 18040 21620 18080
rect 23596 18040 23636 18080
rect 15436 17956 15476 17996
rect 22156 17956 22196 17996
rect 16396 17872 16436 17912
rect 15724 17788 15764 17828
rect 16780 17788 16820 17828
rect 18988 17872 19028 17912
rect 19756 17872 19796 17912
rect 20428 17872 20468 17912
rect 6796 17704 6836 17744
rect 3724 17620 3764 17660
rect 4588 17620 4628 17660
rect 4972 17620 5012 17660
rect 5260 17620 5300 17660
rect 5548 17620 5588 17660
rect 5932 17620 5972 17660
rect 6508 17620 6548 17660
rect 7276 17620 7316 17660
rect 2092 17536 2132 17576
rect 3628 17536 3668 17576
rect 5452 17536 5492 17576
rect 6412 17536 6452 17576
rect 8332 17704 8371 17744
rect 8371 17704 8372 17744
rect 9196 17704 9215 17744
rect 9215 17704 9236 17744
rect 10636 17704 10648 17744
rect 10648 17704 10676 17744
rect 11020 17704 11060 17744
rect 7468 17620 7508 17660
rect 8236 17620 8276 17660
rect 8620 17620 8660 17660
rect 7660 17536 7700 17576
rect 9196 17536 9236 17576
rect 10252 17620 10292 17660
rect 11308 17620 11348 17660
rect 11596 17620 11636 17660
rect 11884 17620 11924 17660
rect 13708 17704 13733 17744
rect 13733 17704 13748 17744
rect 14668 17704 14708 17744
rect 15820 17704 15860 17744
rect 16300 17704 16312 17744
rect 16312 17704 16340 17744
rect 16492 17704 16523 17744
rect 16523 17704 16532 17744
rect 17836 17704 17876 17744
rect 12460 17620 12500 17660
rect 10060 17536 10100 17576
rect 10348 17536 10388 17576
rect 12652 17536 12692 17576
rect 12844 17536 12884 17576
rect 13132 17536 13172 17576
rect 13900 17536 13940 17576
rect 14188 17536 14228 17576
rect 9676 17452 9716 17492
rect 4352 17368 4720 17408
rect 12126 17368 12494 17408
rect 14668 17368 14708 17408
rect 15052 17620 15092 17660
rect 18604 17788 18644 17828
rect 18796 17788 18836 17828
rect 19084 17788 19124 17828
rect 20236 17788 20276 17828
rect 21196 17788 21236 17828
rect 22060 17788 22100 17828
rect 18124 17704 18164 17744
rect 18700 17704 18740 17744
rect 18988 17704 19028 17744
rect 20524 17704 20555 17744
rect 20555 17704 20564 17744
rect 21004 17704 21044 17744
rect 21964 17704 22004 17744
rect 15628 17620 15668 17660
rect 16204 17620 16244 17660
rect 17260 17620 17300 17660
rect 18316 17620 18356 17660
rect 20332 17620 20372 17660
rect 15436 17536 15476 17576
rect 16876 17536 16916 17576
rect 17836 17536 17876 17576
rect 18412 17536 18452 17576
rect 20524 17536 20564 17576
rect 20812 17536 20852 17576
rect 16684 17452 16724 17492
rect 19180 17452 19220 17492
rect 21772 17452 21812 17492
rect 22828 17788 22868 17828
rect 23116 17788 23156 17828
rect 23308 17788 23348 17828
rect 23500 17956 23540 17996
rect 23596 17788 23636 17828
rect 22348 17704 22388 17744
rect 24844 17956 24884 17996
rect 24364 17872 24404 17912
rect 24076 17788 24116 17828
rect 24268 17788 24308 17828
rect 27436 18292 27476 18332
rect 28972 18292 29012 18332
rect 30220 18292 30260 18332
rect 26284 18208 26324 18248
rect 26434 18124 26802 18164
rect 27628 18124 27668 18164
rect 25804 17956 25844 17996
rect 30220 17956 30260 17996
rect 28108 17788 28139 17828
rect 28139 17788 28148 17828
rect 30988 17788 31028 17828
rect 24364 17704 24404 17744
rect 23116 17620 23156 17660
rect 23404 17620 23444 17660
rect 24652 17704 24692 17744
rect 25516 17704 25556 17744
rect 29644 17704 29675 17744
rect 29675 17704 29684 17744
rect 30700 17704 30728 17744
rect 30728 17704 30740 17744
rect 23884 17620 23924 17660
rect 25420 17620 25460 17660
rect 30028 17620 30059 17660
rect 30059 17620 30068 17660
rect 30892 17620 30932 17660
rect 24268 17536 24308 17576
rect 23020 17452 23060 17492
rect 23212 17452 23252 17492
rect 26572 17452 26612 17492
rect 26764 17452 26804 17492
rect 5068 17284 5108 17324
rect 6028 17284 6068 17324
rect 7276 17284 7316 17324
rect 11020 17284 11060 17324
rect 1996 17200 2036 17240
rect 4012 17200 4052 17240
rect 4492 17200 4523 17240
rect 4523 17200 4532 17240
rect 4972 17200 5003 17240
rect 5003 17200 5012 17240
rect 6508 17200 6548 17240
rect 8428 17200 8468 17240
rect 8812 17200 8843 17240
rect 8843 17200 8852 17240
rect 4780 17116 4820 17156
rect 5548 17116 5588 17156
rect 6220 17116 6260 17156
rect 7180 17116 7220 17156
rect 3244 17032 3284 17072
rect 3628 17032 3668 17072
rect 4588 17032 4628 17072
rect 4684 16948 4724 16988
rect 5452 17032 5481 17072
rect 5481 17032 5492 17072
rect 5260 16948 5300 16988
rect 5740 16948 5780 16988
rect 5932 16948 5972 16988
rect 6796 17032 6836 17072
rect 6508 16948 6548 16988
rect 19900 17368 20268 17408
rect 22924 17368 22964 17408
rect 27674 17368 28042 17408
rect 16972 17284 17012 17324
rect 22732 17284 22772 17324
rect 23692 17284 23732 17324
rect 23884 17284 23924 17324
rect 28108 17284 28148 17324
rect 9388 17200 9428 17240
rect 10252 17200 10292 17240
rect 10540 17200 10580 17240
rect 12172 17200 12212 17240
rect 12460 17200 12500 17240
rect 13036 17200 13076 17240
rect 13228 17200 13268 17240
rect 15724 17200 15764 17240
rect 16108 17200 16148 17240
rect 16780 17200 16811 17240
rect 16811 17200 16820 17240
rect 18412 17200 18452 17240
rect 18604 17200 18644 17240
rect 19948 17200 19988 17240
rect 20716 17200 20756 17240
rect 21580 17200 21620 17240
rect 24268 17200 24308 17240
rect 25132 17200 25172 17240
rect 26956 17200 26996 17240
rect 27340 17200 27380 17240
rect 9004 17116 9044 17156
rect 8044 17032 8084 17072
rect 9484 17116 9524 17156
rect 11404 17116 11444 17156
rect 13324 17116 13364 17156
rect 13996 17116 14036 17156
rect 10060 17032 10100 17072
rect 10252 17032 10292 17072
rect 11500 17032 11512 17072
rect 11512 17032 11540 17072
rect 11884 17032 11924 17072
rect 12172 17032 12212 17072
rect 12652 17032 12692 17072
rect 13228 17032 13268 17072
rect 13516 17032 13556 17072
rect 7468 16948 7508 16988
rect 7852 16948 7892 16988
rect 4492 16864 4532 16904
rect 6220 16864 6260 16904
rect 7372 16864 7412 16904
rect 8428 16864 8468 16904
rect 2572 16780 2612 16820
rect 6604 16780 6644 16820
rect 7180 16780 7220 16820
rect 7852 16780 7892 16820
rect 3112 16612 3480 16652
rect 3628 16612 3668 16652
rect 6124 16528 6164 16568
rect 14380 17032 14409 17072
rect 14409 17032 14420 17072
rect 15436 17116 15476 17156
rect 15628 17116 15668 17156
rect 16972 17116 17012 17156
rect 9964 16948 10004 16988
rect 10540 16948 10580 16988
rect 10828 16948 10868 16988
rect 13036 16948 13076 16988
rect 13612 16948 13652 16988
rect 13900 16948 13940 16988
rect 9868 16864 9908 16904
rect 10444 16780 10484 16820
rect 11404 16780 11444 16820
rect 10886 16612 11254 16652
rect 16012 17032 16028 17072
rect 16028 17032 16052 17072
rect 14668 16948 14708 16988
rect 15340 16948 15380 16988
rect 15820 16948 15860 16988
rect 16204 16948 16244 16988
rect 16492 16948 16532 16988
rect 16684 16948 16724 16988
rect 14476 16864 14516 16904
rect 16396 16864 16436 16904
rect 14092 16780 14132 16820
rect 19852 17116 19892 17156
rect 20332 17116 20372 17156
rect 23308 17116 23348 17156
rect 23692 17116 23732 17156
rect 23884 17116 23924 17156
rect 24844 17116 24884 17156
rect 27724 17116 27764 17156
rect 30028 17200 30068 17240
rect 31756 17116 31796 17156
rect 17068 16948 17108 16988
rect 18316 17032 18356 17072
rect 17260 16948 17300 16988
rect 18220 16864 18260 16904
rect 12748 16696 12788 16736
rect 13132 16612 13172 16652
rect 13516 16612 13556 16652
rect 16204 16612 16244 16652
rect 10060 16528 10100 16568
rect 11980 16528 12020 16568
rect 13900 16528 13940 16568
rect 4876 16444 4916 16484
rect 5836 16444 5876 16484
rect 6988 16444 7028 16484
rect 9196 16444 9236 16484
rect 9676 16444 9716 16484
rect 2188 16276 2228 16316
rect 5356 16360 5396 16400
rect 6220 16360 6260 16400
rect 6028 16276 6068 16316
rect 7180 16276 7220 16316
rect 7564 16276 7604 16316
rect 8044 16276 8084 16316
rect 8428 16276 8468 16316
rect 9484 16360 9524 16400
rect 18892 17032 18932 17072
rect 19372 17032 19412 17072
rect 20236 17032 20260 17072
rect 20260 17032 20276 17072
rect 20332 16948 20372 16988
rect 20140 16864 20180 16904
rect 21100 17032 21140 17072
rect 22060 17032 22100 17072
rect 22540 17032 22580 17072
rect 23020 17032 23060 17072
rect 23500 17032 23540 17072
rect 20812 16948 20852 16988
rect 21580 16948 21620 16988
rect 21964 16948 22004 16988
rect 22156 16948 22196 16988
rect 24364 17032 24368 17072
rect 24368 17032 24404 17072
rect 24940 17032 24980 17072
rect 25708 17032 25748 17072
rect 26188 17032 26228 17072
rect 22924 16948 22964 16988
rect 23116 16948 23156 16988
rect 21484 16864 21524 16904
rect 21580 16780 21620 16820
rect 27052 17032 27092 17072
rect 28012 17032 28052 17072
rect 29740 17032 29780 17072
rect 30220 17032 30260 17072
rect 25132 16948 25172 16988
rect 25612 16948 25652 16988
rect 25804 16948 25844 16988
rect 26284 16948 26324 16988
rect 22828 16864 22868 16904
rect 23020 16864 23060 16904
rect 24748 16864 24788 16904
rect 27436 16948 27476 16988
rect 28300 16948 28340 16988
rect 27052 16864 27092 16904
rect 28204 16864 28244 16904
rect 29932 16864 29972 16904
rect 23596 16780 23636 16820
rect 30988 16864 31028 16904
rect 28108 16780 28148 16820
rect 20332 16696 20372 16736
rect 15244 16444 15284 16484
rect 17932 16444 17972 16484
rect 18316 16444 18356 16484
rect 18660 16612 19028 16652
rect 19372 16612 19412 16652
rect 22060 16612 22100 16652
rect 20236 16444 20276 16484
rect 21196 16444 21236 16484
rect 23788 16444 23828 16484
rect 25132 16444 25172 16484
rect 15052 16360 15092 16400
rect 18988 16360 19028 16400
rect 9388 16276 9390 16316
rect 9390 16276 9428 16316
rect 10252 16276 10292 16316
rect 11308 16276 11348 16316
rect 12748 16276 12788 16316
rect 13324 16276 13364 16316
rect 14284 16276 14324 16316
rect 14476 16276 14516 16316
rect 15244 16276 15284 16316
rect 15436 16276 15476 16316
rect 16108 16276 16148 16316
rect 16684 16276 16724 16316
rect 16972 16276 17012 16316
rect 17644 16276 17684 16316
rect 19276 16276 19316 16316
rect 1996 16192 2036 16232
rect 2860 16192 2900 16232
rect 3628 16192 3668 16232
rect 4972 16192 5012 16232
rect 5356 16192 5396 16232
rect 6220 16192 6249 16232
rect 6249 16192 6260 16232
rect 6508 16192 6548 16232
rect 6796 16192 6836 16232
rect 7852 16192 7892 16232
rect 1804 16108 1844 16148
rect 3340 16108 3380 16148
rect 4108 16108 4148 16148
rect 4588 16108 4628 16148
rect 5932 16108 5972 16148
rect 7084 16108 7124 16148
rect 7564 16108 7604 16148
rect 8044 16108 8084 16148
rect 4012 16024 4052 16064
rect 4684 16024 4724 16064
rect 5260 16024 5291 16064
rect 5291 16024 5300 16064
rect 6700 16024 6740 16064
rect 76 15772 116 15812
rect 7948 16024 7988 16064
rect 8428 16108 8468 16148
rect 8716 16108 8756 16148
rect 9100 16108 9140 16148
rect 9676 16108 9716 16148
rect 10924 16192 10964 16232
rect 12076 16192 12116 16232
rect 13228 16192 13268 16232
rect 13900 16192 13940 16232
rect 14572 16192 14612 16232
rect 15148 16192 15188 16232
rect 15628 16192 15668 16232
rect 16204 16192 16244 16232
rect 16876 16192 16916 16232
rect 19756 16276 19796 16316
rect 21484 16276 21524 16316
rect 21868 16276 21908 16316
rect 25132 16276 25172 16316
rect 18316 16192 18356 16232
rect 19180 16192 19220 16232
rect 23308 16192 23348 16232
rect 23788 16192 23828 16232
rect 24268 16192 24308 16232
rect 24652 16192 24692 16232
rect 26284 16696 26324 16736
rect 26434 16612 26802 16652
rect 26956 16612 26996 16652
rect 27532 16528 27572 16568
rect 27052 16360 27092 16400
rect 30220 16360 30260 16400
rect 25516 16276 25556 16316
rect 27340 16276 27380 16316
rect 28204 16276 28235 16316
rect 28235 16276 28244 16316
rect 29932 16276 29972 16316
rect 24940 16192 24971 16203
rect 24971 16192 24980 16203
rect 9964 16108 10004 16148
rect 10252 16108 10292 16148
rect 10828 16108 10868 16148
rect 11308 16108 11348 16148
rect 11500 16108 11540 16148
rect 12460 16108 12500 16148
rect 12748 16108 12788 16148
rect 13804 16108 13844 16148
rect 16396 16108 16436 16148
rect 16972 16108 17012 16148
rect 17932 16108 17972 16148
rect 19564 16108 19604 16148
rect 7276 15940 7316 15980
rect 9484 16024 9524 16064
rect 10444 16024 10484 16064
rect 4352 15856 4720 15896
rect 4012 15772 4052 15812
rect 5164 15772 5204 15812
rect 6892 15856 6932 15896
rect 9292 15856 9332 15896
rect 11404 15856 11444 15896
rect 10924 15772 10964 15812
rect 1996 15688 2036 15728
rect 3532 15688 3572 15728
rect 4876 15688 4916 15728
rect 5068 15688 5108 15728
rect 5356 15688 5396 15728
rect 7564 15688 7604 15728
rect 8812 15688 8852 15728
rect 2860 15604 2900 15644
rect 4492 15604 4532 15644
rect 4684 15604 4724 15644
rect 4972 15604 5012 15644
rect 5452 15604 5492 15644
rect 6220 15604 6260 15644
rect 6892 15604 6932 15644
rect 7660 15604 7700 15644
rect 10060 15688 10100 15728
rect 12748 15940 12788 15980
rect 17260 16024 17300 16064
rect 18604 16024 18644 16064
rect 24940 16163 24980 16192
rect 31084 16276 31124 16316
rect 25804 16192 25844 16232
rect 26284 16192 26324 16232
rect 26668 16223 26708 16232
rect 26668 16192 26699 16223
rect 26699 16192 26708 16223
rect 27436 16192 27476 16232
rect 29644 16192 29684 16232
rect 31756 16192 31796 16232
rect 22060 16108 22100 16148
rect 23116 16108 23156 16148
rect 23404 16108 23444 16148
rect 24172 16108 24212 16148
rect 25420 16108 25460 16148
rect 26188 16108 26228 16148
rect 26764 16108 26804 16148
rect 29164 16108 29204 16148
rect 22732 16024 22772 16064
rect 23596 16024 23636 16064
rect 25612 16024 25652 16064
rect 27052 16024 27092 16064
rect 28012 16024 28052 16064
rect 30508 16108 30548 16148
rect 30796 16108 30836 16148
rect 15340 15940 15380 15980
rect 27148 15940 27188 15980
rect 30700 15940 30740 15980
rect 11980 15856 12020 15896
rect 12126 15856 12494 15896
rect 14764 15856 14804 15896
rect 15628 15856 15668 15896
rect 17452 15856 17492 15896
rect 17932 15856 17972 15896
rect 18316 15856 18356 15896
rect 19900 15856 20268 15896
rect 27674 15856 28042 15896
rect 11788 15688 11819 15728
rect 11819 15688 11828 15728
rect 14476 15772 14516 15812
rect 15244 15772 15284 15812
rect 16876 15772 16916 15812
rect 12172 15688 12212 15728
rect 9580 15604 9620 15644
rect 9868 15604 9908 15644
rect 12364 15604 12404 15644
rect 12940 15604 12980 15644
rect 1708 15520 1748 15560
rect 2572 15551 2612 15560
rect 2572 15520 2612 15551
rect 2956 15520 2996 15560
rect 3340 15520 3380 15560
rect 4012 15520 4052 15560
rect 5548 15520 5588 15560
rect 6604 15520 6644 15560
rect 8140 15520 8180 15560
rect 8620 15520 8660 15560
rect 9484 15520 9524 15560
rect 10732 15520 10741 15560
rect 10741 15520 10772 15560
rect 11020 15520 11060 15560
rect 1612 15436 1652 15476
rect 4588 15436 4628 15476
rect 5164 15436 5204 15476
rect 6700 15436 6739 15476
rect 6739 15436 6740 15476
rect 6796 15352 6836 15392
rect 2956 15268 2996 15308
rect 3724 15184 3764 15224
rect 11884 15520 11900 15560
rect 11900 15520 11924 15560
rect 12748 15520 12788 15560
rect 7948 15436 7988 15476
rect 8428 15436 8468 15476
rect 9196 15436 9236 15476
rect 10060 15436 10100 15476
rect 10636 15436 10676 15476
rect 11116 15436 11156 15476
rect 11404 15436 11444 15476
rect 4204 15268 4244 15308
rect 5932 15268 5972 15308
rect 4588 15184 4628 15224
rect 3112 15100 3480 15140
rect 4972 15100 5012 15140
rect 1612 14932 1652 14972
rect 4204 14932 4235 14972
rect 4235 14932 4244 14972
rect 4876 14848 4916 14888
rect 6028 14848 6068 14888
rect 6892 14848 6932 14888
rect 8524 14848 8564 14888
rect 652 14764 692 14804
rect 2764 14764 2804 14804
rect 2956 14764 2996 14804
rect 3148 14764 3188 14804
rect 4588 14764 4628 14804
rect 1324 14680 1364 14720
rect 1516 14680 1556 14720
rect 2092 14680 2132 14720
rect 3436 14680 3476 14720
rect 3628 14680 3668 14720
rect 4684 14680 4724 14720
rect 6124 14764 6164 14804
rect 6316 14764 6356 14804
rect 5932 14731 5972 14762
rect 5932 14722 5972 14731
rect 5644 14680 5684 14720
rect 6604 14764 6644 14804
rect 7180 14764 7220 14804
rect 7468 14764 7508 14804
rect 8140 14764 8180 14804
rect 8812 14764 8852 14804
rect 8044 14680 8084 14720
rect 1708 14596 1748 14636
rect 2956 14596 2996 14636
rect 4492 14596 4532 14636
rect 6508 14596 6548 14636
rect 2092 14512 2132 14552
rect 4204 14512 4244 14552
rect 4588 14512 4628 14552
rect 4972 14512 5012 14552
rect 5164 14512 5204 14552
rect 5356 14428 5396 14468
rect 11884 15352 11924 15392
rect 10636 15268 10676 15308
rect 11692 15268 11732 15308
rect 21100 15772 21140 15812
rect 28204 15772 28244 15812
rect 13324 15688 13364 15728
rect 13612 15688 13652 15728
rect 18508 15688 18548 15728
rect 13516 15604 13556 15644
rect 13804 15635 13844 15644
rect 13804 15604 13835 15635
rect 13835 15604 13844 15635
rect 14476 15604 14516 15644
rect 14764 15604 14804 15644
rect 15148 15604 15188 15644
rect 16108 15604 16148 15644
rect 17452 15604 17492 15644
rect 19180 15604 19220 15644
rect 20332 15604 20372 15644
rect 22060 15688 22100 15728
rect 24268 15688 24308 15728
rect 25132 15688 25172 15728
rect 27436 15688 27467 15728
rect 27467 15688 27476 15728
rect 13228 15436 13268 15476
rect 13132 15352 13172 15392
rect 12748 15268 12788 15308
rect 13324 15268 13364 15308
rect 12268 15184 12308 15224
rect 10886 15100 11254 15140
rect 9292 15016 9332 15056
rect 10732 15016 10772 15056
rect 12844 15016 12884 15056
rect 10060 14932 10100 14972
rect 11788 14932 11828 14972
rect 12076 14932 12116 14972
rect 14213 15520 14253 15560
rect 15628 15520 15668 15560
rect 13804 15436 13844 15476
rect 14092 15436 14132 15476
rect 15436 15436 15476 15476
rect 16492 15436 16532 15476
rect 16876 15436 16916 15476
rect 14188 15352 14228 15392
rect 14764 15352 14804 15392
rect 15244 15352 15284 15392
rect 14284 15268 14324 15308
rect 13996 15184 14036 15224
rect 22732 15604 22772 15644
rect 24844 15604 24884 15644
rect 26956 15604 26996 15644
rect 29932 15604 29972 15644
rect 18220 15520 18260 15560
rect 19084 15520 19124 15560
rect 19564 15520 19604 15560
rect 20524 15520 20564 15560
rect 21388 15520 21428 15560
rect 21580 15520 21611 15560
rect 21611 15520 21620 15560
rect 22060 15520 22100 15560
rect 22444 15520 22484 15560
rect 17452 15436 17492 15476
rect 17932 15436 17972 15476
rect 18508 15352 18548 15392
rect 18660 15100 19028 15140
rect 17932 15016 17972 15056
rect 20428 15436 20468 15476
rect 24076 15436 24116 15476
rect 21292 15268 21332 15308
rect 22252 15268 22283 15308
rect 22283 15268 22292 15308
rect 24652 15268 24692 15308
rect 25708 15520 25748 15560
rect 27628 15520 27668 15560
rect 28108 15520 28148 15560
rect 25612 15436 25652 15476
rect 25516 15352 25556 15392
rect 25708 15352 25748 15392
rect 26188 15352 26228 15392
rect 26956 15352 26996 15392
rect 28012 15436 28052 15476
rect 30700 15436 30740 15476
rect 31180 15436 31220 15476
rect 30316 15352 30356 15392
rect 27340 15268 27380 15308
rect 19948 15184 19988 15224
rect 24748 15184 24788 15224
rect 26284 15184 26324 15224
rect 26434 15100 26802 15140
rect 23884 15016 23924 15056
rect 27532 15016 27572 15056
rect 19852 14932 19892 14972
rect 11500 14848 11540 14888
rect 9580 14764 9603 14804
rect 9603 14764 9620 14804
rect 11980 14848 12020 14888
rect 12172 14848 12212 14888
rect 15052 14848 15083 14888
rect 15083 14848 15092 14888
rect 16012 14848 16052 14888
rect 17548 14848 17588 14888
rect 20620 14848 20660 14888
rect 10636 14764 10676 14804
rect 14092 14764 14132 14804
rect 15724 14764 15764 14804
rect 16300 14764 16340 14804
rect 18604 14764 18644 14804
rect 21100 14764 21131 14804
rect 21131 14764 21140 14804
rect 8524 14680 8533 14720
rect 8533 14680 8564 14720
rect 9388 14680 9428 14720
rect 9868 14680 9899 14720
rect 9899 14680 9908 14720
rect 10924 14680 10940 14720
rect 10940 14680 10964 14720
rect 12460 14680 12500 14720
rect 13516 14680 13556 14720
rect 13708 14680 13748 14720
rect 9484 14596 9524 14636
rect 9772 14596 9812 14636
rect 10540 14596 10580 14636
rect 10732 14596 10772 14636
rect 12364 14596 12404 14636
rect 6412 14512 6443 14552
rect 6443 14512 6452 14552
rect 7276 14512 7316 14552
rect 9004 14512 9044 14552
rect 10252 14428 10292 14468
rect 10636 14428 10676 14468
rect 12844 14428 12884 14468
rect 3916 14344 3956 14384
rect 4352 14344 4720 14384
rect 5068 14344 5108 14384
rect 6316 14344 6356 14384
rect 6988 14344 7028 14384
rect 9196 14344 9236 14384
rect 11884 14344 11924 14384
rect 12126 14344 12494 14384
rect 1132 14260 1172 14300
rect 652 14176 692 14216
rect 1516 14176 1555 14216
rect 1555 14176 1556 14216
rect 2956 14176 2996 14216
rect 5452 14176 5483 14216
rect 5483 14176 5492 14216
rect 5836 14176 5867 14216
rect 5867 14176 5876 14216
rect 1324 14092 1364 14132
rect 5068 14092 5108 14132
rect 1708 14008 1720 14048
rect 1720 14008 1748 14048
rect 3148 14008 3188 14048
rect 3436 14008 3476 14048
rect 4972 14008 5003 14048
rect 5003 14008 5012 14048
rect 5548 14092 5588 14132
rect 10924 14260 10964 14300
rect 12844 14260 12884 14300
rect 7180 14176 7220 14216
rect 7756 14176 7787 14216
rect 7787 14176 7796 14216
rect 6796 14092 6836 14132
rect 14476 14680 14492 14720
rect 14492 14680 14516 14720
rect 13228 14596 13268 14636
rect 29740 15268 29780 15308
rect 23116 14932 23156 14972
rect 23692 14932 23732 14972
rect 24268 14932 24308 14972
rect 25516 14932 25556 14972
rect 22060 14848 22100 14888
rect 24844 14848 24884 14888
rect 25708 14848 25748 14888
rect 21484 14764 21524 14804
rect 22252 14764 22292 14804
rect 24748 14764 24788 14804
rect 24940 14764 24980 14804
rect 25420 14764 25460 14804
rect 15244 14680 15284 14720
rect 16204 14680 16244 14720
rect 16492 14680 16532 14720
rect 16876 14680 16916 14720
rect 17740 14680 17780 14720
rect 19084 14680 19124 14720
rect 15052 14596 15092 14636
rect 15436 14596 15476 14636
rect 16012 14596 16052 14636
rect 13324 14512 13364 14552
rect 19372 14680 19412 14720
rect 21580 14680 21620 14720
rect 22156 14680 22196 14720
rect 23596 14680 23636 14720
rect 24652 14680 24692 14720
rect 27724 14848 27764 14888
rect 26284 14764 26324 14804
rect 26764 14764 26795 14804
rect 26795 14764 26804 14804
rect 26956 14764 26996 14804
rect 27436 14764 27476 14804
rect 27628 14764 27668 14804
rect 25708 14680 25748 14720
rect 27340 14680 27380 14720
rect 29260 15100 29300 15140
rect 29260 14932 29300 14972
rect 30124 14932 30164 14972
rect 30220 14764 30260 14804
rect 15628 14512 15668 14552
rect 16492 14512 16532 14552
rect 17356 14512 17396 14552
rect 19756 14596 19796 14636
rect 20524 14596 20564 14636
rect 20812 14596 20852 14636
rect 23788 14596 23819 14636
rect 23819 14596 23828 14636
rect 25420 14596 25460 14636
rect 19948 14512 19988 14552
rect 21868 14512 21908 14552
rect 14188 14428 14228 14468
rect 17068 14428 17108 14468
rect 28012 14596 28052 14636
rect 23308 14512 23348 14552
rect 26476 14512 26516 14552
rect 30700 14932 30740 14972
rect 30988 14848 31028 14888
rect 29356 14680 29396 14720
rect 29644 14596 29684 14636
rect 24652 14428 24692 14468
rect 13324 14344 13364 14384
rect 19900 14344 20268 14384
rect 27674 14344 28042 14384
rect 28876 14344 28916 14384
rect 29452 14344 29492 14384
rect 13132 14260 13172 14300
rect 13900 14260 13940 14300
rect 18604 14260 18644 14300
rect 20812 14260 20852 14300
rect 9772 14176 9812 14216
rect 10156 14176 10196 14216
rect 12748 14176 12788 14216
rect 12940 14176 12980 14216
rect 13708 14176 13748 14216
rect 15436 14176 15476 14216
rect 15916 14176 15947 14216
rect 15947 14176 15956 14216
rect 18316 14176 18356 14216
rect 19180 14176 19220 14216
rect 21388 14176 21428 14216
rect 9196 14092 9236 14132
rect 10348 14092 10388 14132
rect 11020 14092 11060 14132
rect 12268 14092 12308 14132
rect 12844 14092 12884 14132
rect 14092 14092 14132 14132
rect 14572 14092 14612 14132
rect 15628 14092 15668 14132
rect 16012 14092 16052 14132
rect 1036 13924 1076 13964
rect 4204 13924 4210 13964
rect 4210 13924 4244 13964
rect 5356 13924 5396 13964
rect 5548 13924 5588 13964
rect 652 13504 692 13544
rect 4396 13840 4436 13880
rect 6412 14008 6452 14048
rect 7468 14008 7508 14048
rect 8620 14008 8660 14048
rect 9772 14008 9812 14048
rect 10060 14008 10100 14048
rect 10444 14008 10484 14048
rect 11308 14008 11348 14048
rect 11692 14008 11713 14048
rect 11713 14008 11732 14048
rect 11980 14008 12005 14048
rect 12005 14008 12020 14048
rect 12364 14008 12404 14048
rect 13132 14008 13172 14048
rect 13804 14008 13844 14048
rect 14284 14008 14324 14048
rect 6796 13924 6836 13964
rect 7564 13924 7604 13964
rect 8524 13840 8564 13880
rect 8716 13840 8756 13880
rect 7372 13756 7403 13796
rect 7403 13756 7412 13796
rect 3112 13588 3480 13628
rect 4972 13588 5012 13628
rect 7756 13588 7796 13628
rect 8812 13588 8852 13628
rect 6796 13504 6836 13544
rect 8044 13504 8084 13544
rect 8140 13420 8171 13460
rect 8171 13420 8180 13460
rect 10540 13924 10580 13964
rect 10732 13924 10772 13964
rect 11020 13924 11060 13964
rect 12076 13924 12116 13964
rect 12940 13924 12980 13964
rect 13612 13924 13652 13964
rect 18604 14092 18644 14132
rect 19564 14092 19604 14132
rect 15052 14008 15077 14048
rect 15077 14008 15092 14048
rect 15724 14008 15764 14048
rect 15916 14008 15956 14048
rect 16492 14008 16532 14048
rect 16876 14008 16916 14048
rect 17452 14008 17492 14048
rect 18508 14008 18548 14048
rect 18700 14008 18731 14048
rect 18731 14008 18740 14048
rect 20236 14008 20276 14048
rect 20524 14008 20564 14048
rect 21484 14008 21524 14048
rect 23116 14260 23156 14300
rect 23692 14176 23732 14216
rect 25708 14176 25748 14216
rect 29644 14176 29684 14216
rect 29356 14092 29396 14132
rect 29740 14092 29780 14132
rect 30124 14092 30164 14132
rect 17740 13924 17780 13964
rect 22540 14008 22580 14048
rect 23020 14008 23060 14048
rect 23596 14008 23636 14048
rect 24268 14008 24308 14048
rect 27148 14008 27188 14048
rect 27436 14008 27476 14048
rect 28300 14008 28340 14048
rect 29164 14008 29204 14048
rect 18316 13924 18356 13964
rect 19756 13924 19796 13964
rect 20620 13924 20660 13964
rect 22636 13924 22676 13964
rect 10252 13840 10292 13880
rect 11788 13840 11828 13880
rect 12844 13840 12884 13880
rect 13516 13840 13556 13880
rect 14476 13840 14516 13880
rect 14668 13840 14708 13880
rect 15532 13840 15572 13880
rect 16396 13840 16436 13880
rect 16972 13840 17012 13880
rect 17548 13840 17588 13880
rect 21580 13840 21620 13880
rect 22156 13840 22196 13880
rect 9388 13756 9428 13796
rect 10924 13756 10964 13796
rect 15148 13756 15188 13796
rect 17740 13756 17780 13796
rect 19084 13756 19124 13796
rect 19756 13756 19796 13796
rect 22636 13756 22676 13796
rect 24364 13924 24404 13964
rect 24652 13924 24683 13964
rect 24683 13924 24692 13964
rect 26188 13924 26228 13964
rect 28876 13924 28916 13964
rect 31084 13924 31124 13964
rect 24652 13756 24692 13796
rect 25612 13756 25652 13796
rect 9772 13672 9812 13712
rect 10060 13672 10100 13712
rect 11404 13672 11444 13712
rect 22156 13672 22196 13712
rect 10886 13588 11254 13628
rect 16492 13588 16532 13628
rect 18660 13588 19028 13628
rect 23884 13588 23924 13628
rect 9100 13504 9140 13544
rect 16108 13504 16148 13544
rect 9964 13420 10004 13460
rect 13516 13420 13556 13460
rect 14380 13420 14420 13460
rect 15244 13420 15284 13460
rect 16012 13420 16052 13460
rect 6892 13336 6932 13376
rect 14572 13336 14612 13376
rect 15820 13336 15860 13376
rect 5164 13252 5204 13292
rect 5740 13252 5780 13292
rect 6028 13252 6068 13292
rect 6220 13252 6260 13292
rect 1612 13168 1652 13208
rect 2092 13168 2132 13208
rect 2572 13168 2612 13208
rect 2764 13168 2804 13208
rect 4300 13168 4340 13208
rect 940 13084 980 13124
rect 2188 13084 2228 13124
rect 1324 13000 1363 13040
rect 1363 13000 1364 13040
rect 2572 13000 2612 13040
rect 3436 13000 3476 13040
rect 4396 13000 4436 13040
rect 6796 13252 6827 13292
rect 6827 13252 6836 13292
rect 6988 13252 7028 13292
rect 9196 13252 9236 13292
rect 11500 13283 11540 13292
rect 11500 13252 11539 13283
rect 11539 13252 11540 13283
rect 8332 13210 8372 13250
rect 4972 13084 5012 13124
rect 5836 13168 5876 13208
rect 6604 13168 6644 13208
rect 7372 13168 7412 13208
rect 7852 13168 7892 13208
rect 10348 13210 10388 13250
rect 12652 13252 12692 13292
rect 15148 13252 15188 13292
rect 15436 13252 15476 13292
rect 8716 13168 8756 13208
rect 9772 13168 9812 13208
rect 10828 13168 10868 13208
rect 11404 13168 11444 13208
rect 12556 13168 12596 13208
rect 13036 13168 13076 13208
rect 14092 13168 14132 13208
rect 14572 13168 14612 13208
rect 15628 13168 15668 13208
rect 5260 13084 5300 13124
rect 4876 13000 4907 13040
rect 4907 13000 4916 13040
rect 5452 13000 5492 13040
rect 7756 13084 7796 13124
rect 8044 13084 8084 13124
rect 9484 13084 9524 13124
rect 9964 13084 10004 13124
rect 11980 13084 12011 13124
rect 12011 13084 12020 13124
rect 6028 13000 6068 13040
rect 6316 13000 6356 13040
rect 14284 13084 14324 13124
rect 8812 13000 8852 13040
rect 9100 13000 9140 13040
rect 9868 13000 9908 13040
rect 10444 13000 10484 13040
rect 11788 13000 11828 13040
rect 12364 13000 12404 13040
rect 17644 13504 17684 13544
rect 19180 13504 19220 13544
rect 19084 13420 19124 13460
rect 19564 13420 19604 13460
rect 16396 13252 16427 13292
rect 16427 13252 16436 13292
rect 26434 13588 26802 13628
rect 21100 13420 21140 13460
rect 21292 13420 21332 13460
rect 23500 13420 23531 13460
rect 23531 13420 23540 13460
rect 24364 13420 24404 13460
rect 27820 13420 27860 13460
rect 18316 13336 18356 13376
rect 18508 13252 18548 13292
rect 16780 13168 16820 13208
rect 17452 13168 17492 13208
rect 17644 13168 17684 13208
rect 18316 13168 18356 13208
rect 19084 13168 19124 13208
rect 22540 13336 22580 13376
rect 22636 13252 22676 13292
rect 20620 13168 20660 13208
rect 24076 13336 24116 13376
rect 24268 13336 24308 13376
rect 26092 13252 26132 13292
rect 26284 13252 26324 13292
rect 27148 13252 27188 13292
rect 30604 13336 30644 13376
rect 31276 13252 31316 13292
rect 22156 13168 22196 13208
rect 22444 13168 22484 13208
rect 23884 13168 23924 13208
rect 26572 13168 26584 13208
rect 26584 13168 26612 13208
rect 29356 13168 29387 13208
rect 29387 13168 29396 13208
rect 31180 13168 31220 13208
rect 15244 13084 15284 13124
rect 15532 13084 15572 13124
rect 22828 13084 22868 13124
rect 16492 13000 16532 13040
rect 20236 13000 20276 13040
rect 23116 13000 23156 13040
rect 25900 13084 25940 13124
rect 24844 13000 24884 13040
rect 25228 13000 25268 13040
rect 29740 13084 29780 13124
rect 26956 13000 26996 13040
rect 6892 12916 6932 12956
rect 8620 12916 8660 12956
rect 9388 12916 9428 12956
rect 12844 12916 12884 12956
rect 13996 12916 14036 12956
rect 14380 12916 14420 12956
rect 16204 12916 16244 12956
rect 17644 12916 17684 12956
rect 20428 12916 20468 12956
rect 23308 12916 23348 12956
rect 28588 12916 28628 12956
rect 4352 12832 4720 12872
rect 11404 12832 11444 12872
rect 12126 12832 12494 12872
rect 12652 12832 12692 12872
rect 1036 12664 1076 12704
rect 5836 12748 5876 12788
rect 6028 12664 6068 12704
rect 6316 12580 6356 12620
rect 7756 12664 7796 12704
rect 9580 12664 9611 12704
rect 9611 12664 9620 12704
rect 9964 12664 10004 12704
rect 8812 12580 8852 12620
rect 10156 12580 10196 12620
rect 1324 12496 1364 12536
rect 1708 12496 1748 12536
rect 2284 12496 2324 12536
rect 3916 12496 3956 12536
rect 5068 12496 5108 12536
rect 5836 12496 5876 12536
rect 6700 12496 6740 12536
rect 7468 12496 7508 12536
rect 8620 12496 8660 12536
rect 9196 12496 9236 12536
rect 9388 12496 9428 12536
rect 1516 12412 1556 12452
rect 2092 12412 2132 12452
rect 4876 12412 4916 12452
rect 6892 12412 6932 12452
rect 8044 12412 8084 12452
rect 8620 12412 8660 12452
rect 8812 12412 8852 12452
rect 9676 12412 9716 12452
rect 9964 12412 10004 12452
rect 5068 12328 5108 12368
rect 5740 12328 5780 12368
rect 6604 12328 6644 12368
rect 8908 12328 8948 12368
rect 14092 12748 14132 12788
rect 19900 12832 20268 12872
rect 21196 12832 21236 12872
rect 24076 12832 24116 12872
rect 27674 12832 28042 12872
rect 28396 12748 28436 12788
rect 30316 12748 30356 12788
rect 10732 12664 10772 12704
rect 11692 12664 11732 12704
rect 13324 12664 13364 12704
rect 14572 12664 14612 12704
rect 16780 12664 16820 12704
rect 18412 12664 18452 12704
rect 11788 12580 11828 12620
rect 12268 12580 12308 12620
rect 12652 12580 12692 12620
rect 15532 12580 15572 12620
rect 16492 12580 16532 12620
rect 17452 12580 17492 12620
rect 18028 12580 18068 12620
rect 10924 12496 10964 12536
rect 11116 12496 11156 12536
rect 12172 12496 12212 12536
rect 12940 12496 12980 12536
rect 13516 12496 13556 12536
rect 13804 12496 13844 12536
rect 13996 12496 14036 12536
rect 14476 12496 14516 12536
rect 15052 12496 15092 12536
rect 15436 12496 15476 12536
rect 4972 12244 5012 12284
rect 9964 12244 10004 12284
rect 8332 12160 8372 12200
rect 9868 12160 9908 12200
rect 11404 12412 11444 12452
rect 11500 12328 11540 12368
rect 15820 12496 15860 12536
rect 16204 12496 16244 12536
rect 17164 12496 17204 12536
rect 18316 12496 18356 12536
rect 13324 12412 13364 12452
rect 14380 12412 14420 12452
rect 16396 12412 16436 12452
rect 16972 12412 17012 12452
rect 17644 12412 17684 12452
rect 18508 12496 18548 12536
rect 22444 12664 22484 12704
rect 29260 12664 29300 12704
rect 22924 12580 22964 12620
rect 21676 12496 21716 12536
rect 23116 12496 23156 12536
rect 18412 12412 18452 12452
rect 19468 12412 19508 12452
rect 20524 12412 20564 12452
rect 15244 12328 15275 12368
rect 15275 12328 15284 12368
rect 16876 12328 16916 12368
rect 17356 12328 17396 12368
rect 20140 12328 20180 12368
rect 11308 12244 11348 12284
rect 15820 12244 15860 12284
rect 20428 12244 20468 12284
rect 21100 12244 21140 12284
rect 11500 12160 11540 12200
rect 3112 12076 3480 12116
rect 5740 12076 5780 12116
rect 6124 12076 6164 12116
rect 9100 12076 9140 12116
rect 10886 12076 11254 12116
rect 13036 12076 13076 12116
rect 17068 12076 17108 12116
rect 18412 12076 18452 12116
rect 18660 12076 19028 12116
rect 19180 12076 19220 12116
rect 21580 12076 21620 12116
rect 9964 11992 10004 12032
rect 13228 11992 13268 12032
rect 13516 11992 13556 12032
rect 2092 11908 2132 11948
rect 3916 11908 3956 11948
rect 4876 11908 4916 11948
rect 5740 11908 5780 11948
rect 6796 11908 6836 11948
rect 7180 11908 7220 11948
rect 9484 11908 9515 11948
rect 9515 11908 9524 11948
rect 11596 11908 11636 11948
rect 1420 11824 1460 11864
rect 5836 11740 5876 11780
rect 7084 11740 7124 11780
rect 7372 11740 7412 11780
rect 2188 11656 2228 11696
rect 2668 11656 2708 11696
rect 3532 11656 3572 11696
rect 4012 11656 4052 11696
rect 10348 11824 10388 11864
rect 11884 11824 11924 11864
rect 13708 11908 13748 11948
rect 14860 11908 14900 11948
rect 9868 11740 9908 11780
rect 4876 11656 4916 11696
rect 5740 11656 5780 11696
rect 6028 11656 6068 11696
rect 6316 11656 6347 11696
rect 6347 11656 6356 11696
rect 8908 11656 8948 11696
rect 9964 11696 10004 11717
rect 13516 11824 13556 11864
rect 14380 11824 14420 11864
rect 11788 11740 11828 11780
rect 13228 11740 13268 11780
rect 14860 11740 14900 11780
rect 15244 11740 15284 11780
rect 15436 11740 15476 11780
rect 9964 11677 10004 11696
rect 10252 11656 10292 11696
rect 11308 11656 11348 11696
rect 12364 11656 12404 11696
rect 12652 11656 12692 11696
rect 13516 11656 13523 11696
rect 13523 11656 13556 11696
rect 16108 11992 16148 12032
rect 16876 11992 16916 12032
rect 19564 11992 19604 12032
rect 16588 11908 16628 11948
rect 17164 11908 17204 11948
rect 18220 11908 18260 11948
rect 18508 11908 18548 11948
rect 16108 11740 16148 11780
rect 16876 11740 16916 11780
rect 15820 11656 15860 11696
rect 17068 11677 17108 11717
rect 19084 11908 19124 11948
rect 20908 11908 20948 11948
rect 20716 11824 20756 11864
rect 19756 11740 19796 11780
rect 20908 11740 20948 11780
rect 21676 11908 21716 11948
rect 22636 12412 22676 12452
rect 22828 12412 22867 12452
rect 22867 12412 22868 12452
rect 23884 12412 23915 12452
rect 23915 12412 23924 12452
rect 26284 12580 26324 12620
rect 28396 12580 28436 12620
rect 28588 12580 28628 12620
rect 29548 12580 29588 12620
rect 25708 12496 25748 12536
rect 27244 12496 27284 12536
rect 31660 12496 31700 12536
rect 25900 12412 25940 12452
rect 26188 12412 26228 12452
rect 28300 12412 28340 12452
rect 28684 12412 28724 12452
rect 29548 12412 29588 12452
rect 29740 12412 29780 12452
rect 30124 12412 30164 12452
rect 31372 12412 31412 12452
rect 30700 12328 30740 12368
rect 28588 12244 28628 12284
rect 30508 12160 30548 12200
rect 26434 12076 26802 12116
rect 26956 12076 26996 12116
rect 28876 12076 28916 12116
rect 24076 11908 24116 11948
rect 24172 11824 24212 11864
rect 21100 11740 21140 11780
rect 24460 11824 24500 11864
rect 25132 11740 25172 11780
rect 29068 11908 29108 11948
rect 29932 11908 29972 11948
rect 30700 11908 30740 11948
rect 27532 11824 27572 11864
rect 29260 11824 29300 11864
rect 29548 11824 29588 11864
rect 30316 11824 30356 11864
rect 30892 11824 30932 11864
rect 25516 11740 25556 11780
rect 26668 11740 26708 11780
rect 28204 11740 28244 11780
rect 29068 11740 29108 11780
rect 29452 11740 29492 11780
rect 30412 11740 30452 11780
rect 17740 11656 17771 11696
rect 17771 11656 17780 11696
rect 18412 11656 18414 11696
rect 18414 11656 18452 11696
rect 19180 11656 19220 11696
rect 20620 11656 20660 11696
rect 22636 11656 22676 11696
rect 23116 11656 23156 11696
rect 23500 11656 23531 11696
rect 23531 11656 23540 11696
rect 24652 11656 24692 11696
rect 26476 11656 26516 11696
rect 27340 11656 27380 11696
rect 27916 11656 27956 11696
rect 28396 11656 28436 11696
rect 31756 11656 31796 11696
rect 1324 11572 1364 11612
rect 1516 11572 1556 11612
rect 1708 11572 1748 11612
rect 2764 11572 2804 11612
rect 5068 11572 5108 11612
rect 5548 11572 5588 11612
rect 5932 11572 5972 11612
rect 7660 11572 7700 11612
rect 8716 11572 8756 11612
rect 9196 11572 9236 11612
rect 10348 11572 10388 11612
rect 10636 11572 10676 11612
rect 11884 11572 11924 11612
rect 12076 11572 12116 11612
rect 1036 11488 1076 11528
rect 1228 11488 1268 11528
rect 3532 11488 3572 11528
rect 4204 11488 4244 11528
rect 2956 11404 2996 11444
rect 4876 11488 4916 11528
rect 6220 11488 6260 11528
rect 7948 11488 7988 11528
rect 8140 11488 8180 11528
rect 9100 11488 9140 11528
rect 10156 11488 10196 11528
rect 10732 11488 10772 11528
rect 10924 11488 10964 11528
rect 11500 11488 11540 11528
rect 12268 11488 12308 11528
rect 13036 11404 13076 11444
rect 13420 11572 13460 11612
rect 14092 11572 14132 11612
rect 15148 11572 15188 11612
rect 15436 11572 15476 11612
rect 16012 11572 16052 11612
rect 16204 11572 16244 11612
rect 16492 11572 16532 11612
rect 13516 11488 13556 11528
rect 18508 11572 18548 11612
rect 23404 11572 23444 11612
rect 25900 11572 25940 11612
rect 28876 11572 28916 11612
rect 31468 11572 31508 11612
rect 16588 11488 16628 11528
rect 16780 11488 16820 11528
rect 18700 11488 18740 11528
rect 26380 11488 26411 11528
rect 26411 11488 26420 11528
rect 27436 11488 27476 11528
rect 29932 11488 29972 11528
rect 24268 11404 24308 11444
rect 25036 11404 25076 11444
rect 1708 11320 1748 11360
rect 4352 11320 4720 11360
rect 6412 11320 6452 11360
rect 12126 11320 12494 11360
rect 12940 11320 12980 11360
rect 19900 11320 20268 11360
rect 21676 11320 21716 11360
rect 25516 11320 25556 11360
rect 27674 11320 28042 11360
rect 652 11236 692 11276
rect 2188 11236 2228 11276
rect 9964 11236 10004 11276
rect 19372 11236 19412 11276
rect 25036 11236 25076 11276
rect 2284 11152 2324 11192
rect 5932 11152 5963 11192
rect 5963 11152 5972 11192
rect 7660 11152 7700 11192
rect 8812 11152 8852 11192
rect 10252 11152 10292 11192
rect 10924 11152 10964 11192
rect 11884 11152 11924 11192
rect 13324 11152 13364 11192
rect 13804 11152 13844 11192
rect 14860 11152 14900 11192
rect 15148 11152 15188 11192
rect 16012 11152 16052 11192
rect 17740 11152 17780 11192
rect 18412 11152 18443 11192
rect 18443 11152 18452 11192
rect 18700 11152 18740 11192
rect 20620 11152 20660 11192
rect 23404 11152 23444 11192
rect 26668 11152 26708 11192
rect 27340 11152 27380 11192
rect 2956 11068 2996 11108
rect 5164 11068 5204 11108
rect 6700 11068 6740 11108
rect 8044 11068 8084 11108
rect 9868 11068 9908 11108
rect 10156 11068 10196 11108
rect 11500 11068 11540 11108
rect 13612 11068 13652 11108
rect 13900 11068 13940 11108
rect 15628 11068 15668 11108
rect 1228 10984 1268 11024
rect 2668 10984 2708 11024
rect 4204 10984 4244 11024
rect 5068 10984 5108 11024
rect 5548 10984 5588 11024
rect 7180 10984 7201 11024
rect 7201 10984 7220 11024
rect 7468 10984 7493 11024
rect 7493 10984 7508 11024
rect 7948 10984 7973 11024
rect 7973 10984 7988 11024
rect 8524 10984 8564 11024
rect 8908 10984 8948 11024
rect 9580 10984 9620 11024
rect 11212 10984 11252 11024
rect 940 10900 980 10940
rect 940 10396 980 10436
rect 11980 10984 12020 11024
rect 12748 10984 12788 11024
rect 2572 10900 2612 10940
rect 4972 10900 5003 10940
rect 5003 10900 5012 10940
rect 5740 10900 5771 10940
rect 5771 10900 5780 10940
rect 6028 10900 6068 10940
rect 6988 10900 7028 10940
rect 7372 10900 7412 10940
rect 7660 10900 7700 10940
rect 8620 10900 8643 10940
rect 8643 10900 8660 10940
rect 12652 10900 12692 10940
rect 18028 11068 18068 11108
rect 21580 11068 21620 11108
rect 13516 10984 13545 11024
rect 13545 10984 13556 11024
rect 5068 10816 5108 10856
rect 8428 10816 8468 10856
rect 14188 10984 14228 11024
rect 15532 10984 15543 11024
rect 15543 10984 15572 11024
rect 16876 10984 16916 11024
rect 17452 10984 17492 11024
rect 13036 10900 13076 10940
rect 13900 10900 13940 10940
rect 16972 10900 17012 10940
rect 3532 10732 3572 10772
rect 7180 10732 7220 10772
rect 12556 10732 12596 10772
rect 7564 10648 7604 10688
rect 12748 10648 12788 10688
rect 3112 10564 3480 10604
rect 5644 10564 5684 10604
rect 9580 10564 9620 10604
rect 10886 10564 11254 10604
rect 8524 10480 8564 10520
rect 940 10228 980 10268
rect 1708 10228 1748 10268
rect 2476 10228 2516 10268
rect 5548 10396 5588 10436
rect 6316 10396 6356 10436
rect 7660 10396 7700 10436
rect 8908 10396 8948 10436
rect 6220 10312 6260 10352
rect 4108 10228 4148 10268
rect 7180 10228 7211 10268
rect 7211 10228 7220 10268
rect 8908 10228 8948 10268
rect 1420 10144 1460 10184
rect 1804 10144 1844 10184
rect 2092 10144 2132 10184
rect 3532 10144 3539 10184
rect 3539 10144 3572 10184
rect 5068 10144 5108 10184
rect 5644 10144 5684 10184
rect 652 10060 692 10100
rect 1036 10060 1076 10100
rect 2476 10060 2516 10100
rect 2092 9976 2132 10016
rect 2860 10060 2891 10100
rect 2891 10060 2900 10100
rect 3436 10060 3476 10100
rect 3052 9892 3092 9932
rect 3820 9892 3860 9932
rect 5260 10060 5300 10100
rect 10156 10396 10187 10436
rect 10187 10396 10196 10436
rect 16780 10396 16820 10436
rect 11980 10228 12019 10268
rect 12019 10228 12020 10268
rect 12652 10228 12692 10268
rect 12940 10228 12980 10268
rect 23020 11068 23060 11108
rect 24556 11068 24596 11108
rect 25132 11068 25172 11108
rect 26380 11068 26420 11108
rect 17836 10984 17876 11024
rect 19564 10984 19604 11024
rect 20716 10984 20756 11024
rect 21196 10984 21236 11024
rect 22060 10984 22100 11024
rect 18220 10900 18260 10940
rect 22540 10984 22580 11024
rect 23212 11015 23252 11024
rect 19468 10900 19508 10940
rect 23212 10984 23243 11015
rect 23243 10984 23252 11015
rect 23596 10984 23636 11024
rect 24460 11015 24500 11024
rect 24460 10984 24500 11015
rect 23980 10900 24020 10940
rect 18124 10816 18164 10856
rect 19084 10816 19124 10856
rect 20140 10816 20180 10856
rect 22540 10732 22580 10772
rect 18412 10648 18452 10688
rect 19180 10648 19220 10688
rect 19372 10648 19412 10688
rect 18660 10564 19028 10604
rect 21580 10564 21620 10604
rect 17740 10480 17780 10520
rect 23692 10480 23732 10520
rect 25612 10984 25652 11024
rect 27820 10984 27860 11024
rect 28588 10984 28628 11024
rect 24364 10816 24404 10856
rect 24844 10816 24884 10856
rect 25132 10816 25172 10856
rect 26284 10900 26324 10940
rect 27436 10900 27476 10940
rect 30124 11320 30164 11360
rect 28972 11236 29012 11276
rect 29452 11152 29492 11192
rect 29836 11152 29876 11192
rect 30124 11152 30164 11192
rect 29548 11068 29588 11108
rect 29260 10984 29300 11024
rect 29644 10900 29684 10940
rect 29836 10900 29876 10940
rect 26860 10816 26900 10856
rect 30412 10816 30452 10856
rect 30796 10816 30836 10856
rect 26092 10732 26132 10772
rect 21580 10396 21620 10436
rect 25036 10396 25076 10436
rect 20236 10312 20276 10352
rect 21004 10312 21044 10352
rect 22732 10312 22772 10352
rect 17164 10228 17204 10268
rect 17548 10228 17588 10268
rect 18220 10228 18260 10268
rect 19468 10228 19508 10268
rect 19660 10228 19700 10268
rect 21196 10228 21236 10268
rect 22540 10228 22580 10268
rect 26434 10564 26802 10604
rect 27820 10396 27851 10436
rect 27851 10396 27860 10436
rect 27532 10312 27572 10352
rect 28492 10312 28532 10352
rect 30412 10312 30452 10352
rect 30796 10312 30836 10352
rect 25900 10228 25940 10268
rect 26764 10228 26804 10268
rect 27052 10228 27092 10268
rect 6604 10144 6644 10184
rect 7276 10144 7316 10184
rect 7948 10144 7988 10184
rect 8140 10144 8180 10184
rect 8428 10144 8468 10184
rect 8812 10144 8852 10184
rect 9004 10144 9044 10184
rect 9868 10144 9908 10184
rect 11308 10144 11348 10184
rect 11884 10144 11924 10184
rect 12748 10144 12788 10184
rect 13420 10144 13460 10184
rect 13708 10144 13736 10184
rect 13736 10144 13748 10184
rect 14476 10144 14516 10184
rect 15148 10144 15188 10184
rect 15628 10144 15668 10184
rect 16012 10144 16052 10184
rect 17644 10144 17684 10184
rect 17836 10144 17861 10184
rect 17861 10144 17876 10184
rect 18508 10144 18548 10184
rect 19372 10144 19403 10184
rect 19403 10144 19412 10184
rect 19756 10144 19796 10184
rect 21292 10144 21332 10184
rect 21676 10144 21716 10184
rect 22444 10144 22484 10184
rect 23116 10144 23156 10184
rect 23500 10144 23540 10184
rect 23788 10144 23828 10184
rect 24076 10144 24116 10184
rect 24364 10144 24368 10184
rect 24368 10144 24404 10184
rect 9388 10060 9428 10100
rect 13036 10060 13076 10100
rect 15820 10060 15860 10100
rect 4972 9976 5012 10016
rect 7660 9976 7700 10016
rect 8140 9976 8180 10016
rect 10156 9976 10196 10016
rect 10828 9976 10868 10016
rect 13996 9976 14036 10016
rect 18124 10060 18164 10100
rect 18316 10060 18356 10100
rect 20620 10060 20660 10100
rect 17836 9976 17876 10016
rect 21676 9976 21716 10016
rect 22348 9976 22388 10016
rect 22636 9976 22676 10016
rect 23788 9976 23828 10016
rect 26764 9976 26804 10016
rect 4876 9892 4916 9932
rect 7180 9892 7220 9932
rect 8524 9892 8564 9932
rect 16396 9892 16436 9932
rect 17548 9892 17588 9932
rect 18412 9892 18452 9932
rect 4352 9808 4720 9848
rect 5452 9808 5492 9848
rect 12126 9808 12494 9848
rect 28108 9976 28148 10016
rect 28684 9976 28724 10016
rect 26956 9892 26996 9932
rect 19900 9808 20268 9848
rect 27674 9808 28042 9848
rect 1516 9724 1556 9764
rect 2476 9724 2516 9764
rect 4108 9724 4148 9764
rect 8812 9724 8852 9764
rect 1804 9640 1844 9680
rect 3148 9640 3188 9680
rect 5164 9640 5204 9680
rect 7276 9640 7316 9680
rect 8620 9640 8660 9680
rect 9004 9640 9044 9680
rect 10444 9640 10484 9680
rect 3820 9556 3860 9596
rect 4108 9556 4148 9596
rect 6604 9556 6644 9596
rect 7180 9556 7220 9596
rect 7948 9556 7988 9596
rect 15916 9724 15956 9764
rect 13708 9640 13739 9680
rect 13739 9640 13748 9680
rect 14476 9640 14516 9680
rect 11980 9556 12020 9596
rect 12364 9556 12404 9596
rect 14188 9556 14228 9596
rect 15148 9640 15188 9680
rect 15628 9640 15668 9680
rect 17644 9640 17684 9680
rect 15532 9556 15572 9596
rect 23116 9724 23156 9764
rect 23692 9724 23732 9764
rect 20908 9640 20939 9680
rect 20939 9640 20948 9680
rect 23404 9640 23444 9680
rect 23596 9640 23636 9680
rect 25804 9640 25843 9680
rect 25843 9640 25844 9680
rect 25996 9640 26036 9680
rect 27532 9640 27572 9680
rect 19372 9556 19412 9596
rect 652 9472 692 9512
rect 1516 9472 1556 9512
rect 2668 9472 2708 9512
rect 3532 9472 3572 9512
rect 4684 9472 4724 9512
rect 5068 9472 5108 9512
rect 5932 9472 5972 9512
rect 6220 9472 6260 9512
rect 6412 9472 6452 9512
rect 6700 9472 6740 9512
rect 6988 9472 7028 9512
rect 7372 9472 7412 9512
rect 7660 9472 7700 9512
rect 8236 9472 8276 9512
rect 8524 9472 8564 9512
rect 9100 9472 9140 9512
rect 9388 9472 9428 9512
rect 10348 9472 10388 9512
rect 11308 9472 11348 9512
rect 11884 9472 11924 9512
rect 13036 9472 13076 9512
rect 13420 9472 13460 9512
rect 13900 9472 13940 9512
rect 14572 9472 14612 9512
rect 15628 9472 15668 9512
rect 16396 9472 16436 9512
rect 18124 9472 18164 9512
rect 1324 9388 1364 9428
rect 2476 9388 2516 9428
rect 2956 9388 2996 9428
rect 3148 9388 3188 9428
rect 2092 9304 2132 9344
rect 2668 9220 2708 9260
rect 5260 9388 5291 9428
rect 5291 9388 5300 9428
rect 7468 9388 7508 9428
rect 9772 9388 9812 9428
rect 4300 9304 4340 9344
rect 4588 9304 4628 9344
rect 5452 9304 5492 9344
rect 9100 9304 9140 9344
rect 9388 9304 9428 9344
rect 10732 9388 10772 9428
rect 12364 9388 12404 9428
rect 13708 9388 13748 9428
rect 3724 9220 3764 9260
rect 6700 9220 6740 9260
rect 6124 9136 6164 9176
rect 3112 9052 3480 9092
rect 9580 8968 9620 9008
rect 556 8884 596 8924
rect 2572 8884 2612 8924
rect 4684 8884 4724 8924
rect 5836 8884 5876 8924
rect 10636 8884 10676 8924
rect 940 8800 980 8840
rect 3724 8800 3764 8840
rect 6988 8800 7028 8840
rect 9100 8800 9140 8840
rect 1996 8716 2036 8756
rect 4588 8716 4628 8756
rect 5260 8716 5300 8756
rect 6604 8716 6644 8756
rect 9676 8716 9716 8756
rect 3052 8632 3092 8672
rect 3340 8632 3369 8672
rect 3369 8632 3380 8672
rect 3628 8632 3668 8672
rect 3916 8632 3956 8672
rect 5452 8632 5492 8672
rect 7180 8632 7220 8672
rect 7372 8639 7376 8679
rect 7376 8639 7412 8679
rect 10886 9052 11254 9092
rect 15148 9388 15188 9428
rect 16108 9388 16148 9428
rect 16780 9388 16820 9428
rect 17260 9388 17300 9428
rect 13900 9304 13940 9344
rect 14572 9304 14612 9344
rect 15820 9304 15860 9344
rect 22636 9556 22676 9596
rect 23788 9556 23828 9596
rect 24940 9556 24980 9596
rect 25900 9556 25940 9596
rect 26284 9556 26324 9596
rect 27340 9556 27380 9596
rect 19468 9472 19508 9512
rect 19852 9472 19892 9512
rect 21196 9472 21236 9512
rect 21964 9472 22004 9512
rect 23212 9472 23243 9512
rect 23243 9472 23252 9512
rect 23500 9472 23540 9512
rect 25420 9472 25460 9512
rect 17452 9388 17492 9428
rect 20332 9388 20372 9428
rect 21868 9388 21874 9428
rect 21874 9388 21908 9428
rect 23020 9388 23060 9428
rect 17260 9220 17300 9260
rect 19468 9220 19508 9260
rect 21676 9136 21716 9176
rect 18660 9052 19028 9092
rect 11884 8968 11924 9008
rect 13132 8968 13172 9008
rect 19180 8968 19220 9008
rect 21868 8968 21908 9008
rect 15916 8884 15956 8924
rect 17260 8884 17291 8924
rect 17291 8884 17300 8924
rect 19756 8884 19796 8924
rect 10828 8800 10868 8840
rect 13036 8800 13076 8840
rect 19660 8800 19700 8840
rect 11308 8716 11348 8756
rect 12364 8716 12404 8756
rect 15052 8716 15092 8756
rect 15436 8716 15476 8756
rect 15820 8716 15860 8756
rect 16780 8716 16820 8756
rect 7660 8632 7700 8672
rect 8236 8632 8276 8672
rect 9484 8632 9524 8672
rect 9868 8632 9908 8672
rect 10444 8632 10484 8672
rect 5068 8548 5108 8588
rect 460 8464 500 8504
rect 4300 8464 4340 8504
rect 4876 8464 4916 8504
rect 5260 8464 5300 8504
rect 4352 8296 4720 8336
rect 8140 8548 8180 8588
rect 9388 8548 9428 8588
rect 9676 8548 9716 8588
rect 9196 8464 9236 8504
rect 11212 8548 11252 8588
rect 3532 8212 3572 8252
rect 7468 8212 7508 8252
rect 9868 8212 9908 8252
rect 652 8128 692 8168
rect 3628 8128 3668 8168
rect 3916 8128 3956 8168
rect 4972 8128 5012 8168
rect 5644 8128 5684 8168
rect 7372 8128 7412 8168
rect 844 8044 884 8084
rect 3820 8044 3860 8084
rect 9100 8128 9131 8168
rect 9131 8128 9140 8168
rect 9676 8128 9716 8168
rect 10732 8464 10772 8504
rect 11692 8464 11723 8504
rect 11723 8464 11732 8504
rect 19468 8716 19508 8756
rect 21772 8884 21812 8924
rect 21964 8884 22004 8924
rect 23020 8884 23060 8924
rect 22828 8800 22868 8840
rect 24652 8800 24692 8840
rect 22732 8716 22772 8756
rect 25708 9472 25748 9512
rect 25996 9472 26008 9512
rect 26008 9472 26036 9512
rect 27052 9472 27092 9512
rect 27532 9472 27572 9512
rect 28684 9472 28724 9512
rect 29356 9472 29387 9512
rect 29387 9472 29396 9512
rect 25324 9304 25364 9344
rect 26956 9388 26996 9428
rect 27244 9388 27284 9428
rect 28492 9388 28532 9428
rect 26860 9220 26900 9260
rect 26434 9052 26802 9092
rect 25612 8716 25652 8756
rect 25996 8716 26036 8756
rect 12268 8632 12299 8672
rect 12299 8632 12308 8672
rect 13708 8632 13748 8672
rect 14764 8632 14804 8672
rect 17932 8632 17972 8672
rect 19180 8632 19220 8672
rect 21676 8632 21716 8672
rect 22924 8632 22964 8672
rect 24556 8632 24596 8672
rect 24844 8632 24884 8672
rect 25420 8632 25460 8672
rect 27436 8632 27476 8672
rect 28108 8632 28148 8672
rect 12844 8464 12884 8504
rect 15916 8548 15956 8588
rect 16204 8548 16244 8588
rect 16684 8548 16724 8588
rect 18220 8548 18260 8588
rect 19756 8548 19796 8588
rect 19948 8548 19988 8588
rect 20620 8548 20660 8588
rect 20908 8548 20919 8588
rect 20919 8548 20948 8588
rect 21100 8548 21131 8588
rect 21131 8548 21140 8588
rect 13996 8464 14036 8504
rect 15436 8464 15476 8504
rect 18796 8464 18836 8504
rect 22156 8464 22196 8504
rect 15052 8380 15092 8420
rect 26860 8548 26900 8588
rect 27148 8548 27188 8588
rect 26092 8464 26132 8504
rect 24652 8380 24692 8420
rect 12126 8296 12494 8336
rect 19372 8296 19412 8336
rect 19900 8296 20268 8336
rect 27674 8296 28042 8336
rect 17548 8212 17588 8252
rect 24844 8212 24884 8252
rect 11404 8128 11444 8168
rect 12652 8128 12692 8168
rect 13132 8128 13172 8168
rect 8236 8044 8276 8084
rect 11596 8044 11636 8084
rect 12268 8044 12308 8084
rect 13324 8044 13364 8084
rect 15916 8128 15956 8168
rect 16204 8128 16235 8168
rect 16235 8128 16244 8168
rect 14764 8044 14804 8084
rect 18028 8128 18068 8168
rect 16780 8044 16820 8084
rect 19756 8128 19796 8168
rect 20428 8128 20468 8168
rect 21100 8128 21140 8168
rect 18796 8044 18836 8084
rect 22156 8044 22187 8084
rect 22187 8044 22196 8084
rect 23980 8044 24020 8084
rect 268 7935 308 7975
rect 940 7960 980 8000
rect 2956 7960 2996 8000
rect 3916 7960 3956 8000
rect 4972 7960 4993 8000
rect 4993 7960 5012 8000
rect 5260 7960 5285 8000
rect 5285 7960 5300 8000
rect 6604 7960 6644 8000
rect 7180 7960 7220 8000
rect 7372 7960 7412 8000
rect 8428 7960 8468 8000
rect 8812 7960 8852 8000
rect 9580 7960 9620 8000
rect 10252 7960 10292 8000
rect 10636 7960 10676 8000
rect 11404 7960 11444 8000
rect 12076 7960 12116 8000
rect 13036 7960 13076 8000
rect 13228 7960 13268 8000
rect 13708 7960 13731 8000
rect 13731 7960 13748 8000
rect 15148 7960 15188 8000
rect 16684 7960 16724 8000
rect 17164 7960 17204 8000
rect 17644 7960 17684 8000
rect 18220 7960 18260 8000
rect 19372 7960 19412 8000
rect 2860 7876 2900 7916
rect 4876 7876 4916 7916
rect 8332 7876 8372 7916
rect 9196 7876 9236 7916
rect 10156 7876 10196 7916
rect 11212 7876 11252 7916
rect 11788 7876 11828 7916
rect 12844 7876 12875 7916
rect 12875 7876 12884 7916
rect 13420 7876 13460 7916
rect 15820 7876 15860 7916
rect 1996 7792 2036 7832
rect 7180 7792 7220 7832
rect 8140 7792 8180 7832
rect 9580 7792 9620 7832
rect 11500 7792 11540 7832
rect 5932 7708 5972 7748
rect 6892 7708 6932 7748
rect 8044 7708 8084 7748
rect 8620 7708 8660 7748
rect 9484 7708 9524 7748
rect 10060 7708 10100 7748
rect 14668 7708 14699 7748
rect 14699 7708 14708 7748
rect 14956 7708 14996 7748
rect 9676 7624 9716 7664
rect 11404 7624 11444 7664
rect 3112 7540 3480 7580
rect 10886 7540 11254 7580
rect 18660 7540 19028 7580
rect 9388 7456 9428 7496
rect 24172 8044 24212 8084
rect 24364 8044 24404 8084
rect 24652 8044 24692 8084
rect 28108 8128 28148 8168
rect 26092 8044 26132 8084
rect 20428 7960 20468 8000
rect 21388 7960 21428 8000
rect 21772 7960 21812 8000
rect 22828 7960 22868 8000
rect 23308 7960 23348 8000
rect 23788 7960 23819 8000
rect 23819 7960 23828 8000
rect 25324 7960 25364 8000
rect 26188 7960 26219 8000
rect 26219 7960 26228 8000
rect 20812 7876 20852 7916
rect 23692 7876 23732 7916
rect 24844 7876 24884 7916
rect 25036 7876 25076 7916
rect 20620 7708 20660 7748
rect 20428 7456 20468 7496
rect 172 7372 212 7412
rect 6028 7372 6068 7412
rect 7180 7372 7220 7412
rect 9196 7372 9236 7412
rect 10252 7372 10292 7412
rect 17164 7372 17204 7412
rect 19276 7372 19316 7412
rect 20812 7372 20852 7412
rect 23404 7792 23444 7832
rect 24940 7792 24980 7832
rect 24364 7708 24404 7748
rect 24556 7708 24596 7748
rect 26764 7708 26804 7748
rect 26434 7540 26802 7580
rect 3628 7288 3668 7328
rect 4204 7288 4244 7328
rect 2476 7204 2516 7244
rect 3916 7204 3956 7244
rect 2860 7120 2900 7160
rect 9388 7288 9428 7328
rect 20908 7288 20948 7328
rect 22348 7319 22388 7328
rect 22348 7288 22380 7319
rect 22380 7288 22388 7319
rect 22732 7288 22772 7328
rect 5644 7204 5684 7244
rect 8044 7204 8084 7244
rect 9484 7204 9524 7244
rect 9772 7204 9812 7244
rect 13420 7204 13460 7244
rect 16012 7204 16052 7244
rect 16300 7204 16340 7244
rect 16684 7204 16724 7244
rect 19660 7204 19700 7244
rect 22252 7204 22292 7244
rect 23596 7204 23636 7244
rect 25516 7204 25556 7244
rect 26860 7204 26900 7244
rect 27340 7204 27380 7244
rect 3628 7120 3668 7160
rect 4012 7120 4052 7160
rect 5068 7120 5108 7160
rect 6892 7193 6932 7202
rect 6892 7162 6932 7193
rect 8332 7120 8363 7160
rect 8363 7120 8372 7160
rect 8620 7120 8631 7160
rect 8631 7120 8660 7160
rect 9100 7120 9140 7160
rect 11116 7120 11156 7160
rect 11692 7120 11732 7160
rect 12652 7120 12692 7160
rect 13324 7120 13364 7160
rect 14668 7120 14708 7160
rect 4108 7036 4148 7076
rect 6124 7036 6164 7076
rect 2572 6952 2612 6992
rect 3916 6952 3956 6992
rect 3340 6868 3380 6908
rect 748 6784 788 6824
rect 4352 6784 4720 6824
rect 3052 6616 3092 6656
rect 5068 6616 5108 6656
rect 2956 6532 2996 6572
rect 6412 6952 6452 6992
rect 6988 6532 7028 6572
rect 2572 6448 2597 6488
rect 2597 6448 2612 6488
rect 4780 6448 4820 6488
rect 5452 6448 5492 6488
rect 5932 6448 5972 6488
rect 6412 6448 6452 6488
rect 6700 6448 6740 6488
rect 7276 6448 7307 6488
rect 7307 6448 7316 6488
rect 1132 6364 1172 6404
rect 2284 6364 2324 6404
rect 2668 6364 2708 6404
rect 4204 6364 4244 6404
rect 5548 6364 5588 6404
rect 5740 6364 5780 6404
rect 8428 6952 8459 6992
rect 8459 6952 8468 6992
rect 10444 6952 10484 6992
rect 9868 6700 9908 6740
rect 9484 6616 9524 6656
rect 9292 6532 9332 6572
rect 14956 7036 14996 7076
rect 11596 6952 11636 6992
rect 12126 6784 12494 6824
rect 16396 7120 16436 7160
rect 17068 7120 17108 7160
rect 19276 7120 19316 7160
rect 20524 7120 20564 7160
rect 21772 7120 21812 7160
rect 22156 7120 22196 7160
rect 23212 7120 23252 7160
rect 24268 7120 24308 7160
rect 25420 7120 25460 7160
rect 25996 7120 26036 7160
rect 26380 7120 26420 7160
rect 27244 7120 27275 7160
rect 27275 7120 27284 7160
rect 15436 7036 15465 7076
rect 15465 7036 15476 7076
rect 17548 7036 17588 7076
rect 16972 6952 17012 6992
rect 17164 6868 17204 6908
rect 14572 6700 14612 6740
rect 13996 6532 14036 6572
rect 14380 6532 14420 6572
rect 8044 6448 8084 6488
rect 8524 6448 8564 6488
rect 9676 6448 9716 6488
rect 9964 6448 10004 6488
rect 10444 6448 10484 6488
rect 11596 6448 11636 6488
rect 11884 6448 11924 6488
rect 12172 6448 12212 6488
rect 19564 7036 19604 7076
rect 16108 6616 16148 6656
rect 16876 6616 16916 6656
rect 18988 6616 19028 6656
rect 15820 6532 15860 6572
rect 16396 6532 16436 6572
rect 21388 7036 21428 7076
rect 21868 7036 21908 7076
rect 22348 7036 22388 7076
rect 23020 7036 23060 7076
rect 23404 7036 23444 7076
rect 27148 7036 27188 7076
rect 27436 7036 27476 7076
rect 22156 6952 22196 6992
rect 23980 6952 24020 6992
rect 21772 6868 21812 6908
rect 19900 6784 20268 6824
rect 21004 6700 21044 6740
rect 12844 6448 12884 6488
rect 13036 6448 13076 6488
rect 14476 6448 14516 6488
rect 9484 6364 9524 6404
rect 10636 6364 10676 6404
rect 9772 6280 9812 6320
rect 15436 6448 15476 6488
rect 16492 6448 16532 6488
rect 16972 6448 17012 6488
rect 17548 6448 17588 6488
rect 15532 6364 15572 6404
rect 3340 6196 3380 6236
rect 5836 6196 5876 6236
rect 6412 6196 6452 6236
rect 6604 6196 6644 6236
rect 7276 6196 7316 6236
rect 9388 6196 9428 6236
rect 9964 6196 10004 6236
rect 11884 6196 11924 6236
rect 12652 6196 12692 6236
rect 14092 6196 14132 6236
rect 16300 6196 16340 6236
rect 7948 6112 7988 6152
rect 10060 6112 10100 6152
rect 3112 6028 3480 6068
rect 6700 6028 6740 6068
rect 9292 6028 9332 6068
rect 10886 6028 11254 6068
rect 15820 6112 15860 6152
rect 17068 6112 17108 6152
rect 24460 6952 24500 6992
rect 25228 6952 25268 6992
rect 27532 6952 27572 6992
rect 27674 6784 28042 6824
rect 21196 6616 21236 6656
rect 21772 6616 21803 6656
rect 21803 6616 21812 6656
rect 22252 6616 22283 6656
rect 22283 6616 22292 6656
rect 23308 6616 23348 6656
rect 23980 6616 24020 6656
rect 20716 6532 20756 6572
rect 21868 6532 21908 6572
rect 22156 6532 22196 6572
rect 23404 6532 23444 6572
rect 20236 6448 20276 6488
rect 20620 6448 20660 6488
rect 20908 6448 20948 6488
rect 22348 6448 22388 6488
rect 23596 6448 23636 6488
rect 24076 6479 24116 6488
rect 24076 6448 24116 6479
rect 24460 6448 24491 6488
rect 24491 6448 24500 6488
rect 19276 6364 19316 6404
rect 21292 6280 21332 6320
rect 460 5944 500 5984
rect 5740 5860 5780 5900
rect 6508 5776 6548 5816
rect 9004 5776 9044 5816
rect 10444 5860 10484 5900
rect 14476 5860 14516 5900
rect 15052 5860 15083 5900
rect 15083 5860 15092 5900
rect 23788 6364 23828 6404
rect 22924 6196 22964 6236
rect 18660 6028 19028 6068
rect 19564 6028 19604 6068
rect 22252 6028 22292 6068
rect 26434 6028 26802 6068
rect 21388 5944 21428 5984
rect 20620 5860 20651 5900
rect 20651 5860 20660 5900
rect 20908 5860 20948 5900
rect 22060 5860 22100 5900
rect 22348 5860 22388 5900
rect 23596 5860 23636 5900
rect 12940 5776 12980 5816
rect 20236 5776 20276 5816
rect 2284 5608 2324 5648
rect 8044 5692 8084 5732
rect 2668 5608 2708 5648
rect 2956 5608 2987 5648
rect 2987 5608 2996 5648
rect 3916 5608 3947 5648
rect 3947 5608 3956 5648
rect 4204 5608 4244 5648
rect 4780 5608 4820 5648
rect 6220 5608 6260 5648
rect 6604 5608 6644 5648
rect 6988 5608 7028 5648
rect 9388 5608 9419 5648
rect 9419 5608 9428 5648
rect 9772 5608 9812 5648
rect 11500 5608 11540 5648
rect 11884 5608 11924 5648
rect 12268 5608 12308 5648
rect 12556 5608 12596 5648
rect 12844 5608 12884 5648
rect 15244 5692 15284 5732
rect 16300 5692 16340 5732
rect 18892 5692 18932 5732
rect 19564 5692 19604 5732
rect 20812 5692 20852 5732
rect 21292 5692 21332 5732
rect 3532 5524 3572 5564
rect 6124 5524 6164 5564
rect 7564 5524 7604 5564
rect 2572 5440 2612 5480
rect 4204 5440 4244 5480
rect 5548 5440 5588 5480
rect 6988 5356 7028 5396
rect 4352 5272 4720 5312
rect 6124 5272 6164 5312
rect 7180 5272 7220 5312
rect 9484 5524 9524 5564
rect 10444 5524 10484 5564
rect 11980 5524 12020 5564
rect 8524 5440 8555 5480
rect 8555 5440 8564 5480
rect 11308 5440 11348 5480
rect 6412 5104 6452 5144
rect 5452 5020 5492 5060
rect 5644 4936 5684 4976
rect 6220 4852 6260 4892
rect 11788 5440 11828 5480
rect 12172 5440 12212 5480
rect 12940 5471 12980 5480
rect 12940 5440 12971 5471
rect 12971 5440 12980 5471
rect 12126 5272 12494 5312
rect 13804 5608 13844 5648
rect 15436 5608 15476 5648
rect 16492 5608 16532 5648
rect 16684 5608 16724 5648
rect 17068 5608 17108 5648
rect 18412 5608 18452 5648
rect 18700 5608 18740 5648
rect 19084 5608 19124 5648
rect 21004 5608 21044 5648
rect 21676 5608 21707 5648
rect 21707 5608 21716 5648
rect 15532 5524 15572 5564
rect 15820 5524 15860 5564
rect 20908 5524 20948 5564
rect 14380 5440 14420 5480
rect 16204 5440 16244 5480
rect 18124 5440 18164 5480
rect 16012 5272 16052 5312
rect 18892 5188 18932 5228
rect 11980 5104 12020 5144
rect 15532 5104 15572 5144
rect 18700 5104 18731 5144
rect 18731 5104 18740 5144
rect 12652 5020 12692 5060
rect 15340 5020 15380 5060
rect 16684 5020 16724 5060
rect 19900 5272 20268 5312
rect 23404 5272 23444 5312
rect 27674 5272 28042 5312
rect 21964 5188 22004 5228
rect 21868 5104 21908 5144
rect 21004 5020 21044 5060
rect 22924 5020 22964 5060
rect 11692 4936 11732 4976
rect 12556 4936 12596 4976
rect 18412 4936 18452 4976
rect 8044 4852 8084 4892
rect 9004 4852 9044 4892
rect 10060 4768 10100 4808
rect 9580 4684 9620 4724
rect 10348 4684 10388 4724
rect 11884 4852 11924 4892
rect 14380 4852 14420 4892
rect 15148 4852 15188 4892
rect 16108 4852 16148 4892
rect 17164 4852 17204 4892
rect 17932 4852 17972 4892
rect 20908 4936 20948 4976
rect 21388 4936 21428 4976
rect 21772 4936 21812 4976
rect 22348 4936 22388 4976
rect 24460 4852 24500 4892
rect 13228 4768 13268 4808
rect 21772 4768 21812 4808
rect 19276 4684 19316 4724
rect 8716 4600 8756 4640
rect 13804 4600 13844 4640
rect 17068 4600 17108 4640
rect 20812 4600 20852 4640
rect 3112 4516 3480 4556
rect 10886 4516 11254 4556
rect 18660 4516 19028 4556
rect 26434 4516 26802 4556
rect 7948 4432 7988 4472
rect 15244 4432 15284 4472
rect 8044 4348 8084 4388
rect 13228 4348 13268 4388
rect 15148 4348 15188 4388
rect 16108 4348 16148 4388
rect 6220 4264 6260 4304
rect 7180 4264 7220 4304
rect 11500 4264 11540 4304
rect 13708 4264 13748 4304
rect 13900 4264 13940 4304
rect 14380 4264 14420 4304
rect 17164 4264 17204 4304
rect 8524 4180 8564 4220
rect 11980 4180 12020 4220
rect 13804 4180 13844 4220
rect 14284 4180 14324 4220
rect 7564 4096 7595 4136
rect 7595 4096 7604 4136
rect 7948 4096 7988 4136
rect 8716 4096 8756 4136
rect 10060 4096 10100 4136
rect 10348 4096 10387 4136
rect 10387 4096 10388 4136
rect 11692 4096 11732 4136
rect 11884 4096 11924 4136
rect 13900 4096 13940 4136
rect 15532 4096 15572 4136
rect 15820 4096 15851 4136
rect 15851 4096 15860 4136
rect 16204 4096 16244 4136
rect 16684 4012 16724 4052
rect 4352 3760 4720 3800
rect 12126 3760 12494 3800
rect 19900 3760 20268 3800
rect 27674 3760 28042 3800
rect 3112 3004 3480 3044
rect 10886 3004 11254 3044
rect 18660 3004 19028 3044
rect 26434 3004 26802 3044
rect 4352 2248 4720 2288
rect 12126 2248 12494 2288
rect 19900 2248 20268 2288
rect 27674 2248 28042 2288
rect 3112 1492 3480 1532
rect 10886 1492 11254 1532
rect 18660 1492 19028 1532
rect 26434 1492 26802 1532
rect 4352 736 4720 776
rect 12126 736 12494 776
rect 19900 736 20268 776
rect 27674 736 28042 776
<< metal3 >>
rect 3128 28600 3208 29000
rect 3896 28600 3976 29000
rect 4664 28600 4744 29000
rect 5432 28600 5512 29000
rect 6200 28600 6280 29000
rect 6968 28600 7048 29000
rect 7736 28600 7816 29000
rect 8504 28600 8584 29000
rect 9272 28600 9352 29000
rect 10040 28600 10120 29000
rect 10808 28600 10888 29000
rect 11576 28600 11656 29000
rect 12344 28600 12424 29000
rect 13112 28600 13192 29000
rect 13880 28600 13960 29000
rect 14648 28600 14728 29000
rect 15416 28600 15496 29000
rect 16184 28600 16264 29000
rect 16396 28664 16436 28673
rect 2956 28496 2996 28505
rect 1804 28412 1844 28421
rect 1516 28160 1556 28169
rect 1516 26648 1556 28120
rect 1804 27656 1844 28372
rect 2764 28160 2804 28169
rect 1900 28076 1940 28085
rect 1900 27740 1940 28036
rect 1900 27691 1940 27700
rect 2188 27992 2228 28001
rect 1804 27607 1844 27616
rect 1516 26599 1556 26608
rect 1900 27572 1940 27581
rect 1900 26648 1940 27532
rect 2188 27572 2228 27952
rect 2188 27523 2228 27532
rect 2476 27740 2516 27749
rect 1900 26599 1940 26608
rect 2092 27488 2132 27497
rect 2092 27068 2132 27448
rect 2380 27488 2420 27497
rect 2380 27353 2420 27448
rect 2092 26480 2132 27028
rect 2092 26431 2132 26440
rect 2476 26228 2516 27700
rect 2668 27656 2708 27665
rect 2668 26816 2708 27616
rect 2764 27488 2804 28120
rect 2956 27992 2996 28456
rect 2956 27572 2996 27952
rect 3148 27824 3188 28600
rect 3148 27775 3188 27784
rect 3532 28160 3572 28169
rect 2956 27523 2996 27532
rect 3148 27656 3188 27665
rect 2764 27439 2804 27448
rect 3148 27404 3188 27616
rect 3532 27488 3572 28120
rect 3532 27439 3572 27448
rect 3628 27824 3668 27833
rect 2956 27364 3188 27404
rect 2860 26984 2900 26993
rect 2956 26984 2996 27364
rect 3112 27236 3480 27245
rect 3112 27187 3480 27196
rect 2900 26944 3092 26984
rect 2860 26935 2900 26944
rect 2668 26767 2708 26776
rect 2860 26816 2900 26825
rect 2900 26776 2996 26816
rect 2860 26767 2900 26776
rect 2956 26396 2996 26776
rect 2956 26347 2996 26356
rect 2476 26179 2516 26188
rect 2956 26228 2996 26237
rect 2860 26144 2900 26153
rect 2188 26060 2228 26069
rect 1132 25976 1172 25985
rect 844 25388 884 25397
rect 556 25220 596 25229
rect 364 24380 404 24389
rect 172 23288 212 23297
rect 76 22532 116 22541
rect 76 15812 116 22492
rect 76 15763 116 15772
rect 172 7412 212 23248
rect 268 22196 308 22205
rect 268 7975 308 22156
rect 364 20768 404 24340
rect 460 22532 500 22541
rect 460 22397 500 22492
rect 556 22364 596 25180
rect 556 22315 596 22324
rect 652 25136 692 25145
rect 460 22028 500 22037
rect 460 21692 500 21988
rect 460 21643 500 21652
rect 556 22028 596 22037
rect 460 21524 500 21533
rect 460 21020 500 21484
rect 460 20971 500 20980
rect 364 20728 500 20768
rect 460 20684 500 20728
rect 460 20635 500 20644
rect 364 20600 404 20609
rect 364 18164 404 20560
rect 460 20348 500 20357
rect 460 19844 500 20308
rect 460 19795 500 19804
rect 364 18124 500 18164
rect 364 14804 404 14813
rect 364 8504 404 14764
rect 460 13796 500 18124
rect 556 14804 596 21988
rect 652 20516 692 25096
rect 652 20467 692 20476
rect 748 23372 788 23381
rect 748 20348 788 23332
rect 844 22784 884 25348
rect 1036 24548 1076 24557
rect 940 23204 980 23213
rect 940 23069 980 23164
rect 1036 22952 1076 24508
rect 1036 22903 1076 22912
rect 844 22735 884 22744
rect 1036 22700 1076 22709
rect 652 20308 788 20348
rect 844 22616 884 22625
rect 652 19424 692 20308
rect 844 20012 884 22576
rect 1036 22028 1076 22660
rect 1036 21979 1076 21988
rect 652 19375 692 19384
rect 748 19972 884 20012
rect 940 20516 980 20525
rect 556 14755 596 14764
rect 652 19088 692 19097
rect 652 14804 692 19048
rect 652 14755 692 14764
rect 748 14636 788 19972
rect 460 13747 500 13756
rect 556 14596 788 14636
rect 844 19844 884 19853
rect 556 8924 596 14596
rect 748 14468 788 14477
rect 652 14216 692 14225
rect 652 13544 692 14176
rect 652 13495 692 13504
rect 556 8875 596 8884
rect 652 11276 692 11285
rect 652 10100 692 11236
rect 652 9512 692 10060
rect 460 8504 500 8513
rect 364 8464 460 8504
rect 460 8455 500 8464
rect 652 8168 692 9472
rect 652 8119 692 8128
rect 268 7926 308 7935
rect 172 7363 212 7372
rect 748 6824 788 14428
rect 844 8084 884 19804
rect 940 19340 980 20476
rect 940 19291 980 19300
rect 1036 20516 1076 20525
rect 940 18752 980 18761
rect 940 13124 980 18712
rect 1036 13964 1076 20476
rect 1132 14300 1172 25936
rect 1516 25976 1556 25985
rect 1228 25388 1268 25397
rect 1228 24128 1268 25348
rect 1228 24079 1268 24088
rect 1324 25220 1364 25229
rect 1228 22364 1268 22373
rect 1228 21020 1268 22324
rect 1324 22112 1364 25180
rect 1516 23876 1556 25936
rect 1900 25976 1940 25985
rect 1900 25841 1940 25936
rect 1612 25472 1652 25481
rect 1612 25337 1652 25432
rect 1516 23827 1556 23836
rect 1612 25220 1652 25229
rect 1612 23708 1652 25180
rect 1996 25136 2036 25145
rect 1708 24800 1748 24809
rect 1708 24665 1748 24760
rect 1996 24632 2036 25096
rect 1996 24583 2036 24592
rect 1612 23659 1652 23668
rect 1996 23708 2036 23717
rect 1420 23372 1460 23381
rect 1420 23288 1460 23332
rect 1420 23237 1460 23248
rect 1612 23120 1652 23129
rect 1612 23060 1652 23080
rect 1516 23020 1652 23060
rect 1900 23036 1940 23045
rect 1324 22063 1364 22072
rect 1420 22196 1460 22205
rect 1324 21524 1364 21533
rect 1324 21272 1364 21484
rect 1420 21440 1460 22156
rect 1516 21575 1556 23020
rect 1708 22868 1748 22877
rect 1708 22280 1748 22828
rect 1708 22231 1748 22240
rect 1804 22196 1844 22205
rect 1516 21526 1556 21535
rect 1612 22028 1652 22037
rect 1612 21776 1652 21988
rect 1420 21391 1460 21400
rect 1612 21440 1652 21736
rect 1324 21232 1460 21272
rect 1228 20971 1268 20980
rect 1324 21104 1364 21113
rect 1228 20600 1268 20609
rect 1228 18752 1268 20560
rect 1228 18703 1268 18712
rect 1324 18584 1364 21064
rect 1420 21020 1460 21232
rect 1420 20971 1460 20980
rect 1420 20852 1460 20861
rect 1420 20717 1460 20812
rect 1612 20600 1652 21400
rect 1612 20551 1652 20560
rect 1708 21860 1748 21869
rect 1132 14251 1172 14260
rect 1228 18544 1364 18584
rect 1420 19844 1460 19853
rect 1036 13915 1076 13924
rect 940 13075 980 13084
rect 1036 13796 1076 13805
rect 1036 12704 1076 13756
rect 1228 12980 1268 18544
rect 1324 14720 1364 14729
rect 1324 14132 1364 14680
rect 1420 14468 1460 19804
rect 1708 18584 1748 21820
rect 1804 21608 1844 22156
rect 1804 20348 1844 21568
rect 1900 21608 1940 22996
rect 1996 21860 2036 23668
rect 2188 23204 2228 26020
rect 2476 26060 2516 26069
rect 2380 25304 2420 25313
rect 2284 25052 2324 25061
rect 2284 24632 2324 25012
rect 2284 23792 2324 24592
rect 2380 24548 2420 25264
rect 2380 24499 2420 24508
rect 2284 23743 2324 23752
rect 2380 24044 2420 24053
rect 2380 23288 2420 24004
rect 2188 23164 2324 23204
rect 2092 23120 2132 23129
rect 2092 22448 2132 23080
rect 2284 23120 2324 23164
rect 2284 23071 2324 23080
rect 2092 22280 2132 22408
rect 2188 23036 2228 23045
rect 2188 22364 2228 22996
rect 2188 22315 2228 22324
rect 2092 22231 2132 22240
rect 2284 22280 2324 22289
rect 2284 22112 2324 22240
rect 2284 22063 2324 22072
rect 1996 21776 2036 21820
rect 1996 21725 2036 21736
rect 2188 21692 2228 21701
rect 2188 21608 2228 21652
rect 1900 20852 1940 21568
rect 1900 20803 1940 20812
rect 1996 21568 2228 21608
rect 1996 20600 2036 21568
rect 2380 21272 2420 23248
rect 1996 20551 2036 20560
rect 2092 21232 2420 21272
rect 2476 23792 2516 26020
rect 2860 26009 2900 26104
rect 2860 25808 2900 25817
rect 2860 25673 2900 25768
rect 2572 25388 2612 25397
rect 2572 25253 2612 25348
rect 2956 25304 2996 26188
rect 3052 25892 3092 26944
rect 3244 26900 3284 26995
rect 3244 26851 3284 26860
rect 3532 26900 3572 26909
rect 3340 26648 3380 26657
rect 3340 26144 3380 26608
rect 3340 26095 3380 26104
rect 3532 25976 3572 26860
rect 3532 25927 3572 25936
rect 3052 25843 3092 25852
rect 3112 25724 3480 25733
rect 3112 25675 3480 25684
rect 3244 25472 3284 25483
rect 3244 25388 3284 25432
rect 3244 25339 3284 25348
rect 2956 25255 2996 25264
rect 3148 25136 3188 25145
rect 2764 25096 3148 25136
rect 2764 24632 2804 25096
rect 3148 25087 3188 25096
rect 2764 24583 2804 24592
rect 3112 24212 3480 24221
rect 3112 24163 3480 24172
rect 2092 20432 2132 21232
rect 2188 20768 2228 20863
rect 2188 20719 2228 20728
rect 2380 20684 2420 20693
rect 2081 20392 2132 20432
rect 2188 20600 2228 20609
rect 2081 20348 2121 20392
rect 2081 20308 2132 20348
rect 1804 20180 1844 20308
rect 1804 20140 1940 20180
rect 1900 20096 1940 20140
rect 1900 20047 1940 20056
rect 1708 18535 1748 18544
rect 1996 18500 2036 18509
rect 1804 17912 1844 17921
rect 1708 16568 1748 16577
rect 1708 15560 1748 16528
rect 1804 16148 1844 17872
rect 1996 17912 2036 18460
rect 2092 18080 2132 20308
rect 2188 20096 2228 20560
rect 2284 20096 2324 20105
rect 2188 20056 2284 20096
rect 2188 19340 2228 20056
rect 2284 20047 2324 20056
rect 2188 19291 2228 19300
rect 2380 19256 2420 20644
rect 2380 19207 2420 19216
rect 2476 19088 2516 23752
rect 3244 23876 3284 23885
rect 2668 23204 2708 23213
rect 2572 22784 2612 22793
rect 2572 21356 2612 22744
rect 2668 22448 2708 23164
rect 3244 23204 3284 23836
rect 3244 23155 3284 23164
rect 2764 22952 2804 22961
rect 2764 22700 2804 22912
rect 2956 22952 2996 22963
rect 2956 22868 2996 22912
rect 2956 22819 2996 22828
rect 3436 22952 3476 22961
rect 3436 22817 3476 22912
rect 2764 22651 2804 22660
rect 3112 22700 3480 22709
rect 3112 22651 3480 22660
rect 2708 22408 2804 22448
rect 2668 22399 2708 22408
rect 2668 22196 2708 22205
rect 2668 22061 2708 22156
rect 2572 21307 2612 21316
rect 2668 21440 2708 21449
rect 2572 20768 2612 20777
rect 2572 20264 2612 20728
rect 2572 20215 2612 20224
rect 2572 19844 2612 19939
rect 2572 19795 2612 19804
rect 2380 19048 2516 19088
rect 2572 19676 2612 19685
rect 2572 19088 2612 19636
rect 2284 18332 2324 18341
rect 2188 18080 2228 18089
rect 2092 18040 2188 18080
rect 1996 17863 2036 17872
rect 2092 17576 2132 17585
rect 1804 16099 1844 16108
rect 1996 17240 2036 17249
rect 1996 16232 2036 17200
rect 1996 15728 2036 16192
rect 1996 15679 2036 15688
rect 1612 15476 1652 15485
rect 1612 14972 1652 15436
rect 1612 14923 1652 14932
rect 1708 14804 1748 15520
rect 1612 14764 1748 14804
rect 1420 14419 1460 14428
rect 1516 14720 1556 14729
rect 1516 14216 1556 14680
rect 1324 14083 1364 14092
rect 1420 14176 1516 14216
rect 1036 12655 1076 12664
rect 1132 12940 1268 12980
rect 1324 13040 1364 13049
rect 1036 11528 1076 11537
rect 940 10940 980 10949
rect 940 10436 980 10900
rect 940 10387 980 10396
rect 844 8035 884 8044
rect 940 10268 980 10277
rect 940 8840 980 10228
rect 1036 10100 1076 11488
rect 1036 10051 1076 10060
rect 940 8000 980 8800
rect 940 7951 980 7960
rect 748 6775 788 6784
rect 1132 6404 1172 12940
rect 1324 12536 1364 13000
rect 1324 11612 1364 12496
rect 1228 11528 1268 11537
rect 1228 11024 1268 11488
rect 1228 10975 1268 10984
rect 1324 11024 1364 11572
rect 1324 10975 1364 10984
rect 1420 11864 1460 14176
rect 1516 14167 1556 14176
rect 1612 13208 1652 14764
rect 2092 14720 2132 17536
rect 2188 16316 2228 18040
rect 2284 17324 2324 18292
rect 2380 17828 2420 19048
rect 2572 19039 2612 19048
rect 2380 17779 2420 17788
rect 2668 17828 2708 21400
rect 2764 20600 2804 22408
rect 3532 22364 3572 22373
rect 3436 22280 3476 22289
rect 3340 22196 3380 22205
rect 3148 22112 3188 22121
rect 3148 21860 3188 22072
rect 3148 21811 3188 21820
rect 3340 21860 3380 22156
rect 3052 21608 3092 21619
rect 3052 21524 3092 21568
rect 3052 21475 3092 21484
rect 3244 21524 3284 21533
rect 3244 21440 3284 21484
rect 3244 21389 3284 21400
rect 3340 21356 3380 21820
rect 3436 21692 3476 22240
rect 3532 21776 3572 22324
rect 3532 21727 3572 21736
rect 3436 21643 3476 21652
rect 3532 21608 3572 21619
rect 3532 21524 3572 21568
rect 3532 21475 3572 21484
rect 3340 21316 3572 21356
rect 2956 21188 2996 21197
rect 2764 20096 2804 20560
rect 2860 20684 2900 20693
rect 2860 20549 2900 20644
rect 2956 20180 2996 21148
rect 3112 21188 3480 21197
rect 3112 21139 3480 21148
rect 3340 21020 3380 21029
rect 3532 21020 3572 21316
rect 3244 20936 3284 20945
rect 2764 19676 2804 20056
rect 2764 19627 2804 19636
rect 2860 20140 2996 20180
rect 3052 20600 3092 20609
rect 3052 20348 3092 20560
rect 2860 19592 2900 20140
rect 3052 20096 3092 20308
rect 3244 20264 3284 20896
rect 3340 20600 3380 20980
rect 3340 20551 3380 20560
rect 3436 20980 3572 21020
rect 3244 20215 3284 20224
rect 3436 20180 3476 20980
rect 3052 20047 3092 20056
rect 3340 20140 3476 20180
rect 3532 20768 3572 20777
rect 3340 20096 3380 20140
rect 3340 20047 3380 20056
rect 2860 19543 2900 19552
rect 2956 19760 2996 19769
rect 2956 19424 2996 19720
rect 3112 19676 3480 19685
rect 3112 19627 3480 19636
rect 2764 19384 2996 19424
rect 3052 19508 3092 19517
rect 2764 19256 2804 19384
rect 3052 19256 3092 19468
rect 3532 19424 3572 20728
rect 2764 19207 2804 19216
rect 2956 19216 3052 19256
rect 2668 17779 2708 17788
rect 2956 17828 2996 19216
rect 3052 19207 3092 19216
rect 3436 19384 3572 19424
rect 3628 19424 3668 27784
rect 3916 27320 3956 28600
rect 4684 28160 4724 28600
rect 4684 28111 4724 28120
rect 4352 27992 4720 28001
rect 4352 27943 4720 27952
rect 5452 27908 5492 28600
rect 5452 27859 5492 27868
rect 5932 28076 5972 28085
rect 3916 27271 3956 27280
rect 4396 27656 4436 27665
rect 4396 26900 4436 27616
rect 4396 26851 4436 26860
rect 5740 27656 5780 27665
rect 4588 26816 4628 26825
rect 4588 26732 4628 26776
rect 5068 26816 5108 26825
rect 4588 26681 4628 26692
rect 4684 26648 4724 26743
rect 4684 26599 4724 26608
rect 4352 26480 4720 26489
rect 4352 26431 4720 26440
rect 5068 26312 5108 26776
rect 5548 26816 5588 26825
rect 5260 26732 5300 26741
rect 5164 26396 5204 26491
rect 5164 26347 5204 26356
rect 5068 26263 5108 26272
rect 4012 26144 4052 26153
rect 3724 25808 3764 25817
rect 3724 25724 3764 25768
rect 3724 25673 3764 25684
rect 3820 23792 3860 23801
rect 3820 23288 3860 23752
rect 4012 23540 4052 26104
rect 4780 26144 4820 26153
rect 4204 25388 4244 25397
rect 4012 23491 4052 23500
rect 4108 24632 4148 24641
rect 3820 23239 3860 23248
rect 4108 23120 4148 24592
rect 4108 23071 4148 23080
rect 4204 23036 4244 25348
rect 4352 24968 4720 24977
rect 4352 24919 4720 24928
rect 4588 24716 4628 24725
rect 4588 24044 4628 24676
rect 4588 23995 4628 24004
rect 4352 23456 4720 23465
rect 4352 23407 4720 23416
rect 4492 23288 4532 23297
rect 4396 23204 4436 23213
rect 4396 23120 4436 23164
rect 4396 23069 4436 23080
rect 3820 22952 3860 22961
rect 3724 22280 3764 22289
rect 3724 22145 3764 22240
rect 3148 19088 3188 19097
rect 3148 18584 3188 19048
rect 3436 18920 3476 19384
rect 3628 19375 3668 19384
rect 3724 21272 3764 21281
rect 3724 19340 3764 21232
rect 3724 19291 3764 19300
rect 3820 20096 3860 22912
rect 3916 22448 3956 22457
rect 4204 22448 4244 22996
rect 4396 22784 4436 22793
rect 3916 22364 3956 22408
rect 3916 22313 3956 22324
rect 4012 22408 4244 22448
rect 4300 22532 4340 22541
rect 4300 22448 4340 22492
rect 3916 21608 3956 21617
rect 3916 21473 3956 21568
rect 4012 21272 4052 22408
rect 4300 22397 4340 22408
rect 4396 22364 4436 22744
rect 4492 22448 4532 23248
rect 4492 22399 4532 22408
rect 4780 22448 4820 26104
rect 5164 26144 5204 26153
rect 5164 25304 5204 26104
rect 5260 25976 5300 26692
rect 5452 26648 5492 26657
rect 5356 26396 5396 26405
rect 5356 26060 5396 26356
rect 5356 26011 5396 26020
rect 5260 25927 5300 25936
rect 5452 25892 5492 26608
rect 5548 26228 5588 26776
rect 5548 26179 5588 26188
rect 5644 26732 5684 26741
rect 5452 25472 5492 25852
rect 5452 25423 5492 25432
rect 5164 25255 5204 25264
rect 5260 25388 5300 25397
rect 4972 24380 5012 24389
rect 4972 23792 5012 24340
rect 4972 23743 5012 23752
rect 5260 23792 5300 25348
rect 5644 25388 5684 26692
rect 5644 25339 5684 25348
rect 5740 26060 5780 27616
rect 5932 26816 5972 28036
rect 5932 26767 5972 26776
rect 5356 25304 5396 25313
rect 5356 25136 5396 25264
rect 5740 25304 5780 26020
rect 5740 25255 5780 25264
rect 5932 25892 5972 25901
rect 5932 25304 5972 25852
rect 5932 25255 5972 25264
rect 5356 25087 5396 25096
rect 5452 25220 5492 25229
rect 5260 23657 5300 23752
rect 5068 23204 5108 23213
rect 5068 23069 5108 23164
rect 5164 23120 5204 23129
rect 5452 23120 5492 25180
rect 6220 24800 6260 28600
rect 6796 28244 6836 28253
rect 6700 27740 6740 27749
rect 6508 27572 6548 27581
rect 6508 26984 6548 27532
rect 6700 27068 6740 27700
rect 6700 27019 6740 27028
rect 6508 26935 6548 26944
rect 6508 26816 6548 26825
rect 6508 26228 6548 26776
rect 6508 26179 6548 26188
rect 6796 26060 6836 28204
rect 6988 27824 7028 28600
rect 6988 27775 7028 27784
rect 7084 28412 7124 28421
rect 6892 27488 6932 27497
rect 6892 26837 6932 27448
rect 6892 26788 6932 26797
rect 7084 26732 7124 28372
rect 7372 27656 7412 27665
rect 6892 26648 6932 26657
rect 6892 26144 6932 26608
rect 6932 26104 7028 26144
rect 6892 26095 6932 26104
rect 6796 26011 6836 26020
rect 6892 25808 6932 25817
rect 6508 25304 6548 25313
rect 6508 25169 6548 25264
rect 6892 25304 6932 25768
rect 6988 25388 7028 26104
rect 7084 25976 7124 26692
rect 7180 26816 7220 26827
rect 7180 26732 7220 26776
rect 7180 26683 7220 26692
rect 7372 26648 7412 27616
rect 7372 26599 7412 26608
rect 7468 27572 7508 27581
rect 7084 25936 7220 25976
rect 6988 25339 7028 25348
rect 7180 25388 7220 25936
rect 7468 25640 7508 27532
rect 7564 26648 7604 26657
rect 7564 25724 7604 26608
rect 7756 26480 7796 28600
rect 8236 28160 8276 28169
rect 7756 26431 7796 26440
rect 7948 26900 7988 26909
rect 7948 26480 7988 26860
rect 7948 26431 7988 26440
rect 8140 26732 8180 26741
rect 7564 25675 7604 25684
rect 8140 26312 8180 26692
rect 7468 25591 7508 25600
rect 8140 25556 8180 26272
rect 8236 26060 8276 28120
rect 8524 27572 8564 28600
rect 8524 27523 8564 27532
rect 9100 28580 9140 28589
rect 8620 27404 8660 27413
rect 8524 27320 8564 27329
rect 8524 26984 8564 27280
rect 8524 26935 8564 26944
rect 8620 26816 8660 27364
rect 8620 26767 8660 26776
rect 8332 26732 8372 26741
rect 8332 26144 8372 26692
rect 8332 26095 8372 26104
rect 8428 26564 8468 26573
rect 8236 26011 8276 26020
rect 8140 25507 8180 25516
rect 8332 25892 8372 25901
rect 6892 25255 6932 25264
rect 6220 24751 6260 24760
rect 5740 24632 5780 24641
rect 5548 24128 5588 24137
rect 5548 23288 5588 24088
rect 5740 24128 5780 24592
rect 5740 23792 5780 24088
rect 5740 23743 5780 23752
rect 6028 24212 6068 24221
rect 6028 23792 6068 24172
rect 7180 23876 7220 25348
rect 8332 25304 8372 25852
rect 7468 24716 7508 24725
rect 7372 23876 7412 23885
rect 7180 23836 7316 23876
rect 6068 23752 6260 23792
rect 6028 23743 6068 23752
rect 5932 23708 5972 23717
rect 5548 23239 5588 23248
rect 5740 23372 5780 23381
rect 5164 22532 5204 23080
rect 5356 23080 5452 23120
rect 5260 23036 5300 23045
rect 5260 22784 5300 22996
rect 5260 22735 5300 22744
rect 5164 22483 5204 22492
rect 4780 22399 4820 22408
rect 4396 22315 4436 22324
rect 5068 22364 5108 22373
rect 4972 22280 5012 22289
rect 4204 22196 4244 22205
rect 4012 21223 4052 21232
rect 4108 21524 4148 21533
rect 4012 20852 4052 20861
rect 4012 20768 4052 20812
rect 4012 20717 4052 20728
rect 3436 18871 3476 18880
rect 3532 19256 3572 19265
rect 3148 18535 3188 18544
rect 3112 18164 3480 18173
rect 3112 18115 3480 18124
rect 2956 17779 2996 17788
rect 3148 17996 3188 18005
rect 2572 17744 2612 17753
rect 2572 17609 2612 17704
rect 3148 17744 3188 17956
rect 2284 17275 2324 17284
rect 2188 16267 2228 16276
rect 2572 16820 2612 16829
rect 3148 16820 3188 17704
rect 3244 17072 3284 17081
rect 3244 16937 3284 17032
rect 2572 15560 2612 16780
rect 2956 16780 3188 16820
rect 2860 16232 2900 16241
rect 2860 15644 2900 16192
rect 2860 15595 2900 15604
rect 2572 15511 2612 15520
rect 2956 15560 2996 16780
rect 3112 16652 3480 16661
rect 3112 16603 3480 16612
rect 2956 15511 2996 15520
rect 3340 16148 3380 16157
rect 3340 15560 3380 16108
rect 3532 15728 3572 19216
rect 3820 19256 3860 20056
rect 3628 19172 3668 19181
rect 3628 18752 3668 19132
rect 3820 19121 3860 19216
rect 3916 20600 3956 20609
rect 3628 17576 3668 18712
rect 3724 18500 3764 18509
rect 3724 17996 3764 18460
rect 3724 17947 3764 17956
rect 3820 17912 3860 17921
rect 3820 17744 3860 17872
rect 3628 17527 3668 17536
rect 3724 17660 3764 17669
rect 3628 17156 3668 17165
rect 3628 17072 3668 17116
rect 3628 17021 3668 17032
rect 3628 16652 3668 16661
rect 3724 16652 3764 17620
rect 3668 16612 3764 16652
rect 3628 16232 3668 16612
rect 3628 16183 3668 16192
rect 3532 15679 3572 15688
rect 3724 15728 3764 15737
rect 3340 15511 3380 15520
rect 3628 15560 3668 15569
rect 2956 15308 2996 15317
rect 2092 14671 2132 14680
rect 2764 14804 2804 14813
rect 1708 14636 1748 14645
rect 1708 14048 1748 14596
rect 1708 13999 1748 14008
rect 2092 14552 2132 14561
rect 1612 13159 1652 13168
rect 2092 13208 2132 14512
rect 2092 13159 2132 13168
rect 2572 13208 2612 13217
rect 2188 13124 2228 13133
rect 1708 12536 1748 12545
rect 1420 10184 1460 11824
rect 1420 10100 1460 10144
rect 1324 10060 1460 10100
rect 1516 12452 1556 12461
rect 1516 11612 1556 12412
rect 1324 9428 1364 10060
rect 1516 9764 1556 11572
rect 1708 11612 1748 12496
rect 2092 12452 2132 12461
rect 2092 11948 2132 12412
rect 2092 11899 2132 11908
rect 1708 11563 1748 11572
rect 2188 11696 2228 13084
rect 2572 13040 2612 13168
rect 2572 12991 2612 13000
rect 2764 13208 2804 14764
rect 2956 14804 2996 15268
rect 3112 15140 3480 15149
rect 3112 15091 3480 15100
rect 2956 14755 2996 14764
rect 3148 14804 3188 14813
rect 2956 14636 2996 14645
rect 2956 14216 2996 14596
rect 2956 14167 2996 14176
rect 3148 14048 3188 14764
rect 3148 13999 3188 14008
rect 3436 14720 3476 14729
rect 3436 14048 3476 14680
rect 3628 14720 3668 15520
rect 3724 15224 3764 15688
rect 3724 15175 3764 15184
rect 3628 14671 3668 14680
rect 3436 13999 3476 14008
rect 3112 13628 3480 13637
rect 3112 13579 3480 13588
rect 2572 12788 2612 12797
rect 1708 11360 1748 11369
rect 1708 10268 1748 11320
rect 2188 11276 2228 11656
rect 2188 11227 2228 11236
rect 2284 12536 2324 12545
rect 2284 11192 2324 12496
rect 2284 11143 2324 11152
rect 2572 10940 2612 12748
rect 2668 11696 2708 11705
rect 2668 11561 2708 11656
rect 2764 11612 2804 13168
rect 3436 13208 3476 13217
rect 3436 13040 3476 13168
rect 3436 12991 3476 13000
rect 3112 12116 3480 12125
rect 3112 12067 3480 12076
rect 2764 11563 2804 11572
rect 3532 11696 3572 11705
rect 3532 11528 3572 11656
rect 3532 11479 3572 11488
rect 2956 11444 2996 11453
rect 2956 11108 2996 11404
rect 2956 11059 2996 11068
rect 1708 10219 1748 10228
rect 2476 10268 2516 10277
rect 1516 9512 1556 9724
rect 1804 10184 1844 10193
rect 1804 9680 1844 10144
rect 1804 9631 1844 9640
rect 2092 10184 2132 10193
rect 2092 10016 2132 10144
rect 2476 10100 2516 10228
rect 2476 10051 2516 10060
rect 1516 9463 1556 9472
rect 1324 9379 1364 9388
rect 2092 9344 2132 9976
rect 2092 9295 2132 9304
rect 2476 9764 2516 9773
rect 2476 9428 2516 9724
rect 1996 8756 2036 8765
rect 1996 7832 2036 8716
rect 1996 7783 2036 7792
rect 2476 7244 2516 9388
rect 2572 9512 2612 10900
rect 2668 11024 2708 11033
rect 2668 10889 2708 10984
rect 3532 10772 3572 10781
rect 3112 10604 3480 10613
rect 3112 10555 3480 10564
rect 3532 10184 3572 10732
rect 3532 10135 3572 10144
rect 2860 10100 2900 10109
rect 3436 10100 3476 10109
rect 2900 10060 2996 10100
rect 2860 10051 2900 10060
rect 2956 9848 2996 10060
rect 3436 10016 3476 10060
rect 3436 9965 3476 9976
rect 3628 10016 3668 10025
rect 2764 9808 2996 9848
rect 3052 9932 3092 9941
rect 2668 9512 2708 9521
rect 2572 9472 2668 9512
rect 2572 8924 2612 9472
rect 2668 9463 2708 9472
rect 2572 8875 2612 8884
rect 2668 9260 2708 9269
rect 2476 7195 2516 7204
rect 2572 6992 2612 7001
rect 2572 6488 2612 6952
rect 1132 6355 1172 6364
rect 2284 6404 2324 6413
rect 460 5984 500 5993
rect 460 5849 500 5944
rect 2284 5648 2324 6364
rect 2284 5599 2324 5608
rect 2572 5480 2612 6448
rect 2668 6404 2708 9220
rect 2764 7916 2804 9808
rect 2956 9428 2996 9437
rect 3052 9428 3092 9892
rect 2996 9388 3092 9428
rect 3148 9680 3188 9689
rect 3148 9428 3188 9640
rect 2956 8000 2996 9388
rect 3148 9379 3188 9388
rect 3532 9512 3572 9521
rect 3112 9092 3480 9101
rect 3112 9043 3480 9052
rect 3340 8840 3380 8849
rect 2956 7951 2996 7960
rect 3052 8672 3092 8681
rect 2860 7916 2900 7925
rect 2764 7876 2860 7916
rect 2764 7160 2804 7876
rect 2860 7848 2900 7876
rect 3052 7832 3092 8632
rect 3340 8672 3380 8800
rect 3340 8623 3380 8632
rect 2956 7792 3092 7832
rect 3532 8252 3572 9472
rect 3628 8840 3668 9976
rect 3820 9932 3860 17704
rect 3916 14384 3956 20560
rect 4012 19172 4052 19181
rect 4012 19088 4052 19132
rect 4108 19088 4148 21484
rect 4204 20768 4244 22156
rect 4876 22196 4916 22205
rect 4876 22061 4916 22156
rect 4352 21944 4720 21953
rect 4352 21895 4720 21904
rect 4972 21776 5012 22240
rect 4972 21727 5012 21736
rect 4492 21692 4532 21701
rect 4204 20719 4244 20728
rect 4396 21020 4436 21029
rect 4396 20852 4436 20980
rect 4492 20936 4532 21652
rect 4780 21524 4820 21619
rect 4780 21475 4820 21484
rect 4876 21608 4916 21617
rect 4492 20887 4532 20896
rect 4588 21356 4628 21365
rect 4396 20600 4436 20812
rect 4588 20768 4628 21316
rect 4588 20719 4628 20728
rect 4780 21272 4820 21281
rect 4396 20551 4436 20560
rect 4352 20432 4720 20441
rect 4352 20383 4720 20392
rect 4588 20264 4628 20273
rect 4300 20012 4340 20021
rect 4300 19877 4340 19972
rect 4396 19844 4436 19853
rect 4396 19508 4436 19804
rect 4396 19459 4436 19468
rect 4300 19256 4340 19351
rect 4588 19340 4628 20224
rect 4684 20096 4724 20105
rect 4684 19961 4724 20056
rect 4588 19291 4628 19300
rect 4300 19207 4340 19216
rect 4300 19088 4340 19097
rect 4012 19048 4300 19088
rect 4300 19039 4340 19048
rect 4352 18920 4720 18929
rect 4352 18871 4720 18880
rect 4780 18752 4820 21232
rect 4876 20264 4916 21568
rect 4972 21524 5012 21533
rect 4972 20768 5012 21484
rect 5068 21104 5108 22324
rect 5068 21055 5108 21064
rect 4972 20633 5012 20728
rect 5068 20936 5108 20945
rect 4876 20215 4916 20224
rect 5068 19844 5108 20896
rect 5164 20852 5204 20861
rect 5164 20264 5204 20812
rect 5260 20684 5300 20693
rect 5356 20684 5396 23080
rect 5452 23071 5492 23080
rect 5644 23204 5684 23213
rect 5452 22448 5492 22543
rect 5452 22399 5492 22408
rect 5548 22364 5588 22373
rect 5452 22280 5492 22289
rect 5452 22145 5492 22240
rect 5548 22112 5588 22324
rect 5548 22063 5588 22072
rect 5644 22028 5684 23164
rect 5740 23120 5780 23332
rect 5740 23071 5780 23080
rect 5836 23036 5876 23045
rect 5836 22364 5876 22996
rect 5836 22315 5876 22324
rect 5740 22280 5780 22291
rect 5740 22196 5780 22240
rect 5740 22112 5780 22156
rect 5740 22032 5780 22072
rect 5644 21979 5684 21988
rect 5932 21692 5972 23668
rect 6124 23540 6164 23549
rect 6124 22532 6164 23500
rect 6124 22483 6164 22492
rect 6124 22196 6164 22205
rect 5740 21652 5972 21692
rect 6028 21776 6068 21785
rect 5300 20644 5396 20684
rect 5452 21608 5492 21617
rect 5260 20635 5300 20644
rect 5452 20432 5492 21568
rect 5548 21608 5588 21648
rect 5740 21608 5780 21652
rect 6028 21641 6068 21736
rect 5548 21524 5588 21568
rect 5548 21020 5588 21484
rect 5548 20971 5588 20980
rect 5644 21568 5780 21608
rect 5548 20852 5588 20861
rect 5548 20717 5588 20812
rect 5452 20383 5492 20392
rect 5164 20096 5204 20224
rect 5164 20047 5204 20056
rect 5356 20264 5396 20273
rect 5356 20096 5396 20224
rect 5356 20047 5396 20056
rect 5068 19795 5108 19804
rect 5260 20012 5300 20021
rect 5644 20012 5684 21568
rect 5932 21524 5972 21533
rect 5740 21440 5780 21449
rect 5740 20936 5780 21400
rect 5740 20887 5780 20896
rect 5836 20852 5876 20861
rect 5740 20600 5780 20609
rect 5740 20180 5780 20560
rect 5836 20264 5876 20812
rect 5836 20215 5876 20224
rect 5740 20131 5780 20140
rect 5836 20096 5876 20105
rect 5644 19972 5780 20012
rect 5260 19340 5300 19972
rect 5260 19291 5300 19300
rect 4588 18712 4820 18752
rect 5068 19256 5108 19265
rect 5068 18752 5108 19216
rect 4108 18584 4148 18593
rect 4012 17240 4052 17249
rect 4012 16064 4052 17200
rect 4108 17156 4148 18544
rect 4204 17912 4244 18007
rect 4204 17863 4244 17872
rect 4396 17828 4436 17837
rect 4204 17744 4244 17753
rect 4204 17609 4244 17704
rect 4396 17744 4436 17788
rect 4396 17693 4436 17704
rect 4588 17660 4628 18712
rect 5068 18703 5108 18712
rect 5164 19172 5204 19181
rect 4588 17611 4628 17620
rect 4684 18584 4724 18593
rect 4684 17576 4724 18544
rect 4972 18584 5012 18593
rect 4876 18500 4916 18509
rect 4684 17527 4724 17536
rect 4780 17744 4820 17753
rect 4352 17408 4720 17417
rect 4352 17359 4720 17368
rect 4108 16316 4148 17116
rect 4492 17240 4532 17249
rect 4492 17105 4532 17200
rect 4780 17156 4820 17704
rect 4780 17107 4820 17116
rect 4588 17072 4628 17081
rect 4492 16904 4532 16913
rect 4492 16769 4532 16864
rect 4108 16148 4148 16276
rect 4108 16099 4148 16108
rect 4588 16148 4628 17032
rect 4684 16988 4724 16997
rect 4724 16948 4820 16988
rect 4684 16939 4724 16948
rect 4588 16099 4628 16108
rect 4012 16015 4052 16024
rect 4684 16064 4724 16159
rect 4684 16015 4724 16024
rect 4352 15896 4720 15905
rect 4352 15847 4720 15856
rect 4012 15812 4052 15821
rect 4052 15772 4148 15812
rect 4012 15763 4052 15772
rect 4012 15560 4052 15655
rect 4012 15511 4052 15520
rect 4108 15476 4148 15772
rect 4492 15644 4532 15653
rect 4492 15509 4532 15604
rect 4684 15644 4724 15653
rect 4108 15427 4148 15436
rect 4588 15476 4628 15485
rect 4588 15341 4628 15436
rect 4204 15308 4244 15317
rect 4204 14972 4244 15268
rect 4204 14923 4244 14932
rect 4588 15224 4628 15233
rect 4588 14804 4628 15184
rect 4588 14755 4628 14764
rect 4684 14720 4724 15604
rect 4780 14720 4820 16948
rect 4876 16484 4916 18460
rect 4972 17912 5012 18544
rect 4972 17863 5012 17872
rect 5068 18500 5108 18509
rect 5068 17828 5108 18460
rect 5068 17779 5108 17788
rect 4972 17660 5012 17669
rect 4972 17240 5012 17620
rect 4972 17072 5012 17200
rect 4972 17023 5012 17032
rect 5068 17408 5108 17417
rect 5068 17324 5108 17368
rect 4876 16435 4916 16444
rect 4972 16232 5012 16241
rect 4876 16064 4916 16073
rect 4876 15728 4916 16024
rect 4876 15679 4916 15688
rect 4972 15644 5012 16192
rect 5068 15728 5108 17284
rect 5164 15812 5204 19132
rect 5356 19172 5396 19181
rect 5260 18752 5300 18761
rect 5260 17660 5300 18712
rect 5356 17996 5396 19132
rect 5548 19172 5588 19181
rect 5356 17828 5396 17956
rect 5356 17779 5396 17788
rect 5452 18584 5492 18593
rect 5260 17611 5300 17620
rect 5452 17576 5492 18544
rect 5548 17660 5588 19132
rect 5740 18668 5780 19972
rect 5836 19424 5876 20056
rect 5836 19375 5876 19384
rect 5740 18628 5876 18668
rect 5548 17611 5588 17620
rect 5740 17744 5780 17753
rect 5356 17536 5452 17576
rect 5260 16988 5300 16997
rect 5260 16853 5300 16948
rect 5356 16400 5396 17536
rect 5452 17527 5492 17536
rect 5452 17240 5492 17249
rect 5452 17072 5492 17200
rect 5740 17240 5780 17704
rect 5452 17023 5492 17032
rect 5548 17156 5588 17165
rect 5740 17156 5780 17200
rect 5356 16351 5396 16360
rect 5356 16232 5396 16241
rect 5164 15763 5204 15772
rect 5260 16064 5300 16073
rect 5068 15679 5108 15688
rect 4972 15140 5012 15604
rect 4972 15091 5012 15100
rect 5164 15476 5204 15485
rect 4876 14888 4916 14897
rect 5164 14888 5204 15436
rect 5260 14972 5300 16024
rect 5356 15896 5396 16192
rect 5356 15847 5396 15856
rect 5260 14923 5300 14932
rect 5356 15728 5396 15737
rect 4916 14848 5204 14888
rect 4876 14839 4916 14848
rect 4780 14680 4916 14720
rect 4492 14636 4532 14645
rect 3916 14335 3956 14344
rect 4204 14552 4244 14561
rect 4204 14216 4244 14512
rect 4492 14501 4532 14596
rect 4588 14552 4628 14647
rect 4684 14636 4724 14680
rect 4684 14596 4820 14636
rect 4588 14503 4628 14512
rect 4352 14384 4720 14393
rect 4352 14335 4720 14344
rect 4204 14176 4340 14216
rect 4204 13964 4244 13973
rect 3916 12536 3956 12545
rect 3916 12401 3956 12496
rect 3820 9883 3860 9892
rect 3916 11948 3956 11957
rect 3820 9596 3860 9605
rect 3628 8791 3668 8800
rect 3724 9260 3764 9269
rect 3724 8840 3764 9220
rect 3724 8791 3764 8800
rect 2860 7160 2900 7169
rect 2764 7120 2860 7160
rect 2860 7092 2900 7120
rect 2956 6572 2996 7792
rect 3112 7580 3480 7589
rect 3112 7531 3480 7540
rect 3340 6908 3380 6917
rect 2956 6523 2996 6532
rect 3052 6656 3092 6665
rect 2668 5648 2708 6364
rect 3052 6236 3092 6616
rect 2668 5599 2708 5608
rect 2956 6196 3092 6236
rect 3340 6236 3380 6868
rect 2956 5648 2996 6196
rect 3340 6187 3380 6196
rect 3112 6068 3480 6077
rect 3112 6019 3480 6028
rect 2956 5599 2996 5608
rect 3532 5564 3572 8212
rect 3628 8672 3668 8681
rect 3628 8168 3668 8632
rect 3628 8119 3668 8128
rect 3820 8084 3860 9556
rect 3916 8672 3956 11908
rect 3916 8168 3956 8632
rect 3916 8119 3956 8128
rect 4012 11696 4052 11705
rect 3820 8035 3860 8044
rect 3916 8000 3956 8009
rect 3628 7328 3668 7337
rect 3628 7160 3668 7288
rect 3628 7111 3668 7120
rect 3916 7244 3956 7960
rect 3916 6992 3956 7204
rect 4012 7160 4052 11656
rect 4204 11528 4244 13924
rect 4300 13208 4340 14176
rect 4300 13159 4340 13168
rect 4396 13880 4436 13889
rect 4396 13040 4436 13840
rect 4780 13292 4820 14596
rect 4780 13243 4820 13252
rect 4396 12991 4436 13000
rect 4876 13040 4916 14680
rect 4972 14552 5012 14561
rect 4972 14048 5012 14512
rect 5164 14552 5204 14848
rect 5164 14503 5204 14512
rect 5356 14468 5396 15688
rect 5068 14384 5108 14393
rect 5068 14132 5108 14344
rect 5068 14083 5108 14092
rect 4972 13999 5012 14008
rect 5356 13964 5396 14428
rect 5452 15644 5492 15653
rect 5452 14216 5492 15604
rect 5452 14167 5492 14176
rect 5548 15560 5588 17116
rect 5548 14132 5588 15520
rect 5548 14083 5588 14092
rect 5644 17116 5780 17156
rect 5644 14720 5684 17116
rect 5740 16988 5780 16999
rect 5740 16904 5780 16948
rect 5740 16855 5780 16864
rect 5836 16652 5876 18628
rect 5932 18164 5972 21484
rect 6028 20348 6068 20357
rect 6028 20096 6068 20308
rect 6028 20012 6068 20056
rect 6124 20096 6164 22156
rect 6220 20852 6260 23752
rect 7180 23708 7220 23717
rect 6700 23624 6740 23633
rect 6316 22532 6356 22541
rect 6316 21776 6356 22492
rect 6316 21727 6356 21736
rect 6412 22280 6452 22320
rect 6412 22196 6452 22240
rect 6220 20600 6260 20812
rect 6220 20551 6260 20560
rect 6316 21608 6356 21617
rect 6316 20264 6356 21568
rect 6316 20215 6356 20224
rect 6124 20047 6164 20056
rect 6412 20096 6452 22156
rect 6604 22196 6644 22205
rect 6604 21860 6644 22156
rect 6604 21811 6644 21820
rect 6604 21608 6644 21617
rect 6604 21473 6644 21568
rect 6700 21356 6740 23584
rect 6796 23204 6836 23213
rect 6796 22364 6836 23164
rect 7180 22532 7220 23668
rect 7276 23624 7316 23836
rect 7276 23575 7316 23584
rect 7180 22483 7220 22492
rect 6796 22315 6836 22324
rect 7084 22028 7124 22037
rect 6988 21608 7028 21617
rect 6796 21524 6836 21533
rect 6796 21389 6836 21484
rect 6988 21440 7028 21568
rect 6700 21307 6740 21316
rect 6796 20768 6836 20777
rect 6412 20047 6452 20056
rect 6508 20684 6548 20693
rect 6028 19172 6068 19972
rect 6508 20012 6548 20644
rect 6604 20600 6644 20609
rect 6604 20264 6644 20560
rect 6604 20215 6644 20224
rect 6700 20264 6740 20273
rect 6700 20180 6740 20224
rect 6796 20264 6836 20728
rect 6796 20215 6836 20224
rect 6700 20100 6740 20140
rect 6508 19963 6548 19972
rect 6892 20096 6932 20105
rect 6892 20012 6932 20056
rect 6604 19928 6644 19937
rect 6220 19760 6260 19769
rect 6220 19340 6260 19720
rect 6604 19508 6644 19888
rect 6604 19459 6644 19468
rect 6220 19291 6260 19300
rect 6028 19123 6068 19132
rect 6124 19256 6164 19265
rect 6124 19121 6164 19216
rect 6604 19256 6644 19265
rect 6316 19172 6356 19181
rect 6124 18920 6164 18929
rect 6124 18584 6164 18880
rect 6124 18535 6164 18544
rect 6220 18500 6260 18509
rect 6316 18500 6356 19132
rect 6508 19172 6548 19181
rect 6508 19037 6548 19132
rect 6260 18460 6356 18500
rect 6412 19004 6452 19013
rect 6412 18500 6452 18964
rect 6604 18752 6644 19216
rect 6892 19256 6932 19972
rect 6892 19121 6932 19216
rect 6988 19088 7028 21400
rect 7084 20600 7124 21988
rect 7084 20551 7124 20560
rect 7180 21524 7220 21533
rect 7180 19592 7220 21484
rect 7276 21440 7316 21449
rect 7276 20936 7316 21400
rect 7372 21020 7412 23836
rect 7468 23288 7508 24676
rect 7660 24380 7700 24389
rect 7660 23792 7700 24340
rect 7660 23743 7700 23752
rect 7852 23708 7892 23717
rect 7468 23120 7508 23248
rect 7564 23540 7604 23549
rect 7564 23204 7604 23500
rect 7564 23155 7604 23164
rect 7468 23071 7508 23080
rect 7852 22952 7892 23668
rect 8044 23708 8084 23717
rect 7852 22903 7892 22912
rect 7948 22868 7988 22963
rect 7948 22819 7988 22828
rect 7756 22784 7796 22793
rect 7468 22364 7508 22373
rect 7468 22196 7508 22324
rect 7468 22147 7508 22156
rect 7564 22364 7604 22373
rect 7564 21944 7604 22324
rect 7660 22280 7700 22289
rect 7660 22145 7700 22240
rect 7564 21895 7604 21904
rect 7660 21860 7700 21869
rect 7660 21776 7700 21820
rect 7660 21725 7700 21736
rect 7372 20971 7412 20980
rect 7468 21692 7508 21701
rect 7276 20887 7316 20896
rect 7468 20852 7508 21652
rect 7564 21524 7604 21533
rect 7564 20936 7604 21484
rect 7564 20887 7604 20896
rect 7468 20803 7508 20812
rect 7660 20852 7700 20861
rect 7276 20768 7316 20777
rect 7276 20633 7316 20728
rect 7276 20432 7316 20441
rect 7276 20180 7316 20392
rect 7276 20131 7316 20140
rect 7180 19543 7220 19552
rect 7372 20096 7412 20105
rect 6988 19039 7028 19048
rect 7276 19172 7316 19181
rect 6604 18703 6644 18712
rect 6892 18920 6932 18929
rect 6892 18752 6932 18880
rect 6892 18703 6932 18712
rect 5932 18124 6164 18164
rect 5932 17912 5972 17921
rect 5932 17660 5972 17872
rect 5932 17611 5972 17620
rect 6028 17324 6068 17333
rect 5740 16612 5876 16652
rect 5932 16988 5972 16997
rect 5740 15728 5780 16612
rect 5740 15679 5780 15688
rect 5836 16484 5876 16493
rect 4972 13628 5012 13637
rect 4972 13124 5012 13588
rect 4972 13075 5012 13084
rect 5164 13292 5204 13301
rect 4876 12991 4916 13000
rect 4352 12872 4720 12881
rect 4352 12823 4720 12832
rect 5068 12536 5108 12545
rect 4876 12452 4916 12461
rect 4876 11948 4916 12412
rect 5068 12368 5108 12496
rect 5068 12319 5108 12328
rect 4876 11696 4916 11908
rect 4876 11647 4916 11656
rect 4972 12284 5012 12293
rect 4204 11479 4244 11488
rect 4876 11528 4916 11537
rect 4352 11360 4720 11369
rect 4352 11311 4720 11320
rect 4780 11192 4820 11201
rect 4204 11024 4244 11033
rect 4204 10889 4244 10984
rect 4108 10268 4148 10277
rect 4108 9764 4148 10228
rect 4352 9848 4720 9857
rect 4352 9799 4720 9808
rect 4108 9596 4148 9724
rect 4108 9547 4148 9556
rect 4684 9512 4724 9521
rect 4300 9344 4340 9353
rect 4300 8504 4340 9304
rect 4588 9344 4628 9353
rect 4588 8756 4628 9304
rect 4684 8924 4724 9472
rect 4684 8875 4724 8884
rect 4588 8707 4628 8716
rect 4300 8455 4340 8464
rect 4352 8336 4720 8345
rect 4352 8287 4720 8296
rect 4012 7111 4052 7120
rect 4204 7328 4244 7337
rect 3916 6943 3956 6952
rect 4108 7076 4148 7085
rect 3532 5515 3572 5524
rect 3916 5648 3956 5657
rect 4108 5648 4148 7036
rect 4204 6404 4244 7288
rect 4352 6824 4720 6833
rect 4352 6775 4720 6784
rect 4780 6488 4820 11152
rect 4876 9932 4916 11488
rect 4972 10940 5012 12244
rect 5068 11612 5108 11621
rect 5068 11024 5108 11572
rect 5164 11108 5204 13252
rect 5164 11059 5204 11068
rect 5260 13124 5300 13133
rect 5068 10975 5108 10984
rect 5260 10940 5300 13084
rect 5356 12788 5396 13924
rect 5548 13964 5588 13973
rect 5644 13964 5684 14680
rect 5588 13924 5684 13964
rect 5740 15560 5780 15569
rect 5548 13915 5588 13924
rect 5740 13292 5780 15520
rect 5836 14216 5876 16444
rect 5932 16148 5972 16948
rect 5932 16013 5972 16108
rect 6028 16652 6068 17284
rect 6028 16316 6068 16612
rect 6124 16568 6164 18124
rect 6220 18080 6260 18460
rect 6412 18451 6452 18460
rect 6700 18584 6740 18593
rect 6220 18031 6260 18040
rect 6604 18248 6644 18257
rect 6220 17912 6260 17923
rect 6220 17828 6260 17872
rect 6220 17779 6260 17788
rect 6604 17828 6644 18208
rect 6604 17779 6644 17788
rect 6508 17660 6548 17669
rect 6412 17576 6452 17585
rect 6220 17240 6260 17249
rect 6220 17156 6260 17200
rect 6220 17105 6260 17116
rect 6124 16519 6164 16528
rect 6220 16904 6260 16913
rect 6220 16484 6260 16864
rect 6220 16400 6260 16444
rect 6220 16349 6260 16360
rect 5932 15308 5972 15317
rect 5932 14762 5972 15268
rect 6028 14888 6068 16276
rect 6220 16232 6260 16241
rect 6220 15644 6260 16192
rect 6220 15595 6260 15604
rect 6412 15140 6452 17536
rect 6508 17240 6548 17620
rect 6508 16988 6548 17200
rect 6508 16232 6548 16948
rect 6508 16183 6548 16192
rect 6604 16820 6644 16829
rect 6412 15091 6452 15100
rect 6508 15896 6548 15905
rect 6028 14839 6068 14848
rect 6124 14804 6164 14813
rect 6316 14804 6356 14813
rect 6164 14764 6260 14804
rect 6124 14755 6164 14764
rect 5932 14713 5972 14722
rect 5836 14167 5876 14176
rect 5740 13243 5780 13252
rect 6028 13292 6068 13301
rect 6220 13292 6260 14764
rect 6316 14384 6356 14764
rect 6508 14636 6548 15856
rect 6604 15560 6644 16780
rect 6700 16400 6740 18544
rect 7084 18584 7124 18593
rect 6892 18332 6932 18341
rect 6796 18164 6836 18173
rect 6796 17744 6836 18124
rect 6796 17072 6836 17704
rect 6796 16568 6836 17032
rect 6796 16519 6836 16528
rect 6700 16351 6740 16360
rect 6796 16232 6836 16241
rect 6700 16064 6740 16073
rect 6700 15980 6740 16024
rect 6700 15929 6740 15940
rect 6796 15812 6836 16192
rect 6796 15763 6836 15772
rect 6892 15896 6932 18292
rect 6892 15644 6932 15856
rect 6892 15595 6932 15604
rect 6988 16568 7028 16577
rect 6988 16484 7028 16528
rect 6604 15511 6644 15520
rect 6700 15476 6740 15485
rect 6508 14587 6548 14596
rect 6604 14804 6644 14813
rect 6316 14335 6356 14344
rect 6412 14552 6452 14561
rect 6412 14216 6452 14512
rect 6412 14167 6452 14176
rect 6068 13252 6164 13292
rect 6028 13243 6068 13252
rect 5836 13208 5876 13217
rect 5356 12739 5396 12748
rect 5452 13040 5492 13049
rect 5452 12620 5492 13000
rect 5836 12788 5876 13168
rect 5836 12739 5876 12748
rect 6028 13040 6068 13049
rect 6028 12704 6068 13000
rect 6028 12655 6068 12664
rect 5452 12571 5492 12580
rect 5836 12620 5876 12629
rect 5836 12536 5876 12580
rect 5836 12485 5876 12496
rect 5740 12368 5780 12377
rect 5780 12328 5876 12368
rect 5740 12319 5780 12328
rect 5740 12116 5780 12125
rect 5740 11948 5780 12076
rect 5740 11899 5780 11908
rect 5836 11780 5876 12328
rect 6124 12116 6164 13252
rect 6220 13157 6260 13252
rect 6412 14048 6452 14057
rect 6316 13040 6356 13049
rect 6316 12620 6356 13000
rect 6316 12571 6356 12580
rect 6124 12067 6164 12076
rect 5740 11696 5780 11705
rect 4972 10891 5012 10900
rect 5164 10900 5300 10940
rect 5548 11612 5588 11621
rect 5548 11024 5588 11572
rect 5068 10856 5108 10865
rect 5068 10184 5108 10816
rect 4876 9883 4916 9892
rect 4972 10016 5012 10025
rect 4972 9881 5012 9976
rect 5068 9512 5108 10144
rect 5164 9680 5204 10900
rect 5548 10436 5588 10984
rect 5740 10940 5780 11656
rect 5740 10891 5780 10900
rect 5548 10387 5588 10396
rect 5644 10604 5684 10613
rect 5644 10184 5684 10564
rect 5164 9631 5204 9640
rect 5260 10100 5300 10109
rect 5068 9463 5108 9472
rect 5260 9428 5300 10060
rect 5260 9379 5300 9388
rect 5452 9848 5492 9857
rect 5452 9344 5492 9808
rect 5260 8756 5300 8765
rect 5452 8756 5492 9304
rect 5300 8716 5492 8756
rect 5260 8707 5300 8716
rect 5452 8672 5492 8716
rect 5452 8623 5492 8632
rect 5068 8588 5108 8597
rect 4876 8504 4916 8513
rect 4876 7916 4916 8464
rect 4972 8168 5012 8177
rect 4972 8000 5012 8128
rect 4972 7951 5012 7960
rect 4876 7867 4916 7876
rect 5068 7160 5108 8548
rect 5260 8504 5300 8513
rect 5260 8000 5300 8464
rect 5260 7951 5300 7960
rect 5644 8168 5684 10144
rect 5836 8924 5876 11740
rect 6028 11696 6068 11705
rect 5932 11612 5972 11621
rect 5932 11192 5972 11572
rect 6028 11561 6068 11656
rect 6316 11696 6356 11705
rect 5932 11143 5972 11152
rect 6220 11528 6260 11537
rect 6028 10940 6068 10949
rect 5836 8875 5876 8884
rect 5932 9512 5972 9521
rect 5068 6656 5108 7120
rect 5068 6607 5108 6616
rect 5644 7244 5684 8128
rect 5932 7916 5972 9472
rect 4780 6439 4820 6448
rect 5452 6488 5492 6497
rect 4204 6355 4244 6364
rect 4204 5648 4244 5657
rect 4108 5608 4204 5648
rect 3916 5513 3956 5608
rect 2572 5431 2612 5440
rect 4204 5480 4244 5608
rect 4780 5648 4820 5657
rect 4780 5513 4820 5608
rect 4204 5431 4244 5440
rect 4352 5312 4720 5321
rect 4352 5263 4720 5272
rect 5452 5060 5492 6448
rect 5548 6404 5588 6413
rect 5548 5480 5588 6364
rect 5548 5431 5588 5440
rect 5452 5011 5492 5020
rect 5644 4976 5684 7204
rect 5836 7876 5972 7916
rect 5740 6404 5780 6413
rect 5740 5900 5780 6364
rect 5836 6236 5876 7876
rect 5932 7748 5972 7757
rect 5932 6488 5972 7708
rect 6028 7412 6068 10900
rect 6220 10352 6260 11488
rect 6316 10436 6356 11656
rect 6412 11696 6452 14008
rect 6604 13208 6644 14764
rect 6604 12536 6644 13168
rect 6604 12368 6644 12496
rect 6604 12319 6644 12328
rect 6700 14552 6740 15436
rect 6796 15392 6836 15401
rect 6988 15392 7028 16444
rect 7084 16148 7124 18544
rect 7180 18584 7220 18593
rect 7276 18584 7316 19132
rect 7220 18544 7316 18584
rect 7180 17996 7220 18544
rect 7180 17947 7220 17956
rect 7276 17660 7316 17669
rect 7276 17525 7316 17620
rect 7276 17324 7316 17333
rect 7180 17156 7220 17165
rect 7180 17021 7220 17116
rect 7180 16820 7220 16829
rect 7180 16316 7220 16780
rect 7180 16267 7220 16276
rect 7084 16099 7124 16108
rect 7276 15980 7316 17284
rect 7372 16904 7412 20056
rect 7468 19844 7508 19853
rect 7468 17828 7508 19804
rect 7660 19340 7700 20812
rect 7756 20348 7796 22744
rect 7852 22784 7892 22793
rect 7852 22700 7892 22744
rect 7852 22448 7892 22660
rect 7948 22532 7988 22560
rect 8044 22532 8084 23668
rect 8332 23708 8372 25264
rect 8428 24380 8468 26524
rect 8620 25892 8660 25901
rect 8620 25304 8660 25852
rect 8620 25255 8660 25264
rect 9004 25724 9044 25733
rect 8524 25220 8564 25229
rect 8524 25085 8564 25180
rect 8812 24968 8852 24977
rect 8428 24331 8468 24340
rect 8524 24632 8564 24641
rect 8236 23624 8276 23633
rect 7988 22492 8084 22532
rect 7948 22483 7988 22492
rect 7852 22399 7892 22408
rect 8044 22112 8084 22492
rect 8044 22063 8084 22072
rect 8140 23288 8180 23297
rect 8044 21524 8084 21533
rect 7948 21188 7988 21197
rect 7948 21020 7988 21148
rect 7948 20971 7988 20980
rect 8044 21020 8084 21484
rect 7852 20684 7892 20693
rect 7852 20549 7892 20644
rect 7756 20299 7796 20308
rect 7948 20516 7988 20525
rect 7852 19844 7892 19853
rect 7852 19709 7892 19804
rect 7660 19291 7700 19300
rect 7756 19256 7796 19265
rect 7756 18752 7796 19216
rect 7756 18703 7796 18712
rect 7756 18584 7796 18595
rect 7468 17779 7508 17788
rect 7564 18500 7604 18509
rect 7468 17660 7508 17669
rect 7468 17324 7508 17620
rect 7468 16988 7508 17284
rect 7468 16939 7508 16948
rect 7372 16855 7412 16864
rect 7564 16316 7604 18460
rect 7756 18500 7796 18544
rect 7756 18451 7796 18460
rect 7852 18416 7892 18425
rect 7756 18332 7796 18341
rect 7660 17576 7700 17585
rect 7660 16652 7700 17536
rect 7660 16603 7700 16612
rect 7564 16267 7604 16276
rect 7276 15931 7316 15940
rect 7564 16148 7604 16157
rect 7564 15728 7604 16108
rect 7564 15679 7604 15688
rect 7660 15644 7700 15653
rect 7660 15392 7700 15604
rect 6988 15352 7124 15392
rect 6796 15257 6836 15352
rect 6700 12536 6740 14512
rect 6796 15140 6836 15149
rect 6796 14132 6836 15100
rect 6796 14083 6836 14092
rect 6892 14888 6932 14897
rect 6796 13964 6836 13973
rect 6796 13544 6836 13924
rect 6796 13495 6836 13504
rect 6892 13880 6932 14848
rect 6892 13376 6932 13840
rect 6892 13327 6932 13336
rect 6988 14384 7028 14393
rect 6412 11647 6452 11656
rect 6316 10387 6356 10396
rect 6412 11360 6452 11369
rect 6412 10940 6452 11320
rect 6220 9512 6260 10312
rect 6220 9463 6260 9472
rect 6412 9512 6452 10900
rect 6700 11108 6740 12496
rect 6796 13292 6836 13301
rect 6796 11948 6836 13252
rect 6988 13292 7028 14344
rect 6988 13243 7028 13252
rect 6892 12956 6932 12965
rect 6892 12452 6932 12916
rect 6892 12403 6932 12412
rect 6796 11899 6836 11908
rect 7084 11780 7124 15352
rect 7660 15343 7700 15352
rect 7468 15056 7508 15065
rect 7180 14804 7220 14813
rect 7180 14216 7220 14764
rect 7468 14804 7508 15016
rect 7468 14755 7508 14764
rect 7180 14167 7220 14176
rect 7276 14552 7316 14561
rect 7084 11731 7124 11740
rect 7180 11948 7220 11957
rect 6604 10184 6644 10193
rect 6604 9596 6644 10144
rect 6604 9547 6644 9556
rect 6412 9463 6452 9472
rect 6700 9512 6740 11068
rect 7180 11024 7220 11908
rect 7276 11192 7316 14512
rect 7756 14216 7796 18292
rect 7852 17576 7892 18376
rect 7852 17527 7892 17536
rect 7852 17240 7892 17249
rect 7852 16988 7892 17200
rect 7852 16939 7892 16948
rect 7852 16820 7892 16829
rect 7852 16685 7892 16780
rect 7852 16400 7892 16409
rect 7852 16232 7892 16360
rect 7852 16148 7892 16192
rect 7852 16068 7892 16108
rect 7948 16064 7988 20476
rect 8044 20432 8084 20980
rect 8044 20383 8084 20392
rect 8140 20096 8180 23248
rect 8236 23120 8276 23584
rect 8236 23071 8276 23080
rect 8236 22112 8276 22121
rect 8236 21977 8276 22072
rect 8236 21692 8276 21701
rect 8236 21440 8276 21652
rect 8236 21391 8276 21400
rect 8236 20936 8276 21031
rect 8236 20887 8276 20896
rect 8236 20768 8276 20777
rect 8236 20600 8276 20728
rect 8236 20264 8276 20560
rect 8236 20215 8276 20224
rect 8140 20047 8180 20056
rect 8140 19928 8180 19937
rect 8044 17828 8084 17837
rect 8044 17408 8084 17788
rect 8044 17359 8084 17368
rect 8044 17072 8084 17081
rect 8044 16736 8084 17032
rect 8140 16820 8180 19888
rect 8236 18584 8276 18593
rect 8236 18449 8276 18544
rect 8332 17744 8372 23668
rect 8524 22952 8564 24592
rect 8716 24548 8756 24557
rect 8716 24413 8756 24508
rect 8620 24044 8660 24053
rect 8812 24044 8852 24928
rect 9004 24548 9044 25684
rect 9100 25388 9140 28540
rect 9100 25339 9140 25348
rect 9196 28496 9236 28505
rect 9196 25220 9236 28456
rect 9292 27740 9332 28600
rect 10060 28244 10100 28600
rect 10060 28204 10292 28244
rect 9292 27691 9332 27700
rect 10060 27740 10100 27749
rect 10060 27605 10100 27700
rect 9580 27572 9620 27581
rect 9580 27068 9620 27532
rect 9580 27019 9620 27028
rect 9580 26648 9620 26657
rect 9580 26228 9620 26608
rect 9580 26179 9620 26188
rect 10156 26648 10196 26657
rect 9388 26144 9428 26153
rect 8660 24004 8852 24044
rect 8908 24508 9004 24548
rect 8620 23995 8660 24004
rect 8524 22903 8564 22912
rect 8620 23792 8660 23801
rect 8428 22868 8468 22877
rect 8428 22616 8468 22828
rect 8428 22567 8468 22576
rect 8524 22532 8564 22541
rect 8428 22448 8468 22457
rect 8428 22313 8468 22408
rect 8524 22397 8564 22492
rect 8620 22364 8660 23752
rect 8812 23624 8852 23633
rect 8812 23540 8852 23584
rect 8812 23489 8852 23500
rect 8908 23120 8948 24508
rect 9004 24499 9044 24508
rect 9100 25180 9236 25220
rect 9292 25304 9332 25313
rect 9100 23876 9140 25180
rect 9292 25136 9332 25264
rect 9100 23827 9140 23836
rect 9196 25096 9332 25136
rect 9196 23792 9236 25096
rect 9388 24716 9428 26104
rect 10060 25640 10100 25668
rect 9964 25600 10060 25640
rect 9388 24667 9428 24676
rect 9772 24716 9812 24725
rect 9196 23708 9236 23752
rect 9292 24632 9332 24641
rect 9292 23792 9332 24592
rect 9484 24632 9524 24641
rect 9484 24548 9524 24592
rect 9292 23743 9332 23752
rect 9388 24508 9524 24548
rect 9100 23668 9196 23708
rect 8908 23071 8948 23080
rect 9004 23204 9044 23213
rect 8812 22952 8852 22961
rect 8620 22315 8660 22324
rect 8716 22868 8756 22877
rect 8524 22280 8564 22289
rect 8524 21860 8564 22240
rect 8524 21811 8564 21820
rect 8428 21608 8468 21617
rect 8428 21473 8468 21568
rect 8428 21272 8468 21281
rect 8428 20432 8468 21232
rect 8524 20852 8564 20861
rect 8524 20768 8564 20812
rect 8524 20717 8564 20728
rect 8620 20852 8660 20861
rect 8620 20768 8660 20812
rect 8620 20717 8660 20728
rect 8428 20383 8468 20392
rect 8620 20180 8660 20189
rect 8524 18836 8564 18845
rect 8524 18701 8564 18796
rect 8620 18668 8660 20140
rect 8716 20096 8756 22828
rect 8812 22616 8852 22912
rect 8908 22952 8948 22961
rect 8908 22868 8948 22912
rect 8908 22817 8948 22828
rect 8812 22567 8852 22576
rect 9004 22196 9044 23164
rect 9004 22147 9044 22156
rect 8908 22028 8948 22037
rect 8812 21944 8852 21953
rect 8812 21104 8852 21904
rect 8812 21055 8852 21064
rect 8716 20047 8756 20056
rect 8812 20936 8852 20945
rect 8236 17660 8276 17669
rect 8236 17156 8276 17620
rect 8236 17107 8276 17116
rect 8140 16780 8276 16820
rect 8044 16687 8084 16696
rect 8044 16400 8084 16409
rect 8044 16316 8084 16360
rect 8044 16265 8084 16276
rect 7948 16015 7988 16024
rect 8044 16148 8084 16157
rect 8044 15980 8084 16108
rect 8044 15931 8084 15940
rect 8140 15560 8180 15569
rect 7948 15476 7988 15485
rect 7948 15341 7988 15436
rect 8140 14804 8180 15520
rect 8044 14720 8084 14729
rect 8044 14585 8084 14680
rect 7756 14167 7796 14176
rect 7468 14048 7508 14057
rect 7372 13796 7412 13805
rect 7372 13208 7412 13756
rect 7372 13159 7412 13168
rect 7468 12980 7508 14008
rect 7372 12940 7508 12980
rect 7564 13964 7604 13973
rect 7372 11948 7412 12940
rect 7372 11899 7412 11908
rect 7468 12536 7508 12545
rect 7564 12536 7604 13924
rect 7756 13628 7796 13637
rect 7756 13124 7796 13588
rect 8044 13544 8084 13553
rect 7756 12989 7796 13084
rect 7852 13208 7892 13217
rect 7852 13073 7892 13168
rect 8044 13124 8084 13504
rect 8140 13460 8180 14764
rect 8236 14636 8276 16780
rect 8332 14720 8372 17704
rect 8428 18500 8468 18509
rect 8428 17240 8468 18460
rect 8428 17191 8468 17200
rect 8524 18332 8564 18341
rect 8428 16904 8468 16913
rect 8428 16820 8468 16864
rect 8428 16769 8468 16780
rect 8428 16400 8468 16409
rect 8428 16316 8468 16360
rect 8428 16265 8468 16276
rect 8428 16148 8468 16157
rect 8428 16013 8468 16108
rect 8332 14671 8372 14680
rect 8428 15476 8468 15485
rect 8236 14587 8276 14596
rect 8428 13880 8468 15436
rect 8524 14888 8564 18292
rect 8620 17828 8660 18628
rect 8716 19088 8756 19097
rect 8716 18416 8756 19048
rect 8716 18367 8756 18376
rect 8620 17779 8660 17788
rect 8716 18080 8756 18089
rect 8716 17912 8756 18040
rect 8620 17660 8660 17669
rect 8620 17525 8660 17620
rect 8716 16148 8756 17872
rect 8812 17240 8852 20896
rect 8908 19844 8948 21988
rect 9100 21104 9140 23668
rect 9196 23657 9236 23668
rect 9196 23372 9236 23381
rect 9196 22028 9236 23332
rect 9388 23372 9428 24508
rect 9676 23792 9716 23801
rect 9388 23323 9428 23332
rect 9484 23456 9524 23465
rect 9196 21979 9236 21988
rect 9100 21055 9140 21064
rect 9196 21860 9236 21869
rect 9196 21020 9236 21820
rect 9004 20852 9044 20861
rect 9004 20768 9044 20812
rect 9004 20717 9044 20728
rect 9196 20684 9236 20980
rect 9196 20635 9236 20644
rect 9292 21776 9332 21785
rect 9196 20516 9236 20525
rect 9196 20264 9236 20476
rect 9196 20215 9236 20224
rect 8908 19795 8948 19804
rect 9196 19340 9236 19349
rect 9004 19256 9044 19265
rect 8908 19172 8948 19181
rect 8908 18920 8948 19132
rect 9004 19121 9044 19216
rect 9196 19004 9236 19300
rect 9196 18955 9236 18964
rect 8908 18871 8948 18880
rect 9196 18836 9236 18845
rect 8812 17191 8852 17200
rect 8908 18668 8948 18677
rect 8716 16099 8756 16108
rect 8812 17072 8852 17081
rect 8812 15896 8852 17032
rect 8716 15856 8852 15896
rect 8620 15560 8660 15569
rect 8620 15425 8660 15520
rect 8524 14839 8564 14848
rect 8428 13831 8468 13840
rect 8524 14720 8564 14729
rect 8524 13880 8564 14680
rect 8524 13831 8564 13840
rect 8620 14048 8660 14057
rect 8140 13411 8180 13420
rect 8044 13075 8084 13084
rect 8332 13250 8372 13259
rect 7756 12704 7796 12713
rect 7756 12620 7796 12664
rect 7756 12569 7796 12580
rect 7508 12496 7604 12536
rect 7276 11143 7316 11152
rect 7372 11780 7412 11789
rect 7180 10975 7220 10984
rect 6700 9463 6740 9472
rect 6988 10940 7028 10949
rect 6988 9512 7028 10900
rect 7372 10940 7412 11740
rect 7372 10891 7412 10900
rect 7468 11024 7508 12496
rect 8044 12452 8084 12461
rect 8332 12452 8372 13210
rect 8620 12956 8660 14008
rect 8716 13880 8756 15856
rect 8716 13831 8756 13840
rect 8812 15728 8852 15737
rect 8812 14804 8852 15688
rect 8812 13796 8852 14764
rect 8812 13747 8852 13756
rect 8812 13628 8852 13637
rect 8812 13493 8852 13588
rect 8716 13208 8756 13217
rect 8716 13073 8756 13168
rect 8620 12907 8660 12916
rect 8812 13040 8852 13049
rect 8812 12620 8852 13000
rect 8812 12571 8852 12580
rect 8084 12412 8372 12452
rect 7468 10889 7508 10984
rect 7564 11948 7604 11957
rect 7180 10772 7220 10781
rect 7180 10268 7220 10732
rect 7564 10688 7604 11908
rect 7660 11612 7700 11621
rect 7660 11192 7700 11572
rect 7660 11143 7700 11152
rect 7948 11528 7988 11537
rect 7948 11024 7988 11488
rect 8044 11108 8084 12412
rect 8332 12200 8372 12412
rect 8620 12536 8660 12545
rect 8620 12452 8660 12496
rect 8620 12401 8660 12412
rect 8812 12452 8852 12461
rect 8332 12151 8372 12160
rect 8716 11612 8756 11621
rect 8044 11059 8084 11068
rect 8140 11528 8180 11537
rect 7948 10975 7988 10984
rect 7564 10639 7604 10648
rect 7660 10940 7700 10949
rect 7660 10436 7700 10900
rect 7660 10387 7700 10396
rect 7180 10219 7220 10228
rect 7276 10184 7316 10193
rect 7180 9932 7220 9941
rect 7180 9596 7220 9892
rect 7276 9680 7316 10144
rect 7948 10184 7988 10193
rect 7276 9631 7316 9640
rect 7660 10016 7700 10025
rect 7180 9547 7220 9556
rect 7372 9512 7412 9521
rect 6700 9260 6740 9269
rect 6028 7363 6068 7372
rect 6124 9176 6164 9185
rect 6124 7076 6164 9136
rect 6124 6992 6164 7036
rect 6604 8756 6644 8765
rect 6604 8000 6644 8716
rect 6412 6992 6452 7001
rect 6124 6952 6412 6992
rect 6412 6943 6452 6952
rect 5932 6439 5972 6448
rect 6412 6488 6452 6497
rect 6452 6448 6548 6488
rect 6412 6439 6452 6448
rect 5836 6187 5876 6196
rect 6412 6236 6452 6245
rect 5740 5851 5780 5860
rect 6220 5648 6260 5657
rect 6124 5564 6164 5573
rect 6124 5312 6164 5524
rect 6220 5513 6260 5608
rect 6124 5263 6164 5272
rect 6412 5144 6452 6196
rect 6508 5816 6548 6448
rect 6508 5767 6548 5776
rect 6604 6236 6644 7960
rect 6604 5648 6644 6196
rect 6700 6488 6740 9220
rect 6988 8840 7028 9472
rect 6892 7748 6932 7757
rect 6892 7202 6932 7708
rect 6892 7153 6932 7162
rect 6700 6068 6740 6448
rect 6700 6019 6740 6028
rect 6988 6572 7028 8800
rect 7276 9472 7372 9512
rect 7180 8672 7220 8681
rect 7180 8000 7220 8632
rect 7180 7951 7220 7960
rect 7180 7832 7220 7841
rect 7276 7832 7316 9472
rect 7372 9463 7412 9472
rect 7660 9512 7700 9976
rect 7948 9596 7988 10144
rect 8140 10184 8180 11488
rect 8524 11024 8564 11033
rect 8140 10135 8180 10144
rect 8428 10856 8468 10865
rect 8428 10184 8468 10816
rect 8524 10520 8564 10984
rect 8524 10471 8564 10480
rect 8620 10940 8660 10949
rect 8428 10135 8468 10144
rect 7948 9547 7988 9556
rect 8140 10016 8180 10025
rect 7468 9428 7508 9437
rect 7372 8679 7412 8688
rect 7372 8168 7412 8639
rect 7468 8252 7508 9388
rect 7660 8672 7700 9472
rect 7660 8623 7700 8632
rect 8140 8588 8180 9976
rect 8524 9932 8564 9941
rect 8236 9512 8276 9521
rect 8236 8672 8276 9472
rect 8236 8623 8276 8632
rect 8524 9512 8564 9892
rect 8620 9680 8660 10900
rect 8620 9631 8660 9640
rect 8140 8539 8180 8548
rect 7468 8203 7508 8212
rect 7372 8119 7412 8128
rect 8236 8084 8276 8093
rect 7220 7792 7316 7832
rect 7372 8000 7412 8009
rect 7180 7412 7220 7792
rect 7180 7363 7220 7372
rect 6604 5599 6644 5608
rect 6988 5648 7028 6532
rect 7276 6488 7316 6497
rect 7276 6236 7316 6448
rect 7276 6187 7316 6196
rect 6988 5396 7028 5608
rect 6988 5347 7028 5356
rect 6412 5095 6452 5104
rect 7180 5312 7220 5321
rect 7372 5312 7412 7960
rect 8140 7832 8180 7841
rect 8236 7832 8276 8044
rect 8428 8000 8468 8009
rect 8180 7792 8276 7832
rect 8332 7916 8372 7925
rect 8140 7783 8180 7792
rect 8044 7748 8084 7757
rect 8044 7244 8084 7708
rect 8044 7195 8084 7204
rect 8332 7160 8372 7876
rect 8332 7111 8372 7120
rect 8428 6992 8468 7960
rect 8428 6943 8468 6952
rect 8044 6488 8084 6497
rect 7948 6152 7988 6161
rect 7220 5272 7412 5312
rect 7564 5564 7604 5573
rect 5644 4927 5684 4936
rect 6220 4892 6260 4901
rect 3112 4556 3480 4565
rect 3112 4507 3480 4516
rect 6220 4304 6260 4852
rect 6220 4255 6260 4264
rect 7180 4304 7220 5272
rect 7180 4255 7220 4264
rect 7564 4136 7604 5524
rect 7564 4087 7604 4096
rect 7948 4472 7988 6112
rect 8044 5732 8084 6448
rect 8044 5683 8084 5692
rect 8524 6488 8564 9472
rect 8716 8000 8756 11572
rect 8812 11192 8852 12412
rect 8908 12368 8948 18628
rect 9100 18584 9140 18593
rect 9196 18584 9236 18796
rect 9292 18668 9332 21736
rect 9388 21524 9428 21533
rect 9388 21389 9428 21484
rect 9388 21020 9428 21029
rect 9388 20768 9428 20980
rect 9388 20719 9428 20728
rect 9388 20600 9428 20609
rect 9388 20096 9428 20560
rect 9388 20047 9428 20056
rect 9388 19256 9428 19296
rect 9388 19172 9428 19216
rect 9388 18836 9428 19132
rect 9388 18787 9428 18796
rect 9292 18628 9428 18668
rect 9196 18544 9332 18584
rect 9004 18332 9044 18341
rect 9004 17156 9044 18292
rect 9100 18080 9140 18544
rect 9196 18248 9236 18257
rect 9196 18113 9236 18208
rect 9100 18031 9140 18040
rect 9004 17107 9044 17116
rect 9100 17912 9140 17921
rect 9100 16988 9140 17872
rect 9196 17744 9236 17753
rect 9196 17576 9236 17704
rect 9196 17441 9236 17536
rect 9004 16948 9140 16988
rect 9196 17240 9236 17249
rect 9004 14552 9044 16948
rect 9100 16820 9140 16829
rect 9100 16148 9140 16780
rect 9196 16484 9236 17200
rect 9196 16435 9236 16444
rect 9100 15896 9140 16108
rect 9100 15476 9140 15856
rect 9196 16316 9236 16325
rect 9196 15644 9236 16276
rect 9292 16064 9332 18544
rect 9388 17660 9428 18628
rect 9484 18080 9524 23416
rect 9676 23204 9716 23752
rect 9676 22532 9716 23164
rect 9676 22483 9716 22492
rect 9676 22196 9716 22205
rect 9580 21776 9620 21785
rect 9580 21641 9620 21736
rect 9676 21188 9716 22156
rect 9676 21139 9716 21148
rect 9676 21020 9716 21029
rect 9580 20852 9620 20861
rect 9580 19256 9620 20812
rect 9676 20348 9716 20980
rect 9676 20299 9716 20308
rect 9772 20180 9812 24676
rect 9964 24380 10004 25600
rect 10060 25591 10100 25600
rect 10060 25472 10100 25481
rect 10060 24548 10100 25432
rect 10060 24499 10100 24508
rect 10060 24380 10100 24389
rect 9964 24340 10060 24380
rect 10060 24312 10100 24340
rect 9964 24044 10004 24053
rect 9964 23456 10004 24004
rect 10156 23876 10196 26608
rect 10252 24632 10292 28204
rect 10636 27908 10676 27917
rect 10540 27572 10580 27581
rect 10348 27320 10388 27329
rect 10348 26648 10388 27280
rect 10444 27152 10484 27161
rect 10444 27017 10484 27112
rect 10348 26599 10388 26608
rect 10444 26816 10484 26825
rect 10444 26480 10484 26776
rect 10444 25304 10484 26440
rect 10444 24884 10484 25264
rect 10444 24835 10484 24844
rect 10252 24592 10388 24632
rect 10156 23827 10196 23836
rect 10252 24464 10292 24473
rect 10060 23708 10100 23717
rect 10252 23708 10292 24424
rect 10060 23624 10100 23668
rect 10060 23573 10100 23584
rect 10156 23668 10292 23708
rect 10060 23456 10100 23465
rect 9964 23416 10060 23456
rect 10060 23388 10100 23416
rect 10060 22868 10100 22877
rect 10060 22733 10100 22828
rect 9964 22280 10004 22289
rect 9868 21860 9908 21869
rect 9868 21020 9908 21820
rect 9964 21860 10004 22240
rect 10156 22280 10196 23668
rect 10252 23204 10292 23299
rect 10252 23155 10292 23164
rect 10348 23120 10388 24592
rect 10444 24380 10484 24389
rect 10444 23876 10484 24340
rect 10540 24296 10580 27532
rect 10636 25472 10676 27868
rect 10732 27404 10772 27413
rect 10732 26732 10772 27364
rect 10828 27404 10868 28600
rect 10828 27355 10868 27364
rect 11308 27656 11348 27665
rect 10886 27236 11254 27245
rect 10886 27187 11254 27196
rect 11212 27068 11252 27077
rect 11212 26933 11252 27028
rect 10924 26900 10964 26909
rect 10924 26765 10964 26860
rect 10732 26683 10772 26692
rect 11116 26648 11156 26657
rect 11116 26312 11156 26608
rect 11116 26263 11156 26272
rect 10886 25724 11254 25733
rect 10886 25675 11254 25684
rect 10636 25423 10676 25432
rect 10732 25388 10772 25397
rect 10540 24247 10580 24256
rect 10636 24884 10676 24893
rect 10444 23827 10484 23836
rect 10540 23960 10580 23971
rect 10540 23876 10580 23920
rect 10540 23827 10580 23836
rect 10636 23708 10676 24844
rect 10444 23540 10484 23549
rect 10444 23456 10484 23500
rect 10444 23405 10484 23416
rect 10636 23372 10676 23668
rect 10636 23323 10676 23332
rect 10732 23204 10772 25348
rect 10828 25304 10868 25313
rect 10828 25169 10868 25264
rect 11020 25136 11060 25145
rect 11020 24884 11060 25096
rect 11020 24835 11060 24844
rect 11308 24800 11348 27616
rect 11596 26816 11636 28600
rect 12364 28160 12404 28600
rect 12364 28111 12404 28120
rect 13036 28160 13076 28169
rect 12126 27992 12494 28001
rect 12126 27943 12494 27952
rect 12940 27740 12980 27749
rect 12172 27656 12212 27665
rect 12172 27521 12212 27616
rect 12076 27320 12116 27329
rect 12076 27068 12116 27280
rect 12076 27019 12116 27028
rect 11596 26767 11636 26776
rect 11692 26984 11732 26993
rect 11596 26648 11636 26657
rect 11596 26228 11636 26608
rect 11596 26179 11636 26188
rect 11404 26060 11444 26069
rect 11404 25304 11444 26020
rect 11692 25556 11732 26944
rect 12172 26900 12212 26911
rect 11980 26816 12020 26825
rect 11788 26564 11828 26573
rect 11788 25976 11828 26524
rect 11884 26396 11924 26405
rect 11884 26261 11924 26356
rect 11788 25927 11828 25936
rect 11692 25507 11732 25516
rect 11788 25472 11828 25481
rect 11404 25052 11444 25264
rect 11692 25304 11732 25315
rect 11692 25220 11732 25264
rect 11692 25171 11732 25180
rect 11596 25052 11636 25061
rect 11404 25003 11444 25012
rect 11500 25012 11596 25052
rect 10886 24212 11254 24221
rect 10886 24163 11254 24172
rect 11308 23792 11348 24760
rect 11308 23743 11348 23752
rect 11020 23708 11060 23717
rect 11020 23573 11060 23668
rect 11500 23456 11540 25012
rect 11596 25003 11636 25012
rect 11788 24464 11828 25432
rect 11788 24415 11828 24424
rect 10732 23155 10772 23164
rect 11116 23288 11156 23297
rect 11116 23204 11156 23248
rect 11116 23153 11156 23164
rect 11404 23204 11444 23213
rect 10252 23036 10292 23045
rect 10252 22448 10292 22996
rect 10348 22448 10388 23080
rect 10540 23036 10580 23045
rect 10444 22784 10484 22793
rect 10444 22649 10484 22744
rect 10444 22448 10484 22457
rect 10348 22408 10444 22448
rect 10252 22399 10292 22408
rect 10444 22399 10484 22408
rect 10156 22196 10196 22240
rect 10156 22145 10196 22156
rect 10444 22196 10484 22205
rect 10060 22112 10100 22121
rect 10060 21977 10100 22072
rect 10252 22112 10292 22121
rect 9964 21811 10004 21820
rect 10156 21692 10196 21701
rect 10156 21524 10196 21652
rect 10156 21475 10196 21484
rect 10252 21440 10292 22072
rect 10348 22028 10388 22037
rect 10348 21893 10388 21988
rect 10444 21776 10484 22156
rect 10444 21727 10484 21736
rect 10060 21356 10100 21365
rect 9868 20971 9908 20980
rect 9964 21272 10004 21281
rect 9964 20180 10004 21232
rect 10060 21188 10100 21316
rect 10060 21139 10100 21148
rect 10252 20516 10292 21400
rect 10252 20467 10292 20476
rect 10348 21608 10388 21617
rect 10348 20180 10388 21568
rect 9772 20131 9812 20140
rect 9868 20140 10004 20180
rect 10156 20140 10388 20180
rect 10444 21524 10484 21533
rect 9772 19256 9812 19265
rect 9580 19216 9772 19256
rect 9676 18668 9716 18677
rect 9580 18500 9620 18509
rect 9580 18164 9620 18460
rect 9580 18115 9620 18124
rect 9484 18031 9524 18040
rect 9676 17912 9716 18628
rect 9772 17996 9812 19216
rect 9772 17947 9812 17956
rect 9676 17863 9716 17872
rect 9388 17620 9620 17660
rect 9388 17240 9428 17249
rect 9388 16904 9428 17200
rect 9484 17156 9524 17165
rect 9484 17021 9524 17116
rect 9388 16864 9524 16904
rect 9484 16400 9524 16864
rect 9388 16316 9428 16327
rect 9388 16232 9428 16276
rect 9484 16316 9524 16360
rect 9484 16265 9524 16276
rect 9388 16183 9428 16192
rect 9484 16064 9524 16073
rect 9292 16024 9484 16064
rect 9484 16015 9524 16024
rect 9292 15896 9332 15907
rect 9292 15812 9332 15856
rect 9292 15763 9332 15772
rect 9580 15644 9620 17620
rect 9676 17492 9716 17501
rect 9676 16484 9716 17452
rect 9868 16904 9908 20140
rect 10156 19676 10196 20140
rect 10156 19627 10196 19636
rect 10156 19256 10196 19265
rect 9868 16855 9908 16864
rect 9964 19088 10004 19097
rect 9964 16988 10004 19048
rect 10156 19004 10196 19216
rect 10196 18964 10292 19004
rect 10156 18955 10196 18964
rect 10156 18584 10196 18593
rect 9676 16435 9716 16444
rect 9868 16736 9908 16745
rect 9196 15604 9428 15644
rect 9100 15427 9140 15436
rect 9196 15476 9236 15485
rect 9004 14503 9044 14512
rect 9196 14384 9236 15436
rect 9196 14132 9236 14344
rect 9196 14083 9236 14092
rect 9292 15056 9332 15065
rect 9196 13796 9236 13805
rect 8908 12319 8948 12328
rect 9004 13628 9044 13637
rect 8908 11780 8948 11789
rect 9004 11780 9044 13588
rect 9100 13544 9140 13553
rect 9100 13040 9140 13504
rect 9196 13292 9236 13756
rect 9196 13243 9236 13252
rect 9100 12991 9140 13000
rect 9196 13124 9236 13133
rect 9196 12620 9236 13084
rect 9196 12536 9236 12580
rect 9196 12456 9236 12496
rect 8948 11740 9044 11780
rect 9100 12116 9140 12125
rect 8908 11696 8948 11740
rect 8908 11645 8948 11656
rect 8812 11143 8852 11152
rect 9100 11528 9140 12076
rect 9196 11612 9236 11621
rect 9292 11612 9332 15016
rect 9388 14720 9428 15604
rect 9580 15595 9620 15604
rect 9676 16148 9716 16157
rect 9388 14671 9428 14680
rect 9484 15560 9524 15569
rect 9484 14636 9524 15520
rect 9484 14587 9524 14596
rect 9580 14804 9620 14813
rect 9388 13796 9428 13805
rect 9388 13292 9428 13756
rect 9388 13243 9428 13252
rect 9484 13124 9524 13133
rect 9388 12956 9428 12965
rect 9388 12536 9428 12916
rect 9388 12487 9428 12496
rect 9484 11948 9524 13084
rect 9580 12704 9620 14764
rect 9676 14216 9716 16108
rect 9868 15644 9908 16696
rect 9964 16400 10004 16948
rect 10060 17576 10100 17585
rect 10060 17072 10100 17536
rect 10060 16568 10100 17032
rect 10060 16519 10100 16528
rect 9964 16351 10004 16360
rect 9868 14720 9908 15604
rect 9868 14671 9908 14680
rect 9964 16148 10004 16157
rect 9676 14167 9716 14176
rect 9772 14636 9812 14645
rect 9772 14216 9812 14596
rect 9772 14167 9812 14176
rect 9772 14048 9812 14057
rect 9772 13712 9812 14008
rect 9772 13663 9812 13672
rect 9964 13460 10004 16108
rect 10060 15728 10100 15737
rect 10060 15593 10100 15688
rect 10060 15476 10100 15485
rect 10060 14972 10100 15436
rect 10060 14048 10100 14932
rect 10156 14216 10196 18544
rect 10252 17912 10292 18964
rect 10348 18752 10388 18763
rect 10348 18668 10388 18712
rect 10348 18619 10388 18628
rect 10252 17863 10292 17872
rect 10252 17660 10292 17669
rect 10252 17240 10292 17620
rect 10252 17072 10292 17200
rect 10252 17023 10292 17032
rect 10348 17576 10388 17585
rect 10252 16400 10292 16409
rect 10252 16316 10292 16360
rect 10252 16265 10292 16276
rect 10252 16148 10292 16157
rect 10252 14468 10292 16108
rect 10348 15392 10388 17536
rect 10444 17156 10484 21484
rect 10540 21272 10580 22996
rect 10828 23036 10868 23045
rect 10636 22952 10676 22961
rect 10636 22532 10676 22912
rect 10828 22868 10868 22996
rect 10828 22819 10868 22828
rect 11308 23036 11348 23045
rect 10886 22700 11254 22709
rect 10886 22651 11254 22660
rect 10636 22483 10676 22492
rect 11308 22532 11348 22996
rect 11308 22483 11348 22492
rect 10540 21223 10580 21232
rect 10636 22280 10676 22289
rect 10636 21188 10676 22240
rect 10924 21776 10964 21871
rect 10924 21727 10964 21736
rect 10732 21608 10772 21617
rect 11045 21608 11085 21617
rect 10732 21473 10772 21568
rect 10924 21568 11045 21608
rect 10924 21356 10964 21568
rect 11045 21559 11085 21568
rect 11404 21440 11444 23164
rect 11500 22364 11540 23416
rect 11500 22315 11540 22324
rect 11596 23624 11636 23633
rect 11596 22280 11636 23584
rect 11692 23540 11732 23549
rect 11692 22532 11732 23500
rect 11788 23372 11828 23383
rect 11788 23288 11828 23332
rect 11788 23239 11828 23248
rect 11884 23204 11924 23213
rect 11788 23036 11828 23131
rect 11788 22987 11828 22996
rect 11692 22483 11732 22492
rect 11788 22784 11828 22793
rect 11596 22231 11636 22240
rect 11788 21692 11828 22744
rect 11788 21643 11828 21652
rect 11404 21391 11444 21400
rect 11596 21608 11636 21617
rect 11596 21440 11636 21568
rect 11884 21608 11924 23164
rect 11980 22280 12020 26776
rect 12172 26816 12212 26860
rect 12172 26767 12212 26776
rect 12556 26816 12596 26825
rect 12460 26648 12500 26743
rect 12460 26599 12500 26608
rect 12126 26480 12494 26489
rect 12126 26431 12494 26440
rect 12460 26144 12500 26155
rect 12460 26060 12500 26104
rect 12460 26011 12500 26020
rect 12460 25388 12500 25397
rect 12172 25304 12212 25313
rect 12172 25220 12212 25264
rect 12172 25169 12212 25180
rect 12460 25220 12500 25348
rect 12556 25388 12596 26776
rect 12652 26732 12692 26741
rect 12652 26396 12692 26692
rect 12940 26648 12980 27700
rect 12940 26599 12980 26608
rect 12844 26564 12884 26573
rect 12844 26429 12884 26524
rect 12652 26347 12692 26356
rect 12844 26228 12884 26237
rect 12556 25339 12596 25348
rect 12652 25892 12692 25901
rect 12460 25171 12500 25180
rect 12126 24968 12494 24977
rect 12126 24919 12494 24928
rect 12556 24464 12596 24473
rect 12172 24380 12212 24389
rect 12172 23792 12212 24340
rect 12172 23657 12212 23752
rect 12556 23792 12596 24424
rect 12652 23792 12692 25852
rect 12748 25220 12788 25229
rect 12748 23960 12788 25180
rect 12844 25136 12884 26188
rect 13036 25388 13076 28120
rect 13132 26480 13172 28600
rect 13900 28496 13940 28600
rect 13900 28447 13940 28456
rect 14092 27992 14132 28001
rect 13516 27152 13556 27161
rect 13324 26984 13364 27079
rect 13324 26935 13364 26944
rect 13420 27068 13460 27077
rect 13420 26900 13460 27028
rect 13420 26851 13460 26860
rect 13132 26431 13172 26440
rect 13324 26816 13364 26825
rect 12844 25087 12884 25096
rect 12940 25348 13076 25388
rect 13132 26228 13172 26237
rect 12748 23911 12788 23920
rect 12844 24380 12884 24389
rect 12652 23752 12788 23792
rect 12556 23743 12596 23752
rect 12126 23456 12494 23465
rect 12126 23407 12494 23416
rect 12556 23372 12596 23381
rect 12076 23120 12116 23129
rect 12076 23036 12116 23080
rect 12076 22985 12116 22996
rect 12268 23036 12308 23045
rect 12172 22784 12212 22793
rect 12172 22649 12212 22744
rect 12268 22448 12308 22996
rect 12268 22399 12308 22408
rect 12364 22868 12404 22877
rect 11980 21692 12020 22240
rect 12364 22112 12404 22828
rect 12364 22063 12404 22072
rect 12126 21944 12494 21953
rect 12126 21895 12494 21904
rect 11980 21643 12020 21652
rect 11884 21524 11924 21568
rect 11884 21444 11924 21484
rect 10636 21139 10676 21148
rect 10732 21316 10964 21356
rect 10732 19508 10772 21316
rect 10886 21188 11254 21197
rect 10886 21139 11254 21148
rect 11596 21104 11636 21400
rect 11596 21055 11636 21064
rect 11884 21020 11924 21029
rect 11788 20768 11828 20777
rect 11404 20600 11444 20609
rect 11404 20348 11444 20560
rect 10886 19676 11254 19685
rect 10886 19627 11254 19636
rect 11404 19508 11444 20308
rect 11788 20264 11828 20728
rect 11884 20684 11924 20980
rect 11884 20635 11924 20644
rect 12556 20768 12596 23332
rect 12748 22280 12788 23752
rect 12844 23540 12884 24340
rect 12844 23120 12884 23500
rect 12844 23071 12884 23080
rect 12940 22280 12980 25348
rect 13036 25220 13076 25229
rect 13036 24464 13076 25180
rect 13132 24548 13172 26188
rect 13324 26228 13364 26776
rect 13516 26732 13556 27112
rect 13516 26597 13556 26692
rect 13708 26816 13748 26825
rect 13708 26648 13748 26776
rect 13708 26599 13748 26608
rect 13804 26816 13844 26825
rect 13804 26648 13844 26776
rect 13996 26732 14036 26741
rect 13804 26599 13844 26608
rect 13900 26648 13940 26657
rect 13324 26179 13364 26188
rect 13516 26228 13556 26237
rect 13420 26144 13460 26153
rect 13324 25388 13364 25397
rect 13132 24499 13172 24508
rect 13228 25304 13268 25313
rect 13036 24415 13076 24424
rect 13228 24044 13268 25264
rect 13324 24716 13364 25348
rect 13420 25220 13460 26104
rect 13420 25171 13460 25180
rect 13516 25304 13556 26188
rect 13900 26228 13940 26608
rect 13900 26179 13940 26188
rect 13804 26144 13844 26153
rect 13804 25976 13844 26104
rect 13804 25388 13844 25936
rect 13804 25339 13844 25348
rect 13324 24667 13364 24676
rect 13516 24716 13556 25264
rect 13516 24581 13556 24676
rect 13708 25220 13748 25229
rect 13612 24548 13652 24557
rect 13516 24464 13556 24473
rect 13228 23995 13268 24004
rect 13324 24212 13364 24221
rect 13132 23876 13172 23885
rect 13132 23288 13172 23836
rect 13324 23708 13364 24172
rect 13324 23659 13364 23668
rect 13420 23960 13460 23969
rect 13132 23239 13172 23248
rect 13228 23624 13268 23633
rect 12748 22240 12884 22280
rect 12652 22112 12692 22121
rect 12652 21608 12692 22072
rect 12748 22112 12788 22121
rect 12748 22028 12788 22072
rect 12748 21977 12788 21988
rect 12652 21473 12692 21568
rect 11500 20180 11540 20189
rect 11500 19676 11540 20140
rect 11500 19627 11540 19636
rect 11692 19760 11732 19769
rect 11404 19468 11540 19508
rect 10732 19459 10772 19468
rect 10636 19340 10676 19349
rect 10540 18668 10580 18677
rect 10540 17996 10580 18628
rect 10540 17947 10580 17956
rect 10636 18332 10676 19300
rect 11308 19256 11348 19265
rect 10444 17107 10484 17116
rect 10540 17828 10580 17837
rect 10540 17240 10580 17788
rect 10636 17744 10676 18292
rect 10732 19172 10772 19181
rect 10732 17828 10772 19132
rect 11308 18752 11348 19216
rect 11308 18703 11348 18712
rect 11404 18584 11444 18593
rect 11308 18500 11348 18509
rect 10886 18164 11254 18173
rect 10886 18115 11254 18124
rect 11020 17996 11060 18005
rect 11212 17996 11252 18005
rect 10732 17779 10772 17788
rect 10828 17912 10868 17921
rect 10636 17695 10676 17704
rect 10540 17105 10580 17200
rect 10636 17576 10676 17585
rect 10540 16988 10580 16997
rect 10444 16820 10484 16829
rect 10444 16064 10484 16780
rect 10540 16316 10580 16948
rect 10636 16736 10676 17536
rect 10828 16988 10868 17872
rect 11020 17744 11060 17956
rect 11020 17324 11060 17704
rect 11020 17275 11060 17284
rect 11116 17956 11212 17996
rect 11116 17072 11156 17956
rect 11212 17947 11252 17956
rect 11116 17023 11156 17032
rect 11308 17660 11348 18460
rect 11404 18449 11444 18544
rect 11500 18164 11540 19468
rect 11500 18115 11540 18124
rect 11596 19172 11636 19181
rect 10828 16939 10868 16948
rect 10636 16687 10676 16696
rect 10886 16652 11254 16661
rect 10886 16603 11254 16612
rect 11308 16316 11348 17620
rect 11404 18080 11444 18089
rect 11404 17996 11444 18040
rect 11404 17156 11444 17956
rect 11404 17107 11444 17116
rect 11500 17912 11540 17921
rect 11500 17072 11540 17872
rect 11596 17660 11636 19132
rect 11596 17525 11636 17620
rect 11500 17023 11540 17032
rect 10540 16276 10676 16316
rect 10444 16015 10484 16024
rect 10636 15476 10676 16276
rect 11308 16267 11348 16276
rect 11404 16820 11444 16829
rect 10924 16232 10964 16241
rect 10828 16148 10868 16157
rect 10636 15427 10676 15436
rect 10732 15560 10772 15569
rect 10348 15343 10388 15352
rect 10252 14419 10292 14428
rect 10444 15308 10484 15317
rect 10156 14167 10196 14176
rect 10060 13999 10100 14008
rect 10348 14132 10388 14141
rect 10252 13964 10292 13973
rect 10252 13880 10292 13924
rect 10060 13712 10100 13807
rect 10060 13663 10100 13672
rect 9964 13411 10004 13420
rect 9580 12655 9620 12664
rect 9772 13208 9812 13217
rect 9484 11899 9524 11908
rect 9676 12452 9716 12461
rect 9236 11572 9332 11612
rect 9196 11563 9236 11572
rect 8908 11024 8948 11033
rect 8908 10436 8948 10984
rect 8908 10268 8948 10396
rect 8908 10219 8948 10228
rect 8812 10184 8852 10193
rect 8812 9764 8852 10144
rect 8812 9715 8852 9724
rect 9004 10184 9044 10193
rect 9004 9680 9044 10144
rect 9004 9631 9044 9640
rect 9100 9512 9140 11488
rect 9580 11024 9620 11033
rect 9580 10604 9620 10984
rect 9100 9344 9140 9472
rect 9388 10100 9428 10109
rect 9388 9512 9428 10060
rect 9388 9463 9428 9472
rect 9100 8840 9140 9304
rect 9100 8791 9140 8800
rect 9388 9344 9428 9353
rect 9388 8588 9428 9304
rect 9580 9008 9620 10564
rect 9580 8959 9620 8968
rect 9676 8756 9716 12412
rect 9772 9596 9812 13168
rect 9964 13124 10004 13133
rect 9868 13040 9908 13049
rect 9868 12452 9908 13000
rect 9964 12704 10004 13084
rect 9964 12655 10004 12664
rect 10156 12620 10196 12629
rect 9868 12200 9908 12412
rect 9964 12536 10004 12545
rect 9964 12452 10004 12496
rect 9964 12401 10004 12412
rect 9868 12151 9908 12160
rect 9964 12284 10004 12293
rect 9964 12032 10004 12244
rect 9964 11983 10004 11992
rect 10060 11948 10100 11957
rect 10060 11864 10100 11908
rect 9868 11824 10100 11864
rect 9868 11780 9908 11824
rect 9868 11731 9908 11740
rect 9964 11717 10004 11726
rect 9964 11276 10004 11677
rect 10156 11528 10196 12580
rect 10252 11864 10292 13840
rect 10348 13250 10388 14092
rect 10444 14048 10484 15268
rect 10636 15308 10676 15317
rect 10636 14804 10676 15268
rect 10636 14755 10676 14764
rect 10732 15056 10772 15520
rect 10828 15308 10868 16108
rect 10924 15812 10964 16192
rect 11308 16148 11348 16157
rect 11404 16148 11444 16780
rect 11348 16108 11444 16148
rect 11500 16148 11540 16157
rect 11308 16099 11348 16108
rect 11404 15896 11444 15905
rect 10924 15763 10964 15772
rect 11020 15812 11060 15821
rect 11020 15560 11060 15772
rect 11404 15761 11444 15856
rect 11020 15511 11060 15520
rect 11404 15560 11444 15571
rect 11116 15476 11156 15485
rect 11116 15341 11156 15436
rect 11404 15476 11444 15520
rect 11404 15427 11444 15436
rect 10828 15259 10868 15268
rect 10886 15140 11254 15149
rect 10886 15091 11254 15100
rect 10540 14636 10580 14645
rect 10540 14501 10580 14596
rect 10732 14636 10772 15016
rect 11116 14972 11156 14981
rect 10732 14587 10772 14596
rect 10924 14720 10964 14729
rect 10924 14585 10964 14680
rect 10636 14468 10676 14477
rect 10444 13999 10484 14008
rect 10540 14216 10580 14225
rect 10540 13964 10580 14176
rect 10540 13915 10580 13924
rect 10348 13201 10388 13210
rect 10444 13040 10484 13049
rect 10252 11815 10292 11824
rect 10348 12368 10388 12377
rect 10348 11864 10388 12328
rect 10348 11815 10388 11824
rect 10156 11479 10196 11488
rect 10252 11696 10292 11705
rect 9964 11227 10004 11236
rect 10252 11192 10292 11656
rect 10252 11143 10292 11152
rect 10348 11612 10388 11621
rect 9868 11108 9908 11117
rect 9868 10184 9908 11068
rect 10156 11108 10196 11117
rect 10156 10436 10196 11068
rect 10156 10387 10196 10396
rect 9868 10135 9908 10144
rect 10156 10016 10196 10025
rect 9772 9556 10004 9596
rect 9676 8707 9716 8716
rect 9772 9428 9812 9437
rect 9484 8672 9524 8681
rect 9524 8632 9620 8672
rect 9484 8623 9524 8632
rect 9388 8539 9428 8548
rect 9196 8504 9236 8513
rect 9100 8168 9140 8177
rect 8812 8000 8852 8009
rect 8716 7960 8812 8000
rect 8620 7748 8660 7757
rect 8620 7160 8660 7708
rect 8620 7111 8660 7120
rect 8524 5480 8564 6448
rect 7948 4136 7988 4432
rect 8044 4892 8084 4901
rect 8044 4388 8084 4852
rect 8044 4339 8084 4348
rect 8524 4220 8564 5440
rect 8524 4171 8564 4180
rect 8716 4640 8756 7960
rect 8812 7951 8852 7960
rect 9100 7160 9140 8128
rect 9196 7916 9236 8464
rect 9196 7412 9236 7876
rect 9388 8420 9428 8429
rect 9388 7496 9428 8380
rect 9580 8000 9620 8632
rect 9676 8588 9716 8597
rect 9676 8420 9716 8548
rect 9676 8168 9716 8380
rect 9676 8119 9716 8128
rect 9580 7832 9620 7960
rect 9388 7447 9428 7456
rect 9484 7748 9524 7757
rect 9196 7363 9236 7372
rect 9100 7111 9140 7120
rect 9388 7328 9428 7337
rect 9292 6572 9332 6581
rect 9292 6068 9332 6532
rect 9292 6019 9332 6028
rect 9388 6236 9428 7288
rect 9484 7244 9524 7708
rect 9484 7195 9524 7204
rect 9004 5816 9044 5825
rect 9004 4892 9044 5776
rect 9388 5648 9428 6196
rect 9388 5599 9428 5608
rect 9484 6656 9524 6665
rect 9484 6404 9524 6616
rect 9484 5564 9524 6364
rect 9484 5515 9524 5524
rect 9004 4843 9044 4852
rect 9580 4724 9620 7792
rect 9676 7664 9716 7673
rect 9676 6488 9716 7624
rect 9676 6439 9716 6448
rect 9772 7244 9812 9388
rect 9868 8672 9908 8681
rect 9868 8252 9908 8632
rect 9868 8203 9908 8212
rect 9772 6320 9812 7204
rect 9868 6740 9908 6749
rect 9964 6740 10004 9556
rect 10156 7916 10196 9976
rect 10348 9512 10388 11572
rect 10444 9680 10484 13000
rect 10444 9631 10484 9640
rect 10540 11864 10580 11873
rect 10348 9463 10388 9472
rect 10540 9008 10580 11824
rect 10636 11612 10676 14428
rect 10924 14300 10964 14309
rect 10732 13964 10772 13973
rect 10732 12704 10772 13924
rect 10924 13796 10964 14260
rect 11020 14132 11060 14227
rect 11020 14083 11060 14092
rect 11116 14048 11156 14932
rect 11500 14888 11540 16108
rect 11500 14839 11540 14848
rect 11596 15896 11636 15905
rect 11308 14048 11348 14057
rect 11116 14008 11308 14048
rect 11348 14008 11444 14048
rect 11308 13999 11348 14008
rect 11020 13964 11060 13975
rect 11020 13880 11060 13924
rect 11020 13831 11060 13840
rect 11308 13880 11348 13889
rect 10924 13747 10964 13756
rect 10886 13628 11254 13637
rect 10886 13579 11254 13588
rect 10732 12655 10772 12664
rect 10828 13208 10868 13217
rect 10828 12284 10868 13168
rect 10924 13124 10964 13133
rect 10924 12536 10964 13084
rect 10924 12487 10964 12496
rect 11116 12620 11156 12629
rect 11116 12536 11156 12580
rect 11116 12485 11156 12496
rect 10636 11563 10676 11572
rect 10732 12244 10868 12284
rect 11308 12284 11348 13840
rect 11404 13712 11444 14008
rect 11404 13663 11444 13672
rect 11500 13292 11540 13301
rect 11404 13208 11444 13217
rect 11404 13073 11444 13168
rect 11404 12872 11444 12881
rect 11404 12620 11444 12832
rect 11404 12571 11444 12580
rect 10732 11528 10772 12244
rect 11308 12235 11348 12244
rect 11404 12452 11444 12461
rect 10886 12116 11254 12125
rect 10886 12067 11254 12076
rect 11308 11864 11348 11873
rect 11212 11696 11252 11705
rect 10732 11479 10772 11488
rect 10924 11528 10964 11537
rect 10924 11192 10964 11488
rect 10924 11143 10964 11152
rect 11212 11024 11252 11656
rect 11308 11696 11348 11824
rect 11308 11647 11348 11656
rect 11252 10984 11348 11024
rect 11212 10975 11252 10984
rect 10886 10604 11254 10613
rect 10886 10555 11254 10564
rect 10828 10268 10868 10277
rect 10828 10016 10868 10228
rect 11308 10184 11348 10984
rect 11308 10135 11348 10144
rect 10828 9967 10868 9976
rect 11308 9512 11348 9521
rect 10444 8968 10580 9008
rect 10732 9428 10772 9437
rect 10444 8840 10484 8968
rect 10444 8672 10484 8800
rect 10444 8623 10484 8632
rect 10636 8924 10676 8933
rect 10156 7867 10196 7876
rect 10252 8000 10292 8009
rect 10060 7748 10100 7757
rect 10060 7613 10100 7708
rect 10252 7412 10292 7960
rect 10252 7363 10292 7372
rect 10636 8000 10676 8884
rect 10732 8504 10772 9388
rect 10886 9092 11254 9101
rect 10886 9043 11254 9052
rect 10828 8840 10868 8849
rect 10828 8705 10868 8800
rect 11308 8756 11348 9472
rect 11308 8707 11348 8716
rect 10732 8455 10772 8464
rect 11212 8588 11252 8597
rect 9908 6700 10004 6740
rect 10444 6992 10484 7001
rect 9868 6691 9908 6700
rect 9772 5648 9812 6280
rect 9964 6488 10004 6497
rect 9964 6236 10004 6448
rect 10444 6488 10484 6952
rect 10444 6439 10484 6448
rect 10636 6404 10676 7960
rect 11212 8084 11252 8548
rect 11404 8168 11444 12412
rect 11500 12368 11540 13252
rect 11500 12200 11540 12328
rect 11500 12151 11540 12160
rect 11596 11948 11636 15856
rect 11692 15308 11732 19720
rect 11788 19256 11828 20224
rect 11788 19207 11828 19216
rect 11884 20432 11924 20441
rect 11884 18920 11924 20392
rect 12126 20432 12494 20441
rect 12126 20383 12494 20392
rect 12556 20264 12596 20728
rect 12556 20215 12596 20224
rect 12844 20768 12884 22240
rect 12940 22231 12980 22240
rect 13036 22868 13076 22877
rect 13036 21944 13076 22828
rect 12940 21904 13076 21944
rect 12940 21776 12980 21904
rect 12940 21727 12980 21736
rect 13228 21524 13268 23584
rect 13324 22868 13364 22877
rect 13324 22733 13364 22828
rect 13132 21484 13268 21524
rect 12844 20264 12884 20728
rect 12940 21188 12980 21197
rect 12940 20684 12980 21148
rect 13132 20768 13172 21484
rect 13132 20719 13172 20728
rect 13228 21356 13268 21365
rect 12940 20635 12980 20644
rect 12844 20096 12884 20224
rect 12844 20047 12884 20056
rect 13132 20264 13172 20273
rect 12748 20012 12788 20021
rect 12652 19424 12692 19433
rect 12556 19256 12596 19265
rect 11788 18880 11924 18920
rect 11980 19088 12020 19097
rect 11788 15896 11828 18880
rect 11884 18752 11924 18761
rect 11884 17660 11924 18712
rect 11884 17240 11924 17620
rect 11884 17191 11924 17200
rect 11884 17072 11924 17081
rect 11884 16937 11924 17032
rect 11980 16568 12020 19048
rect 12126 18920 12494 18929
rect 12126 18871 12494 18880
rect 12556 18752 12596 19216
rect 12652 19004 12692 19384
rect 12652 18955 12692 18964
rect 12748 19340 12788 19972
rect 13036 19844 13076 19853
rect 12556 18703 12596 18712
rect 12460 18584 12500 18593
rect 12748 18584 12788 19300
rect 12940 19424 12980 19433
rect 12940 18836 12980 19384
rect 12940 18787 12980 18796
rect 12500 18544 12788 18584
rect 12460 18535 12500 18544
rect 12172 18500 12212 18509
rect 12172 17996 12212 18460
rect 12652 18416 12692 18425
rect 12652 18332 12692 18376
rect 12652 18281 12692 18292
rect 12460 18164 12500 18173
rect 12172 17947 12212 17956
rect 12364 18080 12404 18091
rect 12364 17996 12404 18040
rect 12364 17947 12404 17956
rect 12460 17660 12500 18124
rect 12460 17611 12500 17620
rect 12556 17996 12596 18005
rect 12126 17408 12494 17417
rect 12126 17359 12494 17368
rect 12172 17240 12212 17249
rect 12172 17072 12212 17200
rect 12172 17023 12212 17032
rect 12460 17240 12500 17249
rect 11980 15896 12020 16528
rect 12076 16232 12116 16241
rect 12076 16097 12116 16192
rect 12460 16148 12500 17200
rect 12460 16099 12500 16108
rect 11788 15856 11924 15896
rect 11692 15259 11732 15268
rect 11788 15728 11828 15737
rect 11884 15728 11924 15856
rect 11980 15847 12020 15856
rect 12126 15896 12494 15905
rect 12126 15847 12494 15856
rect 12172 15728 12212 15737
rect 11884 15688 12116 15728
rect 11788 14972 11828 15688
rect 11884 15560 11924 15569
rect 11884 15392 11924 15520
rect 11884 15308 11924 15352
rect 11884 15257 11924 15268
rect 11788 14923 11828 14932
rect 12076 14972 12116 15688
rect 12172 15476 12212 15688
rect 12172 15427 12212 15436
rect 12364 15644 12404 15653
rect 12364 15392 12404 15604
rect 12268 15224 12308 15233
rect 12268 15089 12308 15184
rect 12076 14923 12116 14932
rect 11980 14888 12020 14897
rect 11788 14552 11828 14561
rect 11692 14048 11732 14057
rect 11692 12704 11732 14008
rect 11788 13880 11828 14512
rect 11788 13831 11828 13840
rect 11884 14384 11924 14395
rect 11884 14300 11924 14344
rect 11692 12655 11732 12664
rect 11788 13040 11828 13049
rect 11596 11899 11636 11908
rect 11788 12620 11828 13000
rect 11788 11780 11828 12580
rect 11884 11864 11924 14260
rect 11980 14048 12020 14848
rect 12172 14888 12212 14897
rect 12172 14552 12212 14848
rect 12364 14636 12404 15352
rect 12460 15644 12500 15653
rect 12460 14720 12500 15604
rect 12460 14671 12500 14680
rect 12364 14587 12404 14596
rect 12172 14503 12212 14512
rect 12126 14384 12494 14393
rect 12126 14335 12494 14344
rect 12268 14216 12308 14227
rect 12268 14132 12308 14176
rect 12268 14083 12308 14092
rect 11980 13999 12020 14008
rect 12076 14048 12116 14057
rect 12076 13964 12116 14008
rect 12076 13913 12116 13924
rect 12364 14048 12404 14057
rect 11980 13124 12020 13133
rect 11980 12284 12020 13084
rect 12364 13040 12404 14008
rect 12556 13208 12596 17956
rect 12652 17576 12692 17585
rect 12652 17072 12692 17536
rect 12652 17023 12692 17032
rect 12748 16904 12788 18544
rect 12844 18584 12884 18593
rect 12844 18449 12884 18544
rect 12940 18248 12980 18257
rect 12844 17576 12884 17585
rect 12844 17408 12884 17536
rect 12844 17359 12884 17368
rect 12652 16864 12788 16904
rect 12844 17240 12884 17249
rect 12940 17240 12980 18208
rect 13036 17660 13076 19804
rect 13132 19256 13172 20224
rect 13228 19340 13268 21316
rect 13228 19291 13268 19300
rect 13324 19928 13364 19937
rect 13132 17912 13172 19216
rect 13132 17863 13172 17872
rect 13228 17828 13268 17837
rect 13036 17620 13172 17660
rect 13132 17576 13172 17620
rect 13132 17527 13172 17536
rect 13036 17240 13076 17249
rect 12940 17200 13036 17240
rect 12652 13292 12692 16864
rect 12748 16736 12788 16745
rect 12748 16316 12788 16696
rect 12748 16148 12788 16276
rect 12748 16099 12788 16108
rect 12748 15980 12788 15989
rect 12748 15812 12788 15940
rect 12748 15560 12788 15772
rect 12748 15511 12788 15520
rect 12844 15392 12884 17200
rect 13036 17105 13076 17200
rect 13228 17240 13268 17788
rect 13228 17191 13268 17200
rect 13324 17156 13364 19888
rect 13420 19928 13460 23920
rect 13516 23204 13556 24424
rect 13612 23624 13652 24508
rect 13612 23575 13652 23584
rect 13708 23624 13748 25180
rect 13900 24800 13940 24809
rect 13900 24665 13940 24760
rect 13996 24716 14036 26692
rect 13996 24667 14036 24676
rect 13708 23575 13748 23584
rect 13996 24380 14036 24389
rect 13516 23155 13556 23164
rect 13804 23372 13844 23381
rect 13804 23204 13844 23332
rect 13804 23155 13844 23164
rect 13996 23204 14036 24340
rect 13996 23155 14036 23164
rect 14092 23060 14132 27952
rect 14188 27572 14228 27581
rect 14188 25472 14228 27532
rect 14188 25423 14228 25432
rect 14284 26480 14324 26489
rect 14668 26480 14708 28600
rect 15340 27656 15380 27665
rect 15052 27572 15092 27581
rect 14860 27488 14900 27497
rect 14188 24632 14228 24641
rect 14188 24212 14228 24592
rect 14188 24163 14228 24172
rect 14188 23876 14228 23885
rect 14188 23741 14228 23836
rect 13612 23036 13652 23045
rect 13612 21860 13652 22996
rect 13996 23020 14132 23060
rect 14188 23120 14228 23129
rect 13996 22952 14036 23020
rect 13996 22903 14036 22912
rect 14188 22952 14228 23080
rect 14092 22868 14132 22877
rect 13708 22280 13748 22289
rect 13708 22112 13748 22240
rect 13996 22280 14036 22289
rect 13708 22063 13748 22072
rect 13804 22196 13844 22205
rect 13516 21608 13556 21617
rect 13516 21188 13556 21568
rect 13612 21524 13652 21820
rect 13612 21475 13652 21484
rect 13708 21776 13748 21785
rect 13516 21139 13556 21148
rect 13612 20684 13652 20693
rect 13516 19928 13556 19956
rect 13420 19888 13516 19928
rect 13420 19508 13460 19888
rect 13516 19879 13556 19888
rect 13420 19459 13460 19468
rect 13516 19004 13556 19013
rect 13516 18248 13556 18964
rect 13228 17072 13268 17081
rect 13036 16988 13076 16997
rect 12940 15644 12980 15655
rect 12940 15560 12980 15604
rect 12940 15511 12980 15520
rect 12844 15352 12980 15392
rect 12748 15308 12788 15317
rect 12748 14216 12788 15268
rect 12844 15056 12884 15151
rect 12844 15007 12884 15016
rect 12844 14552 12884 14561
rect 12844 14468 12884 14512
rect 12940 14468 12980 15352
rect 13036 14636 13076 16948
rect 13132 16652 13172 16661
rect 13132 15392 13172 16612
rect 13228 16232 13268 17032
rect 13324 16316 13364 17116
rect 13324 16267 13364 16276
rect 13420 18208 13556 18248
rect 13228 16183 13268 16192
rect 13324 15728 13364 15737
rect 13132 15343 13172 15352
rect 13228 15476 13268 15485
rect 13036 14587 13076 14596
rect 13132 15140 13172 15149
rect 12940 14428 13076 14468
rect 12844 14417 12884 14428
rect 12748 14167 12788 14176
rect 12844 14300 12884 14309
rect 12844 14132 12884 14260
rect 12844 14083 12884 14092
rect 12940 14216 12980 14225
rect 12844 13964 12884 13975
rect 12844 13880 12884 13924
rect 12940 13964 12980 14176
rect 12940 13915 12980 13924
rect 12844 13831 12884 13840
rect 12652 13243 12692 13252
rect 12748 13796 12788 13805
rect 12556 13073 12596 13168
rect 12364 12991 12404 13000
rect 12126 12872 12494 12881
rect 12126 12823 12494 12832
rect 12652 12872 12692 12881
rect 12268 12620 12308 12629
rect 12172 12536 12212 12545
rect 12172 12401 12212 12496
rect 11980 12235 12020 12244
rect 11924 11824 12020 11864
rect 11884 11815 11924 11824
rect 11788 11731 11828 11740
rect 11884 11612 11924 11621
rect 11500 11528 11540 11537
rect 11500 11108 11540 11488
rect 11884 11192 11924 11572
rect 11884 11143 11924 11152
rect 11500 11059 11540 11068
rect 11980 11024 12020 11824
rect 12076 11612 12116 11707
rect 12076 11563 12116 11572
rect 12268 11528 12308 12580
rect 12652 12620 12692 12832
rect 12652 12571 12692 12580
rect 12364 12284 12404 12293
rect 12364 11696 12404 12244
rect 12364 11561 12404 11656
rect 12652 12032 12692 12041
rect 12652 11696 12692 11992
rect 12268 11479 12308 11488
rect 12126 11360 12494 11369
rect 12126 11311 12494 11320
rect 11980 10975 12020 10984
rect 12652 10940 12692 11656
rect 12748 11192 12788 13756
rect 13036 13208 13076 14428
rect 13132 14300 13172 15100
rect 13132 14251 13172 14260
rect 13228 14636 13268 15436
rect 13324 15308 13364 15688
rect 13324 15259 13364 15268
rect 13132 14048 13172 14143
rect 13132 13999 13172 14008
rect 13228 13796 13268 14596
rect 13324 14636 13364 14645
rect 13324 14552 13364 14596
rect 13324 14501 13364 14512
rect 13228 13747 13268 13756
rect 13324 14384 13364 14393
rect 13036 13159 13076 13168
rect 12844 12956 12884 12965
rect 12844 12536 12884 12916
rect 13324 12704 13364 14344
rect 13324 12655 13364 12664
rect 12940 12536 12980 12545
rect 12844 12496 12940 12536
rect 12940 12487 12980 12496
rect 13036 12452 13076 12461
rect 13036 12116 13076 12412
rect 13036 12067 13076 12076
rect 13324 12452 13364 12461
rect 13228 12032 13268 12041
rect 13228 11780 13268 11992
rect 13228 11731 13268 11740
rect 13036 11444 13076 11453
rect 12940 11360 12980 11369
rect 12748 11152 12884 11192
rect 12652 10891 12692 10900
rect 12748 11024 12788 11033
rect 12556 10772 12596 10781
rect 11980 10268 12020 10277
rect 11884 10184 11924 10193
rect 11884 9512 11924 10144
rect 11980 9596 12020 10228
rect 12126 9848 12494 9857
rect 12126 9799 12494 9808
rect 11980 9547 12020 9556
rect 12364 9596 12404 9605
rect 12556 9596 12596 10732
rect 12748 10688 12788 10984
rect 12404 9556 12596 9596
rect 12652 10268 12692 10277
rect 12364 9547 12404 9556
rect 11884 9008 11924 9472
rect 11884 8959 11924 8968
rect 12364 9428 12404 9437
rect 12364 8756 12404 9388
rect 12364 8707 12404 8716
rect 11692 8672 11732 8681
rect 11692 8504 11732 8632
rect 12268 8672 12308 8681
rect 12268 8537 12308 8632
rect 11404 8119 11444 8128
rect 11500 8464 11692 8504
rect 11212 7916 11252 8044
rect 11212 7867 11252 7876
rect 11404 8000 11444 8009
rect 11404 7664 11444 7960
rect 11404 7615 11444 7624
rect 11500 7832 11540 8464
rect 11692 8455 11732 8464
rect 12126 8336 12494 8345
rect 12652 8336 12692 10228
rect 12748 10184 12788 10648
rect 12748 10135 12788 10144
rect 12844 8672 12884 11152
rect 12940 10268 12980 11320
rect 13036 10940 13076 11404
rect 13324 11192 13364 12412
rect 13420 11612 13460 18208
rect 13612 18164 13652 20644
rect 13708 20012 13748 21736
rect 13804 20180 13844 22156
rect 13900 21440 13940 21449
rect 13900 21020 13940 21400
rect 13900 20971 13940 20980
rect 13804 20131 13844 20140
rect 13900 20768 13940 20777
rect 13708 19172 13748 19972
rect 13900 20096 13940 20728
rect 13900 19961 13940 20056
rect 13900 19844 13940 19853
rect 13900 19256 13940 19804
rect 13900 19207 13940 19216
rect 13708 19123 13748 19132
rect 13900 19088 13940 19097
rect 13900 18920 13940 19048
rect 13516 18124 13652 18164
rect 13708 18752 13748 18761
rect 13708 18584 13748 18712
rect 13516 17324 13556 18124
rect 13708 17744 13748 18544
rect 13900 18500 13940 18880
rect 13900 17912 13940 18460
rect 13996 18416 14036 22240
rect 14092 22280 14132 22828
rect 14092 21440 14132 22240
rect 14188 22280 14228 22912
rect 14284 22364 14324 26440
rect 14572 26440 14708 26480
rect 14764 27320 14804 27329
rect 14476 26060 14516 26069
rect 14380 25136 14420 25145
rect 14380 23288 14420 25096
rect 14476 24548 14516 26020
rect 14476 24499 14516 24508
rect 14380 23239 14420 23248
rect 14572 23060 14612 26440
rect 14668 26312 14708 26321
rect 14668 25388 14708 26272
rect 14764 25388 14804 27280
rect 14860 26060 14900 27448
rect 14956 27320 14996 27329
rect 14956 26984 14996 27280
rect 15052 27152 15092 27532
rect 15052 27103 15092 27112
rect 14956 26935 14996 26944
rect 14860 26011 14900 26020
rect 15052 26732 15092 26741
rect 14764 25348 14900 25388
rect 14668 25339 14708 25348
rect 14860 25304 14900 25348
rect 14764 25136 14804 25145
rect 14668 24884 14708 24893
rect 14668 24044 14708 24844
rect 14764 24716 14804 25096
rect 14764 24667 14804 24676
rect 14860 24632 14900 25264
rect 14956 24632 14996 24641
rect 14860 24592 14956 24632
rect 14956 24583 14996 24592
rect 15052 24464 15092 26692
rect 15340 26144 15380 27616
rect 15340 26095 15380 26104
rect 15244 25808 15284 25817
rect 14668 23708 14708 24004
rect 14668 23204 14708 23668
rect 14668 23155 14708 23164
rect 14860 24424 15092 24464
rect 15148 25304 15188 25313
rect 15148 24464 15188 25264
rect 15244 25052 15284 25768
rect 15244 25003 15284 25012
rect 15340 25136 15380 25145
rect 15340 25001 15380 25096
rect 14860 23060 14900 24424
rect 15148 24415 15188 24424
rect 15436 24380 15476 28600
rect 15628 27656 15668 27665
rect 15628 25388 15668 27616
rect 15724 27572 15764 27581
rect 15724 26984 15764 27532
rect 15724 26935 15764 26944
rect 15820 27404 15860 27413
rect 15628 25339 15668 25348
rect 15436 24331 15476 24340
rect 15820 24632 15860 27364
rect 16108 27404 16148 27413
rect 16108 25556 16148 27364
rect 16204 25976 16244 28600
rect 16300 26564 16340 26573
rect 16300 26312 16340 26524
rect 16300 26263 16340 26272
rect 16204 25927 16244 25936
rect 16396 25892 16436 28624
rect 23096 28600 23176 29000
rect 23864 28600 23944 29000
rect 24632 28600 24712 29000
rect 25400 28600 25480 29000
rect 26168 28600 26248 29000
rect 26936 28600 27016 29000
rect 27704 28600 27784 29000
rect 28472 28600 28552 29000
rect 29240 28600 29320 29000
rect 30008 28600 30088 29000
rect 30776 28600 30856 29000
rect 19900 27992 20268 28001
rect 19900 27943 20268 27952
rect 17068 27740 17108 27749
rect 17068 26816 17108 27700
rect 19180 27656 19220 27665
rect 19084 27488 19124 27497
rect 16108 25388 16148 25516
rect 16108 25339 16148 25348
rect 16300 25852 16436 25892
rect 16972 26228 17012 26237
rect 16204 25304 16244 25313
rect 15724 24212 15764 24221
rect 15436 24128 15476 24137
rect 15340 23792 15380 23801
rect 15244 23372 15284 23381
rect 15244 23204 15284 23332
rect 15244 23155 15284 23164
rect 14284 22315 14324 22324
rect 14380 23036 14420 23045
rect 14572 23020 14804 23060
rect 14860 23020 14996 23060
rect 14188 22231 14228 22240
rect 14380 21776 14420 22996
rect 14764 22616 14804 23020
rect 14764 22567 14804 22576
rect 14188 21608 14228 21619
rect 14188 21524 14228 21568
rect 14188 21475 14228 21484
rect 14092 21391 14132 21400
rect 14380 21272 14420 21736
rect 14476 21608 14516 21617
rect 14476 21473 14516 21568
rect 14380 21223 14420 21232
rect 14860 21272 14900 21281
rect 14860 21104 14900 21232
rect 14860 21055 14900 21064
rect 14092 21020 14132 21029
rect 14092 20852 14132 20980
rect 14092 20803 14132 20812
rect 14860 20852 14900 20861
rect 14572 20768 14612 20777
rect 14476 20516 14516 20525
rect 14476 20432 14516 20476
rect 14188 20264 14228 20273
rect 13996 18367 14036 18376
rect 14092 19256 14132 19265
rect 13900 17863 13940 17872
rect 13708 17695 13748 17704
rect 13996 17828 14036 17837
rect 13516 17275 13556 17284
rect 13900 17576 13940 17585
rect 13516 17072 13556 17081
rect 13516 16652 13556 17032
rect 13516 16603 13556 16612
rect 13612 16988 13652 16997
rect 13612 15728 13652 16948
rect 13900 16988 13940 17536
rect 13996 17156 14036 17788
rect 13996 17107 14036 17116
rect 14092 17051 14132 19216
rect 14188 18752 14228 20224
rect 14476 20180 14516 20392
rect 14476 20131 14516 20140
rect 14188 18703 14228 18712
rect 14284 20096 14324 20105
rect 14284 18920 14324 20056
rect 14380 20012 14420 20021
rect 14380 19760 14420 19972
rect 14380 19711 14420 19720
rect 14476 19844 14516 19853
rect 14476 19256 14516 19804
rect 14572 19508 14612 20728
rect 14860 20717 14900 20812
rect 14668 20684 14708 20693
rect 14668 20264 14708 20644
rect 14668 20215 14708 20224
rect 14860 20096 14900 20105
rect 14572 19459 14612 19468
rect 14668 20012 14708 20021
rect 14668 19340 14708 19972
rect 14860 19844 14900 20056
rect 14860 19795 14900 19804
rect 14668 19291 14708 19300
rect 14476 19207 14516 19216
rect 14764 19256 14804 19267
rect 14764 19172 14804 19216
rect 14284 18668 14324 18880
rect 14284 18619 14324 18628
rect 14476 19004 14516 19013
rect 14284 18500 14324 18509
rect 14188 18416 14228 18425
rect 14188 17912 14228 18376
rect 14284 17996 14324 18460
rect 14380 18416 14420 18425
rect 14380 18248 14420 18376
rect 14380 18199 14420 18208
rect 14284 17947 14324 17956
rect 14476 17996 14516 18964
rect 14764 18752 14804 19132
rect 14764 18703 14804 18712
rect 14860 19172 14900 19181
rect 14572 18584 14612 18593
rect 14572 18416 14612 18544
rect 14572 18367 14612 18376
rect 14668 18416 14708 18427
rect 14668 18332 14708 18376
rect 14668 18283 14708 18292
rect 14764 18332 14804 18341
rect 14188 17576 14228 17872
rect 14188 17527 14228 17536
rect 14380 17912 14420 17921
rect 14380 17240 14420 17872
rect 13900 16939 13940 16948
rect 13996 17011 14132 17051
rect 14284 17200 14420 17240
rect 13900 16568 13940 16577
rect 13612 15679 13652 15688
rect 13708 16232 13748 16241
rect 13516 15644 13556 15653
rect 13516 14720 13556 15604
rect 13708 15224 13748 16192
rect 13900 16232 13940 16528
rect 13900 16183 13940 16192
rect 13804 16148 13844 16157
rect 13804 15644 13844 16108
rect 13804 15595 13844 15604
rect 13804 15476 13844 15485
rect 13804 15341 13844 15436
rect 13900 15308 13940 15317
rect 13708 15184 13844 15224
rect 13516 13880 13556 14680
rect 13708 14720 13748 14729
rect 13708 14216 13748 14680
rect 13708 14167 13748 14176
rect 13804 14048 13844 15184
rect 13516 13831 13556 13840
rect 13612 13964 13652 13973
rect 13612 13829 13652 13924
rect 13516 13460 13556 13469
rect 13516 12536 13556 13420
rect 13804 12956 13844 14008
rect 13516 12032 13556 12496
rect 13516 11983 13556 11992
rect 13708 12916 13804 12956
rect 13708 11948 13748 12916
rect 13804 12907 13844 12916
rect 13900 14300 13940 15268
rect 13996 15224 14036 17011
rect 13996 15175 14036 15184
rect 14092 16820 14132 16829
rect 14092 16232 14132 16780
rect 14284 16316 14324 17200
rect 14284 16267 14324 16276
rect 14380 17072 14420 17081
rect 14092 15476 14132 16192
rect 14213 15560 14253 15569
rect 14092 14804 14132 15436
rect 14092 14755 14132 14764
rect 14188 15520 14213 15560
rect 14188 15511 14253 15520
rect 14188 15392 14228 15511
rect 13708 11899 13748 11908
rect 13804 12536 13844 12545
rect 13516 11864 13556 11873
rect 13516 11696 13556 11824
rect 13516 11647 13556 11656
rect 13708 11696 13748 11705
rect 13420 11563 13460 11572
rect 13324 11143 13364 11152
rect 13516 11528 13556 11537
rect 13516 11024 13556 11488
rect 13612 11192 13652 11203
rect 13612 11108 13652 11152
rect 13612 11059 13652 11068
rect 13516 10975 13556 10984
rect 13036 10891 13076 10900
rect 12940 10219 12980 10228
rect 13420 10184 13460 10193
rect 13036 10100 13076 10109
rect 13036 9512 13076 10060
rect 13036 9463 13076 9472
rect 13420 9512 13460 10144
rect 13708 10184 13748 11656
rect 13804 11192 13844 12496
rect 13900 12536 13940 14260
rect 14188 14468 14228 15352
rect 14284 15308 14324 15317
rect 14284 14636 14324 15268
rect 14284 14587 14324 14596
rect 14092 14132 14132 14141
rect 14092 13208 14132 14092
rect 14188 13544 14228 14428
rect 14284 14300 14324 14309
rect 14284 14048 14324 14260
rect 14284 13999 14324 14008
rect 14188 13495 14228 13504
rect 14380 13460 14420 17032
rect 14476 16904 14516 17956
rect 14668 17996 14708 18005
rect 14572 17828 14612 17837
rect 14572 17660 14612 17788
rect 14572 17611 14612 17620
rect 14668 17744 14708 17956
rect 14668 17576 14708 17704
rect 14668 17527 14708 17536
rect 14668 17408 14708 17417
rect 14668 17156 14708 17368
rect 14764 17240 14804 18292
rect 14764 17191 14804 17200
rect 14668 17107 14708 17116
rect 14476 16855 14516 16864
rect 14668 16988 14708 16997
rect 14668 16820 14708 16948
rect 14668 16771 14708 16780
rect 14476 16316 14516 16325
rect 14476 15812 14516 16276
rect 14476 15763 14516 15772
rect 14572 16232 14612 16241
rect 14476 15644 14516 15653
rect 14476 14720 14516 15604
rect 14476 14671 14516 14680
rect 14572 14468 14612 16192
rect 14764 15896 14804 15905
rect 14764 15644 14804 15856
rect 14764 15595 14804 15604
rect 14476 14428 14612 14468
rect 14764 15392 14804 15401
rect 14476 14048 14516 14428
rect 14476 13999 14516 14008
rect 14572 14132 14612 14141
rect 14572 13997 14612 14092
rect 14476 13880 14516 13889
rect 14476 13745 14516 13840
rect 14668 13880 14708 13889
rect 14668 13712 14708 13840
rect 14380 13411 14420 13420
rect 14572 13672 14708 13712
rect 14572 13376 14612 13672
rect 14572 13327 14612 13336
rect 13900 12487 13940 12496
rect 13996 12956 14036 12965
rect 13996 12536 14036 12916
rect 13996 12487 14036 12496
rect 14092 12788 14132 13168
rect 14572 13208 14612 13217
rect 14092 11864 14132 12748
rect 14284 13124 14324 13133
rect 14284 12704 14324 13084
rect 14284 12655 14324 12664
rect 14380 12956 14420 12965
rect 14380 12452 14420 12916
rect 14380 12403 14420 12412
rect 14476 12704 14516 12713
rect 14476 12536 14516 12664
rect 14572 12704 14612 13168
rect 14572 12655 14612 12664
rect 14092 11612 14132 11824
rect 14380 11864 14420 11873
rect 14476 11864 14516 12496
rect 14420 11824 14516 11864
rect 14572 12536 14612 12545
rect 14380 11815 14420 11824
rect 14092 11563 14132 11572
rect 13804 11143 13844 11152
rect 13900 11192 13940 11201
rect 13900 11108 13940 11152
rect 13900 11057 13940 11068
rect 14188 11024 14228 11033
rect 13900 10940 13940 10949
rect 13940 10900 14132 10940
rect 13900 10891 13940 10900
rect 13708 10135 13748 10144
rect 13996 10016 14036 10025
rect 13420 9463 13460 9472
rect 13708 9680 13748 9689
rect 13708 9428 13748 9640
rect 13612 9388 13708 9428
rect 13132 9008 13172 9017
rect 12844 8623 12884 8632
rect 13036 8840 13076 8849
rect 12126 8287 12494 8296
rect 12556 8296 12692 8336
rect 12844 8504 12884 8513
rect 10886 7580 11254 7589
rect 10886 7531 11254 7540
rect 11116 7160 11156 7169
rect 11116 7025 11156 7120
rect 10636 6355 10676 6364
rect 9964 6187 10004 6196
rect 10060 6152 10100 6161
rect 10060 6017 10100 6112
rect 10886 6068 11254 6077
rect 10886 6019 11254 6028
rect 9772 5599 9812 5608
rect 10444 5900 10484 5909
rect 10444 5564 10484 5860
rect 11500 5648 11540 7792
rect 11596 8084 11636 8093
rect 11596 6992 11636 8044
rect 12268 8084 12308 8093
rect 12076 8000 12116 8009
rect 11788 7916 11828 7925
rect 11596 6943 11636 6952
rect 11692 7160 11732 7169
rect 11596 6488 11636 6497
rect 11596 6353 11636 6448
rect 11500 5599 11540 5608
rect 10444 5515 10484 5524
rect 11308 5480 11348 5489
rect 11308 5312 11348 5440
rect 11308 5272 11540 5312
rect 9580 4675 9620 4684
rect 10060 4808 10100 4817
rect 7948 4087 7988 4096
rect 8716 4136 8756 4600
rect 8716 4087 8756 4096
rect 10060 4136 10100 4768
rect 10060 4087 10100 4096
rect 10348 4724 10388 4733
rect 10348 4136 10388 4684
rect 10886 4556 11254 4565
rect 10886 4507 11254 4516
rect 11500 4304 11540 5272
rect 11500 4255 11540 4264
rect 11692 4976 11732 7120
rect 11788 5480 11828 7876
rect 12076 7748 12116 7960
rect 12268 7949 12308 8044
rect 12076 7699 12116 7708
rect 11884 7160 11924 7169
rect 11884 6488 11924 7120
rect 12126 6824 12494 6833
rect 12126 6775 12494 6784
rect 11884 6439 11924 6448
rect 12172 6488 12212 6497
rect 11884 6236 11924 6245
rect 11884 5648 11924 6196
rect 11884 5599 11924 5608
rect 11788 5431 11828 5440
rect 11980 5564 12020 5573
rect 10348 4087 10388 4096
rect 11692 4136 11732 4936
rect 11980 5144 12020 5524
rect 12172 5480 12212 6448
rect 12268 6488 12308 6497
rect 12268 5648 12308 6448
rect 12268 5599 12308 5608
rect 12556 5648 12596 8296
rect 12652 8168 12692 8177
rect 12652 7160 12692 8128
rect 12844 7916 12884 8464
rect 13036 8000 13076 8800
rect 13132 8168 13172 8968
rect 13132 8000 13172 8128
rect 13324 8084 13364 8093
rect 13228 8000 13268 8009
rect 13132 7960 13228 8000
rect 13036 7951 13076 7960
rect 13228 7951 13268 7960
rect 12844 7867 12884 7876
rect 12652 6236 12692 7120
rect 13324 7160 13364 8044
rect 13420 7916 13460 7925
rect 13420 7244 13460 7876
rect 13420 7195 13460 7204
rect 13324 7111 13364 7120
rect 12652 6187 12692 6196
rect 12844 6488 12884 6497
rect 12172 5431 12212 5440
rect 12126 5312 12494 5321
rect 12126 5263 12494 5272
rect 11692 4087 11732 4096
rect 11884 4892 11924 4901
rect 11884 4136 11924 4852
rect 11980 4220 12020 5104
rect 12556 4976 12596 5608
rect 12844 5648 12884 6448
rect 13036 6488 13076 6497
rect 13036 6152 13076 6448
rect 13612 6488 13652 9388
rect 13708 9379 13748 9388
rect 13900 9512 13940 9521
rect 13900 9344 13940 9472
rect 13900 9295 13940 9304
rect 13612 6439 13652 6448
rect 13708 8672 13748 8681
rect 13708 8000 13748 8632
rect 12940 6112 13076 6152
rect 12940 5816 12980 6112
rect 12940 5767 12980 5776
rect 12844 5599 12884 5608
rect 12940 5480 12980 5489
rect 13036 5480 13076 6112
rect 12980 5440 13076 5480
rect 12940 5412 12980 5440
rect 12556 4927 12596 4936
rect 12652 5060 12692 5069
rect 12652 4925 12692 5020
rect 13228 4808 13268 4817
rect 13228 4388 13268 4768
rect 13228 4339 13268 4348
rect 13708 4304 13748 7960
rect 13996 8504 14036 9976
rect 13996 6572 14036 8464
rect 13996 6523 14036 6532
rect 14092 6236 14132 10900
rect 14188 9596 14228 10984
rect 14476 10184 14516 10193
rect 14476 9680 14516 10144
rect 14476 9631 14516 9640
rect 14188 9547 14228 9556
rect 14572 9512 14612 12496
rect 14572 9344 14612 9472
rect 14572 6740 14612 9304
rect 14764 8672 14804 15352
rect 14860 11948 14900 19132
rect 14860 11899 14900 11908
rect 14956 11864 14996 23020
rect 15148 22280 15188 22289
rect 15148 21776 15188 22240
rect 15148 21727 15188 21736
rect 15052 21608 15092 21617
rect 15052 18668 15092 21568
rect 15148 21356 15188 21365
rect 15148 20600 15188 21316
rect 15148 20551 15188 20560
rect 15244 21188 15284 21197
rect 15244 20348 15284 21148
rect 15148 20264 15188 20273
rect 15148 19508 15188 20224
rect 15244 20012 15284 20308
rect 15244 19963 15284 19972
rect 15148 19459 15188 19468
rect 15148 19340 15188 19349
rect 15148 19205 15188 19300
rect 15244 19172 15284 19181
rect 15148 19004 15188 19013
rect 15148 18920 15188 18964
rect 15148 18869 15188 18880
rect 15052 18619 15092 18628
rect 15244 18836 15284 19132
rect 15244 18584 15284 18796
rect 15244 18535 15284 18544
rect 15148 18500 15188 18509
rect 15052 17660 15092 17669
rect 15052 16400 15092 17620
rect 15148 17660 15188 18460
rect 15148 17611 15188 17620
rect 15244 18416 15284 18425
rect 15244 16484 15284 18376
rect 15244 16435 15284 16444
rect 15340 16988 15380 23752
rect 15436 23036 15476 24088
rect 15436 22987 15476 22996
rect 15724 23372 15764 24172
rect 15532 22280 15572 22289
rect 15532 21692 15572 22240
rect 15532 21524 15572 21652
rect 15436 21440 15476 21449
rect 15436 21020 15476 21400
rect 15436 20971 15476 20980
rect 15532 20852 15572 21484
rect 15436 20812 15572 20852
rect 15628 21188 15668 21197
rect 15436 19844 15476 20812
rect 15628 20768 15668 21148
rect 15628 20719 15668 20728
rect 15628 20600 15668 20609
rect 15532 20071 15572 20107
rect 15532 20012 15572 20031
rect 15532 19963 15572 19972
rect 15436 19804 15572 19844
rect 15436 19256 15476 19265
rect 15436 18752 15476 19216
rect 15436 18703 15476 18712
rect 15532 18584 15572 19804
rect 15436 18544 15572 18584
rect 15436 18248 15476 18544
rect 15628 18416 15668 20560
rect 15628 18367 15668 18376
rect 15724 18584 15764 23332
rect 15436 18199 15476 18208
rect 15532 18164 15572 18173
rect 15436 18080 15476 18091
rect 15436 17996 15476 18040
rect 15436 17947 15476 17956
rect 15436 17576 15476 17585
rect 15436 17441 15476 17536
rect 15436 17156 15476 17165
rect 15436 17021 15476 17116
rect 15052 16351 15092 16360
rect 15244 16316 15284 16325
rect 15148 16232 15188 16241
rect 15148 15644 15188 16192
rect 15244 15812 15284 16276
rect 15244 15763 15284 15772
rect 15340 15980 15380 16948
rect 15148 14972 15188 15604
rect 15244 15644 15284 15653
rect 15244 15392 15284 15604
rect 15244 15343 15284 15352
rect 15148 14923 15188 14932
rect 15052 14888 15092 14897
rect 15052 14753 15092 14848
rect 15244 14720 15284 14729
rect 15052 14636 15092 14645
rect 15052 14048 15092 14596
rect 15052 13999 15092 14008
rect 15148 13796 15188 13891
rect 15148 13747 15188 13756
rect 15244 13460 15284 14680
rect 15244 13411 15284 13420
rect 15148 13292 15188 13301
rect 15148 13157 15188 13252
rect 15244 13124 15284 13133
rect 15052 12536 15092 12545
rect 15052 12401 15092 12496
rect 15244 12368 15284 13084
rect 14956 11824 15092 11864
rect 14860 11780 14900 11789
rect 14860 11192 14900 11740
rect 14860 11143 14900 11152
rect 15052 8924 15092 11824
rect 15244 11780 15284 12328
rect 15244 11731 15284 11740
rect 15148 11612 15188 11621
rect 15148 11192 15188 11572
rect 15148 11143 15188 11152
rect 15148 10184 15188 10193
rect 15148 9680 15188 10144
rect 15148 9428 15188 9640
rect 15148 9379 15188 9388
rect 15052 8884 15284 8924
rect 14764 8084 14804 8632
rect 14764 8035 14804 8044
rect 15052 8756 15092 8765
rect 15052 8420 15092 8716
rect 14668 7748 14708 7757
rect 14668 7160 14708 7708
rect 14668 7111 14708 7120
rect 14956 7748 14996 7757
rect 14956 7076 14996 7708
rect 14956 7027 14996 7036
rect 14572 6691 14612 6700
rect 14092 6187 14132 6196
rect 14380 6572 14420 6581
rect 13708 4255 13748 4264
rect 13804 5648 13844 5657
rect 13804 4640 13844 5608
rect 14380 5480 14420 6532
rect 14476 6488 14516 6497
rect 14476 5900 14516 6448
rect 14476 5851 14516 5860
rect 15052 5900 15092 8380
rect 15052 5851 15092 5860
rect 15148 8000 15188 8009
rect 11980 4171 12020 4180
rect 13804 4220 13844 4600
rect 14284 5440 14380 5480
rect 13804 4171 13844 4180
rect 13900 4304 13940 4313
rect 11884 4087 11924 4096
rect 13900 4136 13940 4264
rect 14284 4220 14324 5440
rect 14380 5431 14420 5440
rect 14380 4892 14420 4901
rect 14380 4304 14420 4852
rect 15148 4892 15188 7960
rect 15148 4388 15188 4852
rect 15244 5732 15284 8884
rect 15244 4472 15284 5692
rect 15340 5060 15380 15940
rect 15436 16316 15476 16325
rect 15436 15476 15476 16276
rect 15436 15427 15476 15436
rect 15436 14636 15476 14645
rect 15436 14216 15476 14596
rect 15436 14167 15476 14176
rect 15532 13880 15572 18124
rect 15724 17828 15764 18544
rect 15820 18500 15860 24592
rect 16108 24884 16148 24893
rect 16012 23876 16052 23885
rect 16012 22952 16052 23836
rect 16108 23060 16148 24844
rect 16204 24800 16244 25264
rect 16204 24751 16244 24760
rect 16204 24212 16244 24221
rect 16204 23204 16244 24172
rect 16204 23155 16244 23164
rect 16108 23020 16244 23060
rect 16012 22903 16052 22912
rect 15916 22280 15956 22289
rect 15916 21356 15956 22240
rect 16108 22196 16148 22205
rect 16108 21776 16148 22156
rect 16012 21692 16052 21701
rect 16012 21557 16052 21652
rect 16108 21608 16148 21736
rect 16108 21559 16148 21568
rect 15916 21307 15956 21316
rect 15916 20936 15956 20945
rect 15916 20801 15956 20896
rect 16108 20852 16148 20861
rect 15916 20684 15956 20693
rect 15916 20264 15956 20644
rect 15916 20215 15956 20224
rect 16012 20600 16052 20609
rect 16012 20012 16052 20560
rect 15916 19844 15956 19853
rect 15916 19709 15956 19804
rect 15820 18451 15860 18460
rect 15916 19340 15956 19349
rect 15916 18164 15956 19300
rect 16012 19088 16052 19972
rect 16012 19039 16052 19048
rect 15916 18115 15956 18124
rect 15628 17660 15668 17669
rect 15628 17156 15668 17620
rect 15724 17240 15764 17788
rect 15820 17912 15860 17921
rect 15820 17744 15860 17872
rect 15820 17695 15860 17704
rect 15724 17191 15764 17200
rect 16108 17240 16148 20812
rect 16204 20012 16244 23020
rect 16204 19963 16244 19972
rect 16204 19256 16244 19265
rect 16204 19121 16244 19216
rect 16204 18836 16244 18845
rect 16204 18668 16244 18796
rect 16204 18619 16244 18628
rect 16204 18500 16244 18509
rect 16204 18365 16244 18460
rect 16300 17744 16340 25852
rect 16876 25640 16916 25649
rect 16396 24044 16436 24053
rect 16396 20768 16436 24004
rect 16684 23876 16724 23885
rect 16684 23741 16724 23836
rect 16684 23288 16724 23299
rect 16684 23204 16724 23248
rect 16876 23288 16916 25600
rect 16876 23239 16916 23248
rect 16972 24716 17012 26188
rect 16684 23155 16724 23164
rect 16876 22616 16916 22625
rect 16876 21608 16916 22576
rect 16876 21559 16916 21568
rect 16396 17912 16436 20728
rect 16684 21524 16724 21533
rect 16684 20348 16724 21484
rect 16972 21020 17012 24676
rect 17068 25304 17108 26776
rect 17548 27404 17588 27413
rect 17548 26732 17588 27364
rect 18660 27236 19028 27245
rect 18660 27187 19028 27196
rect 17548 26683 17588 26692
rect 17740 27068 17780 27077
rect 17740 26732 17780 27028
rect 17740 26683 17780 26692
rect 18316 26900 18356 26909
rect 18220 26648 18260 26657
rect 17068 24716 17108 25264
rect 17356 26564 17396 26573
rect 17068 24667 17108 24676
rect 17260 25220 17300 25229
rect 17068 24380 17108 24389
rect 17068 22280 17108 24340
rect 17260 23960 17300 25180
rect 17260 23911 17300 23920
rect 17260 23792 17300 23801
rect 17260 23204 17300 23752
rect 17260 23155 17300 23164
rect 17068 22231 17108 22240
rect 17260 21860 17300 21869
rect 16972 20971 17012 20980
rect 17164 21356 17204 21365
rect 17068 20852 17108 20861
rect 16972 20684 17012 20693
rect 16588 20264 16628 20273
rect 16492 20096 16532 20105
rect 16492 19928 16532 20056
rect 16492 19879 16532 19888
rect 16588 19844 16628 20224
rect 16684 20180 16724 20308
rect 16684 20131 16724 20140
rect 16876 20516 16916 20525
rect 16780 20012 16820 20021
rect 16588 19804 16724 19844
rect 16396 17863 16436 17872
rect 16492 19172 16532 19181
rect 16492 18332 16532 19132
rect 16588 18584 16628 18679
rect 16588 18535 16628 18544
rect 16492 17744 16532 18292
rect 16300 17695 16340 17704
rect 16396 17704 16492 17744
rect 16108 17191 16148 17200
rect 16204 17660 16244 17669
rect 15628 17107 15668 17116
rect 15724 17072 15764 17081
rect 16012 17072 16052 17081
rect 15628 16232 15668 16241
rect 15628 16097 15668 16192
rect 15628 15896 15668 15905
rect 15628 15560 15668 15856
rect 15628 15511 15668 15520
rect 15724 15560 15764 17032
rect 15916 17032 16012 17072
rect 15724 14804 15764 15520
rect 15724 14755 15764 14764
rect 15820 16988 15860 16997
rect 15724 14636 15764 14645
rect 15628 14552 15668 14561
rect 15628 14132 15668 14512
rect 15628 14083 15668 14092
rect 15724 14048 15764 14596
rect 15724 13999 15764 14008
rect 15532 13831 15572 13840
rect 15532 13544 15572 13553
rect 15436 13292 15476 13301
rect 15436 12704 15476 13252
rect 15436 12655 15476 12664
rect 15532 13124 15572 13504
rect 15628 13376 15668 13385
rect 15628 13208 15668 13336
rect 15820 13376 15860 16948
rect 15916 14216 15956 17032
rect 16012 17023 16052 17032
rect 16204 16988 16244 17620
rect 16204 16939 16244 16948
rect 16396 16904 16436 17704
rect 16492 17695 16532 17704
rect 16588 18416 16628 18425
rect 16396 16855 16436 16864
rect 16492 16988 16532 16997
rect 16204 16652 16244 16661
rect 16108 16316 16148 16325
rect 16012 15644 16052 15653
rect 16012 14888 16052 15604
rect 16108 15644 16148 16276
rect 16204 16232 16244 16612
rect 16244 16192 16340 16232
rect 16204 16183 16244 16192
rect 16108 15595 16148 15604
rect 16012 14839 16052 14848
rect 16108 14888 16148 14897
rect 15916 14167 15956 14176
rect 16012 14636 16052 14645
rect 16012 14132 16052 14596
rect 16012 14083 16052 14092
rect 15820 13327 15860 13336
rect 15916 14048 15956 14057
rect 15628 13159 15668 13168
rect 15532 12620 15572 13084
rect 15532 12571 15572 12580
rect 15628 12704 15668 12713
rect 15436 12536 15476 12545
rect 15436 12401 15476 12496
rect 15436 11864 15476 11873
rect 15436 11780 15476 11824
rect 15436 11729 15476 11740
rect 15436 11612 15476 11621
rect 15436 8756 15476 11572
rect 15628 11108 15668 12664
rect 15820 12536 15860 12545
rect 15820 12284 15860 12496
rect 15820 12235 15860 12244
rect 15820 11696 15860 11705
rect 15820 11561 15860 11656
rect 15628 11059 15668 11068
rect 15532 11024 15572 11033
rect 15532 9596 15572 10984
rect 15532 9547 15572 9556
rect 15628 10184 15668 10193
rect 15628 9680 15668 10144
rect 15628 9512 15668 9640
rect 15628 9463 15668 9472
rect 15820 10100 15860 10109
rect 15820 9344 15860 10060
rect 15916 9764 15956 14008
rect 16108 13544 16148 14848
rect 16300 14804 16340 16192
rect 16300 14755 16340 14764
rect 16396 16148 16436 16157
rect 16204 14720 16244 14729
rect 16396 14720 16436 16108
rect 16492 15476 16532 16948
rect 16492 15427 16532 15436
rect 16492 14720 16532 14815
rect 16396 14680 16492 14720
rect 16204 14585 16244 14680
rect 16492 14671 16532 14680
rect 16492 14552 16532 14561
rect 16492 14048 16532 14512
rect 16492 13999 16532 14008
rect 16396 13880 16436 13889
rect 16012 13460 16052 13469
rect 16012 11948 16052 13420
rect 16108 12032 16148 13504
rect 16204 13796 16244 13805
rect 16204 12956 16244 13756
rect 16204 12536 16244 12916
rect 16204 12487 16244 12496
rect 16300 13292 16340 13301
rect 16108 11983 16148 11992
rect 16012 11899 16052 11908
rect 16108 11864 16148 11873
rect 16108 11780 16148 11824
rect 16108 11729 16148 11740
rect 16012 11612 16052 11621
rect 16012 11192 16052 11572
rect 16012 11143 16052 11152
rect 16204 11612 16244 11621
rect 16204 10856 16244 11572
rect 16204 10807 16244 10816
rect 15916 9715 15956 9724
rect 16012 10184 16052 10193
rect 15820 9295 15860 9304
rect 15916 8924 15956 8933
rect 15436 8707 15476 8716
rect 15820 8756 15860 8765
rect 15436 8504 15476 8513
rect 15436 7076 15476 8464
rect 15820 7916 15860 8716
rect 15916 8588 15956 8884
rect 15916 8168 15956 8548
rect 15916 8119 15956 8128
rect 16012 7916 16052 10144
rect 15820 7867 15860 7876
rect 15916 7876 16052 7916
rect 16108 9428 16148 9437
rect 15436 7027 15476 7036
rect 15820 6572 15860 6581
rect 15916 6572 15956 7876
rect 15860 6532 15956 6572
rect 16012 7244 16052 7253
rect 15436 6488 15476 6497
rect 15436 5648 15476 6448
rect 15436 5599 15476 5608
rect 15532 6404 15572 6413
rect 15340 5011 15380 5020
rect 15532 5564 15572 6364
rect 15820 6152 15860 6532
rect 15820 6103 15860 6112
rect 15532 5144 15572 5524
rect 15244 4423 15284 4432
rect 15148 4339 15188 4348
rect 14380 4255 14420 4264
rect 14284 4171 14324 4180
rect 13900 4087 13940 4096
rect 15532 4136 15572 5104
rect 15532 4087 15572 4096
rect 15820 5564 15860 5573
rect 15820 4136 15860 5524
rect 16012 5312 16052 7204
rect 16108 6656 16148 9388
rect 16204 8588 16244 8597
rect 16204 8168 16244 8548
rect 16204 8119 16244 8128
rect 16300 7244 16340 13252
rect 16396 13292 16436 13840
rect 16396 12452 16436 13252
rect 16492 13628 16532 13637
rect 16492 13040 16532 13588
rect 16492 12991 16532 13000
rect 16396 12403 16436 12412
rect 16492 12788 16532 12797
rect 16492 12620 16532 12748
rect 16492 11612 16532 12580
rect 16588 11948 16628 18376
rect 16684 17492 16724 19804
rect 16684 17408 16724 17452
rect 16684 17359 16724 17368
rect 16780 17828 16820 19972
rect 16876 18668 16916 20476
rect 16972 20180 17012 20644
rect 16972 20131 17012 20140
rect 16972 19256 17012 19265
rect 16972 18752 17012 19216
rect 16972 18703 17012 18712
rect 16876 18619 16916 18628
rect 17068 18584 17108 20812
rect 17164 20768 17204 21316
rect 17164 20719 17204 20728
rect 17260 20852 17300 21820
rect 17260 20717 17300 20812
rect 17164 20180 17204 20189
rect 17164 19928 17204 20140
rect 17164 19088 17204 19888
rect 17260 20012 17300 20021
rect 17260 19760 17300 19972
rect 17260 19711 17300 19720
rect 17164 19039 17204 19048
rect 17068 18535 17108 18544
rect 16780 17240 16820 17788
rect 17260 18416 17300 18425
rect 17260 18248 17300 18376
rect 17260 17660 17300 18208
rect 17260 17611 17300 17620
rect 16780 17191 16820 17200
rect 16876 17576 16916 17585
rect 16876 17156 16916 17536
rect 16972 17324 17012 17419
rect 16972 17275 17012 17284
rect 16876 17072 16916 17116
rect 16780 17032 16916 17072
rect 16588 11899 16628 11908
rect 16684 16988 16724 16997
rect 16684 16316 16724 16948
rect 16492 11563 16532 11572
rect 16588 11528 16628 11537
rect 16588 10100 16628 11488
rect 16588 10051 16628 10060
rect 16396 9932 16436 9941
rect 16396 9512 16436 9892
rect 16396 9463 16436 9472
rect 16300 7195 16340 7204
rect 16684 8588 16724 16276
rect 16780 14132 16820 17032
rect 16876 17021 16916 17032
rect 16972 17156 17012 17165
rect 16972 16316 17012 17116
rect 16972 16267 17012 16276
rect 17068 16988 17108 16997
rect 17260 16988 17300 16997
rect 17108 16948 17260 16988
rect 16876 16232 16916 16241
rect 16876 15812 16916 16192
rect 17068 16232 17108 16948
rect 17260 16939 17300 16948
rect 17260 16820 17300 16829
rect 17260 16232 17300 16780
rect 16876 15763 16916 15772
rect 16972 16148 17012 16157
rect 16972 15644 17012 16108
rect 16972 15595 17012 15604
rect 16876 15476 16916 15485
rect 17068 15476 17108 16192
rect 16916 15436 17108 15476
rect 17164 16192 17300 16232
rect 16876 15427 16916 15436
rect 17068 15308 17108 15317
rect 16876 14720 16916 14729
rect 16876 14300 16916 14680
rect 16876 14251 16916 14260
rect 17068 14468 17108 15268
rect 17164 14636 17204 16192
rect 17260 16064 17300 16073
rect 17260 15644 17300 16024
rect 17260 15595 17300 15604
rect 17164 14596 17300 14636
rect 16780 14083 16820 14092
rect 16972 14216 17012 14225
rect 16876 14048 16916 14057
rect 16876 13913 16916 14008
rect 16972 13880 17012 14176
rect 16972 13831 17012 13840
rect 17068 13880 17108 14428
rect 17068 13831 17108 13840
rect 16780 13208 16820 13217
rect 16780 12704 16820 13168
rect 17260 13040 17300 14596
rect 17356 14552 17396 26524
rect 17740 26564 17780 26573
rect 17452 25976 17492 25985
rect 17452 23120 17492 25936
rect 17548 25976 17588 25985
rect 17548 25388 17588 25936
rect 17548 25339 17588 25348
rect 17644 25808 17684 25817
rect 17548 24884 17588 24893
rect 17548 24800 17588 24844
rect 17548 24749 17588 24760
rect 17644 24548 17684 25768
rect 17740 25388 17780 26524
rect 18028 26396 18068 26405
rect 17740 25348 17876 25388
rect 17452 22532 17492 23080
rect 17452 22483 17492 22492
rect 17548 24508 17684 24548
rect 17740 24548 17780 24557
rect 17452 20012 17492 20021
rect 17452 19340 17492 19972
rect 17452 18332 17492 19300
rect 17452 15896 17492 18292
rect 17452 15847 17492 15856
rect 17452 15728 17492 15737
rect 17452 15644 17492 15688
rect 17452 15593 17492 15604
rect 17452 15476 17492 15485
rect 17452 15341 17492 15436
rect 17548 14888 17588 24508
rect 17740 23792 17780 24508
rect 17740 23743 17780 23752
rect 17644 23624 17684 23633
rect 17836 23624 17876 25348
rect 17644 21608 17684 23584
rect 17740 23584 17876 23624
rect 17740 23120 17780 23584
rect 18028 23372 18068 26356
rect 18220 26060 18260 26608
rect 18220 26011 18260 26020
rect 17932 23332 18068 23372
rect 18124 25640 18164 25649
rect 17740 23071 17780 23080
rect 17836 23288 17876 23297
rect 17836 22952 17876 23248
rect 17836 22903 17876 22912
rect 17644 20348 17684 21568
rect 17644 20299 17684 20308
rect 17740 20684 17780 20693
rect 17644 19844 17684 19853
rect 17644 16316 17684 19804
rect 17644 15140 17684 16276
rect 17644 15091 17684 15100
rect 17548 14839 17588 14848
rect 17644 14972 17684 14981
rect 17356 14503 17396 14512
rect 17452 14048 17492 14057
rect 17452 13376 17492 14008
rect 17452 13208 17492 13336
rect 17548 13880 17588 13889
rect 17548 13208 17588 13840
rect 17644 13544 17684 14932
rect 17740 14888 17780 20644
rect 17836 19256 17876 19265
rect 17836 18836 17876 19216
rect 17836 18787 17876 18796
rect 17836 18584 17876 18593
rect 17836 18449 17876 18544
rect 17836 18248 17876 18257
rect 17836 18080 17876 18208
rect 17836 18031 17876 18040
rect 17836 17912 17876 17921
rect 17836 17744 17876 17872
rect 17836 17695 17876 17704
rect 17740 14839 17780 14848
rect 17836 17576 17876 17585
rect 17740 14720 17780 14729
rect 17740 13964 17780 14680
rect 17740 13915 17780 13924
rect 17644 13495 17684 13504
rect 17740 13796 17780 13805
rect 17644 13208 17684 13217
rect 17548 13168 17644 13208
rect 17452 13159 17492 13168
rect 17644 13159 17684 13168
rect 17260 13000 17588 13040
rect 16780 12655 16820 12664
rect 17356 12620 17396 12629
rect 17164 12536 17204 12545
rect 16972 12452 17012 12461
rect 16876 12368 16916 12377
rect 16876 12032 16916 12328
rect 16876 11780 16916 11992
rect 16876 11731 16916 11740
rect 16780 11528 16820 11537
rect 16780 10436 16820 11488
rect 16780 10387 16820 10396
rect 16876 11024 16916 11033
rect 16684 8000 16724 8548
rect 16780 9428 16820 9437
rect 16780 8756 16820 9388
rect 16780 8084 16820 8716
rect 16780 8035 16820 8044
rect 16684 7244 16724 7960
rect 16684 7195 16724 7204
rect 16108 6607 16148 6616
rect 16396 7160 16436 7169
rect 16396 6572 16436 7120
rect 16876 6656 16916 10984
rect 16972 10940 17012 12412
rect 17068 12116 17108 12125
rect 17068 11717 17108 12076
rect 17068 11668 17108 11677
rect 17164 11948 17204 12496
rect 17356 12368 17396 12580
rect 17356 12319 17396 12328
rect 17452 12620 17492 12629
rect 16972 10891 17012 10900
rect 17164 10268 17204 11908
rect 17452 11024 17492 12580
rect 17452 10975 17492 10984
rect 17164 10219 17204 10228
rect 17548 10268 17588 13000
rect 17644 12956 17684 12965
rect 17644 12821 17684 12916
rect 17644 12452 17684 12461
rect 17644 11528 17684 12412
rect 17740 11696 17780 13756
rect 17740 11647 17780 11656
rect 17836 12536 17876 17536
rect 17932 16484 17972 23332
rect 18028 23120 18068 23129
rect 18028 23036 18068 23080
rect 18028 22985 18068 22996
rect 18124 22448 18164 25600
rect 18220 24464 18260 24473
rect 18220 23624 18260 24424
rect 18220 23575 18260 23584
rect 18220 23288 18260 23297
rect 18220 23036 18260 23248
rect 18220 22987 18260 22996
rect 18316 22952 18356 26860
rect 18508 26900 18548 26909
rect 18412 26648 18452 26657
rect 18412 26228 18452 26608
rect 18508 26564 18548 26860
rect 18508 26515 18548 26524
rect 18892 26648 18932 26659
rect 18892 26564 18932 26608
rect 18412 26093 18452 26188
rect 18892 26228 18932 26524
rect 18988 26480 19028 26489
rect 18988 26345 19028 26440
rect 19084 26312 19124 27448
rect 19180 27068 19220 27616
rect 22348 27656 22388 27665
rect 21100 27572 21140 27581
rect 20428 27404 20468 27413
rect 19180 27019 19220 27028
rect 19372 27068 19412 27077
rect 19372 26900 19412 27028
rect 19372 26851 19412 26860
rect 19660 26816 19700 26825
rect 19084 26263 19124 26272
rect 19276 26480 19316 26489
rect 18892 26179 18932 26188
rect 19084 26144 19124 26153
rect 18508 26060 18548 26069
rect 18412 25976 18452 26004
rect 18508 25976 18548 26020
rect 18452 25936 18548 25976
rect 18412 25927 18452 25936
rect 18412 25808 18452 25817
rect 18412 23060 18452 25768
rect 18508 25220 18548 25936
rect 18660 25724 19028 25733
rect 18660 25675 19028 25684
rect 19084 25472 19124 26104
rect 19084 25423 19124 25432
rect 18508 25171 18548 25180
rect 18988 25304 19028 25313
rect 18988 24716 19028 25264
rect 18988 24667 19028 24676
rect 18508 24632 18548 24641
rect 18508 23288 18548 24592
rect 18604 24548 18644 24557
rect 18604 24413 18644 24508
rect 18660 24212 19028 24221
rect 19180 24212 19220 24221
rect 18660 24163 19028 24172
rect 19084 24172 19180 24212
rect 18508 23239 18548 23248
rect 19084 23120 19124 24172
rect 19180 24163 19220 24172
rect 19180 23792 19220 23801
rect 19180 23288 19220 23752
rect 19180 23239 19220 23248
rect 19084 23071 19124 23080
rect 18412 23020 18548 23060
rect 18124 22399 18164 22408
rect 18220 22868 18260 22908
rect 18316 22903 18356 22912
rect 18220 22784 18260 22828
rect 18508 22784 18548 23020
rect 19276 22952 19316 26440
rect 19468 25976 19508 25985
rect 18220 22744 18548 22784
rect 19180 22912 19276 22952
rect 18028 22280 18068 22289
rect 18220 22280 18260 22744
rect 18660 22700 19028 22709
rect 18660 22651 19028 22660
rect 18604 22364 18644 22373
rect 18028 22145 18068 22240
rect 18124 22240 18260 22280
rect 18508 22280 18548 22289
rect 18028 21776 18068 21785
rect 18028 20600 18068 21736
rect 18028 20551 18068 20560
rect 17932 16435 17972 16444
rect 18028 19088 18068 19097
rect 17932 16148 17972 16157
rect 17932 15896 17972 16108
rect 17932 15847 17972 15856
rect 17932 15476 17972 15485
rect 17932 15308 17972 15436
rect 18028 15308 18068 19048
rect 18124 17912 18164 22240
rect 18316 22196 18356 22205
rect 18508 22196 18548 22240
rect 18356 22156 18548 22196
rect 18316 22147 18356 22156
rect 18220 22112 18260 22121
rect 18220 21524 18260 22072
rect 18220 21475 18260 21484
rect 18316 21608 18356 21617
rect 18124 17863 18164 17872
rect 18220 20768 18260 20777
rect 18124 17744 18164 17753
rect 18124 15392 18164 17704
rect 18220 16904 18260 20728
rect 18316 20600 18356 21568
rect 18508 21608 18548 22156
rect 18604 21776 18644 22324
rect 18988 22364 19028 22373
rect 18988 22112 19028 22324
rect 18988 22063 19028 22072
rect 19180 22196 19220 22912
rect 19276 22903 19316 22912
rect 19372 24968 19412 24977
rect 18604 21727 18644 21736
rect 18508 21559 18548 21568
rect 18988 21608 19028 21617
rect 18988 21473 19028 21568
rect 19180 21608 19220 22156
rect 19276 22700 19316 22709
rect 19276 21692 19316 22660
rect 19372 22448 19412 24928
rect 19468 24632 19508 25936
rect 19660 25808 19700 26776
rect 20332 26816 20372 26825
rect 20140 26648 20180 26743
rect 20140 26599 20180 26608
rect 19900 26480 20268 26489
rect 19900 26431 20268 26440
rect 20044 26228 20084 26237
rect 19660 25759 19700 25768
rect 19756 26060 19796 26069
rect 20044 26060 20084 26188
rect 20140 26060 20180 26069
rect 20044 26020 20140 26060
rect 19468 24583 19508 24592
rect 19660 25136 19700 25145
rect 19468 24296 19508 24305
rect 19468 23456 19508 24256
rect 19660 23792 19700 25096
rect 19756 24548 19796 26020
rect 20140 26011 20180 26020
rect 19900 24968 20268 24977
rect 19900 24919 20268 24928
rect 19756 24499 19796 24508
rect 19852 24800 19892 24809
rect 19852 23792 19892 24760
rect 20332 24548 20372 26776
rect 20428 26648 20468 27364
rect 20428 26599 20468 26608
rect 21004 27152 21044 27161
rect 20812 26144 20852 26153
rect 20812 26009 20852 26104
rect 20620 25220 20660 25229
rect 20620 24884 20660 25180
rect 20620 24835 20660 24844
rect 20716 25136 20756 25145
rect 20524 24800 20564 24809
rect 20428 24632 20468 24641
rect 20524 24632 20564 24760
rect 20468 24592 20564 24632
rect 20428 24583 20468 24592
rect 20236 24464 20276 24473
rect 19660 23743 19700 23752
rect 19756 23752 19852 23792
rect 19468 23407 19508 23416
rect 19660 23204 19700 23213
rect 19372 22399 19412 22408
rect 19564 23120 19604 23129
rect 19276 21643 19316 21652
rect 19180 21559 19220 21568
rect 19468 21524 19508 21533
rect 18508 21356 18548 21365
rect 18316 20516 18356 20560
rect 18316 20436 18356 20476
rect 18412 20852 18452 20861
rect 18412 20516 18452 20812
rect 18412 20467 18452 20476
rect 18508 20768 18548 21316
rect 18660 21188 19028 21197
rect 18660 21139 19028 21148
rect 18700 21020 18740 21029
rect 18508 20012 18548 20728
rect 18508 19963 18548 19972
rect 18604 20936 18644 20945
rect 18604 19844 18644 20896
rect 18700 20852 18740 20980
rect 18892 21020 18932 21029
rect 18740 20812 18836 20852
rect 18700 20803 18740 20812
rect 18604 19795 18644 19804
rect 18700 20432 18740 20441
rect 18700 19844 18740 20392
rect 18796 20348 18836 20812
rect 18796 20299 18836 20308
rect 18892 20264 18932 20980
rect 19468 20936 19508 21484
rect 19468 20887 19508 20896
rect 19084 20852 19124 20861
rect 19084 20717 19124 20812
rect 19372 20852 19412 20861
rect 19180 20684 19220 20693
rect 18892 20215 18932 20224
rect 19084 20600 19124 20609
rect 19084 20012 19124 20560
rect 19084 19963 19124 19972
rect 19180 19928 19220 20644
rect 19372 20684 19412 20812
rect 19372 20180 19412 20644
rect 19372 20131 19412 20140
rect 19468 20600 19508 20609
rect 19180 19879 19220 19888
rect 19276 20096 19316 20105
rect 18700 19795 18740 19804
rect 19084 19844 19124 19853
rect 18508 19760 18548 19769
rect 18316 18920 18356 18929
rect 18316 18416 18356 18880
rect 18316 18367 18356 18376
rect 18412 18752 18452 18761
rect 18412 18332 18452 18712
rect 18508 18584 18548 19720
rect 18660 19676 19028 19685
rect 18660 19627 19028 19636
rect 18604 19256 18644 19265
rect 18604 18752 18644 19216
rect 18604 18703 18644 18712
rect 18508 18535 18548 18544
rect 18604 18584 18644 18593
rect 18604 18332 18644 18544
rect 18988 18500 19028 18509
rect 18988 18365 19028 18460
rect 18412 18283 18452 18292
rect 18508 18292 18644 18332
rect 18316 17660 18356 17755
rect 18316 17611 18356 17620
rect 18412 17576 18452 17585
rect 18412 17240 18452 17536
rect 18412 17191 18452 17200
rect 18316 17072 18356 17081
rect 18316 16937 18356 17032
rect 18220 16855 18260 16864
rect 18412 16904 18452 16913
rect 18316 16484 18356 16493
rect 18316 16232 18356 16444
rect 18316 16183 18356 16192
rect 18316 15896 18356 15905
rect 18220 15560 18260 15655
rect 18220 15511 18260 15520
rect 18124 15352 18260 15392
rect 18028 15268 18164 15308
rect 17932 15259 17972 15268
rect 18028 15140 18068 15149
rect 17836 11696 17876 12496
rect 17836 11647 17876 11656
rect 17932 15056 17972 15065
rect 17644 11488 17780 11528
rect 17740 11192 17780 11488
rect 17740 10520 17780 11152
rect 17740 10471 17780 10480
rect 17836 11024 17876 11033
rect 17548 10219 17588 10228
rect 17644 10184 17684 10279
rect 17644 10135 17684 10144
rect 17836 10268 17876 10984
rect 17836 10184 17876 10228
rect 17836 10135 17876 10144
rect 17836 10016 17876 10025
rect 17548 9932 17588 9941
rect 17260 9428 17300 9437
rect 17452 9428 17492 9437
rect 17300 9388 17452 9428
rect 17260 9379 17300 9388
rect 17452 9379 17492 9388
rect 17260 9260 17300 9269
rect 17260 8924 17300 9220
rect 17260 8875 17300 8884
rect 17548 8252 17588 9892
rect 17644 9680 17684 9689
rect 17836 9680 17876 9976
rect 17684 9640 17876 9680
rect 17644 9631 17684 9640
rect 17164 8000 17204 8009
rect 17164 7412 17204 7960
rect 17068 7160 17108 7169
rect 16876 6607 16916 6616
rect 16972 6992 17012 7001
rect 16396 6523 16436 6532
rect 16492 6488 16532 6497
rect 16300 6236 16340 6245
rect 16300 5732 16340 6196
rect 16300 5683 16340 5692
rect 16492 5648 16532 6448
rect 16972 6488 17012 6952
rect 16972 6439 17012 6448
rect 17068 6152 17108 7120
rect 17164 6908 17204 7372
rect 17164 6859 17204 6868
rect 17548 8000 17588 8212
rect 17932 8672 17972 15016
rect 18028 12620 18068 15100
rect 18028 12571 18068 12580
rect 17644 8000 17684 8009
rect 17548 7960 17644 8000
rect 17548 7076 17588 7960
rect 17644 7951 17684 7960
rect 17548 6488 17588 7036
rect 17548 6439 17588 6448
rect 16492 5599 16532 5608
rect 16684 5648 16724 5657
rect 16012 5263 16052 5272
rect 16204 5480 16244 5489
rect 16108 4892 16148 4901
rect 16108 4388 16148 4852
rect 16108 4339 16148 4348
rect 15820 4087 15860 4096
rect 16204 4136 16244 5440
rect 16204 4087 16244 4096
rect 16684 5060 16724 5608
rect 16684 4052 16724 5020
rect 17068 5648 17108 6112
rect 17068 4640 17108 5608
rect 17068 4591 17108 4600
rect 17164 4892 17204 4901
rect 17164 4304 17204 4852
rect 17932 4892 17972 8632
rect 18028 11108 18068 11117
rect 18028 8168 18068 11068
rect 18124 10856 18164 15268
rect 18220 11948 18260 15352
rect 18316 14216 18356 15856
rect 18316 13964 18356 14176
rect 18316 13915 18356 13924
rect 18316 13712 18356 13721
rect 18316 13376 18356 13672
rect 18316 13327 18356 13336
rect 18316 13208 18356 13219
rect 18316 13124 18356 13168
rect 18316 13075 18356 13084
rect 18412 12704 18452 16864
rect 18508 16148 18548 18292
rect 18660 18164 19028 18173
rect 18660 18115 19028 18124
rect 18988 17912 19028 17921
rect 18604 17828 18644 17837
rect 18604 17240 18644 17788
rect 18796 17828 18836 17837
rect 18604 17191 18644 17200
rect 18700 17744 18740 17753
rect 18700 16904 18740 17704
rect 18700 16855 18740 16864
rect 18796 16820 18836 17788
rect 18988 17744 19028 17872
rect 19084 17828 19124 19804
rect 19276 19760 19316 20056
rect 19084 17779 19124 17788
rect 19180 19720 19316 19760
rect 19372 20012 19412 20021
rect 18988 17695 19028 17704
rect 19180 17660 19220 19720
rect 19372 19676 19412 19972
rect 19276 19636 19412 19676
rect 19276 19256 19316 19636
rect 19276 19207 19316 19216
rect 19372 19340 19412 19349
rect 19276 18752 19316 18847
rect 19276 18703 19316 18712
rect 19276 18584 19316 18593
rect 19276 18164 19316 18544
rect 19276 18115 19316 18124
rect 19372 17828 19412 19300
rect 19372 17779 19412 17788
rect 19084 17620 19220 17660
rect 19276 17660 19316 17669
rect 18892 17156 18932 17165
rect 18892 17072 18932 17116
rect 18892 17021 18932 17032
rect 18796 16771 18836 16780
rect 18660 16652 19028 16661
rect 18660 16603 19028 16612
rect 18988 16400 19028 16409
rect 18988 16265 19028 16360
rect 18508 15728 18548 16108
rect 19084 16148 19124 17620
rect 19180 17492 19220 17501
rect 19180 16652 19220 17452
rect 19180 16603 19220 16612
rect 19276 16316 19316 17620
rect 19276 16267 19316 16276
rect 19372 17072 19412 17081
rect 19372 16652 19412 17032
rect 19084 16099 19124 16108
rect 19180 16232 19220 16241
rect 18508 15679 18548 15688
rect 18604 16064 18644 16073
rect 18604 15560 18644 16024
rect 19180 15644 19220 16192
rect 19180 15595 19220 15604
rect 19276 16148 19316 16157
rect 18508 15520 18644 15560
rect 19084 15560 19124 15569
rect 18508 15392 18548 15520
rect 18508 14048 18548 15352
rect 18660 15140 19028 15149
rect 18660 15091 19028 15100
rect 18604 14972 18644 14981
rect 18604 14804 18644 14932
rect 18604 14755 18644 14764
rect 19084 14720 19124 15520
rect 19084 14468 19124 14680
rect 19276 14636 19316 16108
rect 19372 15224 19412 16612
rect 19372 15175 19412 15184
rect 19276 14587 19316 14596
rect 19372 14720 19412 14729
rect 19372 14468 19412 14680
rect 19084 14428 19412 14468
rect 18604 14300 18644 14309
rect 18604 14132 18644 14260
rect 18604 14083 18644 14092
rect 18508 13964 18548 14008
rect 18508 13292 18548 13924
rect 18700 14048 18740 14057
rect 18700 13913 18740 14008
rect 19084 13796 19124 14428
rect 18660 13628 19028 13637
rect 18660 13579 19028 13588
rect 18508 13243 18548 13252
rect 19084 13460 19124 13756
rect 19180 14216 19220 14225
rect 19180 13544 19220 14176
rect 19180 13495 19220 13504
rect 19372 14216 19412 14225
rect 19084 13208 19124 13420
rect 19084 13159 19124 13168
rect 18412 12655 18452 12664
rect 18316 12536 18356 12545
rect 18316 12401 18356 12496
rect 18508 12536 18548 12545
rect 18412 12452 18452 12461
rect 18412 12116 18452 12412
rect 18412 12067 18452 12076
rect 18220 11899 18260 11908
rect 18508 11948 18548 12496
rect 18660 12116 19028 12125
rect 18660 12067 19028 12076
rect 19180 12116 19220 12125
rect 18508 11899 18548 11908
rect 19084 11948 19124 11957
rect 18412 11696 18452 11705
rect 18412 11192 18452 11656
rect 18508 11696 18548 11705
rect 18508 11612 18548 11656
rect 18508 11561 18548 11572
rect 18412 11143 18452 11152
rect 18700 11528 18740 11537
rect 18700 11192 18740 11488
rect 18700 11143 18740 11152
rect 18124 10807 18164 10816
rect 18220 10940 18260 10949
rect 18220 10268 18260 10900
rect 19084 10856 19124 11908
rect 19180 11696 19220 12076
rect 19180 11561 19220 11656
rect 19276 11948 19316 11957
rect 19084 10807 19124 10816
rect 18220 10219 18260 10228
rect 18412 10688 18452 10697
rect 18124 10184 18164 10195
rect 18124 10100 18164 10144
rect 18124 10051 18164 10060
rect 18316 10100 18356 10109
rect 18316 9965 18356 10060
rect 18412 9932 18452 10648
rect 19180 10688 19220 10697
rect 18660 10604 19028 10613
rect 18660 10555 19028 10564
rect 18412 9883 18452 9892
rect 18508 10184 18548 10193
rect 18508 10016 18548 10144
rect 18028 8119 18068 8128
rect 18124 9512 18164 9521
rect 18124 5480 18164 9472
rect 18220 8588 18260 8597
rect 18220 8000 18260 8548
rect 18508 8588 18548 9976
rect 18660 9092 19028 9101
rect 18660 9043 19028 9052
rect 18508 8539 18548 8548
rect 19180 9008 19220 10648
rect 19180 8672 19220 8968
rect 18796 8504 18836 8513
rect 18796 8084 18836 8464
rect 18796 8035 18836 8044
rect 18220 7951 18260 7960
rect 18660 7580 19028 7589
rect 18660 7531 19028 7540
rect 19180 7160 19220 8632
rect 19276 7412 19316 11908
rect 19372 11276 19412 14176
rect 19468 13292 19508 20560
rect 19564 20264 19604 23080
rect 19564 20215 19604 20224
rect 19564 20096 19604 20105
rect 19660 20096 19700 23164
rect 19756 23120 19796 23752
rect 19852 23743 19892 23752
rect 19948 23960 19988 23969
rect 19948 23624 19988 23920
rect 20236 23876 20276 24424
rect 20236 23827 20276 23836
rect 19948 23575 19988 23584
rect 19900 23456 20268 23465
rect 19900 23407 20268 23416
rect 20236 23288 20276 23297
rect 20236 23153 20276 23248
rect 19756 23071 19796 23080
rect 19756 22364 19796 22373
rect 19756 20852 19796 22324
rect 20332 22280 20372 24508
rect 20524 23792 20564 23801
rect 20428 23624 20468 23633
rect 20428 23204 20468 23584
rect 20524 23372 20564 23752
rect 20524 23323 20564 23332
rect 20620 23624 20660 23633
rect 20620 23204 20660 23584
rect 20428 23155 20468 23164
rect 20524 23164 20660 23204
rect 20332 22240 20468 22280
rect 20332 22112 20372 22121
rect 19900 21944 20268 21953
rect 19900 21895 20268 21904
rect 20332 21608 20372 22072
rect 20332 21559 20372 21568
rect 19756 20803 19796 20812
rect 20044 21440 20084 21449
rect 19756 20684 19796 20693
rect 19756 20549 19796 20644
rect 20044 20600 20084 21400
rect 20428 21020 20468 22240
rect 20428 20971 20468 20980
rect 20044 20551 20084 20560
rect 19900 20432 20268 20441
rect 19900 20383 20268 20392
rect 20044 20264 20084 20273
rect 19660 20056 19796 20096
rect 19564 19508 19604 20056
rect 19564 19459 19604 19468
rect 19660 19928 19700 19937
rect 19570 19256 19610 19265
rect 19564 19216 19570 19256
rect 19564 19207 19610 19216
rect 19564 17156 19604 19207
rect 19660 19172 19700 19888
rect 19660 19123 19700 19132
rect 19564 17107 19604 17116
rect 19660 18500 19700 18509
rect 19756 18500 19796 20056
rect 20044 19088 20084 20224
rect 20140 19340 20180 19349
rect 20140 19205 20180 19300
rect 20524 19256 20564 23164
rect 20716 23060 20756 25096
rect 21004 24548 21044 27112
rect 21004 24499 21044 24508
rect 20908 23708 20948 23717
rect 20908 23060 20948 23668
rect 21100 23060 21140 27532
rect 21964 27572 22004 27581
rect 20620 23020 20756 23060
rect 20812 23020 20948 23060
rect 21004 23020 21140 23060
rect 21196 27404 21236 27413
rect 21196 26816 21236 27364
rect 21964 27068 22004 27532
rect 21964 27019 22004 27028
rect 20620 21440 20660 23020
rect 20716 22868 20756 22877
rect 20716 21608 20756 22828
rect 20716 21559 20756 21568
rect 20812 22112 20852 23020
rect 20908 22952 20948 22963
rect 20908 22868 20948 22912
rect 20908 22819 20948 22828
rect 20620 21400 20756 21440
rect 20428 19216 20564 19256
rect 20620 20768 20660 20777
rect 20044 19039 20084 19048
rect 20332 19172 20372 19181
rect 19900 18920 20268 18929
rect 19900 18871 20268 18880
rect 20332 18752 20372 19132
rect 20332 18703 20372 18712
rect 20428 18584 20468 19216
rect 19700 18460 19796 18500
rect 20332 18500 20372 18509
rect 19564 16232 19604 16241
rect 19564 16148 19604 16192
rect 19564 16097 19604 16108
rect 19564 15560 19604 15569
rect 19564 14132 19604 15520
rect 19564 13460 19604 14092
rect 19564 13411 19604 13420
rect 19660 13292 19700 18460
rect 20236 18080 20276 18089
rect 19756 17912 19796 17921
rect 19756 16316 19796 17872
rect 20236 17828 20276 18040
rect 20236 17779 20276 17788
rect 20332 17660 20372 18460
rect 20428 17912 20468 18544
rect 20428 17863 20468 17872
rect 20524 18668 20564 18677
rect 20524 17744 20564 18628
rect 20524 17695 20564 17704
rect 20620 18080 20660 20728
rect 20716 19340 20756 21400
rect 20812 20768 20852 22072
rect 20908 22280 20948 22289
rect 20908 21776 20948 22240
rect 20908 21727 20948 21736
rect 20812 20719 20852 20728
rect 20908 21440 20948 21449
rect 20812 20180 20852 20189
rect 20812 19760 20852 20140
rect 20812 19711 20852 19720
rect 20716 19291 20756 19300
rect 19900 17408 20268 17417
rect 19900 17359 20268 17368
rect 19948 17240 19988 17249
rect 19852 17156 19892 17165
rect 19852 17021 19892 17116
rect 19756 16267 19796 16276
rect 19948 16148 19988 17200
rect 20332 17156 20372 17620
rect 20332 17107 20372 17116
rect 20524 17576 20564 17585
rect 20236 17072 20276 17081
rect 20140 16904 20180 16913
rect 20140 16769 20180 16864
rect 20236 16484 20276 17032
rect 20236 16435 20276 16444
rect 20332 16988 20372 16997
rect 20332 16736 20372 16948
rect 19756 16108 19988 16148
rect 19756 15728 19796 16108
rect 19900 15896 20268 15905
rect 19900 15847 20268 15856
rect 19756 15679 19796 15688
rect 19852 15644 19892 15653
rect 19852 14972 19892 15604
rect 20332 15644 20372 16696
rect 19948 15560 19988 15569
rect 19948 15224 19988 15520
rect 19948 15175 19988 15184
rect 19852 14923 19892 14932
rect 19948 14720 19988 14729
rect 19756 14636 19796 14645
rect 19756 14300 19796 14596
rect 19948 14552 19988 14680
rect 19948 14503 19988 14512
rect 19900 14384 20268 14393
rect 19900 14335 20268 14344
rect 19756 14251 19796 14260
rect 20140 14216 20180 14225
rect 20332 14216 20372 15604
rect 20524 15560 20564 17536
rect 20620 17072 20660 18040
rect 20716 19172 20756 19181
rect 20716 17240 20756 19132
rect 20812 18584 20852 18593
rect 20812 18080 20852 18544
rect 20812 18031 20852 18040
rect 20716 17191 20756 17200
rect 20812 17576 20852 17585
rect 20620 17032 20756 17072
rect 20524 15511 20564 15520
rect 20180 14176 20372 14216
rect 20428 15476 20468 15485
rect 20140 14167 20180 14176
rect 20236 14048 20276 14059
rect 19756 13964 19796 13973
rect 19756 13796 19796 13924
rect 19756 13747 19796 13756
rect 20236 13964 20276 14008
rect 19468 13252 19604 13292
rect 19468 12788 19508 12797
rect 19468 12452 19508 12748
rect 19468 11780 19508 12412
rect 19468 11731 19508 11740
rect 19564 12032 19604 13252
rect 19660 13243 19700 13252
rect 19756 13544 19796 13553
rect 19372 11227 19412 11236
rect 19564 11024 19604 11992
rect 19756 11780 19796 13504
rect 20236 13040 20276 13924
rect 20236 12991 20276 13000
rect 20428 12956 20468 15436
rect 20620 14888 20660 14897
rect 20524 14636 20564 14645
rect 20524 14468 20564 14596
rect 20524 14419 20564 14428
rect 19900 12872 20268 12881
rect 19900 12823 20268 12832
rect 20140 12368 20180 12377
rect 20140 12233 20180 12328
rect 20428 12284 20468 12916
rect 20524 14300 20564 14309
rect 20524 14048 20564 14260
rect 20524 13040 20564 14008
rect 20620 13964 20660 14848
rect 20620 13208 20660 13924
rect 20620 13159 20660 13168
rect 20524 12452 20564 13000
rect 20716 12980 20756 17032
rect 20812 16988 20852 17536
rect 20812 16939 20852 16948
rect 20812 14636 20852 14645
rect 20812 14300 20852 14596
rect 20812 14251 20852 14260
rect 20716 12940 20852 12980
rect 20524 12403 20564 12412
rect 20428 12235 20468 12244
rect 19756 11731 19796 11740
rect 20716 11864 20756 11873
rect 20620 11696 20660 11705
rect 20428 11612 20468 11621
rect 19900 11360 20268 11369
rect 19900 11311 20268 11320
rect 19564 10975 19604 10984
rect 19468 10940 19508 10949
rect 19372 10688 19412 10697
rect 19372 10184 19412 10648
rect 19372 9596 19412 10144
rect 19372 9547 19412 9556
rect 19468 10268 19508 10900
rect 20140 10856 20180 10865
rect 20140 10721 20180 10816
rect 20236 10352 20276 10361
rect 20276 10312 20372 10352
rect 20236 10303 20276 10312
rect 19468 9512 19508 10228
rect 19468 9463 19508 9472
rect 19660 10268 19700 10277
rect 19468 9260 19508 9269
rect 19468 8756 19508 9220
rect 19660 8840 19700 10228
rect 19756 10184 19796 10193
rect 19756 8924 19796 10144
rect 19900 9848 20268 9857
rect 19900 9799 20268 9808
rect 19756 8875 19796 8884
rect 19852 9512 19892 9521
rect 19660 8791 19700 8800
rect 19468 8707 19508 8716
rect 19660 8588 19700 8597
rect 19372 8336 19412 8345
rect 19372 8000 19412 8296
rect 19372 7951 19412 7960
rect 19276 7363 19316 7372
rect 19660 7244 19700 8548
rect 19756 8588 19796 8628
rect 19756 8504 19796 8548
rect 19852 8504 19892 9472
rect 20332 9428 20372 10312
rect 20332 9379 20372 9388
rect 19948 8588 19988 8683
rect 19948 8539 19988 8548
rect 19756 8464 19892 8504
rect 19756 8168 19796 8464
rect 19900 8336 20268 8345
rect 19900 8287 20268 8296
rect 19756 8119 19796 8128
rect 20428 8168 20468 11572
rect 20620 11192 20660 11656
rect 20620 11143 20660 11152
rect 20716 11024 20756 11824
rect 20716 10975 20756 10984
rect 20428 8119 20468 8128
rect 20620 10100 20660 10109
rect 20620 8588 20660 10060
rect 20812 9680 20852 12940
rect 20908 11948 20948 21400
rect 21004 21188 21044 23020
rect 21196 22196 21236 26776
rect 21484 26816 21524 26825
rect 21388 25976 21428 25985
rect 21292 25724 21332 25733
rect 21292 24632 21332 25684
rect 21292 24583 21332 24592
rect 21292 24464 21332 24473
rect 21292 23288 21332 24424
rect 21292 23239 21332 23248
rect 21196 22147 21236 22156
rect 21292 23120 21332 23129
rect 21004 21139 21044 21148
rect 21292 21020 21332 23080
rect 21292 20971 21332 20980
rect 21004 20684 21044 20693
rect 21004 18332 21044 20644
rect 21292 19256 21332 19265
rect 21292 18836 21332 19216
rect 21292 18787 21332 18796
rect 21292 18668 21332 18708
rect 21292 18584 21332 18628
rect 21004 17744 21044 18292
rect 21196 18500 21236 18509
rect 21196 17828 21236 18460
rect 21196 17779 21236 17788
rect 21004 17695 21044 17704
rect 21100 17072 21140 17081
rect 21100 15812 21140 17032
rect 21100 15763 21140 15772
rect 21196 16484 21236 16493
rect 21100 14804 21140 14813
rect 21100 13460 21140 14764
rect 21100 13411 21140 13420
rect 21196 12872 21236 16444
rect 21292 16232 21332 18544
rect 21388 18416 21428 25936
rect 21484 25808 21524 26776
rect 21484 25304 21524 25768
rect 22348 26144 22388 27616
rect 21772 25640 21812 25649
rect 21484 25255 21524 25264
rect 21580 25556 21620 25565
rect 21580 24716 21620 25516
rect 21772 25388 21812 25600
rect 21772 25339 21812 25348
rect 21676 25304 21716 25313
rect 21676 24800 21716 25264
rect 22348 25304 22388 26104
rect 21676 24751 21716 24760
rect 21868 25220 21908 25229
rect 21868 24800 21908 25180
rect 21868 24751 21908 24760
rect 21580 24667 21620 24676
rect 21964 24548 22004 24557
rect 21676 24464 21716 24473
rect 21484 24380 21524 24389
rect 21484 23876 21524 24340
rect 21484 23120 21524 23836
rect 21676 23792 21716 24424
rect 21484 23071 21524 23080
rect 21580 23752 21676 23792
rect 21484 22028 21524 22037
rect 21484 21356 21524 21988
rect 21484 21307 21524 21316
rect 21580 20852 21620 23752
rect 21676 23657 21716 23752
rect 21772 24380 21812 24389
rect 21772 23288 21812 24340
rect 21772 23239 21812 23248
rect 21868 24128 21908 24137
rect 21772 23036 21812 23045
rect 21772 22532 21812 22996
rect 21676 22364 21716 22373
rect 21676 21524 21716 22324
rect 21772 21692 21812 22492
rect 21772 21643 21812 21652
rect 21676 21475 21716 21484
rect 21868 21440 21908 24088
rect 21868 21391 21908 21400
rect 21964 23792 22004 24508
rect 22156 23960 22196 23969
rect 22156 23876 22196 23920
rect 22156 23825 22196 23836
rect 21580 20803 21620 20812
rect 21868 20936 21908 20945
rect 21868 20012 21908 20896
rect 21964 20852 22004 23752
rect 22156 23708 22196 23717
rect 22156 23204 22196 23668
rect 22156 23155 22196 23164
rect 22348 23204 22388 25264
rect 22540 27572 22580 27581
rect 22444 24380 22484 24389
rect 22444 23708 22484 24340
rect 22444 23659 22484 23668
rect 22348 23155 22388 23164
rect 22060 23120 22100 23129
rect 22060 22616 22100 23080
rect 22060 22567 22100 22576
rect 22156 23036 22196 23045
rect 22156 22532 22196 22996
rect 22540 22784 22580 27532
rect 23116 26984 23156 28600
rect 23404 27404 23444 27413
rect 23116 26935 23156 26944
rect 23308 27320 23348 27329
rect 23116 26816 23156 26825
rect 22540 22735 22580 22744
rect 22636 26312 22676 26321
rect 22636 22868 22676 26272
rect 22828 25892 22868 25901
rect 22732 25136 22772 25145
rect 22732 24548 22772 25096
rect 22828 24632 22868 25852
rect 22924 25220 22964 25229
rect 22924 24716 22964 25180
rect 23116 24800 23156 26776
rect 23116 24751 23156 24760
rect 23308 24716 23348 27280
rect 22924 24676 23060 24716
rect 22828 24592 22964 24632
rect 22732 24499 22772 24508
rect 22828 24464 22868 24473
rect 22828 23792 22868 24424
rect 22828 23743 22868 23752
rect 22924 23624 22964 24592
rect 23020 24548 23060 24676
rect 23308 24667 23348 24676
rect 23404 26900 23444 27364
rect 23020 24499 23060 24508
rect 23116 24632 23156 24641
rect 23116 24296 23156 24592
rect 23116 24247 23156 24256
rect 23212 24632 23252 24641
rect 23212 23876 23252 24592
rect 23308 24464 23348 24473
rect 23308 24044 23348 24424
rect 23308 23995 23348 24004
rect 23212 23827 23252 23836
rect 23308 23792 23348 23801
rect 22924 23575 22964 23584
rect 23212 23708 23252 23717
rect 23212 23204 23252 23668
rect 23308 23372 23348 23752
rect 23308 23323 23348 23332
rect 23212 23155 23252 23164
rect 22156 22483 22196 22492
rect 22636 22448 22676 22828
rect 23404 22952 23444 26860
rect 23596 26648 23636 26657
rect 23500 23876 23540 23885
rect 23500 23741 23540 23836
rect 23020 22616 23060 22625
rect 22636 22399 22676 22408
rect 22924 22576 23020 22616
rect 22252 22364 22292 22373
rect 22060 22280 22100 22289
rect 22060 21860 22100 22240
rect 22060 21811 22100 21820
rect 22252 22196 22292 22324
rect 22252 21608 22292 22156
rect 22732 22364 22772 22373
rect 22540 22112 22580 22121
rect 22540 21692 22580 22072
rect 22732 21776 22772 22324
rect 22828 22280 22868 22289
rect 22828 22145 22868 22240
rect 22732 21727 22772 21736
rect 22540 21643 22580 21652
rect 22252 21559 22292 21568
rect 22828 21608 22868 21617
rect 22060 21524 22100 21533
rect 22060 21389 22100 21484
rect 22828 21272 22868 21568
rect 22924 21524 22964 22576
rect 23020 22548 23060 22576
rect 23116 22364 23156 22373
rect 23116 22229 23156 22324
rect 23404 22364 23444 22912
rect 23404 22315 23444 22324
rect 23500 23624 23540 23633
rect 23212 22280 23252 22291
rect 23212 22196 23252 22240
rect 23212 22147 23252 22156
rect 23308 22280 23348 22289
rect 23308 21860 23348 22240
rect 23308 21811 23348 21820
rect 22924 21475 22964 21484
rect 23308 21440 23348 21449
rect 22828 21223 22868 21232
rect 23116 21356 23156 21365
rect 21964 20803 22004 20812
rect 22156 20768 22196 20777
rect 22156 20096 22196 20728
rect 23116 20768 23156 21316
rect 23116 20719 23156 20728
rect 22156 20047 22196 20056
rect 21868 19963 21908 19972
rect 22828 19844 22868 19853
rect 22636 19592 22676 19601
rect 22348 19424 22388 19433
rect 21772 19256 21812 19265
rect 21388 18367 21428 18376
rect 21676 18584 21716 18593
rect 21580 18080 21620 18089
rect 21580 17240 21620 18040
rect 21580 16988 21620 17200
rect 21580 16939 21620 16948
rect 21484 16904 21524 16913
rect 21484 16316 21524 16864
rect 21484 16267 21524 16276
rect 21580 16820 21620 16829
rect 21292 16183 21332 16192
rect 21580 16148 21620 16780
rect 21388 15560 21428 15569
rect 21292 15308 21332 15317
rect 21292 13460 21332 15268
rect 21388 14216 21428 15520
rect 21580 15560 21620 16108
rect 21580 15511 21620 15520
rect 21388 14167 21428 14176
rect 21484 14804 21524 14813
rect 21484 14048 21524 14764
rect 21484 13999 21524 14008
rect 21580 14720 21620 14729
rect 21580 13880 21620 14680
rect 21580 13831 21620 13840
rect 21292 13411 21332 13420
rect 20908 11899 20948 11908
rect 21100 12284 21140 12293
rect 20428 8000 20468 8009
rect 20428 7496 20468 7960
rect 20620 7748 20660 8548
rect 20620 7699 20660 7708
rect 20716 9640 20852 9680
rect 20908 11780 20948 11789
rect 20908 9680 20948 11740
rect 21100 11780 21140 12244
rect 21100 11731 21140 11740
rect 21196 11024 21236 12832
rect 21676 12536 21716 18544
rect 21772 18500 21812 19216
rect 22156 19256 22196 19265
rect 21772 18451 21812 18460
rect 21868 18500 21908 18509
rect 21772 17576 21812 17585
rect 21772 17492 21812 17536
rect 21772 17441 21812 17452
rect 21868 16316 21908 18460
rect 21964 18248 22004 18343
rect 21964 18199 22004 18208
rect 21964 18080 22004 18089
rect 21964 17744 22004 18040
rect 22156 17996 22196 19216
rect 22252 19172 22292 19181
rect 22252 18332 22292 19132
rect 22348 18668 22388 19384
rect 22636 19256 22676 19552
rect 22636 19207 22676 19216
rect 22348 18619 22388 18628
rect 22252 18283 22292 18292
rect 22444 18500 22484 18509
rect 22156 17947 22196 17956
rect 21964 16988 22004 17704
rect 21964 16939 22004 16948
rect 22060 17828 22100 17837
rect 22060 17072 22100 17788
rect 21868 14552 21908 16276
rect 22060 16652 22100 17032
rect 22348 17744 22388 17753
rect 22060 16148 22100 16612
rect 22060 15728 22100 16108
rect 22060 15679 22100 15688
rect 22156 16988 22196 16997
rect 21868 14503 21908 14512
rect 22060 15560 22100 15569
rect 22060 14888 22100 15520
rect 22060 14552 22100 14848
rect 22156 14720 22196 16948
rect 22252 15308 22292 15317
rect 22252 14804 22292 15268
rect 22252 14755 22292 14764
rect 22156 14671 22196 14680
rect 22060 14503 22100 14512
rect 22156 13880 22196 13889
rect 22156 13712 22196 13840
rect 22156 13208 22196 13672
rect 22156 13159 22196 13168
rect 21580 12116 21620 12125
rect 21580 11108 21620 12076
rect 21676 11948 21716 12496
rect 21676 11899 21716 11908
rect 21580 11059 21620 11068
rect 21676 11360 21716 11369
rect 20428 7447 20468 7456
rect 19660 7195 19700 7204
rect 19276 7160 19316 7169
rect 19180 7120 19276 7160
rect 19276 7111 19316 7120
rect 20524 7160 20564 7169
rect 19564 7076 19604 7085
rect 18988 6908 19028 6917
rect 18988 6656 19028 6868
rect 19028 6616 19124 6656
rect 18988 6607 19028 6616
rect 18660 6068 19028 6077
rect 18660 6019 19028 6028
rect 18892 5732 18932 5741
rect 18124 5431 18164 5440
rect 18412 5648 18452 5657
rect 18412 4976 18452 5608
rect 18700 5648 18740 5657
rect 18700 5144 18740 5608
rect 18892 5228 18932 5692
rect 19084 5648 19124 6616
rect 19084 5599 19124 5608
rect 19276 6404 19316 6413
rect 18892 5179 18932 5188
rect 18700 5095 18740 5104
rect 18412 4927 18452 4936
rect 17932 4843 17972 4852
rect 19276 4724 19316 6364
rect 19564 6068 19604 7036
rect 20524 7025 20564 7120
rect 19900 6824 20268 6833
rect 19900 6775 20268 6784
rect 20716 6572 20756 9640
rect 20908 9631 20948 9640
rect 21004 10352 21044 10361
rect 20908 8588 20948 8597
rect 20812 7916 20852 7925
rect 20812 7412 20852 7876
rect 20812 7363 20852 7372
rect 20908 7328 20948 8548
rect 20908 7279 20948 7288
rect 20716 6523 20756 6532
rect 21004 6740 21044 10312
rect 21196 10268 21236 10984
rect 21580 10604 21620 10613
rect 21580 10436 21620 10564
rect 21580 10387 21620 10396
rect 21196 10219 21236 10228
rect 21292 10184 21332 10279
rect 21292 10135 21332 10144
rect 21676 10184 21716 11320
rect 22060 11024 22100 11033
rect 21676 10135 21716 10144
rect 21868 10184 21908 10193
rect 21676 10016 21716 10025
rect 21196 9512 21236 9521
rect 21100 8588 21140 8597
rect 21100 8168 21140 8548
rect 21100 8119 21140 8128
rect 19564 5732 19604 6028
rect 20236 6488 20276 6497
rect 20236 5816 20276 6448
rect 20620 6488 20660 6497
rect 20620 5900 20660 6448
rect 20620 5851 20660 5860
rect 20908 6488 20948 6497
rect 20908 5900 20948 6448
rect 20908 5851 20948 5860
rect 20236 5767 20276 5776
rect 19564 5683 19604 5692
rect 20812 5732 20852 5741
rect 21004 5732 21044 6700
rect 21196 6656 21236 9472
rect 21676 9176 21716 9976
rect 21868 9428 21908 10144
rect 21868 9379 21908 9388
rect 21964 9512 22004 9521
rect 21676 9127 21716 9136
rect 21868 9008 21908 9017
rect 21772 8924 21812 8933
rect 21676 8672 21716 8681
rect 21388 8000 21428 8009
rect 21388 7076 21428 7960
rect 21388 7027 21428 7036
rect 21196 6607 21236 6616
rect 20852 5692 21044 5732
rect 19900 5312 20268 5321
rect 19900 5263 20268 5272
rect 19276 4675 19316 4684
rect 20812 4640 20852 5692
rect 21004 5648 21044 5692
rect 21292 6320 21332 6329
rect 21292 5732 21332 6280
rect 21292 5683 21332 5692
rect 21388 5984 21428 5993
rect 21004 5599 21044 5608
rect 20908 5564 20948 5573
rect 20908 5060 20948 5524
rect 21004 5060 21044 5088
rect 20908 5020 21004 5060
rect 20908 4976 20948 5020
rect 21004 5011 21044 5020
rect 20908 4927 20948 4936
rect 21388 4976 21428 5944
rect 21676 5648 21716 8632
rect 21772 8000 21812 8884
rect 21772 7951 21812 7960
rect 21772 7244 21812 7255
rect 21772 7160 21812 7204
rect 21772 7111 21812 7120
rect 21868 7076 21908 8968
rect 21964 8924 22004 9472
rect 21964 8875 22004 8884
rect 21908 7036 22004 7076
rect 21868 7027 21908 7036
rect 21772 6908 21812 6917
rect 21772 6656 21812 6868
rect 21772 6607 21812 6616
rect 21676 5599 21716 5608
rect 21868 6572 21908 6581
rect 21868 5144 21908 6532
rect 21964 5228 22004 7036
rect 22060 5900 22100 10984
rect 22348 10016 22388 17704
rect 22444 15560 22484 18460
rect 22636 18332 22676 18341
rect 22540 17072 22580 17081
rect 22540 16937 22580 17032
rect 22636 16232 22676 18292
rect 22828 17828 22868 19804
rect 23020 19760 23060 19769
rect 23060 19720 23252 19760
rect 23020 19711 23060 19720
rect 23116 19340 23156 19349
rect 22924 19256 22964 19265
rect 22924 18752 22964 19216
rect 23020 18752 23060 18761
rect 22924 18712 23020 18752
rect 23020 18684 23060 18712
rect 22732 17492 22772 17501
rect 22732 17324 22772 17452
rect 22732 17275 22772 17284
rect 22828 16904 22868 17788
rect 22924 18248 22964 18257
rect 22924 17408 22964 18208
rect 23020 18248 23060 18257
rect 23020 18164 23060 18208
rect 23020 18113 23060 18124
rect 23116 17828 23156 19300
rect 23212 18920 23252 19720
rect 23308 19592 23348 21400
rect 23308 19543 23348 19552
rect 23404 20516 23444 20525
rect 23404 19256 23444 20476
rect 23500 20348 23540 23584
rect 23596 20768 23636 26608
rect 23884 26396 23924 28600
rect 23884 26347 23924 26356
rect 24076 26816 24116 26825
rect 24076 25976 24116 26776
rect 24556 26648 24596 26657
rect 23788 25892 23828 25901
rect 23692 25388 23732 25397
rect 23692 22532 23732 25348
rect 23788 25052 23828 25852
rect 23788 25003 23828 25012
rect 23884 25640 23924 25649
rect 23788 24800 23828 24809
rect 23788 24296 23828 24760
rect 23884 24632 23924 25600
rect 23884 24583 23924 24592
rect 23980 25556 24020 25565
rect 23980 25472 24020 25516
rect 23980 24548 24020 25432
rect 23980 24499 24020 24508
rect 23788 24247 23828 24256
rect 23692 21776 23732 22492
rect 23788 24128 23828 24137
rect 23788 22280 23828 24088
rect 23980 24044 24020 24053
rect 23980 23876 24020 24004
rect 23980 23827 24020 23836
rect 23788 22028 23828 22240
rect 23788 21979 23828 21988
rect 23980 23708 24020 23717
rect 23692 21727 23732 21736
rect 23980 21020 24020 23668
rect 23980 20971 24020 20980
rect 23596 20728 23924 20768
rect 23500 20299 23540 20308
rect 23596 20600 23636 20609
rect 23596 20096 23636 20560
rect 23596 20047 23636 20056
rect 23404 19207 23444 19216
rect 23212 18871 23252 18880
rect 23404 18920 23444 18929
rect 23212 18668 23252 18677
rect 23212 18248 23252 18628
rect 23212 18199 23252 18208
rect 23116 17779 23156 17788
rect 23308 17828 23348 17837
rect 23404 17828 23444 18880
rect 23788 18668 23828 18677
rect 23692 18628 23788 18668
rect 23596 18584 23636 18595
rect 23500 18500 23540 18509
rect 23500 17996 23540 18460
rect 23596 18500 23636 18544
rect 23596 18080 23636 18460
rect 23596 18031 23636 18040
rect 23500 17947 23540 17956
rect 23596 17828 23636 17837
rect 23404 17788 23540 17828
rect 23020 17660 23060 17669
rect 23020 17492 23060 17620
rect 23020 17443 23060 17452
rect 23116 17660 23156 17669
rect 22924 17359 22964 17368
rect 23020 17156 23060 17165
rect 23020 17072 23060 17116
rect 23020 17021 23060 17032
rect 22828 16855 22868 16864
rect 22924 16988 22964 16997
rect 22924 16853 22964 16948
rect 23116 16988 23156 17620
rect 23212 17576 23252 17587
rect 23212 17492 23252 17536
rect 23212 17443 23252 17452
rect 23308 17324 23348 17788
rect 23116 16939 23156 16948
rect 23212 17284 23348 17324
rect 23404 17660 23444 17669
rect 23020 16904 23060 16913
rect 22636 16192 22868 16232
rect 22732 16064 22772 16073
rect 22732 15644 22772 16024
rect 22732 15595 22772 15604
rect 22444 15511 22484 15520
rect 22540 14048 22580 14057
rect 22540 13376 22580 14008
rect 22540 13327 22580 13336
rect 22636 13964 22676 13973
rect 22636 13796 22676 13924
rect 22636 13292 22676 13756
rect 22636 13243 22676 13252
rect 22444 13208 22484 13217
rect 22444 12704 22484 13168
rect 22444 12655 22484 12664
rect 22828 13124 22868 16192
rect 23020 15728 23060 16864
rect 23212 16232 23252 17284
rect 23308 17156 23348 17165
rect 23308 17072 23348 17116
rect 23404 17072 23444 17620
rect 23500 17240 23540 17788
rect 23596 17576 23636 17788
rect 23596 17527 23636 17536
rect 23692 17324 23732 18628
rect 23788 18619 23828 18628
rect 23884 18248 23924 20728
rect 24076 20684 24116 25936
rect 24364 26144 24404 26153
rect 24172 24800 24212 24809
rect 24172 24548 24212 24760
rect 24172 24499 24212 24508
rect 24268 24716 24308 24725
rect 24172 23876 24212 23887
rect 24172 23792 24212 23836
rect 24172 23743 24212 23752
rect 24268 22532 24308 24676
rect 24364 24716 24404 26104
rect 24364 24667 24404 24676
rect 24460 24632 24500 24641
rect 24460 24497 24500 24592
rect 24460 24044 24500 24053
rect 24364 23960 24404 23969
rect 24364 23825 24404 23920
rect 24460 23876 24500 24004
rect 24460 23827 24500 23836
rect 24364 23708 24404 23717
rect 24364 23624 24404 23668
rect 24364 23573 24404 23584
rect 24460 23540 24500 23549
rect 24364 23372 24404 23381
rect 24364 23036 24404 23332
rect 24364 22987 24404 22996
rect 24268 22483 24308 22492
rect 24364 22196 24404 22205
rect 24364 21944 24404 22156
rect 24172 21524 24212 21533
rect 24172 20852 24212 21484
rect 24364 21524 24404 21904
rect 24460 22112 24500 23500
rect 24556 23204 24596 26608
rect 24652 24884 24692 28600
rect 25228 27992 25268 28001
rect 24940 27572 24980 27581
rect 24652 24835 24692 24844
rect 24748 26732 24788 26741
rect 24748 23876 24788 26692
rect 24844 26144 24884 26153
rect 24844 26060 24884 26104
rect 24844 26009 24884 26020
rect 24844 24716 24884 24811
rect 24844 24667 24884 24676
rect 24748 23827 24788 23836
rect 24844 24548 24884 24557
rect 24556 23155 24596 23164
rect 24748 23456 24788 23465
rect 24652 23036 24692 23131
rect 24652 22987 24692 22996
rect 24460 21608 24500 22072
rect 24460 21559 24500 21568
rect 24556 21776 24596 21785
rect 24364 21475 24404 21484
rect 24460 21356 24500 21365
rect 24172 20803 24212 20812
rect 24364 20936 24404 20945
rect 24172 20684 24212 20693
rect 24076 20644 24172 20684
rect 24172 20264 24212 20644
rect 24172 20215 24212 20224
rect 23980 19256 24020 19265
rect 23980 18752 24020 19216
rect 24364 19256 24404 20896
rect 24364 19207 24404 19216
rect 23980 18703 24020 18712
rect 24172 19088 24212 19097
rect 24076 18668 24116 18677
rect 23980 18584 24020 18593
rect 23980 18449 24020 18544
rect 23884 18208 24020 18248
rect 23500 17200 23636 17240
rect 23500 17072 23540 17081
rect 23308 17032 23500 17072
rect 23500 17023 23540 17032
rect 23596 16820 23636 17200
rect 23692 17156 23732 17284
rect 23692 17107 23732 17116
rect 23788 18164 23828 18173
rect 23596 16771 23636 16780
rect 23788 16484 23828 18124
rect 23884 18080 23924 18089
rect 23884 17660 23924 18040
rect 23884 17611 23924 17620
rect 23884 17492 23924 17501
rect 23884 17324 23924 17452
rect 23884 17275 23924 17284
rect 23884 17156 23924 17167
rect 23884 17072 23924 17116
rect 23884 17023 23924 17032
rect 23788 16435 23828 16444
rect 23308 16232 23348 16241
rect 23212 16192 23308 16232
rect 23308 16183 23348 16192
rect 23788 16232 23828 16243
rect 23980 16232 24020 18208
rect 24076 17996 24116 18628
rect 24076 17947 24116 17956
rect 24076 17828 24116 17837
rect 24076 16316 24116 17788
rect 24076 16267 24116 16276
rect 23020 15679 23060 15688
rect 23116 16148 23156 16157
rect 23116 14972 23156 16108
rect 23116 14923 23156 14932
rect 23404 16148 23444 16157
rect 23404 16064 23444 16108
rect 23788 16148 23828 16192
rect 23116 14636 23156 14645
rect 23020 14468 23060 14477
rect 23020 14048 23060 14428
rect 23116 14300 23156 14596
rect 23116 14251 23156 14260
rect 23308 14552 23348 14561
rect 23020 13913 23060 14008
rect 22636 12452 22676 12461
rect 22636 11696 22676 12412
rect 22828 12452 22868 13084
rect 23212 13208 23252 13217
rect 23116 13040 23156 13049
rect 22828 12403 22868 12412
rect 22924 12620 22964 12629
rect 22636 11647 22676 11656
rect 22924 11108 22964 12580
rect 23116 12536 23156 13000
rect 23116 12487 23156 12496
rect 23116 11780 23156 11791
rect 23116 11696 23156 11740
rect 23116 11647 23156 11656
rect 23020 11108 23060 11117
rect 22924 11068 23020 11108
rect 22540 11024 22580 11033
rect 22540 10772 22580 10984
rect 22540 10268 22580 10732
rect 22540 10219 22580 10228
rect 22732 10352 22772 10361
rect 22732 10217 22772 10312
rect 22348 9967 22388 9976
rect 22444 10184 22484 10193
rect 22444 9512 22484 10144
rect 22636 10016 22676 10025
rect 22636 9596 22676 9976
rect 22636 9547 22676 9556
rect 22444 9463 22484 9472
rect 22828 8840 22868 8849
rect 22732 8756 22772 8765
rect 22156 8504 22196 8513
rect 22156 8084 22196 8464
rect 22156 7160 22196 8044
rect 22348 7328 22388 7337
rect 22156 7111 22196 7120
rect 22252 7244 22292 7253
rect 22156 6992 22196 7001
rect 22156 6572 22196 6952
rect 22156 6523 22196 6532
rect 22252 6656 22292 7204
rect 22252 6068 22292 6616
rect 22348 7076 22388 7288
rect 22732 7328 22772 8716
rect 22828 8000 22868 8800
rect 22924 8672 22964 11068
rect 23020 11040 23060 11068
rect 23212 11024 23252 13168
rect 23212 10975 23252 10984
rect 23308 12956 23348 14512
rect 23116 10184 23156 10193
rect 23116 9764 23156 10144
rect 23116 9715 23156 9724
rect 23212 9512 23252 9521
rect 23020 9428 23060 9437
rect 23020 8924 23060 9388
rect 23212 9377 23252 9472
rect 23020 8875 23060 8884
rect 22924 8168 22964 8632
rect 23308 8168 23348 12916
rect 23404 11612 23444 16024
rect 23596 16064 23636 16073
rect 23596 14720 23636 16024
rect 23596 14048 23636 14680
rect 23692 14972 23732 14981
rect 23692 14216 23732 14932
rect 23788 14804 23828 16108
rect 23884 16192 24020 16232
rect 23884 15056 23924 16192
rect 24172 16148 24212 19048
rect 24364 18584 24404 18593
rect 24268 18332 24308 18341
rect 24268 17828 24308 18292
rect 24364 18248 24404 18544
rect 24364 17912 24404 18208
rect 24364 17863 24404 17872
rect 24268 17779 24308 17788
rect 24364 17744 24404 17753
rect 24268 17576 24308 17585
rect 24268 17240 24308 17536
rect 24364 17576 24404 17704
rect 24364 17527 24404 17536
rect 24268 17191 24308 17200
rect 24364 17072 24404 17083
rect 24364 16988 24404 17032
rect 24364 16939 24404 16948
rect 23884 15007 23924 15016
rect 24076 15476 24116 15485
rect 23788 14755 23828 14764
rect 23788 14636 23828 14645
rect 23788 14501 23828 14596
rect 23692 14167 23732 14176
rect 23596 13999 23636 14008
rect 23884 13628 23924 13637
rect 23500 13460 23540 13469
rect 23500 11696 23540 13420
rect 23884 13208 23924 13588
rect 24076 13376 24116 15436
rect 24076 13327 24116 13336
rect 23884 12452 23924 13168
rect 23884 12403 23924 12412
rect 24076 12872 24116 12881
rect 24076 11948 24116 12832
rect 24076 11899 24116 11908
rect 23500 11647 23540 11656
rect 24172 11864 24212 16108
rect 24268 16232 24308 16241
rect 24268 16097 24308 16192
rect 24268 15728 24308 15737
rect 24268 14972 24308 15688
rect 24268 14923 24308 14932
rect 24268 14048 24308 14057
rect 24268 13376 24308 14008
rect 24364 13964 24404 13973
rect 24364 13460 24404 13924
rect 24364 13411 24404 13420
rect 24268 13327 24308 13336
rect 24172 11696 24212 11824
rect 24460 11864 24500 21316
rect 24556 21020 24596 21736
rect 24556 20971 24596 20980
rect 24652 21692 24692 21701
rect 24652 20096 24692 21652
rect 24748 20180 24788 23416
rect 24844 21608 24884 24508
rect 24844 21272 24884 21568
rect 24844 21223 24884 21232
rect 24748 20131 24788 20140
rect 24652 20047 24692 20056
rect 24844 20096 24884 20105
rect 24748 20012 24788 20021
rect 24556 19340 24596 19349
rect 24556 18416 24596 19300
rect 24556 18367 24596 18376
rect 24652 17744 24692 17753
rect 24652 17576 24692 17704
rect 24652 17527 24692 17536
rect 24748 16904 24788 19972
rect 24844 19256 24884 20056
rect 24844 19207 24884 19216
rect 24844 19088 24884 19097
rect 24844 18953 24884 19048
rect 24940 18920 24980 27532
rect 25036 26984 25076 26993
rect 25036 26144 25076 26944
rect 25228 26228 25268 27952
rect 25420 27824 25460 28600
rect 25420 27775 25460 27784
rect 25516 28496 25556 28505
rect 25516 26312 25556 28456
rect 25900 27404 25940 27413
rect 25900 26816 25940 27364
rect 25516 26263 25556 26272
rect 25804 26648 25844 26657
rect 25228 26179 25268 26188
rect 25420 26228 25460 26237
rect 25036 26095 25076 26104
rect 25324 26060 25364 26069
rect 25132 25976 25172 25985
rect 25036 24212 25076 24221
rect 25036 23204 25076 24172
rect 25036 23155 25076 23164
rect 25132 23120 25172 25936
rect 25036 23036 25076 23045
rect 25036 22280 25076 22996
rect 25132 22985 25172 23080
rect 25228 25472 25268 25481
rect 25228 23876 25268 25432
rect 25324 24800 25364 26020
rect 25420 25556 25460 26188
rect 25612 26144 25652 26153
rect 25420 25516 25556 25556
rect 25420 25388 25460 25397
rect 25420 25304 25460 25348
rect 25420 25253 25460 25264
rect 25420 25136 25460 25147
rect 25420 25052 25460 25096
rect 25420 25003 25460 25012
rect 25516 25136 25556 25516
rect 25324 24751 25364 24760
rect 25516 24716 25556 25096
rect 25516 24667 25556 24676
rect 25420 24632 25460 24641
rect 25324 24296 25364 24305
rect 25324 23960 25364 24256
rect 25420 24044 25460 24592
rect 25420 23995 25460 24004
rect 25324 23911 25364 23920
rect 25516 23960 25556 23969
rect 25036 21524 25076 22240
rect 25132 22196 25172 22205
rect 25132 22061 25172 22156
rect 25132 21944 25172 21953
rect 25132 21692 25172 21904
rect 25132 21643 25172 21652
rect 25132 21524 25172 21533
rect 25076 21484 25132 21524
rect 25036 21389 25076 21484
rect 25132 21475 25172 21484
rect 25132 20684 25172 20693
rect 25132 20096 25172 20644
rect 25132 20047 25172 20056
rect 25132 19928 25172 19937
rect 24940 18880 25076 18920
rect 24940 18752 24980 18761
rect 24844 18500 24884 18509
rect 24844 17996 24884 18460
rect 24940 18500 24980 18712
rect 24940 18451 24980 18460
rect 24844 17947 24884 17956
rect 24748 16855 24788 16864
rect 24844 17156 24884 17165
rect 24652 16232 24692 16241
rect 24652 15308 24692 16192
rect 24652 14720 24692 15268
rect 24844 16232 24884 17116
rect 24940 17072 24980 17081
rect 24940 16937 24980 17032
rect 24844 16203 24980 16232
rect 24844 16192 24940 16203
rect 24844 15644 24884 16192
rect 24940 16154 24980 16163
rect 24748 15224 24788 15233
rect 24748 14804 24788 15184
rect 24748 14755 24788 14764
rect 24844 14888 24884 15604
rect 24652 14671 24692 14680
rect 24652 14468 24692 14477
rect 24652 13964 24692 14428
rect 24652 13915 24692 13924
rect 24652 13796 24692 13805
rect 24500 11824 24596 11864
rect 24460 11815 24500 11824
rect 24172 11647 24212 11656
rect 23404 11563 23444 11572
rect 24268 11444 24308 11453
rect 23404 11192 23444 11201
rect 23404 9680 23444 11152
rect 23596 11024 23636 11033
rect 23404 9631 23444 9640
rect 23500 10184 23540 10193
rect 23500 9512 23540 10144
rect 23596 9680 23636 10984
rect 24076 11024 24116 11033
rect 23980 10940 24020 10949
rect 23980 10805 24020 10900
rect 23692 10520 23732 10529
rect 23692 9764 23732 10480
rect 23692 9715 23732 9724
rect 23788 10184 23828 10193
rect 23788 10016 23828 10144
rect 24076 10184 24116 10984
rect 24076 10135 24116 10144
rect 23596 9631 23636 9640
rect 23788 9596 23828 9976
rect 23788 9547 23828 9556
rect 23500 9463 23540 9472
rect 23308 8128 23444 8168
rect 22924 8119 22964 8128
rect 22828 7951 22868 7960
rect 23308 8000 23348 8009
rect 22732 7279 22772 7288
rect 23212 7160 23252 7169
rect 22348 6488 22388 7036
rect 23020 7076 23060 7085
rect 23020 6941 23060 7036
rect 23212 6908 23252 7120
rect 23212 6859 23252 6868
rect 23308 6656 23348 7960
rect 23404 7832 23444 8128
rect 23980 8084 24020 8093
rect 23404 7076 23444 7792
rect 23404 7027 23444 7036
rect 23596 8000 23636 8009
rect 23596 7244 23636 7960
rect 23788 8000 23828 8009
rect 23308 6607 23348 6616
rect 22348 6439 22388 6448
rect 23404 6572 23444 6581
rect 22252 6019 22292 6028
rect 22924 6236 22964 6245
rect 22060 5851 22100 5860
rect 22348 5900 22388 5909
rect 21964 5179 22004 5188
rect 21868 5095 21908 5104
rect 21388 4927 21428 4936
rect 21772 4976 21812 4985
rect 21772 4808 21812 4936
rect 22348 4976 22388 5860
rect 22924 5060 22964 6196
rect 23404 5312 23444 6532
rect 23596 6488 23636 7204
rect 23596 5900 23636 6448
rect 23692 7916 23732 7925
rect 23692 7160 23732 7876
rect 23692 6488 23732 7120
rect 23692 6439 23732 6448
rect 23788 6404 23828 7960
rect 23980 6992 24020 8044
rect 24172 8084 24212 8095
rect 24172 8000 24212 8044
rect 24172 7951 24212 7960
rect 24268 7160 24308 11404
rect 24556 11108 24596 11824
rect 24652 11696 24692 13756
rect 24844 13040 24884 14848
rect 24940 14804 24980 14813
rect 24940 14669 24980 14764
rect 24844 12991 24884 13000
rect 24652 11647 24692 11656
rect 25036 11444 25076 18880
rect 25132 17240 25172 19888
rect 25132 17191 25172 17200
rect 25132 16988 25172 16997
rect 25132 16484 25172 16948
rect 25132 16435 25172 16444
rect 25132 16316 25172 16325
rect 25132 15728 25172 16276
rect 25132 15593 25172 15688
rect 25036 11395 25076 11404
rect 25132 14720 25172 14729
rect 25132 11780 25172 14680
rect 25228 14552 25268 23836
rect 25324 23792 25364 23801
rect 25324 23372 25364 23752
rect 25516 23792 25556 23920
rect 25516 23743 25556 23752
rect 25324 23323 25364 23332
rect 25420 23708 25460 23717
rect 25324 23120 25364 23129
rect 25324 22364 25364 23080
rect 25420 22952 25460 23668
rect 25516 23624 25556 23633
rect 25516 23120 25556 23584
rect 25612 23456 25652 26104
rect 25708 26144 25748 26153
rect 25708 25976 25748 26104
rect 25708 25927 25748 25936
rect 25708 25472 25748 25481
rect 25708 25337 25748 25432
rect 25708 25136 25748 25145
rect 25708 24716 25748 25096
rect 25708 24632 25748 24676
rect 25708 23876 25748 24592
rect 25804 24044 25844 26608
rect 25900 26060 25940 26776
rect 26188 26396 26228 28600
rect 26956 28076 26996 28600
rect 27724 28160 27764 28600
rect 27724 28111 27764 28120
rect 26956 28027 26996 28036
rect 27674 27992 28042 28001
rect 27674 27943 28042 27952
rect 26956 27908 26996 27917
rect 26860 27656 26900 27665
rect 26434 27236 26802 27245
rect 26434 27187 26802 27196
rect 26860 27068 26900 27616
rect 26956 27572 26996 27868
rect 26956 27523 26996 27532
rect 27340 27572 27380 27581
rect 27340 27437 27380 27532
rect 26860 27019 26900 27028
rect 27916 27404 27956 27413
rect 27052 26816 27092 26825
rect 26092 26356 26228 26396
rect 26284 26732 26324 26741
rect 25900 26011 25940 26020
rect 25996 26312 26036 26321
rect 25996 25388 26036 26272
rect 26092 25724 26132 26356
rect 26092 25675 26132 25684
rect 26188 26228 26228 26237
rect 25996 25339 26036 25348
rect 25804 23995 25844 24004
rect 25996 25052 26036 25061
rect 25996 24380 26036 25012
rect 26188 24884 26228 26188
rect 26284 25388 26324 26692
rect 26764 26144 26804 26153
rect 26380 26060 26420 26069
rect 26380 25925 26420 26020
rect 26764 26009 26804 26104
rect 26860 25976 26900 25985
rect 26434 25724 26802 25733
rect 26434 25675 26802 25684
rect 26284 25339 26324 25348
rect 26860 25388 26900 25936
rect 26956 25976 26996 25985
rect 26956 25472 26996 25936
rect 26956 25423 26996 25432
rect 26860 25339 26900 25348
rect 27052 25388 27092 26776
rect 27916 26816 27956 27364
rect 28492 27404 28532 28600
rect 29260 28580 29300 28600
rect 29260 28531 29300 28540
rect 30028 28580 30068 28600
rect 30028 28531 30068 28540
rect 29260 27740 29300 27749
rect 28492 27355 28532 27364
rect 29164 27404 29204 27413
rect 27916 26767 27956 26776
rect 28300 26648 28340 26657
rect 28204 26564 28244 26573
rect 27674 26480 28042 26489
rect 27674 26431 28042 26440
rect 27820 26312 27860 26321
rect 27820 26177 27860 26272
rect 27052 25339 27092 25348
rect 27340 26144 27380 26153
rect 27244 25304 27284 25313
rect 26380 25220 26420 25231
rect 26380 25136 26420 25180
rect 26668 25220 26708 25229
rect 26380 25087 26420 25096
rect 26476 25136 26516 25145
rect 26476 24968 26516 25096
rect 26188 24835 26228 24844
rect 26284 24928 26516 24968
rect 26092 24800 26132 24809
rect 26092 24665 26132 24760
rect 26188 24716 26228 24727
rect 26188 24632 26228 24676
rect 26188 24583 26228 24592
rect 25708 23836 25940 23876
rect 25804 23624 25844 23633
rect 25612 23416 25748 23456
rect 25516 23071 25556 23080
rect 25612 23120 25652 23129
rect 25516 22952 25556 22961
rect 25420 22912 25516 22952
rect 25324 22315 25364 22324
rect 25420 22280 25460 22289
rect 25420 21776 25460 22240
rect 25516 22196 25556 22912
rect 25516 22147 25556 22156
rect 25420 21727 25460 21736
rect 25612 21692 25652 23080
rect 25708 22532 25748 23416
rect 25708 22483 25748 22492
rect 25804 22364 25844 23584
rect 25804 22315 25844 22324
rect 25708 22280 25748 22289
rect 25708 22196 25748 22240
rect 25708 21860 25748 22156
rect 25708 21811 25748 21820
rect 25804 22196 25844 22205
rect 25652 21652 25748 21692
rect 25612 21643 25652 21652
rect 25420 21608 25460 21617
rect 25324 21356 25364 21365
rect 25324 20852 25364 21316
rect 25324 20803 25364 20812
rect 25324 20600 25364 20609
rect 25324 20096 25364 20560
rect 25324 14720 25364 20056
rect 25420 20264 25460 21568
rect 25708 20936 25748 21652
rect 25804 21020 25844 22156
rect 25804 20971 25844 20980
rect 25420 18752 25460 20224
rect 25612 20852 25652 20861
rect 25612 20600 25652 20812
rect 25708 20801 25748 20896
rect 25516 20096 25556 20107
rect 25516 20012 25556 20056
rect 25516 19963 25556 19972
rect 25420 17660 25460 18712
rect 25612 19256 25652 20560
rect 25612 18920 25652 19216
rect 25420 17611 25460 17620
rect 25516 18668 25556 18677
rect 25516 17744 25556 18628
rect 25612 18500 25652 18880
rect 25708 20516 25748 20525
rect 25708 18584 25748 20476
rect 25804 20012 25844 20021
rect 25804 19877 25844 19972
rect 25708 18535 25748 18544
rect 25804 19088 25844 19097
rect 25804 18668 25844 19048
rect 25612 18451 25652 18460
rect 25804 17996 25844 18628
rect 25804 17947 25844 17956
rect 25516 16316 25556 17704
rect 25708 17576 25748 17585
rect 25708 17072 25748 17536
rect 25420 16148 25460 16157
rect 25420 14804 25460 16108
rect 25516 15392 25556 16276
rect 25612 16988 25652 16997
rect 25612 16064 25652 16948
rect 25612 16015 25652 16024
rect 25708 15644 25748 17032
rect 25708 15560 25748 15604
rect 25708 15509 25748 15520
rect 25804 16988 25844 16997
rect 25804 16232 25844 16948
rect 25516 14972 25556 15352
rect 25516 14923 25556 14932
rect 25612 15476 25652 15485
rect 25420 14755 25460 14764
rect 25516 14804 25556 14813
rect 25324 14671 25364 14680
rect 25420 14636 25460 14645
rect 25516 14636 25556 14764
rect 25460 14596 25556 14636
rect 25228 14512 25364 14552
rect 24460 11024 24500 11033
rect 24460 10889 24500 10984
rect 24364 10856 24404 10865
rect 24364 10184 24404 10816
rect 24556 10856 24596 11068
rect 25036 11276 25076 11285
rect 24556 10807 24596 10816
rect 24844 11024 24884 11033
rect 24844 10856 24884 10984
rect 24844 10807 24884 10816
rect 25036 10436 25076 11236
rect 25132 11108 25172 11740
rect 25132 11059 25172 11068
rect 25228 13040 25268 13049
rect 25132 10856 25172 10865
rect 25132 10721 25172 10816
rect 25036 10387 25076 10396
rect 24364 10135 24404 10144
rect 24940 9596 24980 9605
rect 24652 8840 24692 8849
rect 24692 8800 24884 8840
rect 24652 8791 24692 8800
rect 24556 8672 24596 8681
rect 24364 8084 24404 8093
rect 24364 7748 24404 8044
rect 24364 7699 24404 7708
rect 24556 7748 24596 8632
rect 24844 8672 24884 8800
rect 24844 8623 24884 8632
rect 24652 8420 24692 8429
rect 24652 8084 24692 8380
rect 24652 8035 24692 8044
rect 24844 8252 24884 8261
rect 24844 7916 24884 8212
rect 24844 7867 24884 7876
rect 24940 7832 24980 9556
rect 25036 8000 25076 8011
rect 25036 7916 25076 7960
rect 25036 7867 25076 7876
rect 24940 7783 24980 7792
rect 24556 7699 24596 7708
rect 24268 7111 24308 7120
rect 23980 6656 24020 6952
rect 24460 7076 24500 7087
rect 24460 6992 24500 7036
rect 24460 6943 24500 6952
rect 25228 6992 25268 13000
rect 25324 9344 25364 14512
rect 25420 11780 25460 14596
rect 25612 13796 25652 15436
rect 25708 15392 25748 15401
rect 25708 14888 25748 15352
rect 25708 14839 25748 14848
rect 25708 14720 25748 14729
rect 25708 14468 25748 14680
rect 25708 14419 25748 14428
rect 25612 13747 25652 13756
rect 25708 14216 25748 14225
rect 25708 12536 25748 14176
rect 25708 12487 25748 12496
rect 25420 11731 25460 11740
rect 25516 11780 25556 11789
rect 25516 11360 25556 11740
rect 25324 9295 25364 9304
rect 25420 9512 25460 9521
rect 25420 8672 25460 9472
rect 25324 8084 25364 8093
rect 25324 8000 25364 8044
rect 25324 7949 25364 7960
rect 25420 7160 25460 8632
rect 25516 7244 25556 11320
rect 25612 11024 25652 11033
rect 25612 10889 25652 10984
rect 25804 9680 25844 16192
rect 25900 14300 25940 23836
rect 25900 14251 25940 14260
rect 25900 13124 25940 13133
rect 25900 12452 25940 13084
rect 25900 11612 25940 12412
rect 25900 11563 25940 11572
rect 25708 9512 25748 9521
rect 25804 9512 25844 9640
rect 25900 10268 25940 10277
rect 25900 9596 25940 10228
rect 25996 9680 26036 24340
rect 26092 24464 26132 24473
rect 26092 23120 26132 24424
rect 26284 24296 26324 24928
rect 26668 24800 26708 25180
rect 27052 25220 27092 25229
rect 27052 25085 27092 25180
rect 26956 25052 26996 25061
rect 26380 24632 26420 24643
rect 26380 24548 26420 24592
rect 26380 24499 26420 24508
rect 26668 24380 26708 24760
rect 26764 24968 26804 24977
rect 26764 24464 26804 24928
rect 26956 24716 26996 25012
rect 26956 24667 26996 24676
rect 26764 24415 26804 24424
rect 26860 24548 26900 24557
rect 26668 24331 26708 24340
rect 26284 23624 26324 24256
rect 26434 24212 26802 24221
rect 26434 24163 26802 24172
rect 26284 23575 26324 23584
rect 26476 23792 26516 23801
rect 26380 23540 26420 23549
rect 26092 23071 26132 23080
rect 26188 23204 26228 23213
rect 26092 22364 26132 22459
rect 26092 22315 26132 22324
rect 26092 22196 26132 22236
rect 26092 22112 26132 22156
rect 26092 21608 26132 22072
rect 26092 21559 26132 21568
rect 26092 20768 26132 20777
rect 26092 19004 26132 20728
rect 26092 18955 26132 18964
rect 26092 18500 26132 18509
rect 26092 17744 26132 18460
rect 26092 17695 26132 17704
rect 26188 17240 26228 23164
rect 26380 23120 26420 23500
rect 26380 23036 26420 23080
rect 26284 22952 26324 22961
rect 26380 22956 26420 22996
rect 26284 22532 26324 22912
rect 26476 22868 26516 23752
rect 26668 23792 26708 23887
rect 26668 23743 26708 23752
rect 26764 23876 26804 23885
rect 26668 23624 26708 23633
rect 26668 23489 26708 23584
rect 26764 22868 26804 23836
rect 26860 23036 26900 24508
rect 27052 24548 27092 24557
rect 27052 24413 27092 24508
rect 26956 24380 26996 24389
rect 26956 23204 26996 24340
rect 27244 23960 27284 25264
rect 27340 25136 27380 26104
rect 28108 25976 28148 25985
rect 28108 25841 28148 25936
rect 27340 25087 27380 25096
rect 27436 25388 27476 25397
rect 27340 24548 27380 24557
rect 27340 24044 27380 24508
rect 27340 23995 27380 24004
rect 27244 23911 27284 23920
rect 26956 23155 26996 23164
rect 27052 23792 27092 23801
rect 26860 22987 26900 22996
rect 26956 22952 26996 22961
rect 26764 22828 26900 22868
rect 26476 22819 26516 22828
rect 26434 22700 26802 22709
rect 26434 22651 26802 22660
rect 26860 22616 26900 22828
rect 26860 22567 26900 22576
rect 26284 22483 26324 22492
rect 26668 22448 26708 22457
rect 26572 22408 26668 22448
rect 26380 22196 26420 22205
rect 26284 22112 26324 22121
rect 26284 19088 26324 22072
rect 26380 22061 26420 22156
rect 26572 21692 26612 22408
rect 26668 22399 26708 22408
rect 26572 21643 26612 21652
rect 26668 22196 26708 22205
rect 26668 21776 26708 22156
rect 26860 22196 26900 22205
rect 26860 22028 26900 22156
rect 26860 21944 26900 21988
rect 26860 21895 26900 21904
rect 26668 21356 26708 21736
rect 26668 21307 26708 21316
rect 26860 21776 26900 21785
rect 26434 21188 26802 21197
rect 26434 21139 26802 21148
rect 26476 21020 26516 21029
rect 26380 20768 26420 20777
rect 26380 19928 26420 20728
rect 26380 19879 26420 19888
rect 26476 19928 26516 20980
rect 26860 21020 26900 21736
rect 26860 20971 26900 20980
rect 26860 20852 26900 20863
rect 26860 20768 26900 20812
rect 26860 20719 26900 20728
rect 26572 20684 26612 20693
rect 26572 20549 26612 20644
rect 26860 20600 26900 20609
rect 26764 20516 26804 20525
rect 26572 20264 26612 20359
rect 26668 20348 26708 20443
rect 26668 20299 26708 20308
rect 26572 20215 26612 20224
rect 26668 20180 26708 20189
rect 26476 19879 26516 19888
rect 26572 20096 26612 20105
rect 26572 19844 26612 20056
rect 26668 19928 26708 20140
rect 26764 20180 26804 20476
rect 26860 20465 26900 20560
rect 26764 20131 26804 20140
rect 26860 20096 26900 20105
rect 26860 19961 26900 20056
rect 26956 20012 26996 22912
rect 26956 19963 26996 19972
rect 26668 19879 26708 19888
rect 26572 19795 26612 19804
rect 26860 19760 26900 19769
rect 26434 19676 26802 19685
rect 26434 19627 26802 19636
rect 26860 19508 26900 19720
rect 26764 19468 26900 19508
rect 26572 19340 26612 19349
rect 26284 18668 26324 19048
rect 26284 18619 26324 18628
rect 26380 19256 26420 19265
rect 26380 18584 26420 19216
rect 26572 19205 26612 19300
rect 26380 18535 26420 18544
rect 26476 18668 26516 18677
rect 26476 18533 26516 18628
rect 26764 18584 26804 19468
rect 27052 18584 27092 23752
rect 27340 23708 27380 23717
rect 27148 23204 27188 23213
rect 27148 23069 27188 23164
rect 27244 23036 27284 23131
rect 27244 22987 27284 22996
rect 27148 22952 27188 22961
rect 27148 22784 27188 22912
rect 27148 22735 27188 22744
rect 27244 22868 27284 22877
rect 27148 21860 27188 21869
rect 27148 20348 27188 21820
rect 27244 21608 27284 22828
rect 27244 21524 27284 21568
rect 27244 21475 27284 21484
rect 27244 20684 27284 20693
rect 27340 20684 27380 23668
rect 27436 23624 27476 25348
rect 27628 25388 27668 25397
rect 27628 25253 27668 25348
rect 28108 25220 28148 25229
rect 27674 24968 28042 24977
rect 27674 24919 28042 24928
rect 28108 24968 28148 25180
rect 28108 24919 28148 24928
rect 28012 24800 28052 24809
rect 27820 24760 28012 24800
rect 27436 23575 27476 23584
rect 27532 24716 27572 24725
rect 27436 23120 27476 23129
rect 27436 22985 27476 23080
rect 27436 22112 27476 22121
rect 27436 21692 27476 22072
rect 27436 21643 27476 21652
rect 27532 21608 27572 24676
rect 27820 24632 27860 24760
rect 28012 24751 28052 24760
rect 27820 24583 27860 24592
rect 27628 24296 27668 24305
rect 27628 24161 27668 24256
rect 28204 23792 28244 26524
rect 28300 25052 28340 26608
rect 29164 26648 29204 27364
rect 29164 26599 29204 26608
rect 28780 26228 28820 26237
rect 28300 24917 28340 25012
rect 28588 25220 28628 25229
rect 28492 24800 28532 24809
rect 28204 23743 28244 23752
rect 28300 24716 28340 24725
rect 27628 23708 27668 23717
rect 27628 23573 27668 23668
rect 27724 23624 27764 23719
rect 27724 23575 27764 23584
rect 27674 23456 28042 23465
rect 27674 23407 28042 23416
rect 27820 23288 27860 23297
rect 27628 23036 27668 23047
rect 27628 22952 27668 22996
rect 27628 22903 27668 22912
rect 27724 23036 27764 23045
rect 27628 22784 27668 22793
rect 27628 22649 27668 22744
rect 27724 22532 27764 22996
rect 27724 22483 27764 22492
rect 27820 23036 27860 23248
rect 27724 22280 27764 22289
rect 27820 22280 27860 22996
rect 28204 23036 28244 23045
rect 27764 22240 27860 22280
rect 27916 22868 27956 22877
rect 27916 22280 27956 22828
rect 27724 22231 27764 22240
rect 27916 22231 27956 22240
rect 28108 22700 28148 22709
rect 27674 21944 28042 21953
rect 27674 21895 28042 21904
rect 28108 21776 28148 22660
rect 28204 22280 28244 22996
rect 28204 22231 28244 22240
rect 28012 21736 28108 21776
rect 27916 21692 27956 21701
rect 27628 21608 27668 21617
rect 27532 21568 27628 21608
rect 27628 21559 27668 21568
rect 27916 21608 27956 21652
rect 27916 21557 27956 21568
rect 27532 21440 27572 21449
rect 27284 20644 27476 20684
rect 27244 20635 27284 20644
rect 27148 20299 27188 20308
rect 27244 20516 27284 20525
rect 27244 20348 27284 20476
rect 27244 20299 27284 20308
rect 27340 20264 27380 20273
rect 27244 20012 27284 20021
rect 27148 19928 27188 19937
rect 27148 19424 27188 19888
rect 27148 19375 27188 19384
rect 26764 18416 26804 18544
rect 26764 18367 26804 18376
rect 26860 18544 27092 18584
rect 27148 19256 27188 19265
rect 26284 18248 26324 18257
rect 26284 17660 26324 18208
rect 26434 18164 26802 18173
rect 26434 18115 26802 18124
rect 26284 17611 26324 17620
rect 26572 17492 26612 17501
rect 26764 17492 26804 17501
rect 26612 17452 26764 17492
rect 26572 17443 26612 17452
rect 26764 17443 26804 17452
rect 26092 17200 26228 17240
rect 26092 15392 26132 17200
rect 26188 17072 26228 17081
rect 26188 16148 26228 17032
rect 26284 16988 26324 16997
rect 26284 16853 26324 16948
rect 26284 16736 26324 16745
rect 26284 16316 26324 16696
rect 26434 16652 26802 16661
rect 26434 16603 26802 16612
rect 26284 16232 26324 16276
rect 26284 16181 26324 16192
rect 26668 16232 26708 16243
rect 26188 15560 26228 16108
rect 26668 16148 26708 16192
rect 26668 16099 26708 16108
rect 26764 16148 26804 16159
rect 26764 16064 26804 16108
rect 26764 16015 26804 16024
rect 26188 15511 26228 15520
rect 26092 15343 26132 15352
rect 26188 15392 26228 15401
rect 26092 14552 26132 14561
rect 26092 13292 26132 14512
rect 26188 13964 26228 15352
rect 26188 13915 26228 13924
rect 26284 15224 26324 15233
rect 26284 14804 26324 15184
rect 26434 15140 26802 15149
rect 26434 15091 26802 15100
rect 26092 13243 26132 13252
rect 26188 13796 26228 13805
rect 26188 12452 26228 13756
rect 26284 13292 26324 14764
rect 26764 14804 26804 14813
rect 26764 14636 26804 14764
rect 26764 14587 26804 14596
rect 26476 14552 26516 14561
rect 26476 13796 26516 14512
rect 26476 13747 26516 13756
rect 26434 13628 26802 13637
rect 26434 13579 26802 13588
rect 26284 12620 26324 13252
rect 26572 13208 26612 13217
rect 26572 13073 26612 13168
rect 26284 12571 26324 12580
rect 26188 12403 26228 12412
rect 26434 12116 26802 12125
rect 26860 12116 26900 18544
rect 26956 18416 26996 18425
rect 26956 17240 26996 18376
rect 26956 17191 26996 17200
rect 27052 17072 27092 17081
rect 27052 16904 27092 17032
rect 26956 16652 26996 16661
rect 26956 16232 26996 16612
rect 27052 16400 27092 16864
rect 27052 16351 27092 16360
rect 26956 16183 26996 16192
rect 27052 16064 27092 16073
rect 26956 15644 26996 15653
rect 26956 15509 26996 15604
rect 26956 15392 26996 15401
rect 26956 14804 26996 15352
rect 26956 14636 26996 14764
rect 27052 14804 27092 16024
rect 27148 15980 27188 19216
rect 27148 15931 27188 15940
rect 27052 14755 27092 14764
rect 27148 15644 27188 15653
rect 26956 14587 26996 14596
rect 26956 14468 26996 14477
rect 26956 13040 26996 14428
rect 27148 14048 27188 15604
rect 27148 13292 27188 14008
rect 27148 13243 27188 13252
rect 26996 13000 27092 13040
rect 26956 12991 26996 13000
rect 26956 12116 26996 12125
rect 26860 12076 26956 12116
rect 26434 12067 26802 12076
rect 26956 12067 26996 12076
rect 26668 11780 26708 11789
rect 26476 11696 26516 11705
rect 26476 11561 26516 11656
rect 26380 11528 26420 11537
rect 26380 11108 26420 11488
rect 26668 11192 26708 11740
rect 26668 11143 26708 11152
rect 26380 11059 26420 11068
rect 26284 10940 26324 10949
rect 26284 10805 26324 10900
rect 26860 10856 26900 10865
rect 25996 9631 26036 9640
rect 26092 10772 26132 10781
rect 26092 10352 26132 10732
rect 26434 10604 26802 10613
rect 26434 10555 26802 10564
rect 25900 9547 25940 9556
rect 25748 9472 25844 9512
rect 25996 9512 26036 9521
rect 26092 9512 26132 10312
rect 26764 10268 26804 10277
rect 26764 10016 26804 10228
rect 26764 9967 26804 9976
rect 26036 9472 26132 9512
rect 26284 9596 26324 9605
rect 25612 8756 25652 8765
rect 25708 8756 25748 9472
rect 25996 9463 26036 9472
rect 26284 9461 26324 9556
rect 26284 9344 26324 9353
rect 25652 8716 25748 8756
rect 25996 8756 26036 8765
rect 25612 8707 25652 8716
rect 25516 7195 25556 7204
rect 25420 7111 25460 7120
rect 25996 7160 26036 8716
rect 26092 8504 26132 8513
rect 26092 8084 26132 8464
rect 26092 8035 26132 8044
rect 26188 8168 26228 8177
rect 26188 8000 26228 8128
rect 26188 7951 26228 7960
rect 26284 7244 26324 9304
rect 26860 9260 26900 10816
rect 26956 10268 26996 10279
rect 27052 10268 27092 13000
rect 27244 12536 27284 19972
rect 27340 18668 27380 20224
rect 27436 18752 27476 20644
rect 27532 20348 27572 21400
rect 27628 21356 27668 21365
rect 27628 20768 27668 21316
rect 27724 21104 27764 21113
rect 27724 21020 27764 21064
rect 27724 20969 27764 20980
rect 27916 21020 27956 21029
rect 27628 20719 27668 20728
rect 27916 20768 27956 20980
rect 27916 20719 27956 20728
rect 28012 20684 28052 21736
rect 28108 21727 28148 21736
rect 28012 20635 28052 20644
rect 28108 21608 28148 21617
rect 27674 20432 28042 20441
rect 27674 20383 28042 20392
rect 27532 20299 27572 20308
rect 27820 20264 27860 20273
rect 27436 18703 27476 18712
rect 27532 20096 27572 20105
rect 27340 18619 27380 18628
rect 27340 18500 27380 18509
rect 27340 17240 27380 18460
rect 27436 18500 27476 18509
rect 27436 18332 27476 18460
rect 27436 18283 27476 18292
rect 27340 16316 27380 17200
rect 27436 17156 27476 17165
rect 27436 16988 27476 17116
rect 27436 16400 27476 16948
rect 27532 16568 27572 20056
rect 27724 19928 27764 19937
rect 27628 19844 27668 19853
rect 27628 19709 27668 19804
rect 27724 19592 27764 19888
rect 27724 19543 27764 19552
rect 27820 19340 27860 20224
rect 27820 19291 27860 19300
rect 28012 20264 28052 20273
rect 27628 19088 27668 19183
rect 28012 19088 28052 20224
rect 28108 20180 28148 21568
rect 28204 21608 28244 21617
rect 28204 21020 28244 21568
rect 28204 20971 28244 20980
rect 28300 20852 28340 24676
rect 28396 24464 28436 24473
rect 28396 23204 28436 24424
rect 28396 23155 28436 23164
rect 28300 20803 28340 20812
rect 28396 23036 28436 23045
rect 28396 22364 28436 22996
rect 28108 20131 28148 20140
rect 28204 20684 28244 20693
rect 28108 20012 28148 20040
rect 28204 20012 28244 20644
rect 28148 19972 28244 20012
rect 28108 19963 28148 19972
rect 28204 19508 28244 19972
rect 28204 19459 28244 19468
rect 28300 20684 28340 20693
rect 28204 19340 28244 19349
rect 28012 19048 28148 19088
rect 27628 19039 27668 19048
rect 27674 18920 28042 18929
rect 27674 18871 28042 18880
rect 27628 18668 27668 18677
rect 27628 18164 27668 18628
rect 27628 18115 27668 18124
rect 27724 18416 27764 18425
rect 27724 17576 27764 18376
rect 28108 17996 28148 19048
rect 28108 17947 28148 17956
rect 27724 17527 27764 17536
rect 28108 17828 28148 17837
rect 27674 17408 28042 17417
rect 27674 17359 28042 17368
rect 28108 17324 28148 17788
rect 28108 17275 28148 17284
rect 27724 17156 27764 17165
rect 27724 17021 27764 17116
rect 28012 17072 28052 17081
rect 27532 16519 27572 16528
rect 27436 16360 27572 16400
rect 27340 16267 27380 16276
rect 27436 16232 27476 16241
rect 27436 15728 27476 16192
rect 27436 15679 27476 15688
rect 27340 15308 27380 15317
rect 27340 14720 27380 15268
rect 27532 15056 27572 16360
rect 28012 16064 28052 17032
rect 28204 16904 28244 19300
rect 28300 19088 28340 20644
rect 28300 19039 28340 19048
rect 28396 19256 28436 22324
rect 28492 20684 28532 24760
rect 28588 24128 28628 25180
rect 28684 24884 28724 24893
rect 28684 24548 28724 24844
rect 28684 24499 28724 24508
rect 28588 24079 28628 24088
rect 28780 23288 28820 26188
rect 28972 26060 29012 26069
rect 28972 25976 29012 26020
rect 28972 25925 29012 25936
rect 29164 26060 29204 26069
rect 29164 25925 29204 26020
rect 28876 25304 28916 25313
rect 28876 24800 28916 25264
rect 28876 24632 28916 24760
rect 28876 24583 28916 24592
rect 28972 24548 29012 24643
rect 28972 24499 29012 24508
rect 28972 24380 29012 24389
rect 28972 23876 29012 24340
rect 28972 23827 29012 23836
rect 28780 23239 28820 23248
rect 28876 23792 28916 23801
rect 28588 23204 28628 23213
rect 28588 23036 28628 23164
rect 28588 22987 28628 22996
rect 28492 20635 28532 20644
rect 28588 22364 28628 22373
rect 28300 18584 28340 18593
rect 28300 16988 28340 18544
rect 28396 18500 28436 19216
rect 28396 18451 28436 18460
rect 28492 19508 28532 19517
rect 28300 16939 28340 16948
rect 28396 17996 28436 18005
rect 28204 16855 28244 16864
rect 28012 16015 28052 16024
rect 28108 16820 28148 16829
rect 27674 15896 28042 15905
rect 27674 15847 28042 15856
rect 27724 15728 27764 15737
rect 27532 15007 27572 15016
rect 27628 15560 27668 15569
rect 27340 14671 27380 14680
rect 27436 14804 27476 14813
rect 27436 14048 27476 14764
rect 27628 14804 27668 15520
rect 27724 14888 27764 15688
rect 27724 14839 27764 14848
rect 28012 15560 28052 15569
rect 28012 15476 28052 15520
rect 28108 15560 28148 16780
rect 28204 16316 28244 16325
rect 28204 15812 28244 16276
rect 28204 15763 28244 15772
rect 28108 15511 28148 15520
rect 27628 14755 27668 14764
rect 28012 14636 28052 15436
rect 28012 14587 28052 14596
rect 27674 14384 28042 14393
rect 27674 14335 28042 14344
rect 27436 13999 27476 14008
rect 28204 14300 28244 14309
rect 27820 13964 27860 13973
rect 27820 13460 27860 13924
rect 27820 13411 27860 13420
rect 27674 12872 28042 12881
rect 27674 12823 28042 12832
rect 27244 12487 27284 12496
rect 27532 11864 27572 11873
rect 27340 11696 27380 11705
rect 27340 11192 27380 11656
rect 27340 11143 27380 11152
rect 27436 11528 27476 11537
rect 27436 10940 27476 11488
rect 27436 10891 27476 10900
rect 26956 10228 27052 10268
rect 26956 10184 26996 10228
rect 27052 10219 27092 10228
rect 27532 10352 27572 11824
rect 27916 11780 27956 11789
rect 27916 11696 27956 11740
rect 28204 11780 28244 14260
rect 28300 14048 28340 14057
rect 28300 12452 28340 14008
rect 28396 12788 28436 17956
rect 28396 12739 28436 12748
rect 28300 12403 28340 12412
rect 28396 12620 28436 12629
rect 28204 11731 28244 11740
rect 27916 11645 27956 11656
rect 28396 11696 28436 12580
rect 28492 11780 28532 19468
rect 28588 12956 28628 22324
rect 28684 22280 28724 22289
rect 28684 21608 28724 22240
rect 28684 21473 28724 21568
rect 28684 21104 28724 21113
rect 28684 20852 28724 21064
rect 28684 20803 28724 20812
rect 28588 12620 28628 12916
rect 28588 12571 28628 12580
rect 28684 20600 28724 20609
rect 28684 12452 28724 20560
rect 28876 20600 28916 23752
rect 29068 23792 29108 23801
rect 28972 23204 29012 23213
rect 28972 21692 29012 23164
rect 28972 21643 29012 21652
rect 28876 20551 28916 20560
rect 28972 20768 29012 20777
rect 28972 20264 29012 20728
rect 28972 20215 29012 20224
rect 28876 19424 28916 19433
rect 28876 18920 28916 19384
rect 28876 18871 28916 18880
rect 28780 18752 28820 18761
rect 28820 18712 28916 18740
rect 28780 18700 28916 18712
rect 28876 18668 28916 18700
rect 28876 18619 28916 18628
rect 29068 18500 29108 23752
rect 29260 23792 29300 27700
rect 29356 27656 29396 27665
rect 29356 26816 29396 27616
rect 30124 27656 30164 27665
rect 29356 26228 29396 26776
rect 29356 26179 29396 26188
rect 29644 27404 29684 27413
rect 29164 23120 29204 23129
rect 29164 22448 29204 23080
rect 29164 22399 29204 22408
rect 29260 22196 29300 23752
rect 29356 24632 29396 24641
rect 29356 22364 29396 24592
rect 29548 23708 29588 23717
rect 29548 23288 29588 23668
rect 29548 23239 29588 23248
rect 29548 23120 29588 23129
rect 29548 22952 29588 23080
rect 29548 22903 29588 22912
rect 29356 22324 29492 22364
rect 29452 22280 29492 22324
rect 29356 22196 29396 22205
rect 29260 22156 29356 22196
rect 29260 22028 29300 22037
rect 28876 18460 29108 18500
rect 29164 21524 29204 21533
rect 28876 14384 28916 18460
rect 28876 14335 28916 14344
rect 28972 18332 29012 18341
rect 28876 13964 28916 13973
rect 28876 13829 28916 13924
rect 28684 12403 28724 12412
rect 28492 11731 28532 11740
rect 28588 12284 28628 12293
rect 28396 11647 28436 11656
rect 27674 11360 28042 11369
rect 27674 11311 28042 11320
rect 27820 11024 27860 11033
rect 27820 10436 27860 10984
rect 28588 11024 28628 12244
rect 28876 12116 28916 12125
rect 28876 11612 28916 12076
rect 28876 11563 28916 11572
rect 28972 11276 29012 18292
rect 29164 16316 29204 21484
rect 29068 16276 29204 16316
rect 29068 11948 29108 16276
rect 29164 16148 29204 16157
rect 29164 14132 29204 16108
rect 29260 15140 29300 21988
rect 29356 21608 29396 22156
rect 29356 20852 29396 21568
rect 29356 20803 29396 20812
rect 29452 21776 29492 22240
rect 29452 20096 29492 21736
rect 29548 22028 29588 22037
rect 29548 21356 29588 21988
rect 29548 21307 29588 21316
rect 29452 19256 29492 20056
rect 29452 19207 29492 19216
rect 29548 20180 29588 20189
rect 29452 18836 29492 18845
rect 29452 16484 29492 18796
rect 29548 18584 29588 20140
rect 29644 19844 29684 27364
rect 30124 27068 30164 27616
rect 30124 27019 30164 27028
rect 30412 27656 30452 27665
rect 30124 26900 30164 26909
rect 30124 26765 30164 26860
rect 30028 26648 30068 26657
rect 29932 25304 29972 25313
rect 29836 25136 29876 25145
rect 29836 25001 29876 25096
rect 29836 24716 29876 24725
rect 29740 24548 29780 24557
rect 29740 24413 29780 24508
rect 29644 18836 29684 19804
rect 29644 18787 29684 18796
rect 29740 24296 29780 24305
rect 29548 18535 29588 18544
rect 29644 18668 29684 18677
rect 29644 17744 29684 18628
rect 29740 17996 29780 24256
rect 29836 18416 29876 24676
rect 29932 23624 29972 25264
rect 30028 25052 30068 26608
rect 30028 25003 30068 25012
rect 30124 26396 30164 26405
rect 30028 24800 30068 24809
rect 30028 24296 30068 24760
rect 30028 24247 30068 24256
rect 29932 23372 29972 23584
rect 29932 23323 29972 23332
rect 30028 23876 30068 23885
rect 29932 23204 29972 23213
rect 29932 20432 29972 23164
rect 29932 20348 29972 20392
rect 29932 20299 29972 20308
rect 29932 20180 29972 20189
rect 29932 18836 29972 20140
rect 29932 18787 29972 18796
rect 29836 18367 29876 18376
rect 29932 18668 29972 18677
rect 29740 17956 29876 17996
rect 29452 16444 29588 16484
rect 29260 15091 29300 15100
rect 29164 14048 29204 14092
rect 29164 13997 29204 14008
rect 29260 14972 29300 14981
rect 29260 12704 29300 14932
rect 29260 12655 29300 12664
rect 29356 14720 29396 14729
rect 29356 14132 29396 14680
rect 29356 13208 29396 14092
rect 29068 11899 29108 11908
rect 29260 11864 29300 11873
rect 29068 11780 29108 11789
rect 29068 11645 29108 11740
rect 29260 11729 29300 11824
rect 28972 11227 29012 11236
rect 28588 10975 28628 10984
rect 29260 11024 29300 11033
rect 29260 10889 29300 10984
rect 27820 10387 27860 10396
rect 26956 9932 26996 10144
rect 26956 9883 26996 9892
rect 27052 10100 27092 10109
rect 27052 9512 27092 10060
rect 27532 9680 27572 10312
rect 28492 10352 28532 10361
rect 28108 10016 28148 10025
rect 27674 9848 28042 9857
rect 27674 9799 28042 9808
rect 27532 9631 27572 9640
rect 26434 9092 26802 9101
rect 26434 9043 26802 9052
rect 26860 8924 26900 9220
rect 26764 8884 26900 8924
rect 26956 9428 26996 9437
rect 26764 7748 26804 8884
rect 26764 7699 26804 7708
rect 26860 8588 26900 8597
rect 26956 8588 26996 9388
rect 27052 9344 27092 9472
rect 27340 9596 27380 9605
rect 27052 9295 27092 9304
rect 27244 9428 27284 9437
rect 27148 8588 27188 8597
rect 26956 8548 27148 8588
rect 26434 7580 26802 7589
rect 26434 7531 26802 7540
rect 26380 7244 26420 7253
rect 26284 7204 26380 7244
rect 25996 7111 26036 7120
rect 26380 7160 26420 7204
rect 26860 7244 26900 8548
rect 26860 7195 26900 7204
rect 26380 7109 26420 7120
rect 27148 7076 27188 8548
rect 27244 7160 27284 9388
rect 27340 7244 27380 9556
rect 27532 9512 27572 9521
rect 27340 7195 27380 7204
rect 27436 8672 27476 8681
rect 27244 7111 27284 7120
rect 27148 7027 27188 7036
rect 27436 7076 27476 8632
rect 27436 7027 27476 7036
rect 25228 6943 25268 6952
rect 27532 6992 27572 9472
rect 28108 8672 28148 9976
rect 28492 9428 28532 10312
rect 28684 10016 28724 10025
rect 28684 9512 28724 9976
rect 28684 9463 28724 9472
rect 29356 9512 29396 13168
rect 29452 14384 29492 14393
rect 29452 13124 29492 14344
rect 29452 11780 29492 13084
rect 29548 12620 29588 16444
rect 29644 16232 29684 17704
rect 29740 17072 29780 17081
rect 29740 16937 29780 17032
rect 29644 16183 29684 16192
rect 29740 15308 29780 15317
rect 29644 14636 29684 14645
rect 29644 14216 29684 14596
rect 29644 14167 29684 14176
rect 29740 14132 29780 15268
rect 29740 14083 29780 14092
rect 29548 12571 29588 12580
rect 29644 14048 29684 14057
rect 29548 12452 29588 12461
rect 29548 11864 29588 12412
rect 29548 11815 29588 11824
rect 29452 11731 29492 11740
rect 29452 11192 29492 11201
rect 29452 11057 29492 11152
rect 29548 11108 29588 11117
rect 29548 10973 29588 11068
rect 29644 10940 29684 14008
rect 29740 13124 29780 13133
rect 29740 12989 29780 13084
rect 29740 12452 29780 12461
rect 29836 12452 29876 17956
rect 29932 17072 29972 18628
rect 30028 18668 30068 23836
rect 30124 23060 30164 26356
rect 30412 24968 30452 27616
rect 30604 27572 30644 27581
rect 30604 26312 30644 27532
rect 30796 27404 30836 28600
rect 30988 28160 31028 28169
rect 30796 27355 30836 27364
rect 30892 27572 30932 27581
rect 30604 26263 30644 26272
rect 30700 26732 30740 26741
rect 30412 24919 30452 24928
rect 30220 23876 30260 23885
rect 30220 23741 30260 23836
rect 30316 23120 30356 23129
rect 30124 23020 30260 23060
rect 30028 18619 30068 18628
rect 30124 22616 30164 22625
rect 30028 17660 30068 17669
rect 30028 17240 30068 17620
rect 30028 17191 30068 17200
rect 29932 17032 30068 17072
rect 29932 16904 29972 16913
rect 29932 16316 29972 16864
rect 29932 16267 29972 16276
rect 29932 15644 29972 15653
rect 29932 15509 29972 15604
rect 29780 12412 29876 12452
rect 29932 15392 29972 15401
rect 29740 12403 29780 12412
rect 29836 12284 29876 12293
rect 29836 11192 29876 12244
rect 29932 11948 29972 15352
rect 30028 14048 30068 17032
rect 30124 14972 30164 22576
rect 30220 18332 30260 23020
rect 30316 21104 30356 23080
rect 30412 22364 30452 22373
rect 30412 22229 30452 22324
rect 30316 21055 30356 21064
rect 30412 21524 30452 21533
rect 30316 19592 30356 19601
rect 30316 18752 30356 19552
rect 30316 18703 30356 18712
rect 30220 18283 30260 18292
rect 30316 18500 30356 18509
rect 30220 17996 30260 18005
rect 30220 17072 30260 17956
rect 30220 17023 30260 17032
rect 30124 14923 30164 14932
rect 30220 16400 30260 16409
rect 30220 14804 30260 16360
rect 30316 15392 30356 18460
rect 30412 17492 30452 21484
rect 30508 20768 30548 20777
rect 30508 19508 30548 20728
rect 30508 19004 30548 19468
rect 30508 18955 30548 18964
rect 30604 19340 30644 19349
rect 30412 17443 30452 17452
rect 30508 18836 30548 18845
rect 30508 17324 30548 18796
rect 30316 15343 30356 15352
rect 30412 17284 30548 17324
rect 30220 14755 30260 14764
rect 30028 13999 30068 14008
rect 30124 14132 30164 14141
rect 30124 13997 30164 14092
rect 30316 12788 30356 12797
rect 29932 11528 29972 11908
rect 29932 11479 29972 11488
rect 30124 12452 30164 12461
rect 30124 11360 30164 12412
rect 30316 11864 30356 12748
rect 30316 11815 30356 11824
rect 30412 11780 30452 17284
rect 30508 16148 30548 16157
rect 30508 12200 30548 16108
rect 30604 13376 30644 19300
rect 30700 18668 30740 26692
rect 30892 25892 30932 27532
rect 30892 25843 30932 25852
rect 30700 18619 30740 18628
rect 30796 24884 30836 24893
rect 30796 20768 30836 24844
rect 30988 23060 31028 28120
rect 31084 26648 31124 26657
rect 31084 24380 31124 26608
rect 31084 24331 31124 24340
rect 31468 24968 31508 24977
rect 31180 23624 31220 23633
rect 31180 23372 31220 23584
rect 30700 17744 30740 17753
rect 30700 17609 30740 17704
rect 30796 16148 30836 20728
rect 30892 23020 31028 23060
rect 31084 23120 31124 23129
rect 30892 17660 30932 23020
rect 30988 21356 31028 21365
rect 31084 21356 31124 23080
rect 31028 21316 31124 21356
rect 30988 18836 31028 21316
rect 31180 19424 31220 23332
rect 31276 22868 31316 22877
rect 31276 22364 31316 22828
rect 31276 22315 31316 22324
rect 31372 20012 31412 20021
rect 31180 19384 31316 19424
rect 30988 18787 31028 18796
rect 31084 19088 31124 19097
rect 30892 17611 30932 17620
rect 30988 17828 31028 17837
rect 30796 16099 30836 16108
rect 30892 17492 30932 17501
rect 30700 15980 30740 15989
rect 30700 15476 30740 15940
rect 30700 15427 30740 15436
rect 30700 14972 30740 14981
rect 30700 14837 30740 14932
rect 30604 13327 30644 13336
rect 30700 12368 30740 12377
rect 30700 12233 30740 12328
rect 30508 12151 30548 12160
rect 30700 11948 30740 11957
rect 30700 11813 30740 11908
rect 30892 11864 30932 17452
rect 30988 16904 31028 17788
rect 30988 16855 31028 16864
rect 31084 16316 31124 19048
rect 31084 16267 31124 16276
rect 31180 15476 31220 15485
rect 30988 14888 31028 14897
rect 30988 14753 31028 14848
rect 31084 13964 31124 13973
rect 31084 13829 31124 13924
rect 31180 13208 31220 15436
rect 31276 13292 31316 19384
rect 31276 13243 31316 13252
rect 31180 13159 31220 13168
rect 31372 12452 31412 19972
rect 31372 12403 31412 12412
rect 30892 11815 30932 11824
rect 30412 11731 30452 11740
rect 31468 11612 31508 24928
rect 31660 20684 31700 20693
rect 31660 12536 31700 20644
rect 31660 12487 31700 12496
rect 31756 17156 31796 17165
rect 31756 16232 31796 17116
rect 31756 11696 31796 16192
rect 31756 11647 31796 11656
rect 31468 11563 31508 11572
rect 30124 11311 30164 11320
rect 29836 11143 29876 11152
rect 30124 11192 30164 11201
rect 30124 11057 30164 11152
rect 29644 10891 29684 10900
rect 29836 10940 29876 10949
rect 29836 10805 29876 10900
rect 30412 10856 30452 10865
rect 30412 10721 30452 10816
rect 30796 10856 30836 10865
rect 30796 10721 30836 10816
rect 30412 10604 30452 10613
rect 30412 10352 30452 10564
rect 30412 10303 30452 10312
rect 30796 10352 30836 10361
rect 30796 10217 30836 10312
rect 29356 9463 29396 9472
rect 28492 9379 28532 9388
rect 27674 8336 28042 8345
rect 27674 8287 28042 8296
rect 28108 8168 28148 8632
rect 28108 8119 28148 8128
rect 27532 6943 27572 6952
rect 27674 6824 28042 6833
rect 27674 6775 28042 6784
rect 23980 6607 24020 6616
rect 23788 6355 23828 6364
rect 24076 6488 24116 6497
rect 24076 6353 24116 6448
rect 24460 6488 24500 6497
rect 23596 5851 23636 5860
rect 23404 5263 23444 5272
rect 22924 5011 22964 5020
rect 22348 4927 22388 4936
rect 24460 4892 24500 6448
rect 26434 6068 26802 6077
rect 26434 6019 26802 6028
rect 27674 5312 28042 5321
rect 27674 5263 28042 5272
rect 24460 4843 24500 4852
rect 21772 4759 21812 4768
rect 20812 4591 20852 4600
rect 18660 4556 19028 4565
rect 18660 4507 19028 4516
rect 26434 4556 26802 4565
rect 26434 4507 26802 4516
rect 17164 4255 17204 4264
rect 16684 4003 16724 4012
rect 4352 3800 4720 3809
rect 4352 3751 4720 3760
rect 12126 3800 12494 3809
rect 12126 3751 12494 3760
rect 19900 3800 20268 3809
rect 19900 3751 20268 3760
rect 27674 3800 28042 3809
rect 27674 3751 28042 3760
rect 3112 3044 3480 3053
rect 3112 2995 3480 3004
rect 10886 3044 11254 3053
rect 10886 2995 11254 3004
rect 18660 3044 19028 3053
rect 18660 2995 19028 3004
rect 26434 3044 26802 3053
rect 26434 2995 26802 3004
rect 4352 2288 4720 2297
rect 4352 2239 4720 2248
rect 12126 2288 12494 2297
rect 12126 2239 12494 2248
rect 19900 2288 20268 2297
rect 19900 2239 20268 2248
rect 27674 2288 28042 2297
rect 27674 2239 28042 2248
rect 3112 1532 3480 1541
rect 3112 1483 3480 1492
rect 10886 1532 11254 1541
rect 10886 1483 11254 1492
rect 18660 1532 19028 1541
rect 18660 1483 19028 1492
rect 26434 1532 26802 1541
rect 26434 1483 26802 1492
rect 4352 776 4720 785
rect 4352 727 4720 736
rect 12126 776 12494 785
rect 12126 727 12494 736
rect 19900 776 20268 785
rect 19900 727 20268 736
rect 27674 776 28042 785
rect 27674 727 28042 736
<< via3 >>
rect 1516 28120 1556 28160
rect 1900 27532 1940 27572
rect 2380 27448 2420 27488
rect 3148 27784 3188 27824
rect 3628 27784 3668 27824
rect 3112 27196 3480 27236
rect 2956 26356 2996 26396
rect 2860 26104 2900 26144
rect 556 25180 596 25220
rect 172 23248 212 23288
rect 76 22492 116 22532
rect 460 22492 500 22532
rect 460 21652 500 21692
rect 556 21988 596 22028
rect 364 20560 404 20600
rect 460 20308 500 20348
rect 364 14764 404 14804
rect 652 20476 692 20516
rect 748 23332 788 23372
rect 940 23164 980 23204
rect 844 22744 884 22784
rect 844 22576 884 22616
rect 556 14764 596 14804
rect 460 13756 500 13796
rect 748 14428 788 14468
rect 1036 20476 1076 20516
rect 940 18712 980 18752
rect 1900 25936 1940 25976
rect 1612 25432 1652 25472
rect 1708 24760 1748 24800
rect 1996 24592 2036 24632
rect 1420 23248 1460 23288
rect 1804 22156 1844 22196
rect 1324 21064 1364 21104
rect 1228 20560 1268 20600
rect 1228 18712 1268 18752
rect 1420 20812 1460 20852
rect 1708 21820 1748 21860
rect 1420 19804 1460 19844
rect 1036 13756 1076 13796
rect 2380 24508 2420 24548
rect 2284 22240 2324 22280
rect 1996 21820 2036 21860
rect 1900 21568 1940 21608
rect 2860 25768 2900 25808
rect 2572 25348 2612 25388
rect 3244 26860 3284 26900
rect 3532 25936 3572 25976
rect 3112 25684 3480 25724
rect 3244 25432 3284 25472
rect 3112 24172 3480 24212
rect 2476 23752 2516 23792
rect 2188 20728 2228 20768
rect 2380 20644 2420 20684
rect 1708 18544 1748 18584
rect 1804 17872 1844 17912
rect 1708 16528 1748 16568
rect 2764 22912 2804 22952
rect 2956 22912 2996 22952
rect 3436 22912 3476 22952
rect 3112 22660 3480 22700
rect 2668 22408 2708 22448
rect 2668 22156 2708 22196
rect 2572 21316 2612 21356
rect 2668 21400 2708 21440
rect 2572 19804 2612 19844
rect 2572 19636 2612 19676
rect 2188 18040 2228 18080
rect 1420 14428 1460 14468
rect 940 10900 980 10940
rect 1324 10984 1364 11024
rect 3052 21484 3092 21524
rect 3244 21400 3284 21440
rect 3532 21484 3572 21524
rect 2860 20644 2900 20684
rect 3112 21148 3480 21188
rect 3340 20980 3380 21020
rect 2764 20056 2804 20096
rect 2764 19636 2804 19676
rect 2860 19552 2900 19592
rect 3112 19636 3480 19676
rect 3052 19468 3092 19508
rect 4684 28120 4724 28160
rect 4352 27952 4720 27992
rect 4396 26860 4436 26900
rect 4588 26692 4628 26732
rect 4684 26608 4724 26648
rect 4352 26440 4720 26480
rect 5548 26776 5588 26816
rect 5164 26356 5204 26396
rect 3724 25768 3764 25808
rect 4204 25348 4244 25388
rect 4012 23500 4052 23540
rect 4352 24928 4720 24968
rect 4352 23416 4720 23456
rect 4396 23164 4436 23204
rect 3820 22912 3860 22952
rect 3724 22240 3764 22280
rect 3724 21232 3764 21272
rect 4396 22744 4436 22784
rect 3916 22408 3956 22448
rect 4300 22492 4340 22532
rect 3916 21568 3956 21608
rect 4492 22408 4532 22448
rect 5164 25264 5204 25304
rect 5356 25264 5396 25304
rect 5260 23752 5300 23792
rect 5068 23164 5108 23204
rect 6892 27448 6932 27488
rect 6892 26608 6932 26648
rect 6508 25264 6548 25304
rect 7180 26692 7220 26732
rect 7372 26608 7412 26648
rect 8524 27532 8564 27572
rect 8332 26104 8372 26144
rect 6220 24760 6260 24800
rect 5260 22744 5300 22784
rect 5164 22492 5204 22532
rect 4012 21232 4052 21272
rect 4108 21484 4148 21524
rect 4012 20812 4052 20852
rect 3112 18124 3480 18164
rect 3148 17956 3188 17996
rect 2572 17704 2612 17744
rect 2284 17284 2324 17324
rect 3244 17032 3284 17072
rect 3112 16612 3480 16652
rect 2956 15520 2996 15560
rect 3820 19216 3860 19256
rect 3820 17704 3860 17744
rect 3628 17116 3668 17156
rect 3724 15688 3764 15728
rect 3628 15520 3668 15560
rect 3112 15100 3480 15140
rect 3112 13588 3480 13628
rect 2572 12748 2612 12788
rect 2668 11656 2708 11696
rect 3436 13168 3476 13208
rect 3112 12076 3480 12116
rect 2668 10984 2708 11024
rect 3112 10564 3480 10604
rect 3436 9976 3476 10016
rect 3628 9976 3668 10016
rect 460 5944 500 5984
rect 3112 9052 3480 9092
rect 3340 8800 3380 8840
rect 4876 22156 4916 22196
rect 4352 21904 4720 21944
rect 4204 20728 4244 20768
rect 4396 20980 4436 21020
rect 4780 21484 4820 21524
rect 4492 20896 4532 20936
rect 4588 21316 4628 21356
rect 4352 20392 4720 20432
rect 4588 20224 4628 20264
rect 4300 19972 4340 20012
rect 4684 20056 4724 20096
rect 4300 19216 4340 19256
rect 4352 18880 4720 18920
rect 4972 20728 5012 20768
rect 4876 20224 4916 20264
rect 5452 22408 5492 22448
rect 5452 22240 5492 22280
rect 5548 22072 5588 22112
rect 5740 22156 5780 22196
rect 5644 21988 5684 22028
rect 6124 22156 6164 22196
rect 6028 21736 6068 21776
rect 5548 21568 5588 21608
rect 5548 20812 5588 20852
rect 5452 20392 5492 20432
rect 5356 20056 5396 20096
rect 5932 21484 5972 21524
rect 5740 20140 5780 20180
rect 4204 17872 4244 17912
rect 4396 17788 4436 17828
rect 4204 17704 4244 17744
rect 4972 18544 5012 18584
rect 4684 17536 4724 17576
rect 4352 17368 4720 17408
rect 4108 17116 4148 17156
rect 4492 17200 4532 17240
rect 4492 16864 4532 16904
rect 4108 16276 4148 16316
rect 4684 16024 4724 16064
rect 4352 15856 4720 15896
rect 4012 15520 4052 15560
rect 4492 15604 4532 15644
rect 4108 15436 4148 15476
rect 4588 15436 4628 15476
rect 5068 17788 5108 17828
rect 4972 17032 5012 17072
rect 5068 17368 5108 17408
rect 4876 16024 4916 16064
rect 5356 19132 5396 19172
rect 5356 17956 5396 17996
rect 5260 16948 5300 16988
rect 5452 17200 5492 17240
rect 5740 17200 5780 17240
rect 5356 15856 5396 15896
rect 5260 14932 5300 14972
rect 4492 14596 4532 14636
rect 4588 14512 4628 14552
rect 4352 14344 4720 14384
rect 3916 12496 3956 12536
rect 3628 8800 3668 8840
rect 3112 7540 3480 7580
rect 3112 6028 3480 6068
rect 4780 13252 4820 13292
rect 5740 16864 5780 16904
rect 6028 20056 6068 20096
rect 6412 22240 6452 22280
rect 6316 20224 6356 20264
rect 6604 21568 6644 21608
rect 6796 23164 6836 23204
rect 6796 21484 6836 21524
rect 6700 21316 6740 21356
rect 6412 20056 6452 20096
rect 6700 20224 6740 20264
rect 6508 19972 6548 20012
rect 6892 19972 6932 20012
rect 6124 19216 6164 19256
rect 6124 18880 6164 18920
rect 6508 19132 6548 19172
rect 6892 19216 6932 19256
rect 7084 20560 7124 20600
rect 7180 21484 7220 21524
rect 7852 22912 7892 22952
rect 7948 22828 7988 22868
rect 7468 22324 7508 22364
rect 7660 22240 7700 22280
rect 7660 21820 7700 21860
rect 7276 20728 7316 20768
rect 7276 20392 7316 20432
rect 6892 18880 6932 18920
rect 5932 16948 5972 16988
rect 5740 15688 5780 15728
rect 4352 12832 4720 12872
rect 4352 11320 4720 11360
rect 4780 11152 4820 11192
rect 4204 10984 4244 11024
rect 4352 9808 4720 9848
rect 4352 8296 4720 8336
rect 3916 5608 3956 5648
rect 4352 6784 4720 6824
rect 5740 15520 5780 15560
rect 5932 16108 5972 16148
rect 6028 16612 6068 16652
rect 6220 17788 6260 17828
rect 6412 17536 6452 17576
rect 6220 17200 6260 17240
rect 6220 16444 6260 16484
rect 6412 15100 6452 15140
rect 6508 15856 6548 15896
rect 7084 18544 7124 18584
rect 6796 18124 6836 18164
rect 6796 16528 6836 16568
rect 6700 16360 6740 16400
rect 6700 15940 6740 15980
rect 6796 15772 6836 15812
rect 6988 16528 7028 16568
rect 6412 14176 6452 14216
rect 5356 12748 5396 12788
rect 5452 12580 5492 12620
rect 5836 12580 5876 12620
rect 6220 13252 6260 13292
rect 4972 9976 5012 10016
rect 6028 11656 6068 11696
rect 5932 9472 5972 9512
rect 4780 5608 4820 5648
rect 4352 5272 4720 5312
rect 6604 12496 6644 12536
rect 6796 15352 6836 15392
rect 7276 17620 7316 17660
rect 7180 17116 7220 17156
rect 7852 22744 7892 22784
rect 8620 25264 8660 25304
rect 8524 25180 8564 25220
rect 8332 23668 8372 23708
rect 8236 23584 8276 23624
rect 8044 20980 8084 21020
rect 7852 20644 7892 20684
rect 7756 20308 7796 20348
rect 7852 19804 7892 19844
rect 7468 17284 7508 17324
rect 7756 18460 7796 18500
rect 7852 18376 7892 18416
rect 7660 16612 7700 16652
rect 6700 14512 6740 14552
rect 6796 15100 6836 15140
rect 6892 13840 6932 13880
rect 6412 11656 6452 11696
rect 6412 10900 6452 10940
rect 7660 15352 7700 15392
rect 7468 15016 7508 15056
rect 7852 17536 7892 17576
rect 7852 17200 7892 17240
rect 7852 16948 7892 16988
rect 7852 16780 7892 16820
rect 7852 16360 7892 16400
rect 7852 16108 7892 16148
rect 8044 20392 8084 20432
rect 8236 22072 8276 22112
rect 8236 20896 8276 20936
rect 8236 20224 8276 20264
rect 8044 17368 8084 17408
rect 8236 18544 8276 18584
rect 8716 24508 8756 24548
rect 10060 27700 10100 27740
rect 8428 22828 8468 22868
rect 8524 22492 8564 22532
rect 8428 22408 8468 22448
rect 8812 23584 8852 23624
rect 10060 25600 10100 25640
rect 9196 23752 9236 23792
rect 9292 24592 9332 24632
rect 8620 22324 8660 22364
rect 8524 21820 8564 21860
rect 8428 21568 8468 21608
rect 8524 20812 8564 20852
rect 8620 20728 8660 20768
rect 8524 18796 8564 18836
rect 8908 22912 8948 22952
rect 8812 22576 8852 22616
rect 9004 22156 9044 22196
rect 8908 21988 8948 22028
rect 8812 21064 8852 21104
rect 8812 20896 8852 20936
rect 8236 17116 8276 17156
rect 8044 16696 8084 16736
rect 8044 16360 8084 16400
rect 8044 15940 8084 15980
rect 7948 15436 7988 15476
rect 8044 14680 8084 14720
rect 7372 11908 7412 11948
rect 7756 13084 7796 13124
rect 7852 13168 7892 13208
rect 8428 16780 8468 16820
rect 8428 16360 8468 16400
rect 8428 16108 8468 16148
rect 8332 14680 8372 14720
rect 8236 14596 8276 14636
rect 8716 18040 8756 18080
rect 8620 17620 8660 17660
rect 9196 23332 9236 23372
rect 9388 23332 9428 23372
rect 9196 21988 9236 22028
rect 9196 21820 9236 21860
rect 9004 20812 9044 20852
rect 9196 20644 9236 20684
rect 9292 21736 9332 21776
rect 9196 20224 9236 20264
rect 8908 19804 8948 19844
rect 9004 19216 9044 19256
rect 8908 18880 8948 18920
rect 9196 18796 9236 18836
rect 8812 17032 8852 17072
rect 8620 15520 8660 15560
rect 8428 13840 8468 13880
rect 8620 14008 8660 14048
rect 7756 12580 7796 12620
rect 7276 11152 7316 11192
rect 8812 13756 8852 13796
rect 8812 13588 8852 13628
rect 8716 13168 8756 13208
rect 7468 10984 7508 11024
rect 7564 11908 7604 11948
rect 6220 5608 6260 5648
rect 3112 4516 3480 4556
rect 9388 21484 9428 21524
rect 9388 19216 9428 19256
rect 9196 18208 9236 18248
rect 9100 17872 9140 17912
rect 9196 17536 9236 17576
rect 9196 17200 9236 17240
rect 9100 16780 9140 16820
rect 9100 15856 9140 15896
rect 9196 16276 9236 16316
rect 9580 21736 9620 21776
rect 10060 24340 10100 24380
rect 10444 27112 10484 27152
rect 10252 24424 10292 24464
rect 10060 23584 10100 23624
rect 10060 23416 10100 23456
rect 10060 22828 10100 22868
rect 10252 23164 10292 23204
rect 10828 27364 10868 27404
rect 10886 27196 11254 27236
rect 11212 27028 11252 27068
rect 10924 26860 10964 26900
rect 10886 25684 11254 25724
rect 10540 23836 10580 23876
rect 10444 23500 10484 23540
rect 10828 25264 10868 25304
rect 12364 28120 12404 28160
rect 13036 28120 13076 28160
rect 12126 27952 12494 27992
rect 12172 27616 12212 27656
rect 11596 26776 11636 26816
rect 11596 26188 11636 26228
rect 11980 26776 12020 26816
rect 11884 26356 11924 26396
rect 11692 25180 11732 25220
rect 10886 24172 11254 24212
rect 11020 23668 11060 23708
rect 11116 23164 11156 23204
rect 10348 23080 10388 23120
rect 10444 22744 10484 22784
rect 10156 22240 10196 22280
rect 10060 22072 10100 22112
rect 9964 21820 10004 21860
rect 10156 21484 10196 21524
rect 10348 21988 10388 22028
rect 9868 20980 9908 21020
rect 10060 21148 10100 21188
rect 10348 21568 10388 21608
rect 10444 21484 10484 21524
rect 9580 18124 9620 18164
rect 9484 18040 9524 18080
rect 9676 17872 9716 17912
rect 9484 17116 9524 17156
rect 9484 16276 9524 16316
rect 9388 16192 9428 16232
rect 9292 15772 9332 15812
rect 9868 16696 9908 16736
rect 9100 15436 9140 15476
rect 9196 13756 9236 13796
rect 9004 13588 9044 13628
rect 9196 13084 9236 13124
rect 9196 12580 9236 12620
rect 8908 11740 8948 11780
rect 9388 13252 9428 13292
rect 9964 16360 10004 16400
rect 9676 14176 9716 14216
rect 10060 15688 10100 15728
rect 10348 18712 10388 18752
rect 10252 17872 10292 17912
rect 10252 16360 10292 16400
rect 10886 22660 11254 22700
rect 10924 21736 10964 21776
rect 10732 21568 10772 21608
rect 11788 23332 11828 23372
rect 11788 22996 11828 23036
rect 12172 26776 12212 26816
rect 12460 26608 12500 26648
rect 12126 26440 12494 26480
rect 12460 26020 12500 26060
rect 12460 25348 12500 25388
rect 12172 25264 12212 25304
rect 12844 26524 12884 26564
rect 12126 24928 12494 24968
rect 12172 23752 12212 23792
rect 13324 26944 13364 26984
rect 13420 26860 13460 26900
rect 13132 26440 13172 26480
rect 13324 26776 13364 26816
rect 13132 26188 13172 26228
rect 12844 24340 12884 24380
rect 12126 23416 12494 23456
rect 12556 23332 12596 23372
rect 12076 23080 12116 23120
rect 12172 22744 12212 22784
rect 12364 22072 12404 22112
rect 12126 21904 12494 21944
rect 11884 21484 11924 21524
rect 10636 21148 10676 21188
rect 10886 21148 11254 21188
rect 10886 19636 11254 19676
rect 13516 26692 13556 26732
rect 13708 26776 13748 26816
rect 13804 26608 13844 26648
rect 13036 24424 13076 24464
rect 13420 25180 13460 25220
rect 13516 25264 13556 25304
rect 13516 24676 13556 24716
rect 13708 25180 13748 25220
rect 13228 23584 13268 23624
rect 12652 22072 12692 22112
rect 12748 21988 12788 22028
rect 12652 21568 12692 21608
rect 11500 20140 11540 20180
rect 10540 17956 10580 17996
rect 10444 17116 10484 17156
rect 11404 18544 11444 18584
rect 10886 18124 11254 18164
rect 10828 17872 10868 17912
rect 10540 17200 10580 17240
rect 10636 17536 10676 17576
rect 11116 17032 11156 17072
rect 11596 19132 11636 19172
rect 10636 16696 10676 16736
rect 10886 16612 11254 16652
rect 11404 17956 11444 17996
rect 11596 17620 11636 17660
rect 10828 16108 10868 16148
rect 10732 15520 10772 15560
rect 10348 15352 10388 15392
rect 10444 15268 10484 15308
rect 10252 13924 10292 13964
rect 10060 13672 10100 13712
rect 9868 12412 9908 12452
rect 9964 12496 10004 12536
rect 10060 11908 10100 11948
rect 11404 15856 11444 15896
rect 11020 15772 11060 15812
rect 11404 15520 11444 15560
rect 11116 15436 11156 15476
rect 10828 15268 10868 15308
rect 10886 15100 11254 15140
rect 10540 14596 10580 14636
rect 11116 14932 11156 14972
rect 10924 14680 10964 14720
rect 10540 14176 10580 14216
rect 10252 11824 10292 11864
rect 10348 12328 10388 12368
rect 9388 8380 9428 8420
rect 9676 8380 9716 8420
rect 10540 11824 10580 11864
rect 11020 14092 11060 14132
rect 11596 15856 11636 15896
rect 11020 13840 11060 13880
rect 11308 13840 11348 13880
rect 10886 13588 11254 13628
rect 10924 13084 10964 13124
rect 11116 12580 11156 12620
rect 11404 13168 11444 13208
rect 11404 12580 11444 12620
rect 10886 12076 11254 12116
rect 11308 11824 11348 11864
rect 11212 11656 11252 11696
rect 10886 10564 11254 10604
rect 10828 10228 10868 10268
rect 10444 8800 10484 8840
rect 10060 7708 10100 7748
rect 10886 9052 11254 9092
rect 10828 8800 10868 8840
rect 12126 20392 12494 20432
rect 13324 22828 13364 22868
rect 12940 21148 12980 21188
rect 11884 17200 11924 17240
rect 11884 17032 11924 17072
rect 12126 18880 12494 18920
rect 12652 18964 12692 19004
rect 12940 18796 12980 18836
rect 12652 18292 12692 18332
rect 12364 17956 12404 17996
rect 12126 17368 12494 17408
rect 12076 16192 12116 16232
rect 12126 15856 12494 15896
rect 11884 15268 11924 15308
rect 12172 15436 12212 15476
rect 12364 15352 12404 15392
rect 12268 15184 12308 15224
rect 11788 14512 11828 14552
rect 11884 14260 11924 14300
rect 12460 15604 12500 15644
rect 12172 14512 12212 14552
rect 12126 14344 12494 14384
rect 12268 14176 12308 14216
rect 12076 14008 12116 14048
rect 12844 18544 12884 18584
rect 12940 18208 12980 18248
rect 12844 17368 12884 17408
rect 12844 17200 12884 17240
rect 13132 19216 13172 19256
rect 13036 17200 13076 17240
rect 12748 16696 12788 16736
rect 12748 15772 12788 15812
rect 13612 23584 13652 23624
rect 13900 24760 13940 24800
rect 13804 23332 13844 23372
rect 15340 27616 15380 27656
rect 14284 26440 14324 26480
rect 14188 23836 14228 23876
rect 14188 22912 14228 22952
rect 13996 22240 14036 22280
rect 13516 21148 13556 21188
rect 12940 15520 12980 15560
rect 12844 15016 12884 15056
rect 12844 14512 12884 14552
rect 13228 15436 13268 15476
rect 13036 14596 13076 14636
rect 13132 15100 13172 15140
rect 12844 14092 12884 14132
rect 12844 13924 12884 13964
rect 12748 13756 12788 13796
rect 12556 13168 12596 13208
rect 12126 12832 12494 12872
rect 12172 12496 12212 12536
rect 11980 12244 12020 12284
rect 12076 11572 12116 11612
rect 12364 12244 12404 12284
rect 12364 11656 12404 11696
rect 12652 11992 12692 12032
rect 12126 11320 12494 11360
rect 13132 14008 13172 14048
rect 13324 14596 13364 14636
rect 13228 13756 13268 13796
rect 13036 12412 13076 12452
rect 12126 9808 12494 9848
rect 11692 8632 11732 8672
rect 12268 8632 12308 8672
rect 11212 8044 11252 8084
rect 13708 19972 13748 20012
rect 13900 20056 13940 20096
rect 14476 26020 14516 26060
rect 15052 27112 15092 27152
rect 14956 26944 14996 26984
rect 14764 25096 14804 25136
rect 14668 24844 14708 24884
rect 15340 25096 15380 25136
rect 15628 25348 15668 25388
rect 15436 24340 15476 24380
rect 16300 26524 16340 26564
rect 16204 25936 16244 25976
rect 19900 27952 20268 27992
rect 15436 24088 15476 24128
rect 15244 23164 15284 23204
rect 14188 22240 14228 22280
rect 14380 21736 14420 21776
rect 14188 21484 14228 21524
rect 14476 21568 14516 21608
rect 14860 21232 14900 21272
rect 14092 20980 14132 21020
rect 14860 20812 14900 20852
rect 14476 20476 14516 20516
rect 13516 17284 13556 17324
rect 14476 20140 14516 20180
rect 14476 19804 14516 19844
rect 14860 20056 14900 20096
rect 14764 19132 14804 19172
rect 14284 18880 14324 18920
rect 14188 18376 14228 18416
rect 14380 18208 14420 18248
rect 14572 18376 14612 18416
rect 14668 18292 14708 18332
rect 14476 17956 14516 17996
rect 14188 17872 14228 17912
rect 13708 16192 13748 16232
rect 13804 15436 13844 15476
rect 13900 15268 13940 15308
rect 13612 13924 13652 13964
rect 13516 11992 13556 12032
rect 13804 12916 13844 12956
rect 14092 16192 14132 16232
rect 13708 11656 13748 11696
rect 13612 11152 13652 11192
rect 14284 14596 14324 14636
rect 14284 14260 14324 14300
rect 14188 13504 14228 13544
rect 14572 17620 14612 17660
rect 14668 17536 14708 17576
rect 14764 17200 14804 17240
rect 14668 17116 14708 17156
rect 14668 16780 14708 16820
rect 14476 14008 14516 14048
rect 14572 14092 14612 14132
rect 14476 13840 14516 13880
rect 13900 12496 13940 12536
rect 14284 12664 14324 12704
rect 14476 12664 14516 12704
rect 14092 11824 14132 11864
rect 14572 12496 14612 12536
rect 13900 11152 13940 11192
rect 13996 9976 14036 10016
rect 12844 8632 12884 8672
rect 12126 8296 12494 8336
rect 10886 7540 11254 7580
rect 11116 7120 11156 7160
rect 10060 6112 10100 6152
rect 10886 6028 11254 6068
rect 12268 8044 12308 8084
rect 11596 6448 11636 6488
rect 10886 4516 11254 4556
rect 12076 7708 12116 7748
rect 11884 7120 11924 7160
rect 12126 6784 12494 6824
rect 12268 6448 12308 6488
rect 12126 5272 12494 5312
rect 13612 6448 13652 6488
rect 12652 5020 12692 5060
rect 15148 21316 15188 21356
rect 15244 21148 15284 21188
rect 15244 20308 15284 20348
rect 15148 19300 15188 19340
rect 15148 18964 15188 19004
rect 15148 17620 15188 17660
rect 15532 21484 15572 21524
rect 15532 19972 15572 20012
rect 15724 18544 15764 18584
rect 15532 18124 15572 18164
rect 15436 18040 15476 18080
rect 15436 17536 15476 17576
rect 15436 17116 15476 17156
rect 15244 15604 15284 15644
rect 15148 14932 15188 14972
rect 15052 14848 15092 14888
rect 15148 13756 15188 13796
rect 15148 13252 15188 13292
rect 15052 12496 15092 12536
rect 16108 24844 16148 24884
rect 16108 21736 16148 21776
rect 16012 21652 16052 21692
rect 15916 21316 15956 21356
rect 15916 20896 15956 20936
rect 16108 20812 16148 20852
rect 16012 19972 16052 20012
rect 15916 19804 15956 19844
rect 15820 18460 15860 18500
rect 15916 18124 15956 18164
rect 15628 17620 15668 17660
rect 15820 17872 15860 17912
rect 16204 19216 16244 19256
rect 16204 18460 16244 18500
rect 16684 23836 16724 23876
rect 16684 23248 16724 23288
rect 16876 23248 16916 23288
rect 16972 24676 17012 24716
rect 18660 27196 19028 27236
rect 17740 27028 17780 27068
rect 18220 26608 18260 26648
rect 17068 24340 17108 24380
rect 16684 20308 16724 20348
rect 16492 20056 16532 20096
rect 16588 18544 16628 18584
rect 15724 17032 15764 17072
rect 15628 16192 15668 16232
rect 15724 15520 15764 15560
rect 15724 14596 15764 14636
rect 15532 13504 15572 13544
rect 15436 12664 15476 12704
rect 15628 13336 15668 13376
rect 16012 15604 16052 15644
rect 16108 14848 16148 14888
rect 15916 14008 15956 14048
rect 15628 12664 15668 12704
rect 15436 12496 15476 12536
rect 15436 11824 15476 11864
rect 15820 11656 15860 11696
rect 16204 14680 16244 14720
rect 16492 14680 16532 14720
rect 16204 13756 16244 13796
rect 16300 13252 16340 13292
rect 16012 11908 16052 11948
rect 16108 11824 16148 11864
rect 16204 10816 16244 10856
rect 16492 12748 16532 12788
rect 16684 17368 16724 17408
rect 16972 20140 17012 20180
rect 17260 20812 17300 20852
rect 16972 17284 17012 17324
rect 16876 17116 16916 17156
rect 16588 10060 16628 10100
rect 16972 16276 17012 16316
rect 17260 16780 17300 16820
rect 17068 16192 17108 16232
rect 16972 15604 17012 15644
rect 17068 15268 17108 15308
rect 16876 14680 16916 14720
rect 16876 14260 16916 14300
rect 17260 15604 17300 15644
rect 16780 14092 16820 14132
rect 16972 14176 17012 14216
rect 16876 14008 16916 14048
rect 17068 13840 17108 13880
rect 17740 26524 17780 26564
rect 17452 25936 17492 25976
rect 17548 24760 17588 24800
rect 18028 26356 18068 26396
rect 17452 15688 17492 15728
rect 17452 15436 17492 15476
rect 17836 22912 17876 22952
rect 17644 15100 17684 15140
rect 17644 14932 17684 14972
rect 17452 13336 17492 13376
rect 17836 18796 17876 18836
rect 17836 18544 17876 18584
rect 17836 18208 17876 18248
rect 17836 17872 17876 17912
rect 17740 14848 17780 14888
rect 17740 14680 17780 14720
rect 17356 12580 17396 12620
rect 17644 12916 17684 12956
rect 18028 22996 18068 23036
rect 18220 23248 18260 23288
rect 18892 26524 18932 26564
rect 18412 26188 18452 26228
rect 18988 26440 19028 26480
rect 19276 26440 19316 26480
rect 18412 25768 18452 25808
rect 18660 25684 19028 25724
rect 18604 24508 18644 24548
rect 18660 24172 19028 24212
rect 19084 23080 19124 23120
rect 18660 22660 19028 22700
rect 18028 22240 18068 22280
rect 17932 15268 17972 15308
rect 18316 21568 18356 21608
rect 18124 17872 18164 17912
rect 18988 21568 19028 21608
rect 20332 26776 20372 26816
rect 20140 26608 20180 26648
rect 19900 26440 20268 26480
rect 20044 26188 20084 26228
rect 19660 25768 19700 25808
rect 19900 24928 20268 24968
rect 20812 26104 20852 26144
rect 20524 24760 20564 24800
rect 20332 24508 20372 24548
rect 18316 20476 18356 20516
rect 18660 21148 19028 21188
rect 18700 20980 18740 21020
rect 18604 20896 18644 20936
rect 18796 20308 18836 20348
rect 19084 20812 19124 20852
rect 19372 20812 19412 20852
rect 19180 20644 19220 20684
rect 19276 20056 19316 20096
rect 18700 19804 18740 19844
rect 19084 19804 19124 19844
rect 18316 18880 18356 18920
rect 18412 18712 18452 18752
rect 18660 19636 19028 19676
rect 18508 18544 18548 18584
rect 18988 18460 19028 18500
rect 18316 17620 18356 17660
rect 18316 17032 18356 17072
rect 18412 16864 18452 16904
rect 18220 15520 18260 15560
rect 18028 15100 18068 15140
rect 17836 12496 17876 12536
rect 17836 11656 17876 11696
rect 17644 10144 17684 10184
rect 17836 10228 17876 10268
rect 18316 13672 18356 13712
rect 18316 13084 18356 13124
rect 18660 18124 19028 18164
rect 18700 16864 18740 16904
rect 19372 19300 19412 19340
rect 19276 18712 19316 18752
rect 19372 17788 19412 17828
rect 19276 17620 19316 17660
rect 18892 17116 18932 17156
rect 18796 16780 18836 16820
rect 18660 16612 19028 16652
rect 18988 16360 19028 16400
rect 18508 16108 18548 16148
rect 19180 16612 19220 16652
rect 19084 16108 19124 16148
rect 19276 16108 19316 16148
rect 18660 15100 19028 15140
rect 18604 14932 18644 14972
rect 19372 15184 19412 15224
rect 19276 14596 19316 14636
rect 18508 13924 18548 13964
rect 18700 14008 18740 14048
rect 18660 13588 19028 13628
rect 19372 14176 19412 14216
rect 18316 12496 18356 12536
rect 18660 12076 19028 12116
rect 18508 11656 18548 11696
rect 19180 11656 19220 11696
rect 19276 11908 19316 11948
rect 18124 10144 18164 10184
rect 18316 10060 18356 10100
rect 18660 10564 19028 10604
rect 18508 9976 18548 10016
rect 18660 9052 19028 9092
rect 18508 8548 18548 8588
rect 18660 7540 19028 7580
rect 19564 20224 19604 20264
rect 20236 23836 20276 23876
rect 19900 23416 20268 23456
rect 20236 23248 20276 23288
rect 19900 21904 20268 21944
rect 19756 20644 19796 20684
rect 19900 20392 20268 20432
rect 20044 20224 20084 20264
rect 19564 17116 19604 17156
rect 20140 19300 20180 19340
rect 20908 22828 20948 22868
rect 19900 18880 20268 18920
rect 19564 16192 19604 16232
rect 19900 17368 20268 17408
rect 19948 17200 19988 17240
rect 19852 17116 19892 17156
rect 20140 16864 20180 16904
rect 19900 15856 20268 15896
rect 19756 15688 19796 15728
rect 19852 15604 19892 15644
rect 19948 15520 19988 15560
rect 19948 14680 19988 14720
rect 19900 14344 20268 14384
rect 19756 14260 19796 14300
rect 20140 14176 20180 14216
rect 20236 13924 20276 13964
rect 19468 12748 19508 12788
rect 19468 11740 19508 11780
rect 19660 13252 19700 13292
rect 19756 13504 19796 13544
rect 20524 14428 20564 14468
rect 19900 12832 20268 12872
rect 20140 12328 20180 12368
rect 20524 14260 20564 14300
rect 20524 13000 20564 13040
rect 20428 11572 20468 11612
rect 19900 11320 20268 11360
rect 20140 10816 20180 10856
rect 19900 9808 20268 9848
rect 19660 8548 19700 8588
rect 19948 8548 19988 8588
rect 19900 8296 20268 8336
rect 21292 18628 21332 18668
rect 21004 18292 21044 18332
rect 21484 25768 21524 25808
rect 22156 23836 22196 23876
rect 23116 26944 23156 26984
rect 23212 24592 23252 24632
rect 22636 22828 22676 22868
rect 23500 23836 23540 23876
rect 23404 22912 23444 22952
rect 22252 22324 22292 22364
rect 22828 22240 22868 22280
rect 22060 21484 22100 21524
rect 23116 22324 23156 22364
rect 23212 22240 23252 22280
rect 21676 18544 21716 18584
rect 21292 16192 21332 16232
rect 21580 16108 21620 16148
rect 21772 18460 21812 18500
rect 21772 17536 21812 17576
rect 21964 18208 22004 18248
rect 21964 18040 22004 18080
rect 22444 18460 22484 18500
rect 22060 14512 22100 14552
rect 20524 7120 20564 7160
rect 18988 6868 19028 6908
rect 18660 6028 19028 6068
rect 19900 6784 20268 6824
rect 21292 10144 21332 10184
rect 21868 10144 21908 10184
rect 19900 5272 20268 5312
rect 21772 7204 21812 7244
rect 22540 17032 22580 17072
rect 22732 17452 22772 17492
rect 22924 18208 22964 18248
rect 23020 18124 23060 18164
rect 23980 25432 24020 25472
rect 23788 24256 23828 24296
rect 23788 24088 23828 24128
rect 23980 24004 24020 24044
rect 23980 20980 24020 21020
rect 23596 18460 23636 18500
rect 23020 17620 23060 17660
rect 23020 17116 23060 17156
rect 22924 16948 22964 16988
rect 23212 17536 23252 17576
rect 22636 13924 22676 13964
rect 23596 17788 23636 17828
rect 23596 17536 23636 17576
rect 24172 24760 24212 24800
rect 24172 23752 24212 23792
rect 24364 24676 24404 24716
rect 24460 24592 24500 24632
rect 24364 23920 24404 23960
rect 24460 23836 24500 23876
rect 24364 23668 24404 23708
rect 24364 22996 24404 23036
rect 24844 26104 24884 26144
rect 24844 24676 24884 24716
rect 24556 23164 24596 23204
rect 24652 22996 24692 23036
rect 24364 20896 24404 20936
rect 24172 19048 24212 19088
rect 23980 18544 24020 18584
rect 23788 18124 23828 18164
rect 23884 18040 23924 18080
rect 23884 17452 23924 17492
rect 23884 17032 23924 17072
rect 24076 17956 24116 17996
rect 24076 17788 24116 17828
rect 24076 16276 24116 16316
rect 23020 15688 23060 15728
rect 23788 16108 23828 16148
rect 23404 16024 23444 16064
rect 23116 14596 23156 14636
rect 23020 14428 23060 14468
rect 23308 14512 23348 14552
rect 23020 14008 23060 14048
rect 23212 13168 23252 13208
rect 23116 11740 23156 11780
rect 22732 10312 22772 10352
rect 22444 9472 22484 9512
rect 23212 9472 23252 9512
rect 22924 8128 22964 8168
rect 24364 17536 24404 17576
rect 24364 16948 24404 16988
rect 23788 14764 23828 14804
rect 23788 14596 23828 14636
rect 24268 16192 24308 16232
rect 24844 20056 24884 20096
rect 24652 17536 24692 17576
rect 24844 19048 24884 19088
rect 25036 26944 25076 26984
rect 25324 26020 25364 26060
rect 25132 25936 25172 25976
rect 25132 23080 25172 23120
rect 25036 22996 25076 23036
rect 25612 26104 25652 26144
rect 25420 25348 25460 25388
rect 25420 25012 25460 25052
rect 25516 25096 25556 25136
rect 25420 24592 25460 24632
rect 25324 24256 25364 24296
rect 25132 22156 25172 22196
rect 25036 21484 25076 21524
rect 24940 18460 24980 18500
rect 24844 17116 24884 17156
rect 24940 17032 24980 17072
rect 24172 11656 24212 11696
rect 24076 10984 24116 11024
rect 23980 10900 24020 10940
rect 23020 7036 23060 7076
rect 23212 6868 23252 6908
rect 23596 7960 23636 8000
rect 23692 7120 23732 7160
rect 23692 6448 23732 6488
rect 24172 7960 24212 8000
rect 24940 14764 24980 14804
rect 25132 15688 25172 15728
rect 25132 14680 25172 14720
rect 25516 23752 25556 23792
rect 25324 23332 25364 23372
rect 25708 25936 25748 25976
rect 25708 25432 25748 25472
rect 25708 24676 25748 24716
rect 26956 28036 26996 28076
rect 27674 27952 28042 27992
rect 26434 27196 26802 27236
rect 27340 27532 27380 27572
rect 25996 25348 26036 25388
rect 25804 24004 25844 24044
rect 26764 26104 26804 26144
rect 26380 26020 26420 26060
rect 26860 25936 26900 25976
rect 26434 25684 26802 25724
rect 28492 27364 28532 27404
rect 27674 26440 28042 26480
rect 27820 26272 27860 26312
rect 26380 25096 26420 25136
rect 26188 24844 26228 24884
rect 26092 24760 26132 24800
rect 26188 24592 26228 24632
rect 25612 23080 25652 23120
rect 25324 22324 25364 22364
rect 25708 22156 25748 22196
rect 25708 20896 25748 20936
rect 25420 20224 25460 20264
rect 25516 19972 25556 20012
rect 25516 18628 25556 18668
rect 25804 19972 25844 20012
rect 25708 18544 25748 18584
rect 25708 17536 25748 17576
rect 25612 16948 25652 16988
rect 25708 15604 25748 15644
rect 25516 14764 25556 14804
rect 25324 14680 25364 14720
rect 24460 10984 24500 11024
rect 24556 10816 24596 10856
rect 24844 10984 24884 11024
rect 25132 10816 25172 10856
rect 24364 8044 24404 8084
rect 25036 7960 25076 8000
rect 24460 7036 24500 7076
rect 25708 14428 25748 14468
rect 25420 11740 25460 11780
rect 25324 8044 25364 8084
rect 25612 10984 25652 11024
rect 25900 14260 25940 14300
rect 27052 25180 27092 25220
rect 26956 25012 26996 25052
rect 26380 24508 26420 24548
rect 26668 24340 26708 24380
rect 26284 24256 26324 24296
rect 26434 24172 26802 24212
rect 26380 23500 26420 23540
rect 26092 22324 26132 22364
rect 26092 22156 26132 22196
rect 26092 20728 26132 20768
rect 26092 17704 26132 17744
rect 26380 22996 26420 23036
rect 26668 23752 26708 23792
rect 26668 23584 26708 23624
rect 26476 22828 26516 22868
rect 27052 24508 27092 24548
rect 26956 24340 26996 24380
rect 28108 25936 28148 25976
rect 27436 25348 27476 25388
rect 27244 23920 27284 23960
rect 26860 22996 26900 23036
rect 26956 22912 26996 22952
rect 26434 22660 26802 22700
rect 26380 22156 26420 22196
rect 26860 21988 26900 22028
rect 26434 21148 26802 21188
rect 26476 20980 26516 21020
rect 26860 20812 26900 20852
rect 26572 20644 26612 20684
rect 26860 20560 26900 20600
rect 26764 20476 26804 20516
rect 26668 20308 26708 20348
rect 26572 20224 26612 20264
rect 26476 19888 26516 19928
rect 26764 20140 26804 20180
rect 26860 20056 26900 20096
rect 26668 19888 26708 19928
rect 26572 19804 26612 19844
rect 26434 19636 26802 19676
rect 26572 19300 26612 19340
rect 26476 18628 26516 18668
rect 27148 23164 27188 23204
rect 27244 22996 27284 23036
rect 27148 22744 27188 22784
rect 27244 22828 27284 22868
rect 27244 21484 27284 21524
rect 27628 25348 27668 25388
rect 27674 24928 28042 24968
rect 27436 23080 27476 23120
rect 27628 24256 27668 24296
rect 28300 25012 28340 25052
rect 27628 23668 27668 23708
rect 27724 23584 27764 23624
rect 27674 23416 28042 23456
rect 27820 23248 27860 23288
rect 27628 22912 27668 22952
rect 27724 22996 27764 23036
rect 27628 22744 27668 22784
rect 28108 22660 28148 22700
rect 27674 21904 28042 21944
rect 27916 21568 27956 21608
rect 27244 20308 27284 20348
rect 27340 20224 27380 20264
rect 26764 18376 26804 18416
rect 26434 18124 26802 18164
rect 26284 17620 26324 17660
rect 26284 16948 26324 16988
rect 26434 16612 26802 16652
rect 26284 16276 26324 16316
rect 26668 16108 26708 16148
rect 26764 16024 26804 16064
rect 26188 15520 26228 15560
rect 26092 15352 26132 15392
rect 26092 14512 26132 14552
rect 26434 15100 26802 15140
rect 26188 13756 26228 13796
rect 26764 14596 26804 14636
rect 26476 13756 26516 13796
rect 26434 13588 26802 13628
rect 26572 13168 26612 13208
rect 26434 12076 26802 12116
rect 26956 16192 26996 16232
rect 26956 15604 26996 15644
rect 27052 14764 27092 14804
rect 27148 15604 27188 15644
rect 26956 14596 26996 14636
rect 26956 14428 26996 14468
rect 26476 11656 26516 11696
rect 26284 10900 26324 10940
rect 26434 10564 26802 10604
rect 26092 10312 26132 10352
rect 26284 9556 26324 9596
rect 26284 9304 26324 9344
rect 26188 8128 26228 8168
rect 27724 21064 27764 21104
rect 27916 20980 27956 21020
rect 27628 20728 27668 20768
rect 28012 20644 28052 20684
rect 28108 21568 28148 21608
rect 27674 20392 28042 20432
rect 27532 20308 27572 20348
rect 27820 20224 27860 20264
rect 27340 18628 27380 18668
rect 27436 18460 27476 18500
rect 27436 17116 27476 17156
rect 27724 19888 27764 19928
rect 27628 19804 27668 19844
rect 27628 19048 27668 19088
rect 28396 23164 28436 23204
rect 28396 22996 28436 23036
rect 28396 22324 28436 22364
rect 28300 20644 28340 20684
rect 27674 18880 28042 18920
rect 27628 18628 27668 18668
rect 28108 17956 28148 17996
rect 27724 17536 27764 17576
rect 27674 17368 28042 17408
rect 27724 17116 27764 17156
rect 28300 19048 28340 19088
rect 28972 25936 29012 25976
rect 29164 26020 29204 26060
rect 28876 24592 28916 24632
rect 28972 24508 29012 24548
rect 28780 23248 28820 23288
rect 28588 22996 28628 23036
rect 28300 18544 28340 18584
rect 28396 18460 28436 18500
rect 28396 17956 28436 17996
rect 27674 15856 28042 15896
rect 27724 15688 27764 15728
rect 28012 15520 28052 15560
rect 27674 14344 28042 14384
rect 28204 14260 28244 14300
rect 27820 13924 27860 13964
rect 27674 12832 28042 12872
rect 27916 11740 27956 11780
rect 28300 14008 28340 14048
rect 28684 21568 28724 21608
rect 28684 20812 28724 20852
rect 28972 23164 29012 23204
rect 28876 20560 28916 20600
rect 28972 20728 29012 20768
rect 28780 18712 28820 18752
rect 28876 18628 28916 18668
rect 29548 23248 29588 23288
rect 29548 22912 29588 22952
rect 29164 21484 29204 21524
rect 28876 13924 28916 13964
rect 28492 11740 28532 11780
rect 27674 11320 28042 11360
rect 29548 21988 29588 22028
rect 30124 26860 30164 26900
rect 29836 25096 29876 25136
rect 29740 24508 29780 24548
rect 29644 18796 29684 18836
rect 29740 24256 29780 24296
rect 30028 24256 30068 24296
rect 30028 23836 30068 23876
rect 29932 23164 29972 23204
rect 29932 20308 29972 20348
rect 29932 18628 29972 18668
rect 29164 14092 29204 14132
rect 29260 11824 29300 11864
rect 29068 11740 29108 11780
rect 29260 10984 29300 11024
rect 26956 10144 26996 10184
rect 27052 10060 27092 10100
rect 27674 9808 28042 9848
rect 26434 9052 26802 9092
rect 27052 9304 27092 9344
rect 26434 7540 26802 7580
rect 26380 7204 26420 7244
rect 29452 13084 29492 13124
rect 29740 17032 29780 17072
rect 29644 14008 29684 14048
rect 29452 11152 29492 11192
rect 29548 11068 29588 11108
rect 29740 13084 29780 13124
rect 30796 27364 30836 27404
rect 30220 23836 30260 23876
rect 29932 15604 29972 15644
rect 29932 15352 29972 15392
rect 29836 12244 29876 12284
rect 30412 22324 30452 22364
rect 30412 17452 30452 17492
rect 30508 18796 30548 18836
rect 30028 14008 30068 14048
rect 30124 14092 30164 14132
rect 31084 24340 31124 24380
rect 30700 17704 30740 17744
rect 30988 18796 31028 18836
rect 30892 17452 30932 17492
rect 30700 14932 30740 14972
rect 30700 12328 30740 12368
rect 30700 11908 30740 11948
rect 30988 14848 31028 14888
rect 31084 13924 31124 13964
rect 30124 11152 30164 11192
rect 29836 10900 29876 10940
rect 30412 10816 30452 10856
rect 30796 10816 30836 10856
rect 30412 10564 30452 10604
rect 30796 10312 30836 10352
rect 27674 8296 28042 8336
rect 27674 6784 28042 6824
rect 24076 6448 24116 6488
rect 26434 6028 26802 6068
rect 27674 5272 28042 5312
rect 18660 4516 19028 4556
rect 26434 4516 26802 4556
rect 4352 3760 4720 3800
rect 12126 3760 12494 3800
rect 19900 3760 20268 3800
rect 27674 3760 28042 3800
rect 3112 3004 3480 3044
rect 10886 3004 11254 3044
rect 18660 3004 19028 3044
rect 26434 3004 26802 3044
rect 4352 2248 4720 2288
rect 12126 2248 12494 2288
rect 19900 2248 20268 2288
rect 27674 2248 28042 2288
rect 3112 1492 3480 1532
rect 10886 1492 11254 1532
rect 18660 1492 19028 1532
rect 26434 1492 26802 1532
rect 4352 736 4720 776
rect 12126 736 12494 776
rect 19900 736 20268 776
rect 27674 736 28042 776
<< metal4 >>
rect 1507 28120 1516 28160
rect 1556 28120 4684 28160
rect 4724 28120 4733 28160
rect 12355 28120 12364 28160
rect 12404 28120 13036 28160
rect 13076 28120 13085 28160
rect 26947 28036 26956 28076
rect 26996 28036 27436 28076
rect 27476 28036 27485 28076
rect 4343 27952 4352 27992
rect 4720 27952 4729 27992
rect 12117 27952 12126 27992
rect 12494 27952 12503 27992
rect 19891 27952 19900 27992
rect 20268 27952 20277 27992
rect 27665 27952 27674 27992
rect 28042 27952 28051 27992
rect 3139 27784 3148 27824
rect 3188 27784 3628 27824
rect 3668 27784 3677 27824
rect 10051 27700 10060 27740
rect 10100 27700 10156 27740
rect 10196 27700 10205 27740
rect 12163 27616 12172 27656
rect 12212 27616 15340 27656
rect 15380 27616 15389 27656
rect 1891 27532 1900 27572
rect 1940 27532 8524 27572
rect 8564 27532 8573 27572
rect 27245 27532 27340 27572
rect 27380 27532 27389 27572
rect 2371 27448 2380 27488
rect 2420 27448 6892 27488
rect 6932 27448 6941 27488
rect 10819 27364 10828 27404
rect 10868 27364 11500 27404
rect 11540 27364 11549 27404
rect 28397 27364 28492 27404
rect 28532 27364 28541 27404
rect 30787 27364 30796 27404
rect 30836 27364 31084 27404
rect 31124 27364 31133 27404
rect 3103 27196 3112 27236
rect 3480 27196 3489 27236
rect 10877 27196 10886 27236
rect 11254 27196 11263 27236
rect 18651 27196 18660 27236
rect 19028 27196 19037 27236
rect 26425 27196 26434 27236
rect 26802 27196 26811 27236
rect 10435 27112 10444 27152
rect 10484 27112 15052 27152
rect 15092 27112 15101 27152
rect 11203 27028 11212 27068
rect 11252 27028 17740 27068
rect 17780 27028 17789 27068
rect 13315 26944 13324 26984
rect 13364 26944 14956 26984
rect 14996 26944 15005 26984
rect 23107 26944 23116 26984
rect 23156 26944 25036 26984
rect 25076 26944 25085 26984
rect 3235 26860 3244 26900
rect 3284 26860 4396 26900
rect 4436 26860 4445 26900
rect 10915 26860 10924 26900
rect 10964 26860 13420 26900
rect 13460 26860 13469 26900
rect 30029 26860 30124 26900
rect 30164 26860 30173 26900
rect 5539 26776 5548 26816
rect 5588 26776 10100 26816
rect 11587 26776 11596 26816
rect 11636 26776 11980 26816
rect 12020 26776 12029 26816
rect 12163 26776 12172 26816
rect 12212 26776 13324 26816
rect 13364 26776 13373 26816
rect 13699 26776 13708 26816
rect 13748 26776 20332 26816
rect 20372 26776 20381 26816
rect 10060 26732 10100 26776
rect 4579 26692 4588 26732
rect 4628 26692 7180 26732
rect 7220 26692 7229 26732
rect 10060 26692 13516 26732
rect 13556 26692 13565 26732
rect 4675 26608 4684 26648
rect 4724 26608 6892 26648
rect 6932 26608 7372 26648
rect 7412 26608 7421 26648
rect 12451 26608 12460 26648
rect 12500 26608 13804 26648
rect 13844 26608 13853 26648
rect 18211 26608 18220 26648
rect 18260 26608 20140 26648
rect 20180 26608 20189 26648
rect 12835 26524 12844 26564
rect 12884 26524 16300 26564
rect 16340 26524 16349 26564
rect 17731 26524 17740 26564
rect 17780 26524 18892 26564
rect 18932 26524 18941 26564
rect 4343 26440 4352 26480
rect 4720 26440 4729 26480
rect 12117 26440 12126 26480
rect 12494 26440 12503 26480
rect 13123 26440 13132 26480
rect 13172 26440 14284 26480
rect 14324 26440 14333 26480
rect 18979 26440 18988 26480
rect 19028 26440 19276 26480
rect 19316 26440 19325 26480
rect 19891 26440 19900 26480
rect 20268 26440 20277 26480
rect 27665 26440 27674 26480
rect 28042 26440 28051 26480
rect 2947 26356 2956 26396
rect 2996 26356 5164 26396
rect 5204 26356 5213 26396
rect 11875 26356 11884 26396
rect 11924 26356 18028 26396
rect 18068 26356 18077 26396
rect 27811 26272 27820 26312
rect 27860 26272 28204 26312
rect 28244 26272 28253 26312
rect 11587 26188 11596 26228
rect 11636 26188 13132 26228
rect 13172 26188 13181 26228
rect 18317 26188 18412 26228
rect 18452 26188 20044 26228
rect 20084 26188 20093 26228
rect 2851 26104 2860 26144
rect 2900 26104 8332 26144
rect 8372 26104 8381 26144
rect 20717 26104 20812 26144
rect 20852 26104 20861 26144
rect 24835 26104 24844 26144
rect 24884 26104 25612 26144
rect 25652 26104 26764 26144
rect 26804 26104 26813 26144
rect 12451 26020 12460 26060
rect 12500 26020 14476 26060
rect 14516 26020 14525 26060
rect 25315 26020 25324 26060
rect 25364 26020 26380 26060
rect 26420 26020 26429 26060
rect 29069 26020 29164 26060
rect 29204 26020 29213 26060
rect 1891 25936 1900 25976
rect 1940 25936 3532 25976
rect 3572 25936 3581 25976
rect 16195 25936 16204 25976
rect 16244 25936 17452 25976
rect 17492 25936 17501 25976
rect 25123 25936 25132 25976
rect 25172 25936 25708 25976
rect 25748 25936 26860 25976
rect 26900 25936 26909 25976
rect 27523 25936 27532 25976
rect 27572 25936 28108 25976
rect 28148 25936 28157 25976
rect 28963 25936 28972 25976
rect 29012 25936 30028 25976
rect 30068 25936 30077 25976
rect 2851 25768 2860 25808
rect 2900 25768 3724 25808
rect 3764 25768 3773 25808
rect 18403 25768 18412 25808
rect 18452 25768 19660 25808
rect 19700 25768 21484 25808
rect 21524 25768 21533 25808
rect 3103 25684 3112 25724
rect 3480 25684 3489 25724
rect 10877 25684 10886 25724
rect 11254 25684 11263 25724
rect 18651 25684 18660 25724
rect 19028 25684 19037 25724
rect 26425 25684 26434 25724
rect 26802 25684 26811 25724
rect 10051 25600 10060 25640
rect 10100 25600 10156 25640
rect 10196 25600 10205 25640
rect 1603 25432 1612 25472
rect 1652 25432 3244 25472
rect 3284 25432 3293 25472
rect 23971 25432 23980 25472
rect 24020 25432 25708 25472
rect 25748 25432 25757 25472
rect 2563 25348 2572 25388
rect 2612 25348 4204 25388
rect 4244 25348 4253 25388
rect 12451 25348 12460 25388
rect 12500 25348 15628 25388
rect 15668 25348 15677 25388
rect 25411 25348 25420 25388
rect 25460 25348 25996 25388
rect 26036 25348 26045 25388
rect 27427 25348 27436 25388
rect 27476 25348 27628 25388
rect 27668 25348 27677 25388
rect 5155 25264 5164 25304
rect 5204 25264 5356 25304
rect 5396 25264 6508 25304
rect 6548 25264 8620 25304
rect 8660 25264 8669 25304
rect 10723 25264 10732 25304
rect 10772 25264 10828 25304
rect 10868 25264 10877 25304
rect 12163 25264 12172 25304
rect 12212 25264 13516 25304
rect 13556 25264 13565 25304
rect 547 25180 556 25220
rect 596 25180 8524 25220
rect 8564 25180 8573 25220
rect 11683 25180 11692 25220
rect 11732 25180 13420 25220
rect 13460 25180 13708 25220
rect 13748 25180 13757 25220
rect 26179 25180 26188 25220
rect 26228 25180 27052 25220
rect 27092 25180 27101 25220
rect 14755 25096 14764 25136
rect 14804 25096 15340 25136
rect 15380 25096 15389 25136
rect 25507 25096 25516 25136
rect 25556 25096 26380 25136
rect 26420 25096 26429 25136
rect 29539 25096 29548 25136
rect 29588 25096 29836 25136
rect 29876 25096 29885 25136
rect 20803 25012 20812 25052
rect 20852 25012 25420 25052
rect 25460 25012 26956 25052
rect 26996 25012 28300 25052
rect 28340 25012 28349 25052
rect 4343 24928 4352 24968
rect 4720 24928 4729 24968
rect 12117 24928 12126 24968
rect 12494 24928 12503 24968
rect 19891 24928 19900 24968
rect 20268 24928 20277 24968
rect 27665 24928 27674 24968
rect 28042 24928 28051 24968
rect 14659 24844 14668 24884
rect 14708 24844 16108 24884
rect 16148 24844 26188 24884
rect 26228 24844 26237 24884
rect 1699 24760 1708 24800
rect 1748 24760 6220 24800
rect 6260 24760 6269 24800
rect 13891 24760 13900 24800
rect 13940 24760 17548 24800
rect 17588 24760 17597 24800
rect 20515 24760 20524 24800
rect 20564 24760 24172 24800
rect 24212 24760 26092 24800
rect 26132 24760 26141 24800
rect 13507 24676 13516 24716
rect 13556 24676 16972 24716
rect 17012 24676 17021 24716
rect 24355 24676 24364 24716
rect 24404 24676 24844 24716
rect 24884 24676 25708 24716
rect 25748 24676 25757 24716
rect 1987 24592 1996 24632
rect 2036 24592 9292 24632
rect 9332 24592 9341 24632
rect 23203 24592 23212 24632
rect 23252 24592 24460 24632
rect 24500 24592 25420 24632
rect 25460 24592 25469 24632
rect 26179 24592 26188 24632
rect 26228 24592 28876 24632
rect 28916 24592 28925 24632
rect 2371 24508 2380 24548
rect 2420 24508 8716 24548
rect 8756 24508 8765 24548
rect 18403 24508 18412 24548
rect 18452 24508 18604 24548
rect 18644 24508 18653 24548
rect 20323 24508 20332 24548
rect 20372 24508 26380 24548
rect 26420 24508 27052 24548
rect 27092 24508 27101 24548
rect 28963 24508 28972 24548
rect 29012 24508 29452 24548
rect 29492 24508 29501 24548
rect 29635 24508 29644 24548
rect 29684 24508 29740 24548
rect 29780 24508 29789 24548
rect 8716 24464 8756 24508
rect 8716 24424 10252 24464
rect 10292 24424 13036 24464
rect 13076 24424 13085 24464
rect 10051 24340 10060 24380
rect 10100 24340 12844 24380
rect 12884 24340 12893 24380
rect 15427 24340 15436 24380
rect 15476 24340 17068 24380
rect 17108 24340 17117 24380
rect 26659 24340 26668 24380
rect 26708 24340 26956 24380
rect 26996 24340 27005 24380
rect 27139 24340 27148 24380
rect 27188 24340 31084 24380
rect 31124 24340 31133 24380
rect 23779 24256 23788 24296
rect 23828 24256 25324 24296
rect 25364 24256 26284 24296
rect 26324 24256 26333 24296
rect 27043 24256 27052 24296
rect 27092 24256 27628 24296
rect 27668 24256 27677 24296
rect 29731 24256 29740 24296
rect 29780 24256 30028 24296
rect 30068 24256 30077 24296
rect 3103 24172 3112 24212
rect 3480 24172 3489 24212
rect 10877 24172 10886 24212
rect 11254 24172 11263 24212
rect 18651 24172 18660 24212
rect 19028 24172 19037 24212
rect 26425 24172 26434 24212
rect 26802 24172 26811 24212
rect 15427 24088 15436 24128
rect 15476 24088 23788 24128
rect 23828 24088 23837 24128
rect 23971 24004 23980 24044
rect 24020 24004 25804 24044
rect 25844 24004 25853 24044
rect 24355 23920 24364 23960
rect 24404 23920 27244 23960
rect 27284 23920 27293 23960
rect 10531 23836 10540 23876
rect 10580 23836 10732 23876
rect 10772 23836 12652 23876
rect 12692 23836 14188 23876
rect 14228 23836 16684 23876
rect 16724 23836 16733 23876
rect 20227 23836 20236 23876
rect 20276 23836 20428 23876
rect 20468 23836 20477 23876
rect 22147 23836 22156 23876
rect 22196 23836 23500 23876
rect 23540 23836 23549 23876
rect 24451 23836 24460 23876
rect 24500 23836 30028 23876
rect 30068 23836 30077 23876
rect 30211 23836 30220 23876
rect 30260 23836 30796 23876
rect 30836 23836 30845 23876
rect 2467 23752 2476 23792
rect 2516 23752 5260 23792
rect 5300 23752 9196 23792
rect 9236 23752 9245 23792
rect 12163 23752 12172 23792
rect 12212 23752 16780 23792
rect 16820 23752 16829 23792
rect 24163 23752 24172 23792
rect 24212 23752 25516 23792
rect 25556 23752 25565 23792
rect 26659 23752 26668 23792
rect 26708 23752 29260 23792
rect 29300 23752 29309 23792
rect 8323 23668 8332 23708
rect 8372 23668 11020 23708
rect 11060 23668 11069 23708
rect 24355 23668 24364 23708
rect 24404 23668 27628 23708
rect 27668 23668 27677 23708
rect 8227 23584 8236 23624
rect 8276 23584 8812 23624
rect 8852 23584 8861 23624
rect 10051 23584 10060 23624
rect 10100 23584 13228 23624
rect 13268 23584 13612 23624
rect 13652 23584 13661 23624
rect 26659 23584 26668 23624
rect 26708 23584 26956 23624
rect 26996 23584 27005 23624
rect 27715 23584 27724 23624
rect 27764 23584 27773 23624
rect 27724 23540 27764 23584
rect 4003 23500 4012 23540
rect 4052 23500 10444 23540
rect 10484 23500 10493 23540
rect 26371 23500 26380 23540
rect 26420 23500 27764 23540
rect 4343 23416 4352 23456
rect 4720 23416 4729 23456
rect 10051 23416 10060 23456
rect 10100 23416 12020 23456
rect 12117 23416 12126 23456
rect 12494 23416 12503 23456
rect 19891 23416 19900 23456
rect 20268 23416 20277 23456
rect 27665 23416 27674 23456
rect 28042 23416 28051 23456
rect 11980 23372 12020 23416
rect 739 23332 748 23372
rect 788 23332 2900 23372
rect 9187 23332 9196 23372
rect 9236 23332 9388 23372
rect 9428 23332 11788 23372
rect 11828 23332 11837 23372
rect 11980 23332 12556 23372
rect 12596 23332 12605 23372
rect 13795 23332 13804 23372
rect 13844 23332 23060 23372
rect 25315 23332 25324 23372
rect 25364 23332 30316 23372
rect 30356 23332 30365 23372
rect 2860 23288 2900 23332
rect 23020 23288 23060 23332
rect 163 23248 172 23288
rect 212 23248 1420 23288
rect 1460 23248 1469 23288
rect 2860 23248 16684 23288
rect 16724 23248 16733 23288
rect 16867 23248 16876 23288
rect 16916 23248 18220 23288
rect 18260 23248 18269 23288
rect 20227 23248 20236 23288
rect 20276 23248 20428 23288
rect 20468 23248 20477 23288
rect 23020 23248 27148 23288
rect 27188 23248 27197 23288
rect 27811 23248 27820 23288
rect 27860 23248 28780 23288
rect 28820 23248 28829 23288
rect 29539 23248 29548 23288
rect 29588 23248 29597 23288
rect 29548 23204 29588 23248
rect 931 23164 940 23204
rect 980 23164 4396 23204
rect 4436 23164 4445 23204
rect 5059 23164 5068 23204
rect 5108 23164 6796 23204
rect 6836 23164 6845 23204
rect 10243 23164 10252 23204
rect 10292 23164 11116 23204
rect 11156 23164 11165 23204
rect 15235 23164 15244 23204
rect 15284 23164 24556 23204
rect 24596 23164 24605 23204
rect 27139 23164 27148 23204
rect 27188 23164 27244 23204
rect 27284 23164 27293 23204
rect 28387 23164 28396 23204
rect 28436 23164 28972 23204
rect 29012 23164 29021 23204
rect 29548 23164 29932 23204
rect 29972 23164 29981 23204
rect 10339 23080 10348 23120
rect 10388 23080 12076 23120
rect 12116 23080 19084 23120
rect 19124 23080 19133 23120
rect 25123 23080 25132 23120
rect 25172 23080 25612 23120
rect 25652 23080 25661 23120
rect 27427 23080 27436 23120
rect 27476 23080 30604 23120
rect 30644 23080 30653 23120
rect 11779 22996 11788 23036
rect 11828 22996 11837 23036
rect 18019 22996 18028 23036
rect 18068 22996 20812 23036
rect 20852 22996 20861 23036
rect 24355 22996 24364 23036
rect 24404 22996 24652 23036
rect 24692 22996 24701 23036
rect 25027 22996 25036 23036
rect 25076 22996 26380 23036
rect 26420 22996 26429 23036
rect 26851 22996 26860 23036
rect 26900 22996 27092 23036
rect 27235 22996 27244 23036
rect 27284 22996 27724 23036
rect 27764 22996 27773 23036
rect 28387 22996 28396 23036
rect 28436 22996 28588 23036
rect 28628 22996 28637 23036
rect 11788 22952 11828 22996
rect 27052 22952 27092 22996
rect 2755 22912 2764 22952
rect 2804 22912 2956 22952
rect 2996 22912 3005 22952
rect 3427 22912 3436 22952
rect 3476 22912 3820 22952
rect 3860 22912 3869 22952
rect 7843 22912 7852 22952
rect 7892 22912 8908 22952
rect 8948 22912 8957 22952
rect 11693 22912 11788 22952
rect 11828 22912 14188 22952
rect 14228 22912 14237 22952
rect 17827 22912 17836 22952
rect 17876 22912 23404 22952
rect 23444 22912 23453 22952
rect 26083 22912 26092 22952
rect 26132 22912 26956 22952
rect 26996 22912 27005 22952
rect 27052 22912 27284 22952
rect 27619 22912 27628 22952
rect 27668 22912 29548 22952
rect 29588 22912 29597 22952
rect 27244 22868 27284 22912
rect 7939 22828 7948 22868
rect 7988 22828 8428 22868
rect 8468 22828 8477 22868
rect 10051 22828 10060 22868
rect 10100 22828 13324 22868
rect 13364 22828 13373 22868
rect 20899 22828 20908 22868
rect 20948 22828 22636 22868
rect 22676 22828 22685 22868
rect 26467 22828 26476 22868
rect 26516 22828 26525 22868
rect 27235 22828 27244 22868
rect 27284 22828 27293 22868
rect 26476 22784 26516 22828
rect 835 22744 844 22784
rect 884 22744 4204 22784
rect 4244 22744 4396 22784
rect 4436 22744 5260 22784
rect 5300 22744 7852 22784
rect 7892 22744 7901 22784
rect 10435 22744 10444 22784
rect 10484 22744 12172 22784
rect 12212 22744 12221 22784
rect 26476 22744 27092 22784
rect 27139 22744 27148 22784
rect 27188 22744 27628 22784
rect 27668 22744 27677 22784
rect 27052 22700 27092 22744
rect 3103 22660 3112 22700
rect 3480 22660 3489 22700
rect 10877 22660 10886 22700
rect 11254 22660 11263 22700
rect 18651 22660 18660 22700
rect 19028 22660 19037 22700
rect 26425 22660 26434 22700
rect 26802 22660 26811 22700
rect 27052 22660 28108 22700
rect 28148 22660 28157 22700
rect 835 22576 844 22616
rect 884 22576 8812 22616
rect 8852 22576 8861 22616
rect 67 22492 76 22532
rect 116 22492 460 22532
rect 500 22492 509 22532
rect 4003 22492 4012 22532
rect 4052 22492 4300 22532
rect 4340 22492 5164 22532
rect 5204 22492 8524 22532
rect 8564 22492 11788 22532
rect 11828 22492 11837 22532
rect 2659 22408 2668 22448
rect 2708 22408 3916 22448
rect 3956 22408 4492 22448
rect 4532 22408 4541 22448
rect 5443 22408 5452 22448
rect 5492 22408 8428 22448
rect 8468 22408 8477 22448
rect 3724 22324 7468 22364
rect 7508 22324 8620 22364
rect 8660 22324 8669 22364
rect 22243 22324 22252 22364
rect 22292 22324 23116 22364
rect 23156 22324 23165 22364
rect 25315 22324 25324 22364
rect 25364 22324 26092 22364
rect 26132 22324 28396 22364
rect 28436 22324 28445 22364
rect 30317 22324 30412 22364
rect 30452 22324 30461 22364
rect 3724 22280 3764 22324
rect 2275 22240 2284 22280
rect 2324 22240 3724 22280
rect 3764 22240 3773 22280
rect 5443 22240 5452 22280
rect 5492 22240 6412 22280
rect 6452 22240 6461 22280
rect 7651 22240 7660 22280
rect 7700 22240 10156 22280
rect 10196 22240 13996 22280
rect 14036 22240 14045 22280
rect 14179 22240 14188 22280
rect 14228 22240 18028 22280
rect 18068 22240 18077 22280
rect 22819 22240 22828 22280
rect 22868 22240 23212 22280
rect 23252 22240 23261 22280
rect 1795 22156 1804 22196
rect 1844 22156 2668 22196
rect 2708 22156 2717 22196
rect 4867 22156 4876 22196
rect 4916 22156 5740 22196
rect 5780 22156 5789 22196
rect 6115 22156 6124 22196
rect 6164 22156 9004 22196
rect 9044 22156 9053 22196
rect 25123 22156 25132 22196
rect 25172 22156 25708 22196
rect 25748 22156 25757 22196
rect 26083 22156 26092 22196
rect 26132 22156 26380 22196
rect 26420 22156 26429 22196
rect 5539 22072 5548 22112
rect 5588 22072 8236 22112
rect 8276 22072 8285 22112
rect 8515 22072 8524 22112
rect 8564 22072 10060 22112
rect 10100 22072 10109 22112
rect 12355 22072 12364 22112
rect 12404 22072 12652 22112
rect 12692 22072 12701 22112
rect 547 21988 556 22028
rect 596 21988 5644 22028
rect 5684 21988 5693 22028
rect 8899 21988 8908 22028
rect 8948 21988 9196 22028
rect 9236 21988 9245 22028
rect 10339 21988 10348 22028
rect 10388 21988 12748 22028
rect 12788 21988 12797 22028
rect 26851 21988 26860 22028
rect 26900 21988 29548 22028
rect 29588 21988 29597 22028
rect 4343 21904 4352 21944
rect 4720 21904 4729 21944
rect 12117 21904 12126 21944
rect 12494 21904 12503 21944
rect 19891 21904 19900 21944
rect 20268 21904 20277 21944
rect 27665 21904 27674 21944
rect 28042 21904 28051 21944
rect 1699 21820 1708 21860
rect 1748 21820 1996 21860
rect 2036 21820 2045 21860
rect 7651 21820 7660 21860
rect 7700 21820 8524 21860
rect 8564 21820 8573 21860
rect 9187 21820 9196 21860
rect 9236 21820 9964 21860
rect 10004 21820 10013 21860
rect 67 21736 76 21776
rect 116 21736 2900 21776
rect 6019 21736 6028 21776
rect 6068 21736 9292 21776
rect 9332 21736 9341 21776
rect 9571 21736 9580 21776
rect 9620 21736 10924 21776
rect 10964 21736 10973 21776
rect 14371 21736 14380 21776
rect 14420 21736 16108 21776
rect 16148 21736 16157 21776
rect 2860 21692 2900 21736
rect 365 21652 460 21692
rect 500 21652 509 21692
rect 2860 21652 16012 21692
rect 16052 21652 16061 21692
rect 1891 21568 1900 21608
rect 1940 21568 3916 21608
rect 3956 21568 3965 21608
rect 5539 21568 5548 21608
rect 5588 21568 6604 21608
rect 6644 21568 6653 21608
rect 8419 21568 8428 21608
rect 8468 21568 8524 21608
rect 8564 21568 8573 21608
rect 10339 21568 10348 21608
rect 10388 21568 10732 21608
rect 10772 21568 10781 21608
rect 12643 21568 12652 21608
rect 12692 21568 14476 21608
rect 14516 21568 14525 21608
rect 18307 21568 18316 21608
rect 18356 21568 18988 21608
rect 19028 21568 19037 21608
rect 27907 21568 27916 21608
rect 27956 21568 28108 21608
rect 28148 21568 28157 21608
rect 28589 21568 28684 21608
rect 28724 21568 28733 21608
rect 3043 21484 3052 21524
rect 3092 21484 3532 21524
rect 3572 21484 4108 21524
rect 4148 21484 4157 21524
rect 4771 21484 4780 21524
rect 4820 21484 5932 21524
rect 5972 21484 5981 21524
rect 6787 21484 6796 21524
rect 6836 21484 7180 21524
rect 7220 21484 7229 21524
rect 9379 21484 9388 21524
rect 9428 21484 10156 21524
rect 10196 21484 10444 21524
rect 10484 21484 11884 21524
rect 11924 21484 11933 21524
rect 14179 21484 14188 21524
rect 14228 21484 15532 21524
rect 15572 21484 15581 21524
rect 22051 21484 22060 21524
rect 22100 21484 25036 21524
rect 25076 21484 25085 21524
rect 27235 21484 27244 21524
rect 27284 21484 29164 21524
rect 29204 21484 29213 21524
rect 2659 21400 2668 21440
rect 2708 21400 3244 21440
rect 3284 21400 3293 21440
rect 2563 21316 2572 21356
rect 2612 21316 4588 21356
rect 4628 21316 6700 21356
rect 6740 21316 6749 21356
rect 15139 21316 15148 21356
rect 15188 21316 15916 21356
rect 15956 21316 15965 21356
rect 3715 21232 3724 21272
rect 3764 21232 4012 21272
rect 4052 21232 14860 21272
rect 14900 21232 14909 21272
rect 3103 21148 3112 21188
rect 3480 21148 3489 21188
rect 10051 21148 10060 21188
rect 10100 21148 10636 21188
rect 10676 21148 10685 21188
rect 10877 21148 10886 21188
rect 11254 21148 11263 21188
rect 12931 21148 12940 21188
rect 12980 21148 13516 21188
rect 13556 21148 15244 21188
rect 15284 21148 15293 21188
rect 18651 21148 18660 21188
rect 19028 21148 19037 21188
rect 26425 21148 26434 21188
rect 26802 21148 26811 21188
rect 1315 21064 1324 21104
rect 1364 21064 8812 21104
rect 8852 21064 8861 21104
rect 27235 21064 27244 21104
rect 27284 21064 27724 21104
rect 27764 21064 27773 21104
rect 3331 20980 3340 21020
rect 3380 20980 4204 21020
rect 4244 20980 4396 21020
rect 4436 20980 4445 21020
rect 8035 20980 8044 21020
rect 8084 20980 9868 21020
rect 9908 20980 14092 21020
rect 14132 20980 18700 21020
rect 18740 20980 18749 21020
rect 23971 20980 23980 21020
rect 24020 20980 26476 21020
rect 26516 20980 27916 21020
rect 27956 20980 27965 21020
rect 1420 20896 4492 20936
rect 4532 20896 4541 20936
rect 8227 20896 8236 20936
rect 8276 20896 8812 20936
rect 8852 20896 8861 20936
rect 15907 20896 15916 20936
rect 15956 20896 18604 20936
rect 18644 20896 18653 20936
rect 24355 20896 24364 20936
rect 24404 20896 25708 20936
rect 25748 20896 25757 20936
rect 1420 20852 1460 20896
rect 1411 20812 1420 20852
rect 1460 20812 1469 20852
rect 3917 20812 4012 20852
rect 4052 20812 5548 20852
rect 5588 20812 5597 20852
rect 8429 20812 8524 20852
rect 8564 20812 9004 20852
rect 9044 20812 9053 20852
rect 14851 20812 14860 20852
rect 14900 20812 16108 20852
rect 16148 20812 16157 20852
rect 17251 20812 17260 20852
rect 17300 20812 19084 20852
rect 19124 20812 19372 20852
rect 19412 20812 19421 20852
rect 26851 20812 26860 20852
rect 26900 20812 28684 20852
rect 28724 20812 28733 20852
rect 2179 20728 2188 20768
rect 2228 20728 4204 20768
rect 4244 20728 4253 20768
rect 4963 20728 4972 20768
rect 5012 20728 5021 20768
rect 7267 20728 7276 20768
rect 7316 20728 8620 20768
rect 8660 20728 8669 20768
rect 26083 20728 26092 20768
rect 26132 20728 27628 20768
rect 27668 20728 27677 20768
rect 27724 20728 28972 20768
rect 29012 20728 29021 20768
rect 4972 20684 5012 20728
rect 27724 20684 27764 20728
rect 2371 20644 2380 20684
rect 2420 20644 2860 20684
rect 2900 20644 2909 20684
rect 4972 20644 7852 20684
rect 7892 20644 9196 20684
rect 9236 20644 9245 20684
rect 19171 20644 19180 20684
rect 19220 20644 19756 20684
rect 19796 20644 19805 20684
rect 26563 20644 26572 20684
rect 26612 20644 27764 20684
rect 28003 20644 28012 20684
rect 28052 20644 28300 20684
rect 28340 20644 28349 20684
rect 355 20560 364 20600
rect 404 20560 460 20600
rect 500 20560 509 20600
rect 1219 20560 1228 20600
rect 1268 20560 7084 20600
rect 7124 20560 7133 20600
rect 26851 20560 26860 20600
rect 26900 20560 28876 20600
rect 28916 20560 28925 20600
rect 643 20476 652 20516
rect 692 20476 1036 20516
rect 1076 20476 1085 20516
rect 14467 20476 14476 20516
rect 14516 20476 18316 20516
rect 18356 20476 18365 20516
rect 26755 20476 26764 20516
rect 26804 20476 27052 20516
rect 27092 20476 27101 20516
rect 4343 20392 4352 20432
rect 4720 20392 4729 20432
rect 5443 20392 5452 20432
rect 5492 20392 7276 20432
rect 7316 20392 8044 20432
rect 8084 20392 8093 20432
rect 12117 20392 12126 20432
rect 12494 20392 12503 20432
rect 19891 20392 19900 20432
rect 20268 20392 20277 20432
rect 27665 20392 27674 20432
rect 28042 20392 28051 20432
rect 451 20308 460 20348
rect 500 20308 7756 20348
rect 7796 20308 7805 20348
rect 15235 20308 15244 20348
rect 15284 20308 16684 20348
rect 16724 20308 16733 20348
rect 18787 20308 18796 20348
rect 18836 20308 20084 20348
rect 26659 20308 26668 20348
rect 26708 20308 27244 20348
rect 27284 20308 27293 20348
rect 27523 20308 27532 20348
rect 27572 20308 29932 20348
rect 29972 20308 29981 20348
rect 20044 20264 20084 20308
rect 27820 20264 27860 20308
rect 4579 20224 4588 20264
rect 4628 20224 4876 20264
rect 4916 20224 6316 20264
rect 6356 20224 6700 20264
rect 6740 20224 8236 20264
rect 8276 20224 9196 20264
rect 9236 20224 9245 20264
rect 19276 20224 19564 20264
rect 19604 20224 19613 20264
rect 20035 20224 20044 20264
rect 20084 20224 20093 20264
rect 25411 20224 25420 20264
rect 25460 20224 26572 20264
rect 26612 20224 26621 20264
rect 27331 20224 27340 20264
rect 27380 20224 27436 20264
rect 27476 20224 27485 20264
rect 27811 20224 27820 20264
rect 27860 20224 27869 20264
rect 5731 20140 5740 20180
rect 5780 20140 5789 20180
rect 11405 20140 11500 20180
rect 11540 20140 11549 20180
rect 14381 20140 14476 20180
rect 14516 20140 14525 20180
rect 16877 20140 16972 20180
rect 17012 20140 17021 20180
rect 2755 20056 2764 20096
rect 2804 20056 4684 20096
rect 4724 20056 5356 20096
rect 5396 20056 5405 20096
rect 5740 20012 5780 20140
rect 19276 20096 19316 20224
rect 26755 20140 26764 20180
rect 26804 20140 26813 20180
rect 26764 20096 26804 20140
rect 6019 20056 6028 20096
rect 6068 20056 6412 20096
rect 6452 20056 6461 20096
rect 13891 20056 13900 20096
rect 13940 20056 14860 20096
rect 14900 20056 16492 20096
rect 16532 20056 16541 20096
rect 19267 20056 19276 20096
rect 19316 20056 19325 20096
rect 24835 20056 24844 20096
rect 24884 20056 26804 20096
rect 26851 20056 26860 20096
rect 26900 20056 27532 20096
rect 27572 20056 27581 20096
rect 4291 19972 4300 20012
rect 4340 19972 5780 20012
rect 6499 19972 6508 20012
rect 6548 19972 6892 20012
rect 6932 19972 6941 20012
rect 13699 19972 13708 20012
rect 13748 19972 15532 20012
rect 15572 19972 16012 20012
rect 16052 19972 16061 20012
rect 25421 19972 25516 20012
rect 25556 19972 25565 20012
rect 25795 19972 25804 20012
rect 25844 19972 27148 20012
rect 27188 19972 27197 20012
rect 26275 19888 26284 19928
rect 26324 19888 26476 19928
rect 26516 19888 26525 19928
rect 26659 19888 26668 19928
rect 26708 19888 27724 19928
rect 27764 19888 27773 19928
rect 1411 19804 1420 19844
rect 1460 19804 2572 19844
rect 2612 19804 2621 19844
rect 7843 19804 7852 19844
rect 7892 19804 8908 19844
rect 8948 19804 8957 19844
rect 14467 19804 14476 19844
rect 14516 19804 15916 19844
rect 15956 19804 15965 19844
rect 18691 19804 18700 19844
rect 18740 19804 19084 19844
rect 19124 19804 19133 19844
rect 26563 19804 26572 19844
rect 26612 19804 27628 19844
rect 27668 19804 27677 19844
rect 2563 19636 2572 19676
rect 2612 19636 2764 19676
rect 2804 19636 2813 19676
rect 3103 19636 3112 19676
rect 3480 19636 3489 19676
rect 10877 19636 10886 19676
rect 11254 19636 11263 19676
rect 18651 19636 18660 19676
rect 19028 19636 19037 19676
rect 26425 19636 26434 19676
rect 26802 19636 26811 19676
rect 2851 19552 2860 19592
rect 2900 19552 3092 19592
rect 3052 19508 3092 19552
rect 3043 19468 3052 19508
rect 3092 19468 3101 19508
rect 15043 19300 15052 19340
rect 15092 19300 15148 19340
rect 15188 19300 15197 19340
rect 19363 19300 19372 19340
rect 19412 19300 20140 19340
rect 20180 19300 20189 19340
rect 26275 19300 26284 19340
rect 26324 19300 26572 19340
rect 26612 19300 26621 19340
rect 3811 19216 3820 19256
rect 3860 19216 4300 19256
rect 4340 19216 4349 19256
rect 6115 19216 6124 19256
rect 6164 19216 6892 19256
rect 6932 19216 6941 19256
rect 8995 19216 9004 19256
rect 9044 19216 9388 19256
rect 9428 19216 9437 19256
rect 13123 19216 13132 19256
rect 13172 19216 16204 19256
rect 16244 19216 17836 19256
rect 17876 19216 17885 19256
rect 5347 19132 5356 19172
rect 5396 19132 6508 19172
rect 6548 19132 6557 19172
rect 11587 19132 11596 19172
rect 11636 19132 14764 19172
rect 14804 19132 14813 19172
rect 24163 19048 24172 19088
rect 24212 19048 24844 19088
rect 24884 19048 24893 19088
rect 27523 19048 27532 19088
rect 27572 19048 27628 19088
rect 27668 19048 28300 19088
rect 28340 19048 28349 19088
rect 12643 18964 12652 19004
rect 12692 18964 15148 19004
rect 15188 18964 15197 19004
rect 4343 18880 4352 18920
rect 4720 18880 4729 18920
rect 6115 18880 6124 18920
rect 6164 18880 6892 18920
rect 6932 18880 7948 18920
rect 7988 18880 8908 18920
rect 8948 18880 8957 18920
rect 12117 18880 12126 18920
rect 12494 18880 12503 18920
rect 14275 18880 14284 18920
rect 14324 18880 18316 18920
rect 18356 18880 18365 18920
rect 19891 18880 19900 18920
rect 20268 18880 20277 18920
rect 27665 18880 27674 18920
rect 28042 18880 28051 18920
rect 8515 18796 8524 18836
rect 8564 18796 9196 18836
rect 9236 18796 9245 18836
rect 12931 18796 12940 18836
rect 12980 18796 17836 18836
rect 17876 18796 19316 18836
rect 29635 18796 29644 18836
rect 29684 18796 29972 18836
rect 30499 18796 30508 18836
rect 30548 18796 30988 18836
rect 31028 18796 31037 18836
rect 19276 18752 19316 18796
rect 931 18712 940 18752
rect 980 18712 1228 18752
rect 1268 18712 1277 18752
rect 10339 18712 10348 18752
rect 10388 18712 18412 18752
rect 18452 18712 18461 18752
rect 19181 18712 19276 18752
rect 19316 18712 19325 18752
rect 28675 18712 28684 18752
rect 28724 18712 28780 18752
rect 28820 18712 28829 18752
rect 29932 18668 29972 18796
rect 14572 18628 21292 18668
rect 21332 18628 21341 18668
rect 25507 18628 25516 18668
rect 25556 18628 26476 18668
rect 26516 18628 26525 18668
rect 27331 18628 27340 18668
rect 27380 18628 27628 18668
rect 27668 18628 27677 18668
rect 28867 18628 28876 18668
rect 28916 18628 29011 18668
rect 29923 18628 29932 18668
rect 29972 18628 29981 18668
rect 14572 18584 14612 18628
rect 1699 18544 1708 18584
rect 1748 18544 4972 18584
rect 5012 18544 5021 18584
rect 7075 18544 7084 18584
rect 7124 18544 8236 18584
rect 8276 18544 10636 18584
rect 10676 18544 11404 18584
rect 11444 18544 12844 18584
rect 12884 18544 12893 18584
rect 12940 18544 14612 18584
rect 15715 18544 15724 18584
rect 15764 18544 16588 18584
rect 16628 18544 16637 18584
rect 17827 18544 17836 18584
rect 17876 18544 18508 18584
rect 18548 18544 18557 18584
rect 21667 18544 21676 18584
rect 21716 18544 23980 18584
rect 24020 18544 24076 18584
rect 24116 18544 24144 18584
rect 25699 18544 25708 18584
rect 25748 18544 28300 18584
rect 28340 18544 28349 18584
rect 12940 18500 12980 18544
rect 7747 18460 7756 18500
rect 7796 18460 7805 18500
rect 9676 18460 12980 18500
rect 15811 18460 15820 18500
rect 15860 18460 16204 18500
rect 16244 18460 16253 18500
rect 18979 18460 18988 18500
rect 19028 18460 19180 18500
rect 19220 18460 19229 18500
rect 21763 18460 21772 18500
rect 21812 18460 22444 18500
rect 22484 18460 23596 18500
rect 23636 18460 23645 18500
rect 24931 18460 24940 18500
rect 24980 18460 27436 18500
rect 27476 18460 28396 18500
rect 28436 18460 28445 18500
rect 7756 18332 7796 18460
rect 9676 18416 9716 18460
rect 7843 18376 7852 18416
rect 7892 18376 9716 18416
rect 14179 18376 14188 18416
rect 14228 18376 14476 18416
rect 14516 18376 14572 18416
rect 14612 18376 14621 18416
rect 26275 18376 26284 18416
rect 26324 18376 26764 18416
rect 26804 18376 26813 18416
rect 7756 18292 8620 18332
rect 8660 18292 12652 18332
rect 12692 18292 12701 18332
rect 14659 18292 14668 18332
rect 14708 18292 21004 18332
rect 21044 18292 21053 18332
rect 9187 18208 9196 18248
rect 9236 18208 12940 18248
rect 12980 18208 12989 18248
rect 14371 18208 14380 18248
rect 14420 18208 17836 18248
rect 17876 18208 17885 18248
rect 21955 18208 21964 18248
rect 22004 18208 22924 18248
rect 22964 18208 22973 18248
rect 3103 18124 3112 18164
rect 3480 18124 3489 18164
rect 6787 18124 6796 18164
rect 6836 18124 9580 18164
rect 9620 18124 9629 18164
rect 10877 18124 10886 18164
rect 11254 18124 11263 18164
rect 15523 18124 15532 18164
rect 15572 18124 15916 18164
rect 15956 18124 15965 18164
rect 18651 18124 18660 18164
rect 19028 18124 19037 18164
rect 23011 18124 23020 18164
rect 23060 18124 23788 18164
rect 23828 18124 23837 18164
rect 26425 18124 26434 18164
rect 26802 18124 26811 18164
rect 2179 18040 2188 18080
rect 2228 18040 8716 18080
rect 8756 18040 8765 18080
rect 9475 18040 9484 18080
rect 9524 18040 15436 18080
rect 15476 18040 15485 18080
rect 21955 18040 21964 18080
rect 22004 18040 23884 18080
rect 23924 18040 23933 18080
rect 3139 17956 3148 17996
rect 3188 17956 5356 17996
rect 5396 17956 5405 17996
rect 10531 17956 10540 17996
rect 10580 17956 11404 17996
rect 11444 17956 11453 17996
rect 12355 17956 12364 17996
rect 12404 17956 14476 17996
rect 14516 17956 14525 17996
rect 23596 17956 24076 17996
rect 24116 17956 24125 17996
rect 28099 17956 28108 17996
rect 28148 17956 28396 17996
rect 28436 17956 28445 17996
rect 1795 17872 1804 17912
rect 1844 17872 4204 17912
rect 4244 17872 9100 17912
rect 9140 17872 9676 17912
rect 9716 17872 9725 17912
rect 10243 17872 10252 17912
rect 10292 17872 10828 17912
rect 10868 17872 10877 17912
rect 14179 17872 14188 17912
rect 14228 17872 15820 17912
rect 15860 17872 15869 17912
rect 17741 17872 17836 17912
rect 17876 17872 17885 17912
rect 18029 17872 18124 17912
rect 18164 17872 18173 17912
rect 23596 17828 23636 17956
rect 4387 17788 4396 17828
rect 4436 17788 5068 17828
rect 5108 17788 6220 17828
rect 6260 17788 19372 17828
rect 19412 17788 19421 17828
rect 23299 17788 23308 17828
rect 23348 17788 23596 17828
rect 23636 17788 23645 17828
rect 23981 17788 24076 17828
rect 24116 17788 24125 17828
rect 2563 17704 2572 17744
rect 2612 17704 3820 17744
rect 3860 17704 3869 17744
rect 4195 17704 4204 17744
rect 4244 17704 26092 17744
rect 26132 17704 26141 17744
rect 28483 17704 28492 17744
rect 28532 17704 30700 17744
rect 30740 17704 30749 17744
rect 7267 17620 7276 17660
rect 7316 17620 8620 17660
rect 8660 17620 9388 17660
rect 9428 17620 9437 17660
rect 11501 17620 11596 17660
rect 11636 17620 11645 17660
rect 14563 17620 14572 17660
rect 14612 17620 15148 17660
rect 15188 17620 15628 17660
rect 15668 17620 15677 17660
rect 18307 17620 18316 17660
rect 18356 17620 19276 17660
rect 19316 17620 19325 17660
rect 23011 17620 23020 17660
rect 23060 17620 26284 17660
rect 26324 17620 26333 17660
rect 4675 17536 4684 17576
rect 4724 17536 4733 17576
rect 6403 17536 6412 17576
rect 6452 17536 7852 17576
rect 7892 17536 7901 17576
rect 9187 17536 9196 17576
rect 9236 17536 10636 17576
rect 10676 17536 10685 17576
rect 14659 17536 14668 17576
rect 14708 17536 15436 17576
rect 15476 17536 15485 17576
rect 21763 17536 21772 17576
rect 21812 17536 23212 17576
rect 23252 17536 23261 17576
rect 23587 17536 23596 17576
rect 23636 17536 24364 17576
rect 24404 17536 24413 17576
rect 24643 17536 24652 17576
rect 24692 17536 25708 17576
rect 25748 17536 27724 17576
rect 27764 17536 27773 17576
rect 4684 17492 4724 17536
rect 4684 17452 8852 17492
rect 22723 17452 22732 17492
rect 22772 17452 23884 17492
rect 23924 17452 23933 17492
rect 30403 17452 30412 17492
rect 30452 17452 30892 17492
rect 30932 17452 30941 17492
rect 4343 17368 4352 17408
rect 4720 17368 4729 17408
rect 5059 17368 5068 17408
rect 5108 17368 8044 17408
rect 8084 17368 8093 17408
rect 2275 17284 2284 17324
rect 2324 17284 7468 17324
rect 7508 17284 7517 17324
rect 4483 17200 4492 17240
rect 4532 17200 4876 17240
rect 4916 17200 4925 17240
rect 5443 17200 5452 17240
rect 5492 17200 5740 17240
rect 5780 17200 6220 17240
rect 6260 17200 7852 17240
rect 7892 17200 7901 17240
rect 3619 17116 3628 17156
rect 3668 17116 4108 17156
rect 4148 17116 4157 17156
rect 7085 17116 7180 17156
rect 7220 17116 8236 17156
rect 8276 17116 8285 17156
rect 8812 17072 8852 17452
rect 12117 17368 12126 17408
rect 12494 17368 12503 17408
rect 12835 17368 12844 17408
rect 12884 17368 16684 17408
rect 16724 17368 16733 17408
rect 19891 17368 19900 17408
rect 20268 17368 20277 17408
rect 27665 17368 27674 17408
rect 28042 17368 28051 17408
rect 13507 17284 13516 17324
rect 13556 17284 16972 17324
rect 17012 17284 17021 17324
rect 9187 17200 9196 17240
rect 9236 17200 10540 17240
rect 10580 17200 10589 17240
rect 11875 17200 11884 17240
rect 11924 17200 12844 17240
rect 12884 17200 12893 17240
rect 13027 17200 13036 17240
rect 13076 17200 14764 17240
rect 14804 17200 14813 17240
rect 19171 17200 19180 17240
rect 19220 17200 19948 17240
rect 19988 17200 19997 17240
rect 9475 17116 9484 17156
rect 9524 17116 10156 17156
rect 10196 17116 10444 17156
rect 10484 17116 10493 17156
rect 14659 17116 14668 17156
rect 14708 17116 15436 17156
rect 15476 17116 15485 17156
rect 16867 17116 16876 17156
rect 16916 17116 18892 17156
rect 18932 17116 18941 17156
rect 19555 17116 19564 17156
rect 19604 17116 19852 17156
rect 19892 17116 19901 17156
rect 23011 17116 23020 17156
rect 23060 17116 24844 17156
rect 24884 17116 24893 17156
rect 27427 17116 27436 17156
rect 27476 17116 27724 17156
rect 27764 17116 27773 17156
rect 3235 17032 3244 17072
rect 3284 17032 4972 17072
rect 5012 17032 5021 17072
rect 8803 17032 8812 17072
rect 8852 17032 8861 17072
rect 11107 17032 11116 17072
rect 11156 17032 11884 17072
rect 11924 17032 13132 17072
rect 13172 17032 13181 17072
rect 15715 17032 15724 17072
rect 15764 17032 18316 17072
rect 18356 17032 18365 17072
rect 22531 17032 22540 17072
rect 22580 17032 23884 17072
rect 23924 17032 24940 17072
rect 24980 17032 24989 17072
rect 27523 17032 27532 17072
rect 27572 17032 29740 17072
rect 29780 17032 29789 17072
rect 5251 16948 5260 16988
rect 5300 16948 5932 16988
rect 5972 16948 5981 16988
rect 7843 16948 7852 16988
rect 7892 16948 10732 16988
rect 10772 16948 10781 16988
rect 22915 16948 22924 16988
rect 22964 16948 24364 16988
rect 24404 16948 25612 16988
rect 25652 16948 25661 16988
rect 26189 16948 26284 16988
rect 26324 16948 26333 16988
rect 4483 16864 4492 16904
rect 4532 16864 5740 16904
rect 5780 16864 5789 16904
rect 18403 16864 18412 16904
rect 18452 16864 18700 16904
rect 18740 16864 18749 16904
rect 19747 16864 19756 16904
rect 19796 16864 20140 16904
rect 20180 16864 20189 16904
rect 7171 16780 7180 16820
rect 7220 16780 7852 16820
rect 7892 16780 7901 16820
rect 8419 16780 8428 16820
rect 8468 16780 9100 16820
rect 9140 16780 9149 16820
rect 14659 16780 14668 16820
rect 14708 16780 17260 16820
rect 17300 16780 17309 16820
rect 18307 16780 18316 16820
rect 18356 16780 18796 16820
rect 18836 16780 18845 16820
rect 8035 16696 8044 16736
rect 8084 16696 9868 16736
rect 9908 16696 9917 16736
rect 10627 16696 10636 16736
rect 10676 16696 12748 16736
rect 12788 16696 12797 16736
rect 3103 16612 3112 16652
rect 3480 16612 3489 16652
rect 6019 16612 6028 16652
rect 6068 16612 7660 16652
rect 7700 16612 7709 16652
rect 10877 16612 10886 16652
rect 11254 16612 11263 16652
rect 18651 16612 18660 16652
rect 19028 16612 19037 16652
rect 19171 16612 19180 16652
rect 19220 16612 19229 16652
rect 26425 16612 26434 16652
rect 26802 16612 26811 16652
rect 1699 16528 1708 16568
rect 1748 16528 6796 16568
rect 6836 16528 6988 16568
rect 7028 16528 7037 16568
rect 19180 16484 19220 16612
rect 6211 16444 6220 16484
rect 6260 16444 10252 16484
rect 10292 16444 19220 16484
rect 6691 16360 6700 16400
rect 6740 16360 7852 16400
rect 7892 16360 7901 16400
rect 8035 16360 8044 16400
rect 8084 16360 8428 16400
rect 8468 16360 9964 16400
rect 10004 16360 10013 16400
rect 10147 16360 10156 16400
rect 10196 16360 10252 16400
rect 10292 16360 10301 16400
rect 17347 16360 17356 16400
rect 17396 16360 18988 16400
rect 19028 16360 19276 16400
rect 19316 16360 19325 16400
rect 4099 16276 4108 16316
rect 4148 16276 9196 16316
rect 9236 16276 9484 16316
rect 9524 16276 9533 16316
rect 10723 16276 10732 16316
rect 10772 16276 16972 16316
rect 17012 16276 17021 16316
rect 24067 16276 24076 16316
rect 24116 16276 26284 16316
rect 26324 16276 26333 16316
rect 9293 16192 9388 16232
rect 9428 16192 10964 16232
rect 12067 16192 12076 16232
rect 12116 16192 13708 16232
rect 13748 16192 13757 16232
rect 14083 16192 14092 16232
rect 14132 16192 15628 16232
rect 15668 16192 15677 16232
rect 17059 16192 17068 16232
rect 17108 16192 19564 16232
rect 19604 16192 19613 16232
rect 21283 16192 21292 16232
rect 21332 16192 24268 16232
rect 24308 16192 26956 16232
rect 26996 16192 27005 16232
rect 10924 16148 10964 16192
rect 5837 16108 5932 16148
rect 5972 16108 5981 16148
rect 7843 16108 7852 16148
rect 7892 16108 8428 16148
rect 8468 16108 10156 16148
rect 10196 16108 10205 16148
rect 10627 16108 10636 16148
rect 10676 16108 10828 16148
rect 10868 16108 10877 16148
rect 10924 16108 18508 16148
rect 18548 16108 18557 16148
rect 19075 16108 19084 16148
rect 19124 16108 19276 16148
rect 19316 16108 19325 16148
rect 21571 16108 21580 16148
rect 21620 16108 23788 16148
rect 23828 16108 23837 16148
rect 25507 16108 25516 16148
rect 25556 16108 26668 16148
rect 26708 16108 27052 16148
rect 27092 16108 27101 16148
rect 4675 16024 4684 16064
rect 4724 16024 4876 16064
rect 4916 16024 7948 16064
rect 7988 16024 7997 16064
rect 23395 16024 23404 16064
rect 23444 16024 26764 16064
rect 26804 16024 26813 16064
rect 6691 15940 6700 15980
rect 6740 15940 8044 15980
rect 8084 15940 8093 15980
rect 4343 15856 4352 15896
rect 4720 15856 4729 15896
rect 5347 15856 5356 15896
rect 5396 15856 6508 15896
rect 6548 15856 9100 15896
rect 9140 15856 9149 15896
rect 11395 15856 11404 15896
rect 11444 15856 11596 15896
rect 11636 15856 11645 15896
rect 12117 15856 12126 15896
rect 12494 15856 12503 15896
rect 19891 15856 19900 15896
rect 20268 15856 20277 15896
rect 27665 15856 27674 15896
rect 28042 15856 28051 15896
rect 6787 15772 6796 15812
rect 6836 15772 9292 15812
rect 9332 15772 9341 15812
rect 11011 15772 11020 15812
rect 11060 15772 12748 15812
rect 12788 15772 12797 15812
rect 3715 15688 3724 15728
rect 3764 15688 5740 15728
rect 5780 15688 5789 15728
rect 10051 15688 10060 15728
rect 10100 15688 17452 15728
rect 17492 15688 19756 15728
rect 19796 15688 19805 15728
rect 23011 15688 23020 15728
rect 23060 15688 25132 15728
rect 25172 15688 25181 15728
rect 27523 15688 27532 15728
rect 27572 15688 27724 15728
rect 27764 15688 27773 15728
rect 4483 15604 4492 15644
rect 4532 15604 11596 15644
rect 11636 15604 12460 15644
rect 12500 15604 12509 15644
rect 15235 15604 15244 15644
rect 15284 15604 16012 15644
rect 16052 15604 16972 15644
rect 17012 15604 17021 15644
rect 17251 15604 17260 15644
rect 17300 15604 19852 15644
rect 19892 15604 19901 15644
rect 25699 15604 25708 15644
rect 25748 15604 26956 15644
rect 26996 15604 27148 15644
rect 27188 15604 27197 15644
rect 28867 15604 28876 15644
rect 28916 15604 29932 15644
rect 29972 15604 29981 15644
rect 2947 15520 2956 15560
rect 2996 15520 3628 15560
rect 3668 15520 3677 15560
rect 4003 15520 4012 15560
rect 4052 15520 5740 15560
rect 5780 15520 5789 15560
rect 8611 15520 8620 15560
rect 8660 15520 9388 15560
rect 9428 15520 9437 15560
rect 10723 15520 10732 15560
rect 10772 15520 11404 15560
rect 11444 15520 11453 15560
rect 12931 15520 12940 15560
rect 12980 15520 15724 15560
rect 15764 15520 15773 15560
rect 18125 15520 18220 15560
rect 18260 15520 19948 15560
rect 19988 15520 19997 15560
rect 26179 15520 26188 15560
rect 26228 15520 28012 15560
rect 28052 15520 28061 15560
rect 4099 15436 4108 15476
rect 4148 15436 4588 15476
rect 4628 15436 4637 15476
rect 7853 15436 7948 15476
rect 7988 15436 7997 15476
rect 9091 15436 9100 15476
rect 9140 15436 11116 15476
rect 11156 15436 12172 15476
rect 12212 15436 12221 15476
rect 13219 15436 13228 15476
rect 13268 15436 13804 15476
rect 13844 15436 13853 15476
rect 17357 15436 17452 15476
rect 17492 15436 17501 15476
rect 6787 15352 6796 15392
rect 6836 15352 7660 15392
rect 7700 15352 7709 15392
rect 10339 15352 10348 15392
rect 10388 15352 12364 15392
rect 12404 15352 12413 15392
rect 26083 15352 26092 15392
rect 26132 15352 29932 15392
rect 29972 15352 29981 15392
rect 10435 15268 10444 15308
rect 10484 15268 10828 15308
rect 10868 15268 10877 15308
rect 11875 15268 11884 15308
rect 11924 15268 13900 15308
rect 13940 15268 13949 15308
rect 17059 15268 17068 15308
rect 17108 15268 17932 15308
rect 17972 15268 17981 15308
rect 12259 15184 12268 15224
rect 12308 15184 19372 15224
rect 19412 15184 19421 15224
rect 3103 15100 3112 15140
rect 3480 15100 3489 15140
rect 6403 15100 6412 15140
rect 6452 15100 6796 15140
rect 6836 15100 6845 15140
rect 10877 15100 10886 15140
rect 11254 15100 11263 15140
rect 13037 15100 13132 15140
rect 13172 15100 13181 15140
rect 17635 15100 17644 15140
rect 17684 15100 18028 15140
rect 18068 15100 18077 15140
rect 18651 15100 18660 15140
rect 19028 15100 19037 15140
rect 26425 15100 26434 15140
rect 26802 15100 26811 15140
rect 7171 15016 7180 15056
rect 7220 15016 7468 15056
rect 7508 15016 12844 15056
rect 12884 15016 12893 15056
rect 5251 14932 5260 14972
rect 5300 14932 11116 14972
rect 11156 14932 11165 14972
rect 15139 14932 15148 14972
rect 15188 14932 17644 14972
rect 17684 14932 17693 14972
rect 18115 14932 18124 14972
rect 18164 14932 18604 14972
rect 18644 14932 18653 14972
rect 30307 14932 30316 14972
rect 30356 14932 30700 14972
rect 30740 14932 30749 14972
rect 14957 14848 15052 14888
rect 15092 14848 15101 14888
rect 16099 14848 16108 14888
rect 16148 14848 17740 14888
rect 17780 14848 17789 14888
rect 27331 14848 27340 14888
rect 27380 14848 30988 14888
rect 31028 14848 31037 14888
rect 355 14764 364 14804
rect 404 14764 556 14804
rect 596 14764 605 14804
rect 23779 14764 23788 14804
rect 23828 14764 24940 14804
rect 24980 14764 24989 14804
rect 25507 14764 25516 14804
rect 25556 14764 27052 14804
rect 27092 14764 27101 14804
rect 8035 14680 8044 14720
rect 8084 14680 8332 14720
rect 8372 14680 8381 14720
rect 10723 14680 10732 14720
rect 10772 14680 10924 14720
rect 10964 14680 10973 14720
rect 14284 14680 16204 14720
rect 16244 14680 16253 14720
rect 16483 14680 16492 14720
rect 16532 14680 16541 14720
rect 16867 14680 16876 14720
rect 16916 14680 16972 14720
rect 17012 14680 17021 14720
rect 17731 14680 17740 14720
rect 17780 14680 19948 14720
rect 19988 14680 19997 14720
rect 25123 14680 25132 14720
rect 25172 14680 25324 14720
rect 25364 14680 25373 14720
rect 14284 14636 14324 14680
rect 16492 14636 16532 14680
rect 4483 14596 4492 14636
rect 4532 14596 4876 14636
rect 4916 14596 8236 14636
rect 8276 14596 10540 14636
rect 10580 14596 13036 14636
rect 13076 14596 13324 14636
rect 13364 14596 14284 14636
rect 14324 14596 14333 14636
rect 15715 14596 15724 14636
rect 15764 14596 16532 14636
rect 19267 14596 19276 14636
rect 19316 14596 23116 14636
rect 23156 14596 23165 14636
rect 23779 14596 23788 14636
rect 23828 14596 26764 14636
rect 26804 14596 26956 14636
rect 26996 14596 27005 14636
rect 26092 14552 26132 14596
rect 4579 14512 4588 14552
rect 4628 14512 6700 14552
rect 6740 14512 6749 14552
rect 11779 14512 11788 14552
rect 11828 14512 12172 14552
rect 12212 14512 12221 14552
rect 12835 14512 12844 14552
rect 12884 14512 22060 14552
rect 22100 14512 22109 14552
rect 23213 14512 23308 14552
rect 23348 14512 23357 14552
rect 26083 14512 26092 14552
rect 26132 14512 26172 14552
rect 739 14428 748 14468
rect 788 14428 1420 14468
rect 1460 14428 1469 14468
rect 20515 14428 20524 14468
rect 20564 14428 23020 14468
rect 23060 14428 23069 14468
rect 25699 14428 25708 14468
rect 25748 14428 26956 14468
rect 26996 14428 27005 14468
rect 4343 14344 4352 14384
rect 4720 14344 4729 14384
rect 12117 14344 12126 14384
rect 12494 14344 12503 14384
rect 19891 14344 19900 14384
rect 20268 14344 20277 14384
rect 27665 14344 27674 14384
rect 28042 14344 28051 14384
rect 11875 14260 11884 14300
rect 11924 14260 14284 14300
rect 14324 14260 16876 14300
rect 16916 14260 16925 14300
rect 19747 14260 19756 14300
rect 19796 14260 20524 14300
rect 20564 14260 20573 14300
rect 25891 14260 25900 14300
rect 25940 14260 28204 14300
rect 28244 14260 28253 14300
rect 6403 14176 6412 14216
rect 6452 14176 9676 14216
rect 9716 14176 10540 14216
rect 10580 14176 10589 14216
rect 12259 14176 12268 14216
rect 12308 14176 16972 14216
rect 17012 14176 17021 14216
rect 19363 14176 19372 14216
rect 19412 14176 20140 14216
rect 20180 14176 20189 14216
rect 10147 14092 10156 14132
rect 10196 14092 11020 14132
rect 11060 14092 11069 14132
rect 12835 14092 12844 14132
rect 12884 14092 14572 14132
rect 14612 14092 16780 14132
rect 16820 14092 16829 14132
rect 29155 14092 29164 14132
rect 29204 14092 30124 14132
rect 30164 14092 30173 14132
rect 8525 14008 8620 14048
rect 8660 14008 8669 14048
rect 12067 14008 12076 14048
rect 12116 14008 13132 14048
rect 13172 14008 13181 14048
rect 14467 14008 14476 14048
rect 14516 14008 15916 14048
rect 15956 14008 15965 14048
rect 16771 14008 16780 14048
rect 16820 14008 16876 14048
rect 16916 14008 18700 14048
rect 18740 14008 18749 14048
rect 23011 14008 23020 14048
rect 23060 14008 28300 14048
rect 28340 14008 28349 14048
rect 29635 14008 29644 14048
rect 29684 14008 30028 14048
rect 30068 14008 30077 14048
rect 10157 13924 10252 13964
rect 10292 13924 10301 13964
rect 12835 13924 12844 13964
rect 12884 13924 13612 13964
rect 13652 13924 13661 13964
rect 18499 13924 18508 13964
rect 18548 13924 20236 13964
rect 20276 13924 20285 13964
rect 22627 13924 22636 13964
rect 22676 13924 27820 13964
rect 27860 13924 27869 13964
rect 28867 13924 28876 13964
rect 28916 13924 29011 13964
rect 30989 13924 31084 13964
rect 31124 13924 31133 13964
rect 6883 13840 6892 13880
rect 6932 13840 8428 13880
rect 8468 13840 11020 13880
rect 11060 13840 11308 13880
rect 11348 13840 11357 13880
rect 14467 13840 14476 13880
rect 14516 13840 17068 13880
rect 17108 13840 17117 13880
rect 451 13756 460 13796
rect 500 13756 1036 13796
rect 1076 13756 1085 13796
rect 8803 13756 8812 13796
rect 8852 13756 9196 13796
rect 9236 13756 9245 13796
rect 12739 13756 12748 13796
rect 12788 13756 13228 13796
rect 13268 13756 13277 13796
rect 15139 13756 15148 13796
rect 15188 13756 16204 13796
rect 16244 13756 16253 13796
rect 26179 13756 26188 13796
rect 26228 13756 26476 13796
rect 26516 13756 26525 13796
rect 10051 13672 10060 13712
rect 10100 13672 18220 13712
rect 18260 13672 18316 13712
rect 18356 13672 18365 13712
rect 3103 13588 3112 13628
rect 3480 13588 3489 13628
rect 8803 13588 8812 13628
rect 8852 13588 9004 13628
rect 9044 13588 9053 13628
rect 10877 13588 10886 13628
rect 11254 13588 11263 13628
rect 18651 13588 18660 13628
rect 19028 13588 19037 13628
rect 26425 13588 26434 13628
rect 26802 13588 26811 13628
rect 14179 13504 14188 13544
rect 14228 13504 15532 13544
rect 15572 13504 19756 13544
rect 19796 13504 19805 13544
rect 15619 13336 15628 13376
rect 15668 13336 17452 13376
rect 17492 13336 17501 13376
rect 4771 13252 4780 13292
rect 4820 13252 6220 13292
rect 6260 13252 9388 13292
rect 9428 13252 9437 13292
rect 15139 13252 15148 13292
rect 15188 13252 16300 13292
rect 16340 13252 16349 13292
rect 19651 13252 19660 13292
rect 19700 13252 19756 13292
rect 19796 13252 19805 13292
rect 3427 13168 3436 13208
rect 3476 13168 7852 13208
rect 7892 13168 8716 13208
rect 8756 13168 8765 13208
rect 11395 13168 11404 13208
rect 11444 13168 12556 13208
rect 12596 13168 12605 13208
rect 23203 13168 23212 13208
rect 23252 13168 26572 13208
rect 26612 13168 28876 13208
rect 28916 13168 28925 13208
rect 7747 13084 7756 13124
rect 7796 13084 9196 13124
rect 9236 13084 9245 13124
rect 10915 13084 10924 13124
rect 10964 13084 17452 13124
rect 17492 13084 18316 13124
rect 18356 13084 18365 13124
rect 29443 13084 29452 13124
rect 29492 13084 29740 13124
rect 29780 13084 29789 13124
rect 18316 13040 18356 13084
rect 18316 13000 20524 13040
rect 20564 13000 20573 13040
rect 13795 12916 13804 12956
rect 13844 12916 17644 12956
rect 17684 12916 17693 12956
rect 4343 12832 4352 12872
rect 4720 12832 4729 12872
rect 12117 12832 12126 12872
rect 12494 12832 12503 12872
rect 19891 12832 19900 12872
rect 20268 12832 20277 12872
rect 27665 12832 27674 12872
rect 28042 12832 28051 12872
rect 2563 12748 2572 12788
rect 2612 12748 5356 12788
rect 5396 12748 5405 12788
rect 14284 12748 16492 12788
rect 16532 12748 16541 12788
rect 19459 12748 19468 12788
rect 19508 12748 19756 12788
rect 19796 12748 19805 12788
rect 14284 12704 14324 12748
rect 11116 12664 14284 12704
rect 14324 12664 14333 12704
rect 14467 12664 14476 12704
rect 14516 12664 15436 12704
rect 15476 12664 15628 12704
rect 15668 12664 15677 12704
rect 11116 12620 11156 12664
rect 5443 12580 5452 12620
rect 5492 12580 5836 12620
rect 5876 12580 7756 12620
rect 7796 12580 7805 12620
rect 9187 12580 9196 12620
rect 9236 12580 11116 12620
rect 11156 12580 11165 12620
rect 11395 12580 11404 12620
rect 11444 12580 17356 12620
rect 17396 12580 17405 12620
rect 9964 12536 10004 12580
rect 3907 12496 3916 12536
rect 3956 12496 6604 12536
rect 6644 12496 6653 12536
rect 9955 12496 9964 12536
rect 10004 12496 10013 12536
rect 12163 12496 12172 12536
rect 12212 12496 13900 12536
rect 13940 12496 13949 12536
rect 14563 12496 14572 12536
rect 14612 12496 15052 12536
rect 15092 12496 15101 12536
rect 15427 12496 15436 12536
rect 15476 12496 17836 12536
rect 17876 12496 17885 12536
rect 18221 12496 18316 12536
rect 18356 12496 18365 12536
rect 9859 12412 9868 12452
rect 9908 12412 13036 12452
rect 13076 12412 13085 12452
rect 10339 12328 10348 12368
rect 10388 12328 20140 12368
rect 20180 12328 20189 12368
rect 30115 12328 30124 12368
rect 30164 12328 30700 12368
rect 30740 12328 30749 12368
rect 11971 12244 11980 12284
rect 12020 12244 12364 12284
rect 12404 12244 12413 12284
rect 27139 12244 27148 12284
rect 27188 12244 29836 12284
rect 29876 12244 29885 12284
rect 3103 12076 3112 12116
rect 3480 12076 3489 12116
rect 10877 12076 10886 12116
rect 11254 12076 11263 12116
rect 18651 12076 18660 12116
rect 19028 12076 19037 12116
rect 26425 12076 26434 12116
rect 26802 12076 26811 12116
rect 12643 11992 12652 12032
rect 12692 11992 13516 12032
rect 13556 11992 13565 12032
rect 7363 11908 7372 11948
rect 7412 11908 7564 11948
rect 7604 11908 7613 11948
rect 10051 11908 10060 11948
rect 10100 11908 10156 11948
rect 10196 11908 10205 11948
rect 16003 11908 16012 11948
rect 16052 11908 19276 11948
rect 19316 11908 19325 11948
rect 30595 11908 30604 11948
rect 30644 11908 30700 11948
rect 30740 11908 30749 11948
rect 10243 11824 10252 11864
rect 10292 11824 10540 11864
rect 10580 11824 11308 11864
rect 11348 11824 11357 11864
rect 14083 11824 14092 11864
rect 14132 11824 15436 11864
rect 15476 11824 16108 11864
rect 16148 11824 16157 11864
rect 29165 11824 29260 11864
rect 29300 11824 29309 11864
rect 8899 11740 8908 11780
rect 8948 11740 19468 11780
rect 19508 11740 19517 11780
rect 23107 11740 23116 11780
rect 23156 11740 25420 11780
rect 25460 11740 27916 11780
rect 27956 11740 27965 11780
rect 28483 11740 28492 11780
rect 28532 11740 29068 11780
rect 29108 11740 29117 11780
rect 2659 11656 2668 11696
rect 2708 11656 6028 11696
rect 6068 11656 6412 11696
rect 6452 11656 6461 11696
rect 11203 11656 11212 11696
rect 11252 11656 12364 11696
rect 12404 11656 13708 11696
rect 13748 11656 15820 11696
rect 15860 11656 15869 11696
rect 17827 11656 17836 11696
rect 17876 11656 18508 11696
rect 18548 11656 19180 11696
rect 19220 11656 19229 11696
rect 24163 11656 24172 11696
rect 24212 11656 26476 11696
rect 26516 11656 26525 11696
rect 12067 11572 12076 11612
rect 12116 11572 20428 11612
rect 20468 11572 20477 11612
rect 4343 11320 4352 11360
rect 4720 11320 4729 11360
rect 12117 11320 12126 11360
rect 12494 11320 12503 11360
rect 19891 11320 19900 11360
rect 20268 11320 20277 11360
rect 27665 11320 27674 11360
rect 28042 11320 28051 11360
rect 4771 11152 4780 11192
rect 4820 11152 7276 11192
rect 7316 11152 7325 11192
rect 13603 11152 13612 11192
rect 13652 11152 13900 11192
rect 13940 11152 13949 11192
rect 29357 11152 29452 11192
rect 29492 11152 29501 11192
rect 30019 11152 30028 11192
rect 30068 11152 30124 11192
rect 30164 11152 30173 11192
rect 29453 11068 29548 11108
rect 29588 11068 29597 11108
rect 1315 10984 1324 11024
rect 1364 10984 2668 11024
rect 2708 10984 4204 11024
rect 4244 10984 7468 11024
rect 7508 10984 7517 11024
rect 24067 10984 24076 11024
rect 24116 10984 24460 11024
rect 24500 10984 24509 11024
rect 24835 10984 24844 11024
rect 24884 10984 25612 11024
rect 25652 10984 25661 11024
rect 26947 10984 26956 11024
rect 26996 10984 29260 11024
rect 29300 10984 29309 11024
rect 931 10900 940 10940
rect 980 10900 6412 10940
rect 6452 10900 6461 10940
rect 23971 10900 23980 10940
rect 24020 10900 26284 10940
rect 26324 10900 26333 10940
rect 28195 10900 28204 10940
rect 28244 10900 29836 10940
rect 29876 10900 29885 10940
rect 16195 10816 16204 10856
rect 16244 10816 20140 10856
rect 20180 10816 20189 10856
rect 24547 10816 24556 10856
rect 24596 10816 25132 10856
rect 25172 10816 25181 10856
rect 30317 10816 30412 10856
rect 30452 10816 30461 10856
rect 30701 10816 30796 10856
rect 30836 10816 30845 10856
rect 3103 10564 3112 10604
rect 3480 10564 3489 10604
rect 10877 10564 10886 10604
rect 11254 10564 11263 10604
rect 18651 10564 18660 10604
rect 19028 10564 19037 10604
rect 26425 10564 26434 10604
rect 26802 10564 26811 10604
rect 29155 10564 29164 10604
rect 29204 10564 30412 10604
rect 30452 10564 30461 10604
rect 22723 10312 22732 10352
rect 22772 10312 26092 10352
rect 26132 10312 26141 10352
rect 29635 10312 29644 10352
rect 29684 10312 30796 10352
rect 30836 10312 30845 10352
rect 10819 10228 10828 10268
rect 10868 10228 17836 10268
rect 17876 10228 17885 10268
rect 17635 10144 17644 10184
rect 17684 10144 18124 10184
rect 18164 10144 18173 10184
rect 21283 10144 21292 10184
rect 21332 10144 21868 10184
rect 21908 10144 26956 10184
rect 26996 10144 27005 10184
rect 16579 10060 16588 10100
rect 16628 10060 18316 10100
rect 18356 10060 18365 10100
rect 26957 10060 27052 10100
rect 27092 10060 27101 10100
rect 3427 9976 3436 10016
rect 3476 9976 3628 10016
rect 3668 9976 4972 10016
rect 5012 9976 5021 10016
rect 13987 9976 13996 10016
rect 14036 9976 18508 10016
rect 18548 9976 18557 10016
rect 4343 9808 4352 9848
rect 4720 9808 4729 9848
rect 12117 9808 12126 9848
rect 12494 9808 12503 9848
rect 19891 9808 19900 9848
rect 20268 9808 20277 9848
rect 27665 9808 27674 9848
rect 28042 9808 28051 9848
rect 26179 9556 26188 9596
rect 26228 9556 26284 9596
rect 26324 9556 26333 9596
rect 5837 9472 5932 9512
rect 5972 9472 5981 9512
rect 22435 9472 22444 9512
rect 22484 9472 23212 9512
rect 23252 9472 23261 9512
rect 26275 9304 26284 9344
rect 26324 9304 27052 9344
rect 27092 9304 27101 9344
rect 3103 9052 3112 9092
rect 3480 9052 3489 9092
rect 10877 9052 10886 9092
rect 11254 9052 11263 9092
rect 18651 9052 18660 9092
rect 19028 9052 19037 9092
rect 26425 9052 26434 9092
rect 26802 9052 26811 9092
rect 3331 8800 3340 8840
rect 3380 8800 3628 8840
rect 3668 8800 3677 8840
rect 10435 8800 10444 8840
rect 10484 8800 10828 8840
rect 10868 8800 10877 8840
rect 11683 8632 11692 8672
rect 11732 8632 12268 8672
rect 12308 8632 12844 8672
rect 12884 8632 12893 8672
rect 18499 8548 18508 8588
rect 18548 8548 19660 8588
rect 19700 8548 19948 8588
rect 19988 8548 19997 8588
rect 9379 8380 9388 8420
rect 9428 8380 9676 8420
rect 9716 8380 9725 8420
rect 4343 8296 4352 8336
rect 4720 8296 4729 8336
rect 12117 8296 12126 8336
rect 12494 8296 12503 8336
rect 19891 8296 19900 8336
rect 20268 8296 20277 8336
rect 27665 8296 27674 8336
rect 28042 8296 28051 8336
rect 22915 8128 22924 8168
rect 22964 8128 26188 8168
rect 26228 8128 26237 8168
rect 11203 8044 11212 8084
rect 11252 8044 12268 8084
rect 12308 8044 12317 8084
rect 24355 8044 24364 8084
rect 24404 8044 25324 8084
rect 25364 8044 25373 8084
rect 23587 7960 23596 8000
rect 23636 7960 24172 8000
rect 24212 7960 25036 8000
rect 25076 7960 25085 8000
rect 10051 7708 10060 7748
rect 10100 7708 12076 7748
rect 12116 7708 12125 7748
rect 3103 7540 3112 7580
rect 3480 7540 3489 7580
rect 10877 7540 10886 7580
rect 11254 7540 11263 7580
rect 18651 7540 18660 7580
rect 19028 7540 19037 7580
rect 26425 7540 26434 7580
rect 26802 7540 26811 7580
rect 21763 7204 21772 7244
rect 21812 7204 26380 7244
rect 26420 7204 26429 7244
rect 11107 7120 11116 7160
rect 11156 7120 11884 7160
rect 11924 7120 11933 7160
rect 20515 7120 20524 7160
rect 20564 7120 23692 7160
rect 23732 7120 23741 7160
rect 23011 7036 23020 7076
rect 23060 7036 24460 7076
rect 24500 7036 24509 7076
rect 18979 6868 18988 6908
rect 19028 6868 23212 6908
rect 23252 6868 23261 6908
rect 4343 6784 4352 6824
rect 4720 6784 4729 6824
rect 12117 6784 12126 6824
rect 12494 6784 12503 6824
rect 19891 6784 19900 6824
rect 20268 6784 20277 6824
rect 27665 6784 27674 6824
rect 28042 6784 28051 6824
rect 11587 6448 11596 6488
rect 11636 6448 12268 6488
rect 12308 6448 13612 6488
rect 13652 6448 13661 6488
rect 23683 6448 23692 6488
rect 23732 6448 24076 6488
rect 24116 6448 24125 6488
rect 10051 6112 10060 6152
rect 10100 6112 12652 6152
rect 12692 6112 12701 6152
rect 3103 6028 3112 6068
rect 3480 6028 3489 6068
rect 10877 6028 10886 6068
rect 11254 6028 11263 6068
rect 18651 6028 18660 6068
rect 19028 6028 19037 6068
rect 26425 6028 26434 6068
rect 26802 6028 26811 6068
rect 67 5944 76 5984
rect 116 5944 460 5984
rect 500 5944 509 5984
rect 3907 5608 3916 5648
rect 3956 5608 4780 5648
rect 4820 5608 6220 5648
rect 6260 5608 6269 5648
rect 4343 5272 4352 5312
rect 4720 5272 4729 5312
rect 12117 5272 12126 5312
rect 12494 5272 12503 5312
rect 19891 5272 19900 5312
rect 20268 5272 20277 5312
rect 27665 5272 27674 5312
rect 28042 5272 28051 5312
rect 12557 5020 12652 5060
rect 12692 5020 12701 5060
rect 3103 4516 3112 4556
rect 3480 4516 3489 4556
rect 10877 4516 10886 4556
rect 11254 4516 11263 4556
rect 18651 4516 18660 4556
rect 19028 4516 19037 4556
rect 26425 4516 26434 4556
rect 26802 4516 26811 4556
rect 4343 3760 4352 3800
rect 4720 3760 4729 3800
rect 12117 3760 12126 3800
rect 12494 3760 12503 3800
rect 19891 3760 19900 3800
rect 20268 3760 20277 3800
rect 27665 3760 27674 3800
rect 28042 3760 28051 3800
rect 3103 3004 3112 3044
rect 3480 3004 3489 3044
rect 10877 3004 10886 3044
rect 11254 3004 11263 3044
rect 18651 3004 18660 3044
rect 19028 3004 19037 3044
rect 26425 3004 26434 3044
rect 26802 3004 26811 3044
rect 4343 2248 4352 2288
rect 4720 2248 4729 2288
rect 12117 2248 12126 2288
rect 12494 2248 12503 2288
rect 19891 2248 19900 2288
rect 20268 2248 20277 2288
rect 27665 2248 27674 2288
rect 28042 2248 28051 2288
rect 3103 1492 3112 1532
rect 3480 1492 3489 1532
rect 10877 1492 10886 1532
rect 11254 1492 11263 1532
rect 18651 1492 18660 1532
rect 19028 1492 19037 1532
rect 26425 1492 26434 1532
rect 26802 1492 26811 1532
rect 4343 736 4352 776
rect 4720 736 4729 776
rect 12117 736 12126 776
rect 12494 736 12503 776
rect 19891 736 19900 776
rect 20268 736 20277 776
rect 27665 736 27674 776
rect 28042 736 28051 776
<< via4 >>
rect 27436 28036 27476 28076
rect 4352 27952 4720 27992
rect 12126 27952 12494 27992
rect 19900 27952 20268 27992
rect 27674 27952 28042 27992
rect 10156 27700 10196 27740
rect 27340 27532 27380 27572
rect 11500 27364 11540 27404
rect 28492 27364 28532 27404
rect 31084 27364 31124 27404
rect 3112 27196 3480 27236
rect 10886 27196 11254 27236
rect 18660 27196 19028 27236
rect 26434 27196 26802 27236
rect 30124 26860 30164 26900
rect 4352 26440 4720 26480
rect 12126 26440 12494 26480
rect 19900 26440 20268 26480
rect 27674 26440 28042 26480
rect 28204 26272 28244 26312
rect 18412 26188 18452 26228
rect 20812 26104 20852 26144
rect 29164 26020 29204 26060
rect 27532 25936 27572 25976
rect 30028 25936 30068 25976
rect 3112 25684 3480 25724
rect 10886 25684 11254 25724
rect 18660 25684 19028 25724
rect 26434 25684 26802 25724
rect 10156 25600 10196 25640
rect 10732 25264 10772 25304
rect 26188 25180 26228 25220
rect 29548 25096 29588 25136
rect 20812 25012 20852 25052
rect 4352 24928 4720 24968
rect 12126 24928 12494 24968
rect 19900 24928 20268 24968
rect 27674 24928 28042 24968
rect 26092 24760 26132 24800
rect 18412 24508 18452 24548
rect 29452 24508 29492 24548
rect 29644 24508 29684 24548
rect 27148 24340 27188 24380
rect 27052 24256 27092 24296
rect 3112 24172 3480 24212
rect 10886 24172 11254 24212
rect 18660 24172 19028 24212
rect 26434 24172 26802 24212
rect 10732 23836 10772 23876
rect 12652 23836 12692 23876
rect 20428 23836 20468 23876
rect 30796 23836 30836 23876
rect 16780 23752 16820 23792
rect 29260 23752 29300 23792
rect 26956 23584 26996 23624
rect 4352 23416 4720 23456
rect 12126 23416 12494 23456
rect 19900 23416 20268 23456
rect 27674 23416 28042 23456
rect 30316 23332 30356 23372
rect 20428 23248 20468 23288
rect 27148 23248 27188 23288
rect 27244 23164 27284 23204
rect 30604 23080 30644 23120
rect 20812 22996 20852 23036
rect 11788 22912 11828 22952
rect 26092 22912 26132 22952
rect 4204 22744 4244 22784
rect 3112 22660 3480 22700
rect 10886 22660 11254 22700
rect 18660 22660 19028 22700
rect 26434 22660 26802 22700
rect 4012 22492 4052 22532
rect 11788 22492 11828 22532
rect 30412 22324 30452 22364
rect 8524 22072 8564 22112
rect 4352 21904 4720 21944
rect 12126 21904 12494 21944
rect 19900 21904 20268 21944
rect 27674 21904 28042 21944
rect 76 21736 116 21776
rect 460 21652 500 21692
rect 8524 21568 8564 21608
rect 28684 21568 28724 21608
rect 3112 21148 3480 21188
rect 10886 21148 11254 21188
rect 18660 21148 19028 21188
rect 26434 21148 26802 21188
rect 27244 21064 27284 21104
rect 4204 20980 4244 21020
rect 4012 20812 4052 20852
rect 8524 20812 8564 20852
rect 460 20560 500 20600
rect 27052 20476 27092 20516
rect 4352 20392 4720 20432
rect 12126 20392 12494 20432
rect 19900 20392 20268 20432
rect 27674 20392 28042 20432
rect 27436 20224 27476 20264
rect 11500 20140 11540 20180
rect 14476 20140 14516 20180
rect 16972 20140 17012 20180
rect 27532 20056 27572 20096
rect 25516 19972 25556 20012
rect 27148 19972 27188 20012
rect 26284 19888 26324 19928
rect 3112 19636 3480 19676
rect 10886 19636 11254 19676
rect 18660 19636 19028 19676
rect 26434 19636 26802 19676
rect 15052 19300 15092 19340
rect 26284 19300 26324 19340
rect 17836 19216 17876 19256
rect 27532 19048 27572 19088
rect 4352 18880 4720 18920
rect 7948 18880 7988 18920
rect 12126 18880 12494 18920
rect 19900 18880 20268 18920
rect 27674 18880 28042 18920
rect 19276 18712 19316 18752
rect 28684 18712 28724 18752
rect 28876 18628 28916 18668
rect 10636 18544 10676 18584
rect 24076 18544 24116 18584
rect 19180 18460 19220 18500
rect 14476 18376 14516 18416
rect 26284 18376 26324 18416
rect 8620 18292 8660 18332
rect 3112 18124 3480 18164
rect 10886 18124 11254 18164
rect 18660 18124 19028 18164
rect 26434 18124 26802 18164
rect 17836 17872 17876 17912
rect 18124 17872 18164 17912
rect 23308 17788 23348 17828
rect 24076 17788 24116 17828
rect 28492 17704 28532 17744
rect 9388 17620 9428 17660
rect 11596 17620 11636 17660
rect 4352 17368 4720 17408
rect 4876 17200 4916 17240
rect 7180 17116 7220 17156
rect 12126 17368 12494 17408
rect 19900 17368 20268 17408
rect 27674 17368 28042 17408
rect 19180 17200 19220 17240
rect 10156 17116 10196 17156
rect 13132 17032 13172 17072
rect 27532 17032 27572 17072
rect 10732 16948 10772 16988
rect 26284 16948 26324 16988
rect 19756 16864 19796 16904
rect 7180 16780 7220 16820
rect 18316 16780 18356 16820
rect 3112 16612 3480 16652
rect 10886 16612 11254 16652
rect 18660 16612 19028 16652
rect 26434 16612 26802 16652
rect 10252 16444 10292 16484
rect 10156 16360 10196 16400
rect 17356 16360 17396 16400
rect 19276 16360 19316 16400
rect 10732 16276 10772 16316
rect 9388 16192 9428 16232
rect 5932 16108 5972 16148
rect 10156 16108 10196 16148
rect 10636 16108 10676 16148
rect 25516 16108 25556 16148
rect 27052 16108 27092 16148
rect 7948 16024 7988 16064
rect 4352 15856 4720 15896
rect 12126 15856 12494 15896
rect 19900 15856 20268 15896
rect 27674 15856 28042 15896
rect 27532 15688 27572 15728
rect 11596 15604 11636 15644
rect 28876 15604 28916 15644
rect 9388 15520 9428 15560
rect 18220 15520 18260 15560
rect 7948 15436 7988 15476
rect 17452 15436 17492 15476
rect 3112 15100 3480 15140
rect 10886 15100 11254 15140
rect 13132 15100 13172 15140
rect 18660 15100 19028 15140
rect 26434 15100 26802 15140
rect 7180 15016 7220 15056
rect 18124 14932 18164 14972
rect 30316 14932 30356 14972
rect 15052 14848 15092 14888
rect 27340 14848 27380 14888
rect 10732 14680 10772 14720
rect 16972 14680 17012 14720
rect 4876 14596 4916 14636
rect 23308 14512 23348 14552
rect 4352 14344 4720 14384
rect 12126 14344 12494 14384
rect 19900 14344 20268 14384
rect 27674 14344 28042 14384
rect 10156 14092 10196 14132
rect 8620 14008 8660 14048
rect 16780 14008 16820 14048
rect 10252 13924 10292 13964
rect 28876 13924 28916 13964
rect 31084 13924 31124 13964
rect 18220 13672 18260 13712
rect 3112 13588 3480 13628
rect 10886 13588 11254 13628
rect 18660 13588 19028 13628
rect 26434 13588 26802 13628
rect 19756 13504 19796 13544
rect 19756 13252 19796 13292
rect 28876 13168 28916 13208
rect 17452 13084 17492 13124
rect 4352 12832 4720 12872
rect 12126 12832 12494 12872
rect 19900 12832 20268 12872
rect 27674 12832 28042 12872
rect 19756 12748 19796 12788
rect 17356 12580 17396 12620
rect 18316 12496 18356 12536
rect 30124 12328 30164 12368
rect 27148 12244 27188 12284
rect 3112 12076 3480 12116
rect 10886 12076 11254 12116
rect 18660 12076 19028 12116
rect 26434 12076 26802 12116
rect 10156 11908 10196 11948
rect 30604 11908 30644 11948
rect 29260 11824 29300 11864
rect 4352 11320 4720 11360
rect 12126 11320 12494 11360
rect 19900 11320 20268 11360
rect 27674 11320 28042 11360
rect 29452 11152 29492 11192
rect 30028 11152 30068 11192
rect 29548 11068 29588 11108
rect 26956 10984 26996 11024
rect 28204 10900 28244 10940
rect 30412 10816 30452 10856
rect 30796 10816 30836 10856
rect 3112 10564 3480 10604
rect 10886 10564 11254 10604
rect 18660 10564 19028 10604
rect 26434 10564 26802 10604
rect 29164 10564 29204 10604
rect 29644 10312 29684 10352
rect 27052 10060 27092 10100
rect 4352 9808 4720 9848
rect 12126 9808 12494 9848
rect 19900 9808 20268 9848
rect 27674 9808 28042 9848
rect 26188 9556 26228 9596
rect 5932 9472 5972 9512
rect 3112 9052 3480 9092
rect 10886 9052 11254 9092
rect 18660 9052 19028 9092
rect 26434 9052 26802 9092
rect 4352 8296 4720 8336
rect 12126 8296 12494 8336
rect 19900 8296 20268 8336
rect 27674 8296 28042 8336
rect 3112 7540 3480 7580
rect 10886 7540 11254 7580
rect 18660 7540 19028 7580
rect 26434 7540 26802 7580
rect 4352 6784 4720 6824
rect 12126 6784 12494 6824
rect 19900 6784 20268 6824
rect 27674 6784 28042 6824
rect 12652 6112 12692 6152
rect 3112 6028 3480 6068
rect 10886 6028 11254 6068
rect 18660 6028 19028 6068
rect 26434 6028 26802 6068
rect 76 5944 116 5984
rect 4352 5272 4720 5312
rect 12126 5272 12494 5312
rect 19900 5272 20268 5312
rect 27674 5272 28042 5312
rect 12652 5020 12692 5060
rect 3112 4516 3480 4556
rect 10886 4516 11254 4556
rect 18660 4516 19028 4556
rect 26434 4516 26802 4556
rect 4352 3760 4720 3800
rect 12126 3760 12494 3800
rect 19900 3760 20268 3800
rect 27674 3760 28042 3800
rect 3112 3004 3480 3044
rect 10886 3004 11254 3044
rect 18660 3004 19028 3044
rect 26434 3004 26802 3044
rect 4352 2248 4720 2288
rect 12126 2248 12494 2288
rect 19900 2248 20268 2288
rect 27674 2248 28042 2288
rect 3112 1492 3480 1532
rect 10886 1492 11254 1532
rect 18660 1492 19028 1532
rect 26434 1492 26802 1532
rect 4352 736 4720 776
rect 12126 736 12494 776
rect 19900 736 20268 776
rect 27674 736 28042 776
<< metal5 >>
rect 27436 28076 27476 28085
rect 3076 27236 3516 28016
rect 3076 27196 3112 27236
rect 3480 27196 3516 27236
rect 3076 25724 3516 27196
rect 3076 25684 3112 25724
rect 3480 25684 3516 25724
rect 3076 24212 3516 25684
rect 3076 24172 3112 24212
rect 3480 24172 3516 24212
rect 3076 22700 3516 24172
rect 4316 27992 4756 28016
rect 4316 27952 4352 27992
rect 4720 27952 4756 27992
rect 4316 26480 4756 27952
rect 4316 26440 4352 26480
rect 4720 26440 4756 26480
rect 4316 24968 4756 26440
rect 10156 27740 10196 27749
rect 10156 25640 10196 27700
rect 10156 25591 10196 25600
rect 10850 27236 11290 28016
rect 12090 27992 12530 28016
rect 12090 27952 12126 27992
rect 12494 27952 12530 27992
rect 10850 27196 10886 27236
rect 11254 27196 11290 27236
rect 10850 25724 11290 27196
rect 10850 25684 10886 25724
rect 11254 25684 11290 25724
rect 4316 24928 4352 24968
rect 4720 24928 4756 24968
rect 4316 23456 4756 24928
rect 10732 25304 10772 25313
rect 10732 23876 10772 25264
rect 10732 23827 10772 23836
rect 10850 24212 11290 25684
rect 10850 24172 10886 24212
rect 11254 24172 11290 24212
rect 4316 23416 4352 23456
rect 4720 23416 4756 23456
rect 3076 22660 3112 22700
rect 3480 22660 3516 22700
rect 76 21776 116 21785
rect 76 5984 116 21736
rect 460 21692 500 21701
rect 460 20600 500 21652
rect 460 20551 500 20560
rect 3076 21188 3516 22660
rect 4204 22784 4244 22793
rect 3076 21148 3112 21188
rect 3480 21148 3516 21188
rect 76 5935 116 5944
rect 3076 19676 3516 21148
rect 4012 22532 4052 22541
rect 4012 20852 4052 22492
rect 4204 21020 4244 22744
rect 4204 20971 4244 20980
rect 4316 21944 4756 23416
rect 10850 22700 11290 24172
rect 10850 22660 10886 22700
rect 11254 22660 11290 22700
rect 4316 21904 4352 21944
rect 4720 21904 4756 21944
rect 4012 20803 4052 20812
rect 3076 19636 3112 19676
rect 3480 19636 3516 19676
rect 3076 18164 3516 19636
rect 3076 18124 3112 18164
rect 3480 18124 3516 18164
rect 3076 16652 3516 18124
rect 3076 16612 3112 16652
rect 3480 16612 3516 16652
rect 3076 15140 3516 16612
rect 3076 15100 3112 15140
rect 3480 15100 3516 15140
rect 3076 13628 3516 15100
rect 3076 13588 3112 13628
rect 3480 13588 3516 13628
rect 3076 12116 3516 13588
rect 3076 12076 3112 12116
rect 3480 12076 3516 12116
rect 3076 10604 3516 12076
rect 3076 10564 3112 10604
rect 3480 10564 3516 10604
rect 3076 9092 3516 10564
rect 3076 9052 3112 9092
rect 3480 9052 3516 9092
rect 3076 7580 3516 9052
rect 3076 7540 3112 7580
rect 3480 7540 3516 7580
rect 3076 6068 3516 7540
rect 3076 6028 3112 6068
rect 3480 6028 3516 6068
rect 3076 4556 3516 6028
rect 3076 4516 3112 4556
rect 3480 4516 3516 4556
rect 3076 3044 3516 4516
rect 3076 3004 3112 3044
rect 3480 3004 3516 3044
rect 3076 1532 3516 3004
rect 3076 1492 3112 1532
rect 3480 1492 3516 1532
rect 3076 712 3516 1492
rect 4316 20432 4756 21904
rect 8524 22112 8564 22121
rect 8524 21608 8564 22072
rect 8524 20852 8564 21568
rect 8524 20803 8564 20812
rect 10850 21188 11290 22660
rect 10850 21148 10886 21188
rect 11254 21148 11290 21188
rect 4316 20392 4352 20432
rect 4720 20392 4756 20432
rect 4316 18920 4756 20392
rect 10850 19676 11290 21148
rect 11500 27404 11540 27413
rect 11500 20180 11540 27364
rect 12090 26480 12530 27952
rect 12090 26440 12126 26480
rect 12494 26440 12530 26480
rect 12090 24968 12530 26440
rect 18624 27236 19064 28016
rect 18624 27196 18660 27236
rect 19028 27196 19064 27236
rect 12090 24928 12126 24968
rect 12494 24928 12530 24968
rect 12090 23456 12530 24928
rect 18412 26228 18452 26237
rect 18412 24548 18452 26188
rect 18412 24499 18452 24508
rect 18624 25724 19064 27196
rect 18624 25684 18660 25724
rect 19028 25684 19064 25724
rect 18624 24212 19064 25684
rect 18624 24172 18660 24212
rect 19028 24172 19064 24212
rect 12090 23416 12126 23456
rect 12494 23416 12530 23456
rect 11788 22952 11828 22961
rect 11788 22532 11828 22912
rect 11788 22483 11828 22492
rect 11500 20131 11540 20140
rect 12090 21944 12530 23416
rect 12090 21904 12126 21944
rect 12494 21904 12530 21944
rect 12090 20432 12530 21904
rect 12090 20392 12126 20432
rect 12494 20392 12530 20432
rect 10850 19636 10886 19676
rect 11254 19636 11290 19676
rect 4316 18880 4352 18920
rect 4720 18880 4756 18920
rect 4316 17408 4756 18880
rect 4316 17368 4352 17408
rect 4720 17368 4756 17408
rect 4316 15896 4756 17368
rect 7948 18920 7988 18929
rect 4316 15856 4352 15896
rect 4720 15856 4756 15896
rect 4316 14384 4756 15856
rect 4876 17240 4916 17249
rect 4876 14636 4916 17200
rect 7180 17156 7220 17165
rect 7180 16820 7220 17116
rect 4876 14587 4916 14596
rect 5932 16148 5972 16157
rect 4316 14344 4352 14384
rect 4720 14344 4756 14384
rect 4316 12872 4756 14344
rect 4316 12832 4352 12872
rect 4720 12832 4756 12872
rect 4316 11360 4756 12832
rect 4316 11320 4352 11360
rect 4720 11320 4756 11360
rect 4316 9848 4756 11320
rect 4316 9808 4352 9848
rect 4720 9808 4756 9848
rect 4316 8336 4756 9808
rect 5932 9512 5972 16108
rect 7180 15056 7220 16780
rect 7948 16064 7988 18880
rect 10636 18584 10676 18593
rect 7948 15476 7988 16024
rect 7948 15427 7988 15436
rect 8620 18332 8660 18341
rect 7180 15007 7220 15016
rect 8620 14048 8660 18292
rect 9388 17660 9428 17669
rect 9388 16232 9428 17620
rect 9388 15560 9428 16192
rect 10156 17156 10196 17165
rect 10156 16400 10196 17116
rect 10156 16148 10196 16360
rect 10156 16099 10196 16108
rect 10252 16484 10292 16493
rect 9388 15511 9428 15520
rect 8620 13999 8660 14008
rect 10156 14132 10196 14141
rect 10156 11948 10196 14092
rect 10252 13964 10292 16444
rect 10636 16148 10676 18544
rect 10850 18164 11290 19636
rect 10850 18124 10886 18164
rect 11254 18124 11290 18164
rect 10636 16099 10676 16108
rect 10732 16988 10772 16997
rect 10732 16316 10772 16948
rect 10732 14720 10772 16276
rect 10732 14671 10772 14680
rect 10850 16652 11290 18124
rect 12090 18920 12530 20392
rect 12090 18880 12126 18920
rect 12494 18880 12530 18920
rect 10850 16612 10886 16652
rect 11254 16612 11290 16652
rect 10850 15140 11290 16612
rect 11596 17660 11636 17669
rect 11596 15644 11636 17620
rect 11596 15595 11636 15604
rect 12090 17408 12530 18880
rect 12090 17368 12126 17408
rect 12494 17368 12530 17408
rect 12090 15896 12530 17368
rect 12090 15856 12126 15896
rect 12494 15856 12530 15896
rect 10850 15100 10886 15140
rect 11254 15100 11290 15140
rect 10252 13915 10292 13924
rect 10156 11899 10196 11908
rect 10850 13628 11290 15100
rect 10850 13588 10886 13628
rect 11254 13588 11290 13628
rect 10850 12116 11290 13588
rect 10850 12076 10886 12116
rect 11254 12076 11290 12116
rect 5932 9463 5972 9472
rect 10850 10604 11290 12076
rect 10850 10564 10886 10604
rect 11254 10564 11290 10604
rect 4316 8296 4352 8336
rect 4720 8296 4756 8336
rect 4316 6824 4756 8296
rect 4316 6784 4352 6824
rect 4720 6784 4756 6824
rect 4316 5312 4756 6784
rect 4316 5272 4352 5312
rect 4720 5272 4756 5312
rect 4316 3800 4756 5272
rect 4316 3760 4352 3800
rect 4720 3760 4756 3800
rect 4316 2288 4756 3760
rect 4316 2248 4352 2288
rect 4720 2248 4756 2288
rect 4316 776 4756 2248
rect 4316 736 4352 776
rect 4720 736 4756 776
rect 4316 712 4756 736
rect 10850 9092 11290 10564
rect 10850 9052 10886 9092
rect 11254 9052 11290 9092
rect 10850 7580 11290 9052
rect 10850 7540 10886 7580
rect 11254 7540 11290 7580
rect 10850 6068 11290 7540
rect 10850 6028 10886 6068
rect 11254 6028 11290 6068
rect 10850 4556 11290 6028
rect 10850 4516 10886 4556
rect 11254 4516 11290 4556
rect 10850 3044 11290 4516
rect 10850 3004 10886 3044
rect 11254 3004 11290 3044
rect 10850 1532 11290 3004
rect 10850 1492 10886 1532
rect 11254 1492 11290 1532
rect 10850 712 11290 1492
rect 12090 14384 12530 15856
rect 12090 14344 12126 14384
rect 12494 14344 12530 14384
rect 12090 12872 12530 14344
rect 12090 12832 12126 12872
rect 12494 12832 12530 12872
rect 12090 11360 12530 12832
rect 12090 11320 12126 11360
rect 12494 11320 12530 11360
rect 12090 9848 12530 11320
rect 12090 9808 12126 9848
rect 12494 9808 12530 9848
rect 12090 8336 12530 9808
rect 12090 8296 12126 8336
rect 12494 8296 12530 8336
rect 12090 6824 12530 8296
rect 12090 6784 12126 6824
rect 12494 6784 12530 6824
rect 12090 5312 12530 6784
rect 12090 5272 12126 5312
rect 12494 5272 12530 5312
rect 12090 3800 12530 5272
rect 12652 23876 12692 23885
rect 12652 6152 12692 23836
rect 16780 23792 16820 23801
rect 14476 20180 14516 20189
rect 14476 18416 14516 20140
rect 14476 18367 14516 18376
rect 15052 19340 15092 19349
rect 13132 17072 13172 17081
rect 13132 15140 13172 17032
rect 13132 15091 13172 15100
rect 15052 14888 15092 19300
rect 15052 14839 15092 14848
rect 16780 14048 16820 23752
rect 18624 22700 19064 24172
rect 18624 22660 18660 22700
rect 19028 22660 19064 22700
rect 18624 21188 19064 22660
rect 18624 21148 18660 21188
rect 19028 21148 19064 21188
rect 16972 20180 17012 20189
rect 16972 14720 17012 20140
rect 18624 19676 19064 21148
rect 18624 19636 18660 19676
rect 19028 19636 19064 19676
rect 17836 19256 17876 19265
rect 17836 17912 17876 19216
rect 18624 18164 19064 19636
rect 19864 27992 20304 28016
rect 19864 27952 19900 27992
rect 20268 27952 20304 27992
rect 19864 26480 20304 27952
rect 19864 26440 19900 26480
rect 20268 26440 20304 26480
rect 19864 24968 20304 26440
rect 26398 27236 26838 28016
rect 26398 27196 26434 27236
rect 26802 27196 26838 27236
rect 19864 24928 19900 24968
rect 20268 24928 20304 24968
rect 19864 23456 20304 24928
rect 20812 26144 20852 26153
rect 20812 25052 20852 26104
rect 26398 25724 26838 27196
rect 26398 25684 26434 25724
rect 26802 25684 26838 25724
rect 19864 23416 19900 23456
rect 20268 23416 20304 23456
rect 19864 21944 20304 23416
rect 20428 23876 20468 23885
rect 20428 23288 20468 23836
rect 20428 23239 20468 23248
rect 20812 23036 20852 25012
rect 26188 25220 26228 25229
rect 20812 22987 20852 22996
rect 26092 24800 26132 24809
rect 26092 22952 26132 24760
rect 26092 22903 26132 22912
rect 19864 21904 19900 21944
rect 20268 21904 20304 21944
rect 19864 20432 20304 21904
rect 19864 20392 19900 20432
rect 20268 20392 20304 20432
rect 19864 18920 20304 20392
rect 19864 18880 19900 18920
rect 20268 18880 20304 18920
rect 19276 18752 19316 18761
rect 18624 18124 18660 18164
rect 19028 18124 19064 18164
rect 17836 17863 17876 17872
rect 18124 17912 18164 17921
rect 16972 14671 17012 14680
rect 17356 16400 17396 16409
rect 16780 13999 16820 14008
rect 17356 12620 17396 16360
rect 17452 15476 17492 15485
rect 17452 13124 17492 15436
rect 18124 14972 18164 17872
rect 18316 16820 18356 16829
rect 18124 14923 18164 14932
rect 18220 15560 18260 15569
rect 18220 13712 18260 15520
rect 18220 13663 18260 13672
rect 17452 13075 17492 13084
rect 17356 12571 17396 12580
rect 18316 12536 18356 16780
rect 18316 12487 18356 12496
rect 18624 16652 19064 18124
rect 19180 18500 19220 18509
rect 19180 17240 19220 18460
rect 19180 17191 19220 17200
rect 18624 16612 18660 16652
rect 19028 16612 19064 16652
rect 18624 15140 19064 16612
rect 19276 16400 19316 18712
rect 19864 17408 20304 18880
rect 25516 20012 25556 20021
rect 24076 18584 24116 18593
rect 19864 17368 19900 17408
rect 20268 17368 20304 17408
rect 19276 16351 19316 16360
rect 19756 16904 19796 16913
rect 18624 15100 18660 15140
rect 19028 15100 19064 15140
rect 18624 13628 19064 15100
rect 18624 13588 18660 13628
rect 19028 13588 19064 13628
rect 12652 5060 12692 6112
rect 12652 5011 12692 5020
rect 18624 12116 19064 13588
rect 19756 13544 19796 16864
rect 19756 13495 19796 13504
rect 19864 15896 20304 17368
rect 19864 15856 19900 15896
rect 20268 15856 20304 15896
rect 19864 14384 20304 15856
rect 23308 17828 23348 17837
rect 23308 14552 23348 17788
rect 24076 17828 24116 18544
rect 24076 17779 24116 17788
rect 25516 16148 25556 19972
rect 25516 16099 25556 16108
rect 23308 14503 23348 14512
rect 19864 14344 19900 14384
rect 20268 14344 20304 14384
rect 19756 13292 19796 13301
rect 19756 12788 19796 13252
rect 19756 12739 19796 12748
rect 19864 12872 20304 14344
rect 19864 12832 19900 12872
rect 20268 12832 20304 12872
rect 18624 12076 18660 12116
rect 19028 12076 19064 12116
rect 18624 10604 19064 12076
rect 18624 10564 18660 10604
rect 19028 10564 19064 10604
rect 18624 9092 19064 10564
rect 18624 9052 18660 9092
rect 19028 9052 19064 9092
rect 18624 7580 19064 9052
rect 18624 7540 18660 7580
rect 19028 7540 19064 7580
rect 18624 6068 19064 7540
rect 18624 6028 18660 6068
rect 19028 6028 19064 6068
rect 12090 3760 12126 3800
rect 12494 3760 12530 3800
rect 12090 2288 12530 3760
rect 12090 2248 12126 2288
rect 12494 2248 12530 2288
rect 12090 776 12530 2248
rect 12090 736 12126 776
rect 12494 736 12530 776
rect 12090 712 12530 736
rect 18624 4556 19064 6028
rect 18624 4516 18660 4556
rect 19028 4516 19064 4556
rect 18624 3044 19064 4516
rect 18624 3004 18660 3044
rect 19028 3004 19064 3044
rect 18624 1532 19064 3004
rect 18624 1492 18660 1532
rect 19028 1492 19064 1532
rect 18624 712 19064 1492
rect 19864 11360 20304 12832
rect 19864 11320 19900 11360
rect 20268 11320 20304 11360
rect 19864 9848 20304 11320
rect 19864 9808 19900 9848
rect 20268 9808 20304 9848
rect 19864 8336 20304 9808
rect 26188 9596 26228 25180
rect 26398 24212 26838 25684
rect 27340 27572 27380 27581
rect 27148 24380 27188 24389
rect 26398 24172 26434 24212
rect 26802 24172 26838 24212
rect 26398 22700 26838 24172
rect 27052 24296 27092 24305
rect 26398 22660 26434 22700
rect 26802 22660 26838 22700
rect 26398 21188 26838 22660
rect 26398 21148 26434 21188
rect 26802 21148 26838 21188
rect 26284 19928 26324 19937
rect 26284 19340 26324 19888
rect 26284 19291 26324 19300
rect 26398 19676 26838 21148
rect 26398 19636 26434 19676
rect 26802 19636 26838 19676
rect 26284 18416 26324 18425
rect 26284 16988 26324 18376
rect 26284 16939 26324 16948
rect 26398 18164 26838 19636
rect 26398 18124 26434 18164
rect 26802 18124 26838 18164
rect 26188 9547 26228 9556
rect 26398 16652 26838 18124
rect 26398 16612 26434 16652
rect 26802 16612 26838 16652
rect 26398 15140 26838 16612
rect 26398 15100 26434 15140
rect 26802 15100 26838 15140
rect 26398 13628 26838 15100
rect 26398 13588 26434 13628
rect 26802 13588 26838 13628
rect 26398 12116 26838 13588
rect 26398 12076 26434 12116
rect 26802 12076 26838 12116
rect 26398 10604 26838 12076
rect 26956 23624 26996 23633
rect 26956 11024 26996 23584
rect 27052 20516 27092 24256
rect 27052 20467 27092 20476
rect 27148 23288 27188 24340
rect 27148 20012 27188 23248
rect 27244 23204 27284 23213
rect 27244 21104 27284 23164
rect 27244 21055 27284 21064
rect 26956 10975 26996 10984
rect 27052 16148 27092 16157
rect 26398 10564 26434 10604
rect 26802 10564 26838 10604
rect 19864 8296 19900 8336
rect 20268 8296 20304 8336
rect 19864 6824 20304 8296
rect 19864 6784 19900 6824
rect 20268 6784 20304 6824
rect 19864 5312 20304 6784
rect 19864 5272 19900 5312
rect 20268 5272 20304 5312
rect 19864 3800 20304 5272
rect 19864 3760 19900 3800
rect 20268 3760 20304 3800
rect 19864 2288 20304 3760
rect 19864 2248 19900 2288
rect 20268 2248 20304 2288
rect 19864 776 20304 2248
rect 19864 736 19900 776
rect 20268 736 20304 776
rect 19864 712 20304 736
rect 26398 9092 26838 10564
rect 27052 10100 27092 16108
rect 27148 12284 27188 19972
rect 27340 14888 27380 27532
rect 27436 20264 27476 28036
rect 27638 27992 28078 28016
rect 27638 27952 27674 27992
rect 28042 27952 28078 27992
rect 27638 26480 28078 27952
rect 27638 26440 27674 26480
rect 28042 26440 28078 26480
rect 27436 20215 27476 20224
rect 27532 25976 27572 25985
rect 27532 20096 27572 25936
rect 27532 20047 27572 20056
rect 27638 24968 28078 26440
rect 28492 27404 28532 27413
rect 27638 24928 27674 24968
rect 28042 24928 28078 24968
rect 27638 23456 28078 24928
rect 27638 23416 27674 23456
rect 28042 23416 28078 23456
rect 27638 21944 28078 23416
rect 27638 21904 27674 21944
rect 28042 21904 28078 21944
rect 27638 20432 28078 21904
rect 27638 20392 27674 20432
rect 28042 20392 28078 20432
rect 27532 19088 27572 19097
rect 27532 17072 27572 19048
rect 27532 15728 27572 17032
rect 27532 15679 27572 15688
rect 27638 18920 28078 20392
rect 27638 18880 27674 18920
rect 28042 18880 28078 18920
rect 27638 17408 28078 18880
rect 27638 17368 27674 17408
rect 28042 17368 28078 17408
rect 27638 15896 28078 17368
rect 27638 15856 27674 15896
rect 28042 15856 28078 15896
rect 27340 14839 27380 14848
rect 27148 12235 27188 12244
rect 27638 14384 28078 15856
rect 27638 14344 27674 14384
rect 28042 14344 28078 14384
rect 27638 12872 28078 14344
rect 27638 12832 27674 12872
rect 28042 12832 28078 12872
rect 27052 10051 27092 10060
rect 27638 11360 28078 12832
rect 27638 11320 27674 11360
rect 28042 11320 28078 11360
rect 26398 9052 26434 9092
rect 26802 9052 26838 9092
rect 26398 7580 26838 9052
rect 26398 7540 26434 7580
rect 26802 7540 26838 7580
rect 26398 6068 26838 7540
rect 26398 6028 26434 6068
rect 26802 6028 26838 6068
rect 26398 4556 26838 6028
rect 26398 4516 26434 4556
rect 26802 4516 26838 4556
rect 26398 3044 26838 4516
rect 26398 3004 26434 3044
rect 26802 3004 26838 3044
rect 26398 1532 26838 3004
rect 26398 1492 26434 1532
rect 26802 1492 26838 1532
rect 26398 712 26838 1492
rect 27638 9848 28078 11320
rect 28204 26312 28244 26321
rect 28204 10940 28244 26272
rect 28492 17744 28532 27364
rect 31084 27404 31124 27413
rect 30124 26900 30164 26909
rect 29164 26060 29204 26069
rect 28684 21608 28724 21617
rect 28684 18752 28724 21568
rect 28684 18703 28724 18712
rect 28492 17695 28532 17704
rect 28876 18668 28916 18677
rect 28876 15644 28916 18628
rect 28876 13964 28916 15604
rect 28876 13208 28916 13924
rect 28876 13159 28916 13168
rect 28204 10891 28244 10900
rect 29164 10604 29204 26020
rect 30028 25976 30068 25985
rect 29548 25136 29588 25145
rect 29452 24548 29492 24557
rect 29260 23792 29300 23801
rect 29260 11864 29300 23752
rect 29260 11815 29300 11824
rect 29452 11192 29492 24508
rect 29452 11143 29492 11152
rect 29548 11108 29588 25096
rect 29548 11059 29588 11068
rect 29644 24548 29684 24557
rect 29164 10555 29204 10564
rect 29644 10352 29684 24508
rect 30028 11192 30068 25936
rect 30124 12368 30164 26860
rect 30796 23876 30836 23885
rect 30316 23372 30356 23381
rect 30316 14972 30356 23332
rect 30604 23120 30644 23129
rect 30316 14923 30356 14932
rect 30412 22364 30452 22373
rect 30124 12319 30164 12328
rect 30028 11143 30068 11152
rect 30412 10856 30452 22324
rect 30604 11948 30644 23080
rect 30604 11899 30644 11908
rect 30412 10807 30452 10816
rect 30796 10856 30836 23836
rect 31084 13964 31124 27364
rect 31084 13915 31124 13924
rect 30796 10807 30836 10816
rect 29644 10303 29684 10312
rect 27638 9808 27674 9848
rect 28042 9808 28078 9848
rect 27638 8336 28078 9808
rect 27638 8296 27674 8336
rect 28042 8296 28078 8336
rect 27638 6824 28078 8296
rect 27638 6784 27674 6824
rect 28042 6784 28078 6824
rect 27638 5312 28078 6784
rect 27638 5272 27674 5312
rect 28042 5272 28078 5312
rect 27638 3800 28078 5272
rect 27638 3760 27674 3800
rect 28042 3760 28078 3800
rect 27638 2288 28078 3760
rect 27638 2248 27674 2288
rect 28042 2248 28078 2288
rect 27638 776 28078 2248
rect 27638 736 27674 776
rect 28042 736 28078 776
rect 27638 712 28078 736
use sg13g2_inv_1  _1039_
timestamp 1746816402
transform -1 0 25728 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1040_
timestamp 1746816402
transform -1 0 27072 0 -1 24948
box -48 -56 336 834
use sg13g2_inv_1  _1041_
timestamp 1746816402
transform 1 0 25728 0 1 8316
box -48 -56 336 834
use sg13g2_inv_1  _1042_
timestamp 1746816402
transform 1 0 21216 0 -1 5292
box -48 -56 336 834
use sg13g2_inv_1  _1043_
timestamp 1746816402
transform 1 0 12096 0 -1 11340
box -48 -56 336 834
use sg13g2_inv_1  _1044_
timestamp 1746816402
transform -1 0 4512 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1045_
timestamp 1746816402
transform 1 0 9408 0 1 23436
box -48 -56 336 834
use sg13g2_inv_2  _1046_
timestamp 1746816402
transform 1 0 30144 0 -1 17388
box -48 -56 432 834
use sg13g2_inv_2  _1047_
timestamp 1746816402
transform -1 0 21888 0 1 11340
box -48 -56 432 834
use sg13g2_inv_1  _1048_
timestamp 1746816402
transform -1 0 25824 0 -1 21924
box -48 -56 336 834
use sg13g2_inv_2  _1049_
timestamp 1746816402
transform 1 0 21504 0 1 9828
box -48 -56 432 834
use sg13g2_inv_2  _1050_
timestamp 1746816402
transform 1 0 7680 0 -1 20412
box -48 -56 432 834
use sg13g2_inv_1  _1051_
timestamp 1746816402
transform -1 0 13344 0 1 20412
box -48 -56 336 834
use sg13g2_inv_1  _1052_
timestamp 1746816402
transform -1 0 23520 0 -1 24948
box -48 -56 336 834
use sg13g2_inv_1  _1053_
timestamp 1746816402
transform -1 0 19776 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1054_
timestamp 1746816402
transform -1 0 18240 0 -1 27972
box -48 -56 336 834
use sg13g2_inv_1  _1055_
timestamp 1746816402
transform -1 0 16608 0 -1 26460
box -48 -56 336 834
use sg13g2_inv_1  _1056_
timestamp 1746816402
transform -1 0 8736 0 1 3780
box -48 -56 336 834
use sg13g2_inv_2  _1057_
timestamp 1746816402
transform -1 0 13920 0 1 3780
box -48 -56 432 834
use sg13g2_o21ai_1  _1058_
timestamp 1746816402
transform -1 0 25536 0 -1 17388
box -48 -56 538 834
use sg13g2_nand3b_1  _1059_
timestamp 1746816402
transform -1 0 25824 0 -1 15876
box -48 -56 720 834
use sg13g2_nor3_1  _1060_
timestamp 1746816402
transform 1 0 24672 0 1 15876
box -48 -56 528 834
use sg13g2_nor2b_1  _1061_
timestamp 1746816402
transform -1 0 26304 0 1 14364
box -54 -56 528 834
use sg13g2_o21ai_1  _1062_
timestamp 1746816402
transform -1 0 25824 0 1 14364
box -48 -56 538 834
use sg13g2_nor2_1  _1063_
timestamp 1746816402
transform 1 0 25152 0 1 15876
box -48 -56 432 834
use sg13g2_nor2_2  _1064_
timestamp 1746816402
transform 1 0 21792 0 1 17388
box -48 -56 624 834
use sg13g2_nor2b_1  _1065_
timestamp 1746816402
transform -1 0 22944 0 -1 17388
box -54 -56 528 834
use sg13g2_nand2_1  _1066_
timestamp 1746816402
transform 1 0 23520 0 -1 17388
box -48 -56 432 834
use sg13g2_nand2_1  _1067_
timestamp 1746816402
transform -1 0 24288 0 1 17388
box -48 -56 432 834
use sg13g2_nor4_1  _1068_
timestamp 1746816402
transform 1 0 22944 0 -1 17388
box -48 -56 624 834
use sg13g2_nor3_1  _1069_
timestamp 1746816402
transform -1 0 25056 0 -1 17388
box -48 -56 528 834
use sg13g2_a21oi_2  _1070_
timestamp 1746816402
transform 1 0 24192 0 -1 20412
box -48 -56 816 834
use sg13g2_inv_1  _1071_
timestamp 1746816402
transform 1 0 12672 0 -1 23436
box -48 -56 336 834
use sg13g2_and2_2  _1072_
timestamp 1746816402
transform 1 0 25440 0 1 20412
box -48 -56 624 834
use sg13g2_nor2_1  _1073_
timestamp 1746816402
transform -1 0 29952 0 -1 12852
box -48 -56 432 834
use sg13g2_nor3_1  _1074_
timestamp 1746816402
transform 1 0 24576 0 1 21924
box -48 -56 528 834
use sg13g2_nand2_1  _1075_
timestamp 1746816402
transform -1 0 30912 0 1 14364
box -48 -56 432 834
use sg13g2_nand3_1  _1076_
timestamp 1746816402
transform -1 0 25440 0 1 23436
box -48 -56 528 834
use sg13g2_nand2_1  _1077_
timestamp 1746816402
transform -1 0 30528 0 1 11340
box -48 -56 432 834
use sg13g2_nand2b_1  _1078_
timestamp 1746816402
transform 1 0 28128 0 -1 23436
box -48 -56 528 834
use sg13g2_nor3_2  _1079_
timestamp 1746816402
transform 1 0 26304 0 -1 23436
box -48 -56 912 834
use sg13g2_or2_1  _1080_
timestamp 1746816402
transform 1 0 25536 0 1 24948
box -48 -56 528 834
use sg13g2_nor3_1  _1081_
timestamp 1746816402
transform -1 0 26304 0 -1 24948
box -48 -56 528 834
use sg13g2_nor2b_1  _1082_
timestamp 1746816402
transform 1 0 26784 0 1 21924
box -54 -56 528 834
use sg13g2_a221oi_1  _1083_
timestamp 1746816402
transform 1 0 25440 0 -1 23436
box -48 -56 816 834
use sg13g2_a21oi_2  _1084_
timestamp 1746816402
transform 1 0 24576 0 -1 23436
box -48 -56 816 834
use sg13g2_and2_1  _1085_
timestamp 1746816402
transform 1 0 18144 0 -1 23436
box -48 -56 528 834
use sg13g2_nand2_1  _1086_
timestamp 1746816402
transform -1 0 19488 0 -1 23436
box -48 -56 432 834
use sg13g2_nor2_1  _1087_
timestamp 1746816402
transform -1 0 13728 0 -1 23436
box -48 -56 432 834
use sg13g2_a21oi_1  _1088_
timestamp 1746816402
transform -1 0 7392 0 1 23436
box -48 -56 528 834
use sg13g2_nand2_1  _1089_
timestamp 1746816402
transform 1 0 1728 0 1 24948
box -48 -56 432 834
use sg13g2_nor2_1  _1090_
timestamp 1746816402
transform 1 0 8256 0 -1 23436
box -48 -56 432 834
use sg13g2_a21oi_1  _1091_
timestamp 1746816402
transform 1 0 8640 0 -1 24948
box -48 -56 528 834
use sg13g2_o21ai_1  _1092_
timestamp 1746816402
transform 1 0 8928 0 1 23436
box -48 -56 538 834
use sg13g2_nor2_1  _1093_
timestamp 1746816402
transform 1 0 2016 0 -1 26460
box -48 -56 432 834
use sg13g2_a21oi_1  _1094_
timestamp 1746816402
transform 1 0 5280 0 1 26460
box -48 -56 528 834
use sg13g2_nor2_1  _1095_
timestamp 1746816402
transform 1 0 2880 0 -1 27972
box -48 -56 432 834
use sg13g2_or2_1  _1096_
timestamp 1746816402
transform 1 0 7488 0 1 24948
box -48 -56 528 834
use sg13g2_inv_1  _1097_
timestamp 1746816402
transform 1 0 10560 0 1 24948
box -48 -56 336 834
use sg13g2_nor2_1  _1098_
timestamp 1746816402
transform 1 0 2112 0 -1 27972
box -48 -56 432 834
use sg13g2_nor2_1  _1099_
timestamp 1746816402
transform -1 0 2400 0 1 26460
box -48 -56 432 834
use sg13g2_a21oi_1  _1100_
timestamp 1746816402
transform 1 0 7872 0 1 26460
box -48 -56 528 834
use sg13g2_nor2_1  _1101_
timestamp 1746816402
transform 1 0 1728 0 -1 27972
box -48 -56 432 834
use sg13g2_xnor2_1  _1102_
timestamp 1746816402
transform -1 0 26208 0 -1 26460
box -48 -56 816 834
use sg13g2_nor2_2  _1103_
timestamp 1746816402
transform 1 0 12480 0 1 20412
box -48 -56 624 834
use sg13g2_and2_1  _1104_
timestamp 1746816402
transform -1 0 13728 0 -1 21924
box -48 -56 528 834
use sg13g2_nand2_1  _1105_
timestamp 1746816402
transform 1 0 15264 0 -1 20412
box -48 -56 432 834
use sg13g2_nor2_2  _1106_
timestamp 1746816402
transform 1 0 13536 0 -1 20412
box -48 -56 624 834
use sg13g2_nand2_1  _1107_
timestamp 1746816402
transform 1 0 12288 0 -1 23436
box -48 -56 432 834
use sg13g2_nand2_1  _1108_
timestamp 1746816402
transform 1 0 9696 0 1 23436
box -48 -56 432 834
use sg13g2_nand3b_1  _1109_
timestamp 1746816402
transform -1 0 24576 0 -1 17388
box -48 -56 720 834
use sg13g2_nor2_1  _1110_
timestamp 1746816402
transform 1 0 19200 0 1 18900
box -48 -56 432 834
use sg13g2_or2_1  _1111_
timestamp 1746816402
transform -1 0 20448 0 -1 20412
box -48 -56 528 834
use sg13g2_xnor2_1  _1112_
timestamp 1746816402
transform 1 0 23904 0 1 20412
box -48 -56 816 834
use sg13g2_nand2_1  _1113_
timestamp 1746816402
transform 1 0 15168 0 -1 23436
box -48 -56 432 834
use sg13g2_xnor2_1  _1114_
timestamp 1746816402
transform 1 0 23424 0 1 21924
box -48 -56 816 834
use sg13g2_inv_1  _1115_
timestamp 1746816402
transform 1 0 24576 0 -1 24948
box -48 -56 336 834
use sg13g2_nor2_1  _1116_
timestamp 1746816402
transform -1 0 21600 0 1 20412
box -48 -56 432 834
use sg13g2_nand2_1  _1117_
timestamp 1746816402
transform 1 0 17760 0 -1 23436
box -48 -56 432 834
use sg13g2_nand2_1  _1118_
timestamp 1746816402
transform 1 0 18432 0 -1 26460
box -48 -56 432 834
use sg13g2_xnor2_1  _1119_
timestamp 1746816402
transform -1 0 21216 0 -1 26460
box -48 -56 816 834
use sg13g2_o21ai_1  _1120_
timestamp 1746816402
transform -1 0 19584 0 -1 24948
box -48 -56 538 834
use sg13g2_and2_1  _1121_
timestamp 1746816402
transform 1 0 20448 0 -1 24948
box -48 -56 528 834
use sg13g2_xor2_1  _1122_
timestamp 1746816402
transform -1 0 20448 0 -1 24948
box -48 -56 816 834
use sg13g2_nand2_1  _1123_
timestamp 1746816402
transform 1 0 18048 0 -1 24948
box -48 -56 432 834
use sg13g2_a21oi_1  _1124_
timestamp 1746816402
transform 1 0 22272 0 -1 24948
box -48 -56 528 834
use sg13g2_a21o_1  _1125_
timestamp 1746816402
transform 1 0 21024 0 -1 23436
box -48 -56 720 834
use sg13g2_nand2_1  _1126_
timestamp 1746816402
transform 1 0 21600 0 -1 21924
box -48 -56 432 834
use sg13g2_xnor2_1  _1127_
timestamp 1746816402
transform -1 0 20832 0 1 21924
box -48 -56 816 834
use sg13g2_nand2_1  _1128_
timestamp 1746816402
transform 1 0 23040 0 1 21924
box -48 -56 432 834
use sg13g2_nor2_1  _1129_
timestamp 1746816402
transform 1 0 21984 0 -1 21924
box -48 -56 432 834
use sg13g2_xnor2_1  _1130_
timestamp 1746816402
transform -1 0 21696 0 1 21924
box -48 -56 816 834
use sg13g2_nor2_1  _1131_
timestamp 1746816402
transform -1 0 22080 0 -1 23436
box -48 -56 432 834
use sg13g2_inv_1  _1132_
timestamp 1746816402
transform 1 0 20736 0 -1 23436
box -48 -56 336 834
use sg13g2_a221oi_1  _1133_
timestamp 1746816402
transform 1 0 22272 0 1 23436
box -48 -56 816 834
use sg13g2_o21ai_1  _1134_
timestamp 1746816402
transform 1 0 22560 0 1 21924
box -48 -56 538 834
use sg13g2_nor2_1  _1135_
timestamp 1746816402
transform -1 0 24576 0 1 21924
box -48 -56 432 834
use sg13g2_o21ai_1  _1136_
timestamp 1746816402
transform 1 0 24576 0 -1 21924
box -48 -56 538 834
use sg13g2_a21oi_2  _1137_
timestamp 1746816402
transform -1 0 25440 0 1 20412
box -48 -56 816 834
use sg13g2_a21o_1  _1138_
timestamp 1746816402
transform -1 0 25632 0 -1 20412
box -48 -56 720 834
use sg13g2_and2_1  _1139_
timestamp 1746816402
transform -1 0 26208 0 1 18900
box -48 -56 528 834
use sg13g2_a21oi_1  _1140_
timestamp 1746816402
transform -1 0 26016 0 -1 18900
box -48 -56 528 834
use sg13g2_o21ai_1  _1141_
timestamp 1746816402
transform -1 0 26016 0 1 17388
box -48 -56 538 834
use sg13g2_xor2_1  _1142_
timestamp 1746816402
transform -1 0 25728 0 1 18900
box -48 -56 816 834
use sg13g2_nor2_1  _1143_
timestamp 1746816402
transform -1 0 24384 0 1 15876
box -48 -56 432 834
use sg13g2_nor3_1  _1144_
timestamp 1746816402
transform 1 0 21696 0 -1 18900
box -48 -56 528 834
use sg13g2_a21oi_1  _1145_
timestamp 1746816402
transform -1 0 22656 0 -1 18900
box -48 -56 528 834
use sg13g2_nand2_1  _1146_
timestamp 1746816402
transform -1 0 22080 0 1 18900
box -48 -56 432 834
use sg13g2_xnor2_1  _1147_
timestamp 1746816402
transform -1 0 22272 0 1 23436
box -48 -56 816 834
use sg13g2_a21oi_1  _1148_
timestamp 1746816402
transform -1 0 20736 0 -1 23436
box -48 -56 528 834
use sg13g2_xnor2_1  _1149_
timestamp 1746816402
transform -1 0 21312 0 1 23436
box -48 -56 816 834
use sg13g2_nor2b_1  _1150_
timestamp 1746816402
transform -1 0 22272 0 -1 17388
box -54 -56 528 834
use sg13g2_xor2_1  _1151_
timestamp 1746816402
transform 1 0 19680 0 -1 26460
box -48 -56 816 834
use sg13g2_nand2b_1  _1152_
timestamp 1746816402
transform 1 0 20544 0 -1 18900
box -48 -56 528 834
use sg13g2_and2_1  _1153_
timestamp 1746816402
transform 1 0 20832 0 -1 15876
box -48 -56 528 834
use sg13g2_nand2_2  _1154_
timestamp 1746816402
transform 1 0 19296 0 -1 17388
box -48 -56 624 834
use sg13g2_xor2_1  _1155_
timestamp 1746816402
transform 1 0 19776 0 1 24948
box -48 -56 816 834
use sg13g2_o21ai_1  _1156_
timestamp 1746816402
transform 1 0 19584 0 1 18900
box -48 -56 538 834
use sg13g2_nor2_1  _1157_
timestamp 1746816402
transform -1 0 21408 0 -1 18900
box -48 -56 432 834
use sg13g2_xnor2_1  _1158_
timestamp 1746816402
transform 1 0 19776 0 1 23436
box -48 -56 816 834
use sg13g2_inv_1  _1159_
timestamp 1746816402
transform -1 0 5568 0 1 8316
box -48 -56 336 834
use sg13g2_a221oi_1  _1160_
timestamp 1746816402
transform 1 0 19776 0 -1 18900
box -48 -56 816 834
use sg13g2_nor2_1  _1161_
timestamp 1746816402
transform -1 0 21600 0 1 18900
box -48 -56 432 834
use sg13g2_and3_1  _1162_
timestamp 1746816402
transform 1 0 23904 0 -1 21924
box -48 -56 720 834
use sg13g2_or2_2  _1163_
timestamp 1746816402
transform -1 0 24480 0 1 11340
box -48 -56 624 834
use sg13g2_xnor2_1  _1164_
timestamp 1746816402
transform 1 0 22464 0 -1 21924
box -48 -56 816 834
use sg13g2_nor2b_1  _1165_
timestamp 1746816402
transform 1 0 20448 0 1 17388
box -54 -56 528 834
use sg13g2_xor2_1  _1166_
timestamp 1746816402
transform -1 0 20832 0 -1 21924
box -48 -56 816 834
use sg13g2_nand2b_1  _1167_
timestamp 1746816402
transform 1 0 20160 0 -1 15876
box -48 -56 528 834
use sg13g2_o21ai_1  _1168_
timestamp 1746816402
transform -1 0 20064 0 -1 21924
box -48 -56 538 834
use sg13g2_xor2_1  _1169_
timestamp 1746816402
transform -1 0 21600 0 -1 21924
box -48 -56 816 834
use sg13g2_a221oi_1  _1170_
timestamp 1746816402
transform -1 0 20928 0 -1 17388
box -48 -56 816 834
use sg13g2_a21oi_1  _1171_
timestamp 1746816402
transform -1 0 21408 0 -1 17388
box -48 -56 528 834
use sg13g2_nor2_2  _1172_
timestamp 1746816402
transform 1 0 23424 0 1 15876
box -48 -56 624 834
use sg13g2_nor3_2  _1173_
timestamp 1746816402
transform -1 0 21216 0 1 18900
box -48 -56 912 834
use sg13g2_nand2_1  _1174_
timestamp 1746816402
transform 1 0 9216 0 -1 21924
box -48 -56 432 834
use sg13g2_a21oi_1  _1175_
timestamp 1746816402
transform -1 0 10080 0 -1 21924
box -48 -56 528 834
use sg13g2_or4_1  _1176_
timestamp 1746816402
transform 1 0 10752 0 1 21924
box -48 -56 816 834
use sg13g2_mux4_1  _1177_
timestamp 1746816402
transform 1 0 17088 0 -1 15876
box -48 -56 2064 834
use sg13g2_nor2_1  _1178_
timestamp 1746816402
transform -1 0 7488 0 1 17388
box -48 -56 432 834
use sg13g2_nor2_1  _1179_
timestamp 1746816402
transform -1 0 16320 0 1 14364
box -48 -56 432 834
use sg13g2_or2_2  _1180_
timestamp 1746816402
transform 1 0 12384 0 -1 17388
box -48 -56 624 834
use sg13g2_nor2b_1  _1181_
timestamp 1746816402
transform -1 0 14016 0 1 15876
box -54 -56 528 834
use sg13g2_a221oi_1  _1182_
timestamp 1746816402
transform -1 0 6432 0 1 17388
box -48 -56 816 834
use sg13g2_nor2b_2  _1183_
timestamp 1746816402
transform -1 0 12864 0 -1 20412
box -54 -56 720 834
use sg13g2_and2_1  _1184_
timestamp 1746816402
transform 1 0 12096 0 -1 18900
box -48 -56 528 834
use sg13g2_nand2_2  _1185_
timestamp 1746816402
transform -1 0 13152 0 1 18900
box -48 -56 624 834
use sg13g2_nor2_1  _1186_
timestamp 1746816402
transform 1 0 25152 0 -1 18900
box -48 -56 432 834
use sg13g2_mux2_1  _1187_
timestamp 1746816402
transform -1 0 19392 0 -1 18900
box -48 -56 1008 834
use sg13g2_and2_1  _1188_
timestamp 1746816402
transform 1 0 14112 0 -1 20412
box -48 -56 528 834
use sg13g2_nor2b_2  _1189_
timestamp 1746816402
transform 1 0 12864 0 -1 20412
box -54 -56 720 834
use sg13g2_and2_1  _1190_
timestamp 1746816402
transform 1 0 16128 0 1 18900
box -48 -56 528 834
use sg13g2_nand2_1  _1191_
timestamp 1746816402
transform -1 0 12192 0 1 17388
box -48 -56 432 834
use sg13g2_nor2_1  _1192_
timestamp 1746816402
transform -1 0 11808 0 1 17388
box -48 -56 432 834
use sg13g2_nand2b_2  _1193_
timestamp 1746816402
transform -1 0 11136 0 -1 17388
box -48 -56 816 834
use sg13g2_nor2_1  _1194_
timestamp 1746816402
transform -1 0 19776 0 -1 18900
box -48 -56 432 834
use sg13g2_nand2b_1  _1195_
timestamp 1746816402
transform -1 0 14208 0 -1 18900
box -48 -56 528 834
use sg13g2_xnor2_1  _1196_
timestamp 1746816402
transform 1 0 4608 0 -1 18900
box -48 -56 816 834
use sg13g2_nor2_2  _1197_
timestamp 1746816402
transform -1 0 5664 0 1 17388
box -48 -56 624 834
use sg13g2_nand2_1  _1198_
timestamp 1746816402
transform 1 0 4992 0 1 18900
box -48 -56 432 834
use sg13g2_and2_1  _1199_
timestamp 1746816402
transform 1 0 16512 0 -1 20412
box -48 -56 528 834
use sg13g2_nand2_1  _1200_
timestamp 1746816402
transform 1 0 16992 0 -1 21924
box -48 -56 432 834
use sg13g2_nor2_1  _1201_
timestamp 1746816402
transform 1 0 5664 0 -1 18900
box -48 -56 432 834
use sg13g2_a221oi_1  _1202_
timestamp 1746816402
transform -1 0 6816 0 -1 18900
box -48 -56 816 834
use sg13g2_o21ai_1  _1203_
timestamp 1746816402
transform 1 0 6336 0 1 18900
box -48 -56 538 834
use sg13g2_a21oi_1  _1204_
timestamp 1746816402
transform -1 0 11040 0 -1 21924
box -48 -56 528 834
use sg13g2_o21ai_1  _1205_
timestamp 1746816402
transform 1 0 11136 0 -1 23436
box -48 -56 538 834
use sg13g2_o21ai_1  _1206_
timestamp 1746816402
transform -1 0 12192 0 -1 23436
box -48 -56 538 834
use sg13g2_o21ai_1  _1207_
timestamp 1746816402
transform 1 0 7680 0 1 21924
box -48 -56 538 834
use sg13g2_nor2_1  _1208_
timestamp 1746816402
transform -1 0 10272 0 1 21924
box -48 -56 432 834
use sg13g2_nand2b_1  _1209_
timestamp 1746816402
transform -1 0 8544 0 -1 21924
box -48 -56 528 834
use sg13g2_nand2_1  _1210_
timestamp 1746816402
transform -1 0 8064 0 -1 21924
box -48 -56 432 834
use sg13g2_nand2_1  _1211_
timestamp 1746816402
transform -1 0 2400 0 1 14364
box -48 -56 432 834
use sg13g2_nor2_1  _1212_
timestamp 1746816402
transform 1 0 960 0 -1 14364
box -48 -56 432 834
use sg13g2_xor2_1  _1213_
timestamp 1746816402
transform 1 0 1248 0 1 14364
box -48 -56 816 834
use sg13g2_xnor2_1  _1214_
timestamp 1746816402
transform 1 0 1344 0 -1 15876
box -48 -56 816 834
use sg13g2_nand2_1  _1215_
timestamp 1746816402
transform -1 0 1728 0 1 15876
box -48 -56 432 834
use sg13g2_and2_1  _1216_
timestamp 1746816402
transform 1 0 2112 0 -1 17388
box -48 -56 528 834
use sg13g2_xor2_1  _1217_
timestamp 1746816402
transform 1 0 1728 0 1 15876
box -48 -56 816 834
use sg13g2_xnor2_1  _1218_
timestamp 1746816402
transform 1 0 2496 0 1 15876
box -48 -56 816 834
use sg13g2_xnor2_1  _1219_
timestamp 1746816402
transform 1 0 2784 0 1 12852
box -48 -56 816 834
use sg13g2_xnor2_1  _1220_
timestamp 1746816402
transform 1 0 6816 0 -1 14364
box -48 -56 816 834
use sg13g2_and2_2  _1221_
timestamp 1746816402
transform 1 0 17664 0 1 17388
box -48 -56 624 834
use sg13g2_nand2_1  _1222_
timestamp 1746816402
transform 1 0 12576 0 1 17388
box -48 -56 432 834
use sg13g2_a21oi_1  _1223_
timestamp 1746816402
transform -1 0 8064 0 1 12852
box -48 -56 528 834
use sg13g2_o21ai_1  _1224_
timestamp 1746816402
transform 1 0 8736 0 1 12852
box -48 -56 538 834
use sg13g2_nor2b_2  _1225_
timestamp 1746816402
transform 1 0 13344 0 1 12852
box -54 -56 720 834
use sg13g2_nand2b_2  _1226_
timestamp 1746816402
transform -1 0 13344 0 1 12852
box -48 -56 816 834
use sg13g2_a21o_1  _1227_
timestamp 1746816402
transform 1 0 8064 0 1 12852
box -48 -56 720 834
use sg13g2_nor2b_1  _1228_
timestamp 1746816402
transform 1 0 6432 0 -1 17388
box -54 -56 528 834
use sg13g2_mux2_1  _1229_
timestamp 1746816402
transform 1 0 19008 0 1 12852
box -48 -56 1008 834
use sg13g2_mux2_1  _1230_
timestamp 1746816402
transform 1 0 18816 0 1 14364
box -48 -56 1008 834
use sg13g2_mux2_2  _1231_
timestamp 1746816402
transform -1 0 20160 0 -1 15876
box -48 -56 1104 834
use sg13g2_a221oi_1  _1232_
timestamp 1746816402
transform 1 0 7008 0 -1 17388
box -48 -56 816 834
use sg13g2_inv_1  _1233_
timestamp 1746816402
transform 1 0 6240 0 -1 15876
box -48 -56 336 834
use sg13g2_a22oi_1  _1234_
timestamp 1746816402
transform 1 0 7584 0 -1 15876
box -48 -56 624 834
use sg13g2_o21ai_1  _1235_
timestamp 1746816402
transform 1 0 7008 0 -1 15876
box -48 -56 538 834
use sg13g2_a221oi_1  _1236_
timestamp 1746816402
transform -1 0 7872 0 1 15876
box -48 -56 816 834
use sg13g2_o21ai_1  _1237_
timestamp 1746816402
transform -1 0 9024 0 1 20412
box -48 -56 538 834
use sg13g2_nand2_1  _1238_
timestamp 1746816402
transform 1 0 7200 0 1 20412
box -48 -56 432 834
use sg13g2_a21oi_1  _1239_
timestamp 1746816402
transform 1 0 8448 0 1 23436
box -48 -56 528 834
use sg13g2_o21ai_1  _1240_
timestamp 1746816402
transform -1 0 4512 0 1 20412
box -48 -56 538 834
use sg13g2_nor2_1  _1241_
timestamp 1746816402
transform 1 0 1152 0 -1 23436
box -48 -56 432 834
use sg13g2_nand2b_1  _1242_
timestamp 1746816402
transform -1 0 3648 0 -1 20412
box -48 -56 528 834
use sg13g2_nand2_1  _1243_
timestamp 1746816402
transform -1 0 1824 0 1 20412
box -48 -56 432 834
use sg13g2_mux4_1  _1244_
timestamp 1746816402
transform -1 0 18720 0 1 12852
box -48 -56 2064 834
use sg13g2_and2_1  _1245_
timestamp 1746816402
transform 1 0 4416 0 1 14364
box -48 -56 528 834
use sg13g2_a221oi_1  _1246_
timestamp 1746816402
transform 1 0 4896 0 -1 14364
box -48 -56 816 834
use sg13g2_and2_1  _1247_
timestamp 1746816402
transform -1 0 4704 0 1 15876
box -48 -56 528 834
use sg13g2_a21o_1  _1248_
timestamp 1746816402
transform -1 0 2976 0 -1 15876
box -48 -56 720 834
use sg13g2_and2_1  _1249_
timestamp 1746816402
transform 1 0 2976 0 1 11340
box -48 -56 528 834
use sg13g2_xor2_1  _1250_
timestamp 1746816402
transform 1 0 3456 0 1 11340
box -48 -56 816 834
use sg13g2_xnor2_1  _1251_
timestamp 1746816402
transform -1 0 4704 0 -1 14364
box -48 -56 816 834
use sg13g2_o21ai_1  _1252_
timestamp 1746816402
transform 1 0 1920 0 1 12852
box -48 -56 538 834
use sg13g2_nor2b_1  _1253_
timestamp 1746816402
transform 1 0 1824 0 -1 14364
box -54 -56 528 834
use sg13g2_xnor2_1  _1254_
timestamp 1746816402
transform 1 0 2304 0 -1 14364
box -48 -56 816 834
use sg13g2_xor2_1  _1255_
timestamp 1746816402
transform 1 0 3072 0 -1 14364
box -48 -56 816 834
use sg13g2_xor2_1  _1256_
timestamp 1746816402
transform 1 0 7008 0 -1 12852
box -48 -56 816 834
use sg13g2_a21oi_2  _1257_
timestamp 1746816402
transform -1 0 8640 0 -1 12852
box -48 -56 816 834
use sg13g2_nand2_1  _1258_
timestamp 1746816402
transform 1 0 768 0 -1 11340
box -48 -56 432 834
use sg13g2_nand2_1  _1259_
timestamp 1746816402
transform -1 0 1248 0 -1 9828
box -48 -56 432 834
use sg13g2_nor2_1  _1260_
timestamp 1746816402
transform 1 0 864 0 1 11340
box -48 -56 432 834
use sg13g2_xor2_1  _1261_
timestamp 1746816402
transform 1 0 960 0 1 9828
box -48 -56 816 834
use sg13g2_xnor2_1  _1262_
timestamp 1746816402
transform 1 0 1152 0 -1 11340
box -48 -56 816 834
use sg13g2_nand2_1  _1263_
timestamp 1746816402
transform 1 0 1248 0 1 11340
box -48 -56 432 834
use sg13g2_xnor2_1  _1264_
timestamp 1746816402
transform 1 0 576 0 -1 12852
box -48 -56 816 834
use sg13g2_nand2_1  _1265_
timestamp 1746816402
transform -1 0 2496 0 1 11340
box -48 -56 432 834
use sg13g2_xnor2_1  _1266_
timestamp 1746816402
transform 1 0 1344 0 -1 12852
box -48 -56 816 834
use sg13g2_o21ai_1  _1267_
timestamp 1746816402
transform 1 0 2592 0 -1 12852
box -48 -56 538 834
use sg13g2_a21oi_1  _1268_
timestamp 1746816402
transform -1 0 2592 0 -1 12852
box -48 -56 528 834
use sg13g2_o21ai_1  _1269_
timestamp 1746816402
transform 1 0 3936 0 -1 12852
box -48 -56 538 834
use sg13g2_a21oi_1  _1270_
timestamp 1746816402
transform 1 0 5664 0 -1 14364
box -48 -56 528 834
use sg13g2_o21ai_1  _1271_
timestamp 1746816402
transform -1 0 4224 0 1 15876
box -48 -56 538 834
use sg13g2_o21ai_1  _1272_
timestamp 1746816402
transform 1 0 3072 0 -1 15876
box -48 -56 538 834
use sg13g2_a21oi_1  _1273_
timestamp 1746816402
transform -1 0 3840 0 1 18900
box -48 -56 528 834
use sg13g2_o21ai_1  _1274_
timestamp 1746816402
transform 1 0 2112 0 -1 20412
box -48 -56 538 834
use sg13g2_a21oi_1  _1275_
timestamp 1746816402
transform 1 0 2112 0 1 18900
box -48 -56 528 834
use sg13g2_o21ai_1  _1276_
timestamp 1746816402
transform -1 0 4512 0 1 21924
box -48 -56 538 834
use sg13g2_nor2_1  _1277_
timestamp 1746816402
transform -1 0 2208 0 1 20412
box -48 -56 432 834
use sg13g2_nand2b_1  _1278_
timestamp 1746816402
transform -1 0 3552 0 1 21924
box -48 -56 528 834
use sg13g2_nand2_1  _1279_
timestamp 1746816402
transform 1 0 1056 0 -1 21924
box -48 -56 432 834
use sg13g2_mux2_1  _1280_
timestamp 1746816402
transform 1 0 19776 0 1 14364
box -48 -56 1008 834
use sg13g2_mux2_2  _1281_
timestamp 1746816402
transform -1 0 20448 0 -1 14364
box -48 -56 1104 834
use sg13g2_and2_1  _1282_
timestamp 1746816402
transform 1 0 4416 0 -1 17388
box -48 -56 528 834
use sg13g2_a221oi_1  _1283_
timestamp 1746816402
transform 1 0 4896 0 -1 17388
box -48 -56 816 834
use sg13g2_and2_1  _1284_
timestamp 1746816402
transform -1 0 3456 0 -1 17388
box -48 -56 528 834
use sg13g2_a21oi_1  _1285_
timestamp 1746816402
transform 1 0 2976 0 1 14364
box -48 -56 528 834
use sg13g2_and2_1  _1286_
timestamp 1746816402
transform 1 0 6240 0 -1 8316
box -48 -56 528 834
use sg13g2_xor2_1  _1287_
timestamp 1746816402
transform 1 0 5568 0 1 8316
box -48 -56 816 834
use sg13g2_xor2_1  _1288_
timestamp 1746816402
transform -1 0 7104 0 1 8316
box -48 -56 816 834
use sg13g2_a21o_1  _1289_
timestamp 1746816402
transform -1 0 4896 0 1 11340
box -48 -56 720 834
use sg13g2_nand2_1  _1290_
timestamp 1746816402
transform 1 0 4896 0 1 11340
box -48 -56 432 834
use sg13g2_nor2_1  _1291_
timestamp 1746816402
transform -1 0 5568 0 -1 12852
box -48 -56 432 834
use sg13g2_xor2_1  _1292_
timestamp 1746816402
transform -1 0 5184 0 -1 12852
box -48 -56 816 834
use sg13g2_xnor2_1  _1293_
timestamp 1746816402
transform 1 0 3936 0 1 12852
box -48 -56 816 834
use sg13g2_xnor2_1  _1294_
timestamp 1746816402
transform -1 0 20064 0 -1 12852
box -48 -56 816 834
use sg13g2_o21ai_1  _1295_
timestamp 1746816402
transform -1 0 11712 0 1 12852
box -48 -56 538 834
use sg13g2_o21ai_1  _1296_
timestamp 1746816402
transform 1 0 1632 0 1 11340
box -48 -56 538 834
use sg13g2_xnor2_1  _1297_
timestamp 1746816402
transform -1 0 5280 0 1 8316
box -48 -56 816 834
use sg13g2_xor2_1  _1298_
timestamp 1746816402
transform 1 0 3744 0 1 8316
box -48 -56 816 834
use sg13g2_and2_1  _1299_
timestamp 1746816402
transform 1 0 2400 0 1 6804
box -48 -56 528 834
use sg13g2_xor2_1  _1300_
timestamp 1746816402
transform 1 0 3360 0 1 6804
box -48 -56 816 834
use sg13g2_o21ai_1  _1301_
timestamp 1746816402
transform 1 0 2496 0 1 9828
box -48 -56 538 834
use sg13g2_xnor2_1  _1302_
timestamp 1746816402
transform -1 0 4512 0 -1 8316
box -48 -56 816 834
use sg13g2_a21oi_1  _1303_
timestamp 1746816402
transform 1 0 3264 0 1 8316
box -48 -56 528 834
use sg13g2_o21ai_1  _1304_
timestamp 1746816402
transform 1 0 4416 0 -1 9828
box -48 -56 538 834
use sg13g2_a221oi_1  _1305_
timestamp 1746816402
transform -1 0 5472 0 1 12852
box -48 -56 816 834
use sg13g2_o21ai_1  _1306_
timestamp 1746816402
transform 1 0 3456 0 -1 17388
box -48 -56 538 834
use sg13g2_o21ai_1  _1307_
timestamp 1746816402
transform -1 0 5088 0 1 17388
box -48 -56 538 834
use sg13g2_a21oi_1  _1308_
timestamp 1746816402
transform 1 0 2784 0 -1 21924
box -48 -56 528 834
use sg13g2_o21ai_1  _1309_
timestamp 1746816402
transform -1 0 1920 0 -1 21924
box -48 -56 538 834
use sg13g2_a21oi_1  _1310_
timestamp 1746816402
transform -1 0 2016 0 -1 23436
box -48 -56 528 834
use sg13g2_o21ai_1  _1311_
timestamp 1746816402
transform -1 0 5472 0 -1 23436
box -48 -56 538 834
use sg13g2_nor2_1  _1312_
timestamp 1746816402
transform 1 0 4704 0 1 20412
box -48 -56 432 834
use sg13g2_nand2b_1  _1313_
timestamp 1746816402
transform -1 0 5760 0 -1 21924
box -48 -56 528 834
use sg13g2_nand2_1  _1314_
timestamp 1746816402
transform -1 0 5088 0 1 21924
box -48 -56 432 834
use sg13g2_nor2b_1  _1315_
timestamp 1746816402
transform 1 0 9792 0 1 14364
box -54 -56 528 834
use sg13g2_mux4_1  _1316_
timestamp 1746816402
transform -1 0 18528 0 -1 14364
box -48 -56 2064 834
use sg13g2_a221oi_1  _1317_
timestamp 1746816402
transform 1 0 10272 0 1 14364
box -48 -56 816 834
use sg13g2_and2_1  _1318_
timestamp 1746816402
transform -1 0 10176 0 -1 14364
box -48 -56 528 834
use sg13g2_o21ai_1  _1319_
timestamp 1746816402
transform 1 0 4800 0 -1 11340
box -48 -56 538 834
use sg13g2_xor2_1  _1320_
timestamp 1746816402
transform -1 0 12768 0 1 9828
box -48 -56 816 834
use sg13g2_nand2b_1  _1321_
timestamp 1746816402
transform 1 0 11904 0 -1 9828
box -48 -56 528 834
use sg13g2_xnor2_1  _1322_
timestamp 1746816402
transform -1 0 12000 0 1 9828
box -48 -56 816 834
use sg13g2_a21o_1  _1323_
timestamp 1746816402
transform -1 0 7776 0 1 8316
box -48 -56 720 834
use sg13g2_and2_1  _1324_
timestamp 1746816402
transform 1 0 9408 0 -1 11340
box -48 -56 528 834
use sg13g2_or2_1  _1325_
timestamp 1746816402
transform 1 0 9792 0 1 9828
box -48 -56 528 834
use sg13g2_nand2b_1  _1326_
timestamp 1746816402
transform 1 0 10368 0 -1 11340
box -48 -56 528 834
use sg13g2_xnor2_1  _1327_
timestamp 1746816402
transform 1 0 9600 0 1 11340
box -48 -56 816 834
use sg13g2_xor2_1  _1328_
timestamp 1746816402
transform 1 0 10944 0 1 11340
box -48 -56 816 834
use sg13g2_o21ai_1  _1329_
timestamp 1746816402
transform -1 0 11712 0 -1 11340
box -48 -56 538 834
use sg13g2_a22oi_1  _1330_
timestamp 1746816402
transform 1 0 4800 0 -1 8316
box -48 -56 624 834
use sg13g2_or2_1  _1331_
timestamp 1746816402
transform 1 0 12096 0 1 8316
box -48 -56 528 834
use sg13g2_and2_1  _1332_
timestamp 1746816402
transform 1 0 11616 0 1 8316
box -48 -56 528 834
use sg13g2_xor2_1  _1333_
timestamp 1746816402
transform -1 0 9696 0 -1 8316
box -48 -56 816 834
use sg13g2_xnor2_1  _1334_
timestamp 1746816402
transform 1 0 8928 0 1 6804
box -48 -56 816 834
use sg13g2_nand2_1  _1335_
timestamp 1746816402
transform 1 0 6528 0 1 5292
box -48 -56 432 834
use sg13g2_xnor2_1  _1336_
timestamp 1746816402
transform 1 0 7008 0 -1 6804
box -48 -56 816 834
use sg13g2_a21oi_1  _1337_
timestamp 1746816402
transform 1 0 2880 0 1 6804
box -48 -56 528 834
use sg13g2_xnor2_1  _1338_
timestamp 1746816402
transform 1 0 7488 0 1 6804
box -48 -56 816 834
use sg13g2_a21oi_1  _1339_
timestamp 1746816402
transform -1 0 10176 0 -1 8316
box -48 -56 528 834
use sg13g2_o21ai_1  _1340_
timestamp 1746816402
transform 1 0 9600 0 1 8316
box -48 -56 538 834
use sg13g2_a221oi_1  _1341_
timestamp 1746816402
transform 1 0 9504 0 -1 12852
box -48 -56 816 834
use sg13g2_o21ai_1  _1342_
timestamp 1746816402
transform -1 0 9792 0 1 14364
box -48 -56 538 834
use sg13g2_o21ai_1  _1343_
timestamp 1746816402
transform -1 0 10080 0 -1 15876
box -48 -56 538 834
use sg13g2_a21oi_1  _1344_
timestamp 1746816402
transform 1 0 5760 0 -1 21924
box -48 -56 528 834
use sg13g2_o21ai_1  _1345_
timestamp 1746816402
transform 1 0 6432 0 1 21924
box -48 -56 538 834
use sg13g2_a21oi_1  _1346_
timestamp 1746816402
transform 1 0 4512 0 -1 23436
box -48 -56 528 834
use sg13g2_o21ai_1  _1347_
timestamp 1746816402
transform -1 0 5568 0 1 20412
box -48 -56 538 834
use sg13g2_nor2_1  _1348_
timestamp 1746816402
transform -1 0 6336 0 1 20412
box -48 -56 432 834
use sg13g2_nand2b_1  _1349_
timestamp 1746816402
transform 1 0 7008 0 -1 20412
box -48 -56 528 834
use sg13g2_nand2_1  _1350_
timestamp 1746816402
transform -1 0 6720 0 1 20412
box -48 -56 432 834
use sg13g2_mux2_1  _1351_
timestamp 1746816402
transform -1 0 22368 0 1 12852
box -48 -56 1008 834
use sg13g2_mux2_2  _1352_
timestamp 1746816402
transform -1 0 21024 0 1 12852
box -48 -56 1104 834
use sg13g2_and2_1  _1353_
timestamp 1746816402
transform 1 0 13152 0 1 14364
box -48 -56 528 834
use sg13g2_a221oi_1  _1354_
timestamp 1746816402
transform 1 0 13440 0 -1 15876
box -48 -56 816 834
use sg13g2_nand2_1  _1355_
timestamp 1746816402
transform 1 0 12672 0 -1 14364
box -48 -56 432 834
use sg13g2_a21oi_1  _1356_
timestamp 1746816402
transform -1 0 10368 0 -1 11340
box -48 -56 528 834
use sg13g2_and2_1  _1357_
timestamp 1746816402
transform 1 0 13632 0 -1 9828
box -48 -56 528 834
use sg13g2_xor2_1  _1358_
timestamp 1746816402
transform 1 0 14112 0 -1 9828
box -48 -56 816 834
use sg13g2_xor2_1  _1359_
timestamp 1746816402
transform -1 0 14880 0 1 9828
box -48 -56 816 834
use sg13g2_o21ai_1  _1360_
timestamp 1746816402
transform 1 0 12384 0 -1 9828
box -48 -56 538 834
use sg13g2_nand2_1  _1361_
timestamp 1746816402
transform 1 0 13152 0 -1 9828
box -48 -56 432 834
use sg13g2_xnor2_1  _1362_
timestamp 1746816402
transform 1 0 12768 0 1 9828
box -48 -56 816 834
use sg13g2_xnor2_1  _1363_
timestamp 1746816402
transform 1 0 12672 0 -1 11340
box -48 -56 816 834
use sg13g2_xnor2_1  _1364_
timestamp 1746816402
transform -1 0 13440 0 1 11340
box -48 -56 816 834
use sg13g2_o21ai_1  _1365_
timestamp 1746816402
transform -1 0 12672 0 1 11340
box -48 -56 538 834
use sg13g2_o21ai_1  _1366_
timestamp 1746816402
transform 1 0 12672 0 -1 8316
box -48 -56 538 834
use sg13g2_xor2_1  _1367_
timestamp 1746816402
transform 1 0 12192 0 1 6804
box -48 -56 816 834
use sg13g2_xnor2_1  _1368_
timestamp 1746816402
transform 1 0 12960 0 1 6804
box -48 -56 816 834
use sg13g2_and2_1  _1369_
timestamp 1746816402
transform 1 0 12192 0 -1 5292
box -48 -56 528 834
use sg13g2_xor2_1  _1370_
timestamp 1746816402
transform 1 0 12096 0 1 5292
box -48 -56 816 834
use sg13g2_o21ai_1  _1371_
timestamp 1746816402
transform 1 0 7776 0 -1 6804
box -48 -56 538 834
use sg13g2_xor2_1  _1372_
timestamp 1746816402
transform 1 0 12768 0 -1 6804
box -48 -56 816 834
use sg13g2_a21oi_1  _1373_
timestamp 1746816402
transform -1 0 14016 0 -1 6804
box -48 -56 528 834
use sg13g2_o21ai_1  _1374_
timestamp 1746816402
transform 1 0 14016 0 -1 6804
box -48 -56 538 834
use sg13g2_a21oi_1  _1375_
timestamp 1746816402
transform 1 0 13440 0 -1 11340
box -48 -56 528 834
use sg13g2_o21ai_1  _1376_
timestamp 1746816402
transform -1 0 14112 0 -1 12852
box -48 -56 538 834
use sg13g2_a21o_1  _1377_
timestamp 1746816402
transform 1 0 12480 0 1 14364
box -48 -56 720 834
use sg13g2_o21ai_1  _1378_
timestamp 1746816402
transform -1 0 12672 0 -1 15876
box -48 -56 538 834
use sg13g2_a21oi_1  _1379_
timestamp 1746816402
transform 1 0 5856 0 1 18900
box -48 -56 528 834
use sg13g2_o21ai_1  _1380_
timestamp 1746816402
transform -1 0 5856 0 1 18900
box -48 -56 538 834
use sg13g2_a21oi_1  _1381_
timestamp 1746816402
transform 1 0 4608 0 -1 20412
box -48 -56 528 834
use sg13g2_o21ai_1  _1382_
timestamp 1746816402
transform -1 0 14592 0 -1 23436
box -48 -56 538 834
use sg13g2_nor2_1  _1383_
timestamp 1746816402
transform -1 0 16416 0 -1 20412
box -48 -56 432 834
use sg13g2_nand2b_1  _1384_
timestamp 1746816402
transform -1 0 14304 0 1 20412
box -48 -56 528 834
use sg13g2_nand2_1  _1385_
timestamp 1746816402
transform 1 0 16800 0 -1 18900
box -48 -56 432 834
use sg13g2_o21ai_1  _1386_
timestamp 1746816402
transform 1 0 13920 0 -1 11340
box -48 -56 538 834
use sg13g2_nand2_1  _1387_
timestamp 1746816402
transform -1 0 16704 0 1 6804
box -48 -56 432 834
use sg13g2_xnor2_1  _1388_
timestamp 1746816402
transform 1 0 15456 0 -1 6804
box -48 -56 816 834
use sg13g2_xnor2_1  _1389_
timestamp 1746816402
transform -1 0 16512 0 -1 9828
box -48 -56 816 834
use sg13g2_a21oi_1  _1390_
timestamp 1746816402
transform -1 0 15360 0 -1 9828
box -48 -56 528 834
use sg13g2_nor2_1  _1391_
timestamp 1746816402
transform -1 0 15744 0 -1 9828
box -48 -56 432 834
use sg13g2_xor2_1  _1392_
timestamp 1746816402
transform -1 0 15648 0 1 9828
box -48 -56 816 834
use sg13g2_nor2_1  _1393_
timestamp 1746816402
transform 1 0 14784 0 -1 11340
box -48 -56 432 834
use sg13g2_nand2_1  _1394_
timestamp 1746816402
transform -1 0 14784 0 -1 11340
box -48 -56 432 834
use sg13g2_nor2_1  _1395_
timestamp 1746816402
transform -1 0 16032 0 -1 11340
box -48 -56 432 834
use sg13g2_xnor2_1  _1396_
timestamp 1746816402
transform 1 0 14400 0 -1 12852
box -48 -56 816 834
use sg13g2_a21o_1  _1397_
timestamp 1746816402
transform 1 0 15168 0 -1 12852
box -48 -56 720 834
use sg13g2_a22oi_1  _1398_
timestamp 1746816402
transform -1 0 13824 0 -1 8316
box -48 -56 624 834
use sg13g2_nor2_1  _1399_
timestamp 1746816402
transform 1 0 16608 0 1 8316
box -48 -56 432 834
use sg13g2_xor2_1  _1400_
timestamp 1746816402
transform -1 0 16800 0 -1 8316
box -48 -56 816 834
use sg13g2_nor2b_1  _1401_
timestamp 1746816402
transform 1 0 16128 0 1 8316
box -54 -56 528 834
use sg13g2_xor2_1  _1402_
timestamp 1746816402
transform 1 0 15264 0 -1 8316
box -48 -56 816 834
use sg13g2_xnor2_1  _1403_
timestamp 1746816402
transform -1 0 16032 0 1 5292
box -48 -56 816 834
use sg13g2_a21o_1  _1404_
timestamp 1746816402
transform -1 0 13536 0 1 5292
box -48 -56 720 834
use sg13g2_nor2b_1  _1405_
timestamp 1746816402
transform 1 0 14016 0 1 5292
box -54 -56 528 834
use sg13g2_xnor2_1  _1406_
timestamp 1746816402
transform 1 0 14496 0 1 5292
box -48 -56 816 834
use sg13g2_a21oi_1  _1407_
timestamp 1746816402
transform -1 0 15456 0 1 8316
box -48 -56 528 834
use sg13g2_o21ai_1  _1408_
timestamp 1746816402
transform -1 0 15936 0 1 8316
box -48 -56 538 834
use sg13g2_a221oi_1  _1409_
timestamp 1746816402
transform -1 0 15456 0 1 11340
box -48 -56 816 834
use sg13g2_nor2b_1  _1410_
timestamp 1746816402
transform 1 0 14208 0 1 15876
box -54 -56 528 834
use sg13g2_mux4_1  _1411_
timestamp 1746816402
transform -1 0 23328 0 -1 14364
box -48 -56 2064 834
use sg13g2_a221oi_1  _1412_
timestamp 1746816402
transform 1 0 14592 0 -1 15876
box -48 -56 816 834
use sg13g2_nor2_1  _1413_
timestamp 1746816402
transform -1 0 16032 0 -1 20412
box -48 -56 432 834
use sg13g2_a21oi_1  _1414_
timestamp 1746816402
transform -1 0 14496 0 1 18900
box -48 -56 528 834
use sg13g2_or3_1  _1415_
timestamp 1746816402
transform -1 0 15168 0 1 18900
box -48 -56 720 834
use sg13g2_a21oi_1  _1416_
timestamp 1746816402
transform 1 0 14688 0 -1 20412
box -48 -56 528 834
use sg13g2_a21oi_1  _1417_
timestamp 1746816402
transform 1 0 14304 0 1 20412
box -48 -56 528 834
use sg13g2_o21ai_1  _1418_
timestamp 1746816402
transform 1 0 13728 0 -1 21924
box -48 -56 538 834
use sg13g2_a21oi_2  _1419_
timestamp 1746816402
transform 1 0 14208 0 -1 21924
box -48 -56 816 834
use sg13g2_o21ai_1  _1420_
timestamp 1746816402
transform -1 0 18336 0 1 21924
box -48 -56 538 834
use sg13g2_nor2_1  _1421_
timestamp 1746816402
transform -1 0 19296 0 -1 21924
box -48 -56 432 834
use sg13g2_nand2b_1  _1422_
timestamp 1746816402
transform 1 0 18624 0 1 20412
box -48 -56 528 834
use sg13g2_nand2_1  _1423_
timestamp 1746816402
transform 1 0 19008 0 -1 20412
box -48 -56 432 834
use sg13g2_xor2_1  _1424_
timestamp 1746816402
transform 1 0 15936 0 1 9828
box -48 -56 816 834
use sg13g2_a21o_1  _1425_
timestamp 1746816402
transform -1 0 17472 0 1 11340
box -48 -56 720 834
use sg13g2_inv_1  _1426_
timestamp 1746816402
transform -1 0 17280 0 -1 12852
box -48 -56 336 834
use sg13g2_nor2_1  _1427_
timestamp 1746816402
transform 1 0 16992 0 1 8316
box -48 -56 432 834
use sg13g2_a21oi_1  _1428_
timestamp 1746816402
transform 1 0 14976 0 -1 6804
box -48 -56 528 834
use sg13g2_xor2_1  _1429_
timestamp 1746816402
transform 1 0 16608 0 1 5292
box -48 -56 816 834
use sg13g2_xnor2_1  _1430_
timestamp 1746816402
transform 1 0 17376 0 1 5292
box -48 -56 816 834
use sg13g2_xor2_1  _1431_
timestamp 1746816402
transform -1 0 19296 0 -1 9828
box -48 -56 816 834
use sg13g2_xnor2_1  _1432_
timestamp 1746816402
transform -1 0 18528 0 -1 9828
box -48 -56 816 834
use sg13g2_xnor2_1  _1433_
timestamp 1746816402
transform 1 0 16992 0 -1 9828
box -48 -56 816 834
use sg13g2_o21ai_1  _1434_
timestamp 1746816402
transform -1 0 18432 0 1 9828
box -48 -56 538 834
use sg13g2_a21oi_1  _1435_
timestamp 1746816402
transform -1 0 15648 0 -1 11340
box -48 -56 528 834
use sg13g2_o21ai_1  _1436_
timestamp 1746816402
transform -1 0 17472 0 -1 6804
box -48 -56 538 834
use sg13g2_xor2_1  _1437_
timestamp 1746816402
transform 1 0 16224 0 -1 6804
box -48 -56 816 834
use sg13g2_xor2_1  _1438_
timestamp 1746816402
transform -1 0 21408 0 1 9828
box -48 -56 816 834
use sg13g2_xnor2_1  _1439_
timestamp 1746816402
transform 1 0 16512 0 -1 11340
box -48 -56 816 834
use sg13g2_xnor2_1  _1440_
timestamp 1746816402
transform 1 0 16704 0 1 9828
box -48 -56 816 834
use sg13g2_mux2_1  _1441_
timestamp 1746816402
transform 1 0 17280 0 -1 11340
box -48 -56 1008 834
use sg13g2_nor2b_1  _1442_
timestamp 1746816402
transform -1 0 22272 0 1 14364
box -54 -56 528 834
use sg13g2_nor2_1  _1443_
timestamp 1746816402
transform -1 0 21408 0 1 12852
box -48 -56 432 834
use sg13g2_a21oi_2  _1444_
timestamp 1746816402
transform -1 0 21792 0 1 14364
box -48 -56 816 834
use sg13g2_and2_1  _1445_
timestamp 1746816402
transform 1 0 16320 0 1 14364
box -48 -56 528 834
use sg13g2_a221oi_1  _1446_
timestamp 1746816402
transform -1 0 17088 0 -1 15876
box -48 -56 816 834
use sg13g2_a21oi_1  _1447_
timestamp 1746816402
transform 1 0 17184 0 -1 18900
box -48 -56 528 834
use sg13g2_nand2b_1  _1448_
timestamp 1746816402
transform 1 0 17088 0 1 18900
box -48 -56 528 834
use sg13g2_nand2_1  _1449_
timestamp 1746816402
transform -1 0 18912 0 1 18900
box -48 -56 432 834
use sg13g2_a21o_1  _1450_
timestamp 1746816402
transform -1 0 18528 0 1 18900
box -48 -56 720 834
use sg13g2_a21oi_1  _1451_
timestamp 1746816402
transform -1 0 17952 0 -1 20412
box -48 -56 528 834
use sg13g2_a21oi_1  _1452_
timestamp 1746816402
transform -1 0 18528 0 -1 20412
box -48 -56 528 834
use sg13g2_o21ai_1  _1453_
timestamp 1746816402
transform 1 0 19584 0 1 20412
box -48 -56 538 834
use sg13g2_a21oi_2  _1454_
timestamp 1746816402
transform -1 0 18912 0 -1 21924
box -48 -56 816 834
use sg13g2_nor2_1  _1455_
timestamp 1746816402
transform 1 0 12192 0 1 17388
box -48 -56 432 834
use sg13g2_nand2b_2  _1456_
timestamp 1746816402
transform 1 0 11616 0 -1 17388
box -48 -56 816 834
use sg13g2_a22oi_1  _1457_
timestamp 1746816402
transform -1 0 9408 0 1 17388
box -48 -56 624 834
use sg13g2_o21ai_1  _1458_
timestamp 1746816402
transform 1 0 8832 0 -1 18900
box -48 -56 538 834
use sg13g2_nand2_1  _1459_
timestamp 1746816402
transform -1 0 9024 0 1 18900
box -48 -56 432 834
use sg13g2_nor2_1  _1460_
timestamp 1746816402
transform -1 0 9408 0 -1 15876
box -48 -56 432 834
use sg13g2_nand2_2  _1461_
timestamp 1746816402
transform -1 0 13632 0 -1 12852
box -48 -56 624 834
use sg13g2_nor2_1  _1462_
timestamp 1746816402
transform -1 0 8640 0 -1 15876
box -48 -56 432 834
use sg13g2_or2_1  _1463_
timestamp 1746816402
transform 1 0 7968 0 1 14364
box -48 -56 528 834
use sg13g2_a22oi_1  _1464_
timestamp 1746816402
transform 1 0 8448 0 1 14364
box -48 -56 624 834
use sg13g2_o21ai_1  _1465_
timestamp 1746816402
transform 1 0 7776 0 -1 18900
box -48 -56 538 834
use sg13g2_o21ai_1  _1466_
timestamp 1746816402
transform -1 0 10176 0 1 18900
box -48 -56 538 834
use sg13g2_a21o_1  _1467_
timestamp 1746816402
transform -1 0 9696 0 1 18900
box -48 -56 720 834
use sg13g2_a21oi_1  _1468_
timestamp 1746816402
transform -1 0 11520 0 -1 21924
box -48 -56 528 834
use sg13g2_o21ai_1  _1469_
timestamp 1746816402
transform -1 0 10656 0 -1 23436
box -48 -56 538 834
use sg13g2_nor2_1  _1470_
timestamp 1746816402
transform 1 0 6720 0 1 17388
box -48 -56 432 834
use sg13g2_a221oi_1  _1471_
timestamp 1746816402
transform 1 0 7488 0 1 17388
box -48 -56 816 834
use sg13g2_and2_1  _1472_
timestamp 1746816402
transform 1 0 6816 0 -1 18900
box -48 -56 528 834
use sg13g2_o21ai_1  _1473_
timestamp 1746816402
transform -1 0 7488 0 1 14364
box -48 -56 538 834
use sg13g2_and2_1  _1474_
timestamp 1746816402
transform 1 0 2496 0 1 11340
box -48 -56 528 834
use sg13g2_xnor2_1  _1475_
timestamp 1746816402
transform 1 0 2112 0 -1 11340
box -48 -56 816 834
use sg13g2_xnor2_1  _1476_
timestamp 1746816402
transform 1 0 2880 0 -1 11340
box -48 -56 816 834
use sg13g2_nand2_1  _1477_
timestamp 1746816402
transform 1 0 576 0 1 9828
box -48 -56 432 834
use sg13g2_nand2_1  _1478_
timestamp 1746816402
transform 1 0 2208 0 -1 9828
box -48 -56 432 834
use sg13g2_nor2_1  _1479_
timestamp 1746816402
transform -1 0 4416 0 -1 9828
box -48 -56 432 834
use sg13g2_xor2_1  _1480_
timestamp 1746816402
transform 1 0 1248 0 -1 9828
box -48 -56 816 834
use sg13g2_xnor2_1  _1481_
timestamp 1746816402
transform 1 0 1728 0 1 9828
box -48 -56 816 834
use sg13g2_a21oi_1  _1482_
timestamp 1746816402
transform -1 0 3456 0 1 9828
box -48 -56 528 834
use sg13g2_o21ai_1  _1483_
timestamp 1746816402
transform 1 0 3456 0 1 9828
box -48 -56 538 834
use sg13g2_nor2_1  _1484_
timestamp 1746816402
transform -1 0 14592 0 -1 14364
box -48 -56 432 834
use sg13g2_a221oi_1  _1485_
timestamp 1746816402
transform -1 0 8352 0 -1 14364
box -48 -56 816 834
use sg13g2_o21ai_1  _1486_
timestamp 1746816402
transform 1 0 7296 0 -1 18900
box -48 -56 538 834
use sg13g2_o21ai_1  _1487_
timestamp 1746816402
transform -1 0 8160 0 1 18900
box -48 -56 538 834
use sg13g2_a21oi_1  _1488_
timestamp 1746816402
transform -1 0 8064 0 1 20412
box -48 -56 528 834
use sg13g2_o21ai_1  _1489_
timestamp 1746816402
transform -1 0 9024 0 -1 21924
box -48 -56 538 834
use sg13g2_a21oi_1  _1490_
timestamp 1746816402
transform 1 0 7200 0 1 21924
box -48 -56 528 834
use sg13g2_and2_1  _1491_
timestamp 1746816402
transform -1 0 5376 0 -1 15876
box -48 -56 528 834
use sg13g2_a221oi_1  _1492_
timestamp 1746816402
transform 1 0 4896 0 1 14364
box -48 -56 816 834
use sg13g2_or2_1  _1493_
timestamp 1746816402
transform 1 0 3840 0 1 14364
box -48 -56 528 834
use sg13g2_nand2_1  _1494_
timestamp 1746816402
transform -1 0 4896 0 -1 15876
box -48 -56 432 834
use sg13g2_nor2_1  _1495_
timestamp 1746816402
transform 1 0 6144 0 1 12852
box -48 -56 432 834
use sg13g2_nor2_1  _1496_
timestamp 1746816402
transform 1 0 5760 0 -1 12852
box -48 -56 432 834
use sg13g2_a22oi_1  _1497_
timestamp 1746816402
transform 1 0 3648 0 -1 11340
box -48 -56 624 834
use sg13g2_xor2_1  _1498_
timestamp 1746816402
transform 1 0 3936 0 1 9828
box -48 -56 816 834
use sg13g2_xnor2_1  _1499_
timestamp 1746816402
transform 1 0 4704 0 1 9828
box -48 -56 816 834
use sg13g2_and2_1  _1500_
timestamp 1746816402
transform 1 0 5760 0 -1 8316
box -48 -56 528 834
use sg13g2_or2_1  _1501_
timestamp 1746816402
transform 1 0 4512 0 1 6804
box -48 -56 528 834
use sg13g2_nand2b_1  _1502_
timestamp 1746816402
transform 1 0 5856 0 -1 6804
box -48 -56 528 834
use sg13g2_o21ai_1  _1503_
timestamp 1746816402
transform 1 0 3072 0 -1 9828
box -48 -56 538 834
use sg13g2_xnor2_1  _1504_
timestamp 1746816402
transform -1 0 6624 0 1 6804
box -48 -56 816 834
use sg13g2_o21ai_1  _1505_
timestamp 1746816402
transform 1 0 5568 0 -1 11340
box -48 -56 538 834
use sg13g2_a21oi_1  _1506_
timestamp 1746816402
transform -1 0 5760 0 1 11340
box -48 -56 528 834
use sg13g2_nor3_1  _1507_
timestamp 1746816402
transform -1 0 10752 0 -1 12852
box -48 -56 528 834
use sg13g2_nor2_1  _1508_
timestamp 1746816402
transform 1 0 6144 0 -1 12852
box -48 -56 432 834
use sg13g2_o21ai_1  _1509_
timestamp 1746816402
transform -1 0 6144 0 1 12852
box -48 -56 538 834
use sg13g2_and2_1  _1510_
timestamp 1746816402
transform -1 0 4032 0 -1 15876
box -48 -56 528 834
use sg13g2_o21ai_1  _1511_
timestamp 1746816402
transform -1 0 4512 0 -1 15876
box -48 -56 538 834
use sg13g2_a21oi_1  _1512_
timestamp 1746816402
transform 1 0 4320 0 1 18900
box -48 -56 528 834
use sg13g2_o21ai_1  _1513_
timestamp 1746816402
transform -1 0 3072 0 -1 20412
box -48 -56 538 834
use sg13g2_a21oi_1  _1514_
timestamp 1746816402
transform 1 0 2208 0 1 20412
box -48 -56 528 834
use sg13g2_and2_1  _1515_
timestamp 1746816402
transform -1 0 4416 0 -1 17388
box -48 -56 528 834
use sg13g2_a221oi_1  _1516_
timestamp 1746816402
transform 1 0 5664 0 -1 17388
box -48 -56 816 834
use sg13g2_nor2_1  _1517_
timestamp 1746816402
transform -1 0 11328 0 -1 14364
box -48 -56 432 834
use sg13g2_nor2_1  _1518_
timestamp 1746816402
transform 1 0 9216 0 1 11340
box -48 -56 432 834
use sg13g2_and2_1  _1519_
timestamp 1746816402
transform -1 0 10272 0 1 5292
box -48 -56 528 834
use sg13g2_xor2_1  _1520_
timestamp 1746816402
transform 1 0 8256 0 -1 6804
box -48 -56 816 834
use sg13g2_a21o_1  _1521_
timestamp 1746816402
transform -1 0 7296 0 1 6804
box -48 -56 720 834
use sg13g2_xnor2_1  _1522_
timestamp 1746816402
transform -1 0 10560 0 -1 6804
box -48 -56 816 834
use sg13g2_or2_1  _1523_
timestamp 1746816402
transform -1 0 6048 0 -1 9828
box -48 -56 528 834
use sg13g2_o21ai_1  _1524_
timestamp 1746816402
transform 1 0 5088 0 -1 9828
box -48 -56 538 834
use sg13g2_nor2_1  _1525_
timestamp 1746816402
transform -1 0 8928 0 -1 8316
box -48 -56 432 834
use sg13g2_xnor2_1  _1526_
timestamp 1746816402
transform 1 0 7008 0 -1 8316
box -48 -56 816 834
use sg13g2_xnor2_1  _1527_
timestamp 1746816402
transform 1 0 7776 0 -1 8316
box -48 -56 816 834
use sg13g2_xnor2_1  _1528_
timestamp 1746816402
transform 1 0 9024 0 -1 6804
box -48 -56 816 834
use sg13g2_a21oi_1  _1529_
timestamp 1746816402
transform 1 0 9504 0 1 12852
box -48 -56 528 834
use sg13g2_nor3_1  _1530_
timestamp 1746816402
transform -1 0 9696 0 -1 14364
box -48 -56 528 834
use sg13g2_nor3_1  _1531_
timestamp 1746816402
transform 1 0 8736 0 -1 14364
box -48 -56 528 834
use sg13g2_and2_1  _1532_
timestamp 1746816402
transform 1 0 3264 0 1 15876
box -48 -56 528 834
use sg13g2_o21ai_1  _1533_
timestamp 1746816402
transform -1 0 4512 0 -1 18900
box -48 -56 538 834
use sg13g2_o21ai_1  _1534_
timestamp 1746816402
transform -1 0 3168 0 1 17388
box -48 -56 538 834
use sg13g2_a21oi_1  _1535_
timestamp 1746816402
transform -1 0 3744 0 -1 21924
box -48 -56 528 834
use sg13g2_o21ai_1  _1536_
timestamp 1746816402
transform -1 0 2784 0 1 21924
box -48 -56 538 834
use sg13g2_a21oi_1  _1537_
timestamp 1746816402
transform 1 0 2016 0 -1 23436
box -48 -56 528 834
use sg13g2_nor2_1  _1538_
timestamp 1746816402
transform -1 0 11904 0 1 15876
box -48 -56 432 834
use sg13g2_a221oi_1  _1539_
timestamp 1746816402
transform 1 0 11232 0 -1 15876
box -48 -56 816 834
use sg13g2_or2_1  _1540_
timestamp 1746816402
transform 1 0 11520 0 1 14364
box -48 -56 528 834
use sg13g2_nor2_1  _1541_
timestamp 1746816402
transform -1 0 12288 0 -1 12852
box -48 -56 432 834
use sg13g2_a21oi_1  _1542_
timestamp 1746816402
transform -1 0 8736 0 1 6804
box -48 -56 528 834
use sg13g2_xnor2_1  _1543_
timestamp 1746816402
transform 1 0 11136 0 -1 6804
box -48 -56 816 834
use sg13g2_xor2_1  _1544_
timestamp 1746816402
transform 1 0 11040 0 1 6804
box -48 -56 816 834
use sg13g2_nand2_1  _1545_
timestamp 1746816402
transform -1 0 12000 0 1 3780
box -48 -56 432 834
use sg13g2_xnor2_1  _1546_
timestamp 1746816402
transform -1 0 12096 0 -1 5292
box -48 -56 816 834
use sg13g2_a21oi_1  _1547_
timestamp 1746816402
transform -1 0 9792 0 1 5292
box -48 -56 528 834
use sg13g2_xnor2_1  _1548_
timestamp 1746816402
transform 1 0 10848 0 1 5292
box -48 -56 816 834
use sg13g2_a21oi_1  _1549_
timestamp 1746816402
transform -1 0 12288 0 -1 8316
box -48 -56 528 834
use sg13g2_o21ai_1  _1550_
timestamp 1746816402
transform -1 0 11808 0 -1 8316
box -48 -56 538 834
use sg13g2_o21ai_1  _1551_
timestamp 1746816402
transform -1 0 11904 0 -1 12852
box -48 -56 538 834
use sg13g2_nor2_1  _1552_
timestamp 1746816402
transform -1 0 12672 0 -1 14364
box -48 -56 432 834
use sg13g2_a21oi_1  _1553_
timestamp 1746816402
transform -1 0 14112 0 -1 14364
box -48 -56 528 834
use sg13g2_a22oi_1  _1554_
timestamp 1746816402
transform 1 0 11520 0 -1 14364
box -48 -56 624 834
use sg13g2_o21ai_1  _1555_
timestamp 1746816402
transform -1 0 12480 0 1 14364
box -48 -56 538 834
use sg13g2_a21oi_1  _1556_
timestamp 1746816402
transform 1 0 6720 0 -1 21924
box -48 -56 528 834
use sg13g2_o21ai_1  _1557_
timestamp 1746816402
transform 1 0 5472 0 1 21924
box -48 -56 538 834
use sg13g2_a21oi_1  _1558_
timestamp 1746816402
transform 1 0 5472 0 -1 23436
box -48 -56 528 834
use sg13g2_and2_1  _1559_
timestamp 1746816402
transform 1 0 13152 0 -1 14364
box -48 -56 528 834
use sg13g2_a221oi_1  _1560_
timestamp 1746816402
transform 1 0 13824 0 1 14364
box -48 -56 816 834
use sg13g2_or2_1  _1561_
timestamp 1746816402
transform 1 0 14688 0 1 14364
box -48 -56 528 834
use sg13g2_nor2_1  _1562_
timestamp 1746816402
transform -1 0 16224 0 -1 12852
box -48 -56 432 834
use sg13g2_nand2b_1  _1563_
timestamp 1746816402
transform 1 0 11616 0 1 5292
box -48 -56 528 834
use sg13g2_o21ai_1  _1564_
timestamp 1746816402
transform 1 0 11904 0 -1 6804
box -48 -56 538 834
use sg13g2_nor2_1  _1565_
timestamp 1746816402
transform -1 0 15264 0 -1 8316
box -48 -56 432 834
use sg13g2_xnor2_1  _1566_
timestamp 1746816402
transform 1 0 14112 0 -1 8316
box -48 -56 816 834
use sg13g2_xnor2_1  _1567_
timestamp 1746816402
transform 1 0 14592 0 1 6804
box -48 -56 816 834
use sg13g2_and2_1  _1568_
timestamp 1746816402
transform -1 0 19392 0 1 5292
box -48 -56 528 834
use sg13g2_xor2_1  _1569_
timestamp 1746816402
transform 1 0 17856 0 -1 6804
box -48 -56 816 834
use sg13g2_o21ai_1  _1570_
timestamp 1746816402
transform -1 0 10848 0 1 5292
box -48 -56 538 834
use sg13g2_xor2_1  _1571_
timestamp 1746816402
transform -1 0 18912 0 1 5292
box -48 -56 816 834
use sg13g2_a21oi_1  _1572_
timestamp 1746816402
transform 1 0 15360 0 1 6804
box -48 -56 528 834
use sg13g2_o21ai_1  _1573_
timestamp 1746816402
transform 1 0 15840 0 1 6804
box -48 -56 538 834
use sg13g2_o21ai_1  _1574_
timestamp 1746816402
transform -1 0 15168 0 1 12852
box -48 -56 538 834
use sg13g2_nor3_1  _1575_
timestamp 1746816402
transform -1 0 15648 0 1 12852
box -48 -56 528 834
use sg13g2_nor2_1  _1576_
timestamp 1746816402
transform -1 0 15552 0 1 14364
box -48 -56 432 834
use sg13g2_a22oi_1  _1577_
timestamp 1746816402
transform 1 0 14592 0 -1 14364
box -48 -56 624 834
use sg13g2_o21ai_1  _1578_
timestamp 1746816402
transform -1 0 16128 0 1 18900
box -48 -56 538 834
use sg13g2_a21oi_1  _1579_
timestamp 1746816402
transform 1 0 6816 0 1 18900
box -48 -56 528 834
use sg13g2_o21ai_1  _1580_
timestamp 1746816402
transform -1 0 6048 0 -1 20412
box -48 -56 538 834
use sg13g2_a21oi_1  _1581_
timestamp 1746816402
transform 1 0 5088 0 -1 20412
box -48 -56 528 834
use sg13g2_o21ai_1  _1582_
timestamp 1746816402
transform 1 0 16224 0 1 12852
box -48 -56 538 834
use sg13g2_nand2_1  _1583_
timestamp 1746816402
transform -1 0 21120 0 1 5292
box -48 -56 432 834
use sg13g2_nor2_1  _1584_
timestamp 1746816402
transform 1 0 20352 0 1 5292
box -48 -56 432 834
use sg13g2_xnor2_1  _1585_
timestamp 1746816402
transform -1 0 20640 0 -1 6804
box -48 -56 816 834
use sg13g2_a21oi_1  _1586_
timestamp 1746816402
transform -1 0 19008 0 -1 5292
box -48 -56 528 834
use sg13g2_xnor2_1  _1587_
timestamp 1746816402
transform -1 0 19872 0 -1 6804
box -48 -56 816 834
use sg13g2_a21oi_1  _1588_
timestamp 1746816402
transform -1 0 14592 0 1 6804
box -48 -56 528 834
use sg13g2_nand2b_1  _1589_
timestamp 1746816402
transform -1 0 18624 0 -1 8316
box -48 -56 528 834
use sg13g2_nor2b_1  _1590_
timestamp 1746816402
transform -1 0 18144 0 -1 8316
box -54 -56 528 834
use sg13g2_xnor2_1  _1591_
timestamp 1746816402
transform 1 0 17184 0 1 6804
box -48 -56 816 834
use sg13g2_xnor2_1  _1592_
timestamp 1746816402
transform 1 0 17952 0 1 6804
box -48 -56 816 834
use sg13g2_xnor2_1  _1593_
timestamp 1746816402
transform -1 0 19488 0 1 6804
box -48 -56 816 834
use sg13g2_o21ai_1  _1594_
timestamp 1746816402
transform -1 0 16224 0 1 12852
box -48 -56 538 834
use sg13g2_nor2_1  _1595_
timestamp 1746816402
transform -1 0 17184 0 1 14364
box -48 -56 432 834
use sg13g2_a21oi_1  _1596_
timestamp 1746816402
transform 1 0 15744 0 -1 14364
box -48 -56 528 834
use sg13g2_a22oi_1  _1597_
timestamp 1746816402
transform -1 0 16032 0 1 15876
box -48 -56 624 834
use sg13g2_o21ai_1  _1598_
timestamp 1746816402
transform 1 0 14784 0 -1 18900
box -48 -56 538 834
use sg13g2_o21ai_1  _1599_
timestamp 1746816402
transform 1 0 14304 0 1 17388
box -48 -56 538 834
use sg13g2_a221oi_1  _1600_
timestamp 1746816402
transform 1 0 15360 0 -1 17388
box -48 -56 816 834
use sg13g2_o21ai_1  _1601_
timestamp 1746816402
transform 1 0 15456 0 1 17388
box -48 -56 538 834
use sg13g2_nor2_1  _1602_
timestamp 1746816402
transform -1 0 16512 0 -1 17388
box -48 -56 432 834
use sg13g2_o21ai_1  _1603_
timestamp 1746816402
transform 1 0 14784 0 1 20412
box -48 -56 538 834
use sg13g2_a21oi_1  _1604_
timestamp 1746816402
transform 1 0 15456 0 1 21924
box -48 -56 528 834
use sg13g2_nor2_2  _1605_
timestamp 1746816402
transform -1 0 14208 0 1 21924
box -48 -56 624 834
use sg13g2_nand2_1  _1606_
timestamp 1746816402
transform 1 0 17280 0 -1 17388
box -48 -56 432 834
use sg13g2_a22oi_1  _1607_
timestamp 1746816402
transform 1 0 16128 0 1 15876
box -48 -56 624 834
use sg13g2_a21oi_1  _1608_
timestamp 1746816402
transform 1 0 18336 0 -1 17388
box -48 -56 528 834
use sg13g2_nand3_1  _1609_
timestamp 1746816402
transform -1 0 19296 0 -1 17388
box -48 -56 528 834
use sg13g2_o21ai_1  _1610_
timestamp 1746816402
transform 1 0 15552 0 1 11340
box -48 -56 538 834
use sg13g2_nor2_1  _1611_
timestamp 1746816402
transform -1 0 15744 0 -1 14364
box -48 -56 432 834
use sg13g2_nor2_1  _1612_
timestamp 1746816402
transform 1 0 17472 0 1 11340
box -48 -56 432 834
use sg13g2_o21ai_1  _1613_
timestamp 1746816402
transform 1 0 17184 0 -1 8316
box -48 -56 538 834
use sg13g2_xor2_1  _1614_
timestamp 1746816402
transform -1 0 21696 0 -1 11340
box -48 -56 816 834
use sg13g2_o21ai_1  _1615_
timestamp 1746816402
transform 1 0 20640 0 -1 6804
box -48 -56 538 834
use sg13g2_xnor2_1  _1616_
timestamp 1746816402
transform -1 0 22368 0 -1 9828
box -48 -56 816 834
use sg13g2_xnor2_1  _1617_
timestamp 1746816402
transform -1 0 21600 0 -1 9828
box -48 -56 816 834
use sg13g2_xnor2_1  _1618_
timestamp 1746816402
transform -1 0 21024 0 1 11340
box -48 -56 816 834
use sg13g2_or2_1  _1619_
timestamp 1746816402
transform -1 0 19200 0 -1 11340
box -48 -56 528 834
use sg13g2_a21oi_1  _1620_
timestamp 1746816402
transform 1 0 18240 0 -1 11340
box -48 -56 528 834
use sg13g2_a21oi_1  _1621_
timestamp 1746816402
transform 1 0 18048 0 1 11340
box -48 -56 528 834
use sg13g2_nand2b_1  _1622_
timestamp 1746816402
transform 1 0 17760 0 1 15876
box -48 -56 528 834
use sg13g2_o21ai_1  _1623_
timestamp 1746816402
transform -1 0 19680 0 1 15876
box -48 -56 538 834
use sg13g2_o21ai_1  _1624_
timestamp 1746816402
transform 1 0 18240 0 1 17388
box -48 -56 538 834
use sg13g2_a21o_1  _1625_
timestamp 1746816402
transform -1 0 18336 0 -1 17388
box -48 -56 720 834
use sg13g2_a21oi_1  _1626_
timestamp 1746816402
transform -1 0 18624 0 1 20412
box -48 -56 528 834
use sg13g2_o21ai_1  _1627_
timestamp 1746816402
transform 1 0 17664 0 1 20412
box -48 -56 538 834
use sg13g2_a21oi_2  _1628_
timestamp 1746816402
transform 1 0 18336 0 1 21924
box -48 -56 816 834
use sg13g2_nor2_2  _1629_
timestamp 1746816402
transform 1 0 15744 0 -1 15876
box -48 -56 624 834
use sg13g2_a22oi_1  _1630_
timestamp 1746816402
transform 1 0 9024 0 1 15876
box -48 -56 624 834
use sg13g2_o21ai_1  _1631_
timestamp 1746816402
transform 1 0 9408 0 1 17388
box -48 -56 538 834
use sg13g2_and2_1  _1632_
timestamp 1746816402
transform 1 0 5760 0 1 11340
box -48 -56 528 834
use sg13g2_xnor2_1  _1633_
timestamp 1746816402
transform 1 0 6720 0 1 11340
box -48 -56 816 834
use sg13g2_xnor2_1  _1634_
timestamp 1746816402
transform -1 0 8256 0 1 11340
box -48 -56 816 834
use sg13g2_nand2_1  _1635_
timestamp 1746816402
transform -1 0 6528 0 -1 9828
box -48 -56 432 834
use sg13g2_nand2_1  _1636_
timestamp 1746816402
transform 1 0 6720 0 -1 9828
box -48 -56 432 834
use sg13g2_nor2_1  _1637_
timestamp 1746816402
transform 1 0 6624 0 -1 11340
box -48 -56 432 834
use sg13g2_xor2_1  _1638_
timestamp 1746816402
transform 1 0 5472 0 1 9828
box -48 -56 816 834
use sg13g2_xnor2_1  _1639_
timestamp 1746816402
transform -1 0 7008 0 1 9828
box -48 -56 816 834
use sg13g2_o21ai_1  _1640_
timestamp 1746816402
transform -1 0 8064 0 -1 11340
box -48 -56 538 834
use sg13g2_a21oi_1  _1641_
timestamp 1746816402
transform -1 0 6720 0 1 11340
box -48 -56 528 834
use sg13g2_a21oi_1  _1642_
timestamp 1746816402
transform 1 0 7104 0 1 12852
box -48 -56 528 834
use sg13g2_o21ai_1  _1643_
timestamp 1746816402
transform 1 0 6624 0 1 12852
box -48 -56 538 834
use sg13g2_o21ai_1  _1644_
timestamp 1746816402
transform -1 0 10848 0 1 15876
box -48 -56 538 834
use sg13g2_a22oi_1  _1645_
timestamp 1746816402
transform 1 0 9504 0 -1 17388
box -48 -56 624 834
use sg13g2_o21ai_1  _1646_
timestamp 1746816402
transform 1 0 10080 0 -1 21924
box -48 -56 538 834
use sg13g2_and2_1  _1647_
timestamp 1746816402
transform 1 0 10272 0 1 21924
box -48 -56 528 834
use sg13g2_o21ai_1  _1648_
timestamp 1746816402
transform -1 0 11136 0 -1 23436
box -48 -56 538 834
use sg13g2_a22oi_1  _1649_
timestamp 1746816402
transform 1 0 7008 0 -1 11340
box -48 -56 624 834
use sg13g2_xor2_1  _1650_
timestamp 1746816402
transform 1 0 8640 0 -1 9828
box -48 -56 816 834
use sg13g2_xor2_1  _1651_
timestamp 1746816402
transform 1 0 8352 0 1 9828
box -48 -56 816 834
use sg13g2_and2_1  _1652_
timestamp 1746816402
transform 1 0 7776 0 1 9828
box -48 -56 528 834
use sg13g2_xor2_1  _1653_
timestamp 1746816402
transform 1 0 7104 0 -1 9828
box -48 -56 816 834
use sg13g2_o21ai_1  _1654_
timestamp 1746816402
transform 1 0 7008 0 1 9828
box -48 -56 538 834
use sg13g2_xnor2_1  _1655_
timestamp 1746816402
transform 1 0 7872 0 -1 9828
box -48 -56 816 834
use sg13g2_a21oi_1  _1656_
timestamp 1746816402
transform -1 0 9600 0 1 9828
box -48 -56 528 834
use sg13g2_o21ai_1  _1657_
timestamp 1746816402
transform -1 0 8832 0 -1 11340
box -48 -56 538 834
use sg13g2_nor2_1  _1658_
timestamp 1746816402
transform 1 0 8640 0 1 15876
box -48 -56 432 834
use sg13g2_a221oi_1  _1659_
timestamp 1746816402
transform -1 0 8640 0 -1 17388
box -48 -56 816 834
use sg13g2_a22oi_1  _1660_
timestamp 1746816402
transform -1 0 9216 0 -1 12852
box -48 -56 624 834
use sg13g2_o21ai_1  _1661_
timestamp 1746816402
transform 1 0 8256 0 -1 18900
box -48 -56 538 834
use sg13g2_a221oi_1  _1662_
timestamp 1746816402
transform -1 0 9408 0 -1 17388
box -48 -56 816 834
use sg13g2_o21ai_1  _1663_
timestamp 1746816402
transform -1 0 8544 0 1 20412
box -48 -56 538 834
use sg13g2_nand2_1  _1664_
timestamp 1746816402
transform -1 0 7680 0 -1 21924
box -48 -56 432 834
use sg13g2_a21oi_1  _1665_
timestamp 1746816402
transform 1 0 8160 0 1 21924
box -48 -56 528 834
use sg13g2_nand2_1  _1666_
timestamp 1746816402
transform 1 0 9696 0 1 6804
box -48 -56 432 834
use sg13g2_xnor2_1  _1667_
timestamp 1746816402
transform -1 0 10848 0 1 6804
box -48 -56 816 834
use sg13g2_a21oi_1  _1668_
timestamp 1746816402
transform -1 0 8544 0 1 8316
box -48 -56 528 834
use sg13g2_xor2_1  _1669_
timestamp 1746816402
transform 1 0 10176 0 -1 8316
box -48 -56 816 834
use sg13g2_or2_1  _1670_
timestamp 1746816402
transform 1 0 9120 0 1 8316
box -48 -56 528 834
use sg13g2_o21ai_1  _1671_
timestamp 1746816402
transform 1 0 9408 0 -1 9828
box -48 -56 538 834
use sg13g2_nor2_1  _1672_
timestamp 1746816402
transform -1 0 14496 0 1 8316
box -48 -56 432 834
use sg13g2_xnor2_1  _1673_
timestamp 1746816402
transform -1 0 14112 0 1 8316
box -48 -56 816 834
use sg13g2_xnor2_1  _1674_
timestamp 1746816402
transform -1 0 11616 0 -1 9828
box -48 -56 816 834
use sg13g2_a21oi_1  _1675_
timestamp 1746816402
transform -1 0 11232 0 1 8316
box -48 -56 528 834
use sg13g2_o21ai_1  _1676_
timestamp 1746816402
transform -1 0 10848 0 -1 9828
box -48 -56 538 834
use sg13g2_nand2b_1  _1677_
timestamp 1746816402
transform -1 0 11424 0 -1 12852
box -48 -56 528 834
use sg13g2_and2_1  _1678_
timestamp 1746816402
transform 1 0 5376 0 -1 15876
box -48 -56 528 834
use sg13g2_a221oi_1  _1679_
timestamp 1746816402
transform 1 0 5856 0 1 14364
box -48 -56 816 834
use sg13g2_o21ai_1  _1680_
timestamp 1746816402
transform 1 0 10464 0 -1 14364
box -48 -56 538 834
use sg13g2_a21o_1  _1681_
timestamp 1746816402
transform 1 0 10272 0 1 12852
box -48 -56 720 834
use sg13g2_a221oi_1  _1682_
timestamp 1746816402
transform -1 0 10368 0 1 15876
box -48 -56 816 834
use sg13g2_o21ai_1  _1683_
timestamp 1746816402
transform -1 0 4320 0 1 18900
box -48 -56 538 834
use sg13g2_nand2_1  _1684_
timestamp 1746816402
transform -1 0 2112 0 1 18900
box -48 -56 432 834
use sg13g2_a21oi_1  _1685_
timestamp 1746816402
transform -1 0 3648 0 1 20412
box -48 -56 528 834
use sg13g2_a21oi_2  _1686_
timestamp 1746816402
transform 1 0 12576 0 1 8316
box -48 -56 816 834
use sg13g2_xnor2_1  _1687_
timestamp 1746816402
transform -1 0 20256 0 1 6804
box -48 -56 816 834
use sg13g2_xnor2_1  _1688_
timestamp 1746816402
transform 1 0 19008 0 -1 8316
box -48 -56 816 834
use sg13g2_and2_1  _1689_
timestamp 1746816402
transform 1 0 22176 0 -1 6804
box -48 -56 528 834
use sg13g2_or2_1  _1690_
timestamp 1746816402
transform -1 0 22560 0 1 6804
box -48 -56 528 834
use sg13g2_nand2b_1  _1691_
timestamp 1746816402
transform -1 0 22176 0 -1 6804
box -48 -56 528 834
use sg13g2_o21ai_1  _1692_
timestamp 1746816402
transform 1 0 10560 0 -1 6804
box -48 -56 538 834
use sg13g2_xnor2_1  _1693_
timestamp 1746816402
transform 1 0 20352 0 1 6804
box -48 -56 816 834
use sg13g2_a21oi_1  _1694_
timestamp 1746816402
transform 1 0 21120 0 1 6804
box -48 -56 528 834
use sg13g2_o21ai_1  _1695_
timestamp 1746816402
transform -1 0 20736 0 -1 8316
box -48 -56 538 834
use sg13g2_and2_1  _1696_
timestamp 1746816402
transform 1 0 5184 0 1 15876
box -48 -56 528 834
use sg13g2_a221oi_1  _1697_
timestamp 1746816402
transform 1 0 5664 0 1 15876
box -48 -56 816 834
use sg13g2_nor2_1  _1698_
timestamp 1746816402
transform -1 0 12096 0 -1 11340
box -48 -56 432 834
use sg13g2_a21oi_1  _1699_
timestamp 1746816402
transform 1 0 11712 0 1 11340
box -48 -56 528 834
use sg13g2_o21ai_1  _1700_
timestamp 1746816402
transform -1 0 7104 0 1 15876
box -48 -56 538 834
use sg13g2_a221oi_1  _1701_
timestamp 1746816402
transform -1 0 8640 0 1 15876
box -48 -56 816 834
use sg13g2_o21ai_1  _1702_
timestamp 1746816402
transform 1 0 4416 0 -1 21924
box -48 -56 538 834
use sg13g2_nand2_1  _1703_
timestamp 1746816402
transform -1 0 1440 0 1 20412
box -48 -56 432 834
use sg13g2_a21oi_1  _1704_
timestamp 1746816402
transform -1 0 2304 0 1 21924
box -48 -56 528 834
use sg13g2_nand2b_1  _1705_
timestamp 1746816402
transform 1 0 18432 0 1 8316
box -48 -56 528 834
use sg13g2_o21ai_1  _1706_
timestamp 1746816402
transform 1 0 19776 0 -1 8316
box -48 -56 538 834
use sg13g2_nor2_1  _1707_
timestamp 1746816402
transform 1 0 19104 0 1 9828
box -48 -56 432 834
use sg13g2_xor2_1  _1708_
timestamp 1746816402
transform 1 0 19296 0 -1 9828
box -48 -56 816 834
use sg13g2_xnor2_1  _1709_
timestamp 1746816402
transform 1 0 19200 0 1 8316
box -48 -56 816 834
use sg13g2_a21oi_1  _1710_
timestamp 1746816402
transform 1 0 23712 0 -1 6804
box -48 -56 528 834
use sg13g2_nor2_1  _1711_
timestamp 1746816402
transform 1 0 24960 0 -1 8316
box -48 -56 432 834
use sg13g2_xor2_1  _1712_
timestamp 1746816402
transform 1 0 22656 0 1 6804
box -48 -56 816 834
use sg13g2_xnor2_1  _1713_
timestamp 1746816402
transform -1 0 23712 0 -1 8316
box -48 -56 816 834
use sg13g2_a21oi_1  _1714_
timestamp 1746816402
transform 1 0 19968 0 1 8316
box -48 -56 528 834
use sg13g2_o21ai_1  _1715_
timestamp 1746816402
transform -1 0 20064 0 1 9828
box -48 -56 538 834
use sg13g2_a21oi_1  _1716_
timestamp 1746816402
transform 1 0 14208 0 1 11340
box -48 -56 528 834
use sg13g2_o21ai_1  _1717_
timestamp 1746816402
transform 1 0 13440 0 1 11340
box -48 -56 538 834
use sg13g2_a22oi_1  _1718_
timestamp 1746816402
transform 1 0 10656 0 -1 15876
box -48 -56 624 834
use sg13g2_o21ai_1  _1719_
timestamp 1746816402
transform -1 0 11520 0 1 15876
box -48 -56 538 834
use sg13g2_o21ai_1  _1720_
timestamp 1746816402
transform -1 0 11424 0 -1 18900
box -48 -56 538 834
use sg13g2_a21oi_1  _1721_
timestamp 1746816402
transform -1 0 10944 0 -1 18900
box -48 -56 528 834
use sg13g2_o21ai_1  _1722_
timestamp 1746816402
transform 1 0 10752 0 1 17388
box -48 -56 538 834
use sg13g2_a21oi_1  _1723_
timestamp 1746816402
transform 1 0 10944 0 1 18900
box -48 -56 528 834
use sg13g2_o21ai_1  _1724_
timestamp 1746816402
transform -1 0 6720 0 -1 21924
box -48 -56 538 834
use sg13g2_a21oi_1  _1725_
timestamp 1746816402
transform 1 0 5952 0 1 21924
box -48 -56 528 834
use sg13g2_nor2_1  _1726_
timestamp 1746816402
transform 1 0 768 0 -1 23436
box -48 -56 432 834
use sg13g2_xnor2_1  _1727_
timestamp 1746816402
transform -1 0 25632 0 1 8316
box -48 -56 816 834
use sg13g2_a221oi_1  _1728_
timestamp 1746816402
transform 1 0 23712 0 -1 8316
box -48 -56 816 834
use sg13g2_nor2_1  _1729_
timestamp 1746816402
transform -1 0 25728 0 -1 8316
box -48 -56 432 834
use sg13g2_nor3_1  _1730_
timestamp 1746816402
transform -1 0 24960 0 -1 8316
box -48 -56 528 834
use sg13g2_xor2_1  _1731_
timestamp 1746816402
transform 1 0 24096 0 1 8316
box -48 -56 816 834
use sg13g2_a21oi_2  _1732_
timestamp 1746816402
transform -1 0 20832 0 -1 9828
box -48 -56 816 834
use sg13g2_nor2b_1  _1733_
timestamp 1746816402
transform 1 0 23136 0 -1 9828
box -54 -56 528 834
use sg13g2_nand2b_1  _1734_
timestamp 1746816402
transform -1 0 23616 0 1 9828
box -48 -56 528 834
use sg13g2_xnor2_1  _1735_
timestamp 1746816402
transform 1 0 22368 0 -1 9828
box -48 -56 816 834
use sg13g2_inv_1  _1736_
timestamp 1746816402
transform -1 0 23904 0 1 9828
box -48 -56 336 834
use sg13g2_xnor2_1  _1737_
timestamp 1746816402
transform 1 0 23616 0 -1 9828
box -48 -56 816 834
use sg13g2_xnor2_1  _1738_
timestamp 1746816402
transform -1 0 25152 0 -1 9828
box -48 -56 816 834
use sg13g2_o21ai_1  _1739_
timestamp 1746816402
transform -1 0 17952 0 1 9828
box -48 -56 538 834
use sg13g2_a21oi_1  _1740_
timestamp 1746816402
transform 1 0 14208 0 1 12852
box -48 -56 528 834
use sg13g2_nand2_1  _1741_
timestamp 1746816402
transform -1 0 14592 0 -1 15876
box -48 -56 432 834
use sg13g2_a22oi_1  _1742_
timestamp 1746816402
transform -1 0 13440 0 -1 15876
box -48 -56 624 834
use sg13g2_nand2_1  _1743_
timestamp 1746816402
transform 1 0 13440 0 -1 17388
box -48 -56 432 834
use sg13g2_o21ai_1  _1744_
timestamp 1746816402
transform -1 0 13824 0 1 17388
box -48 -56 538 834
use sg13g2_a221oi_1  _1745_
timestamp 1746816402
transform 1 0 13824 0 -1 17388
box -48 -56 816 834
use sg13g2_o21ai_1  _1746_
timestamp 1746816402
transform -1 0 14304 0 1 17388
box -48 -56 538 834
use sg13g2_nor2_1  _1747_
timestamp 1746816402
transform -1 0 13344 0 1 17388
box -48 -56 432 834
use sg13g2_o21ai_1  _1748_
timestamp 1746816402
transform -1 0 7008 0 -1 20412
box -48 -56 538 834
use sg13g2_a21oi_1  _1749_
timestamp 1746816402
transform 1 0 6048 0 -1 20412
box -48 -56 528 834
use sg13g2_nor2_1  _1750_
timestamp 1746816402
transform 1 0 5568 0 1 20412
box -48 -56 432 834
use sg13g2_o21ai_1  _1751_
timestamp 1746816402
transform -1 0 23136 0 1 9828
box -48 -56 538 834
use sg13g2_xor2_1  _1752_
timestamp 1746816402
transform -1 0 27264 0 1 9828
box -48 -56 816 834
use sg13g2_a21oi_1  _1753_
timestamp 1746816402
transform 1 0 25152 0 -1 9828
box -48 -56 528 834
use sg13g2_nor2b_1  _1754_
timestamp 1746816402
transform 1 0 27264 0 1 9828
box -54 -56 528 834
use sg13g2_xnor2_1  _1755_
timestamp 1746816402
transform -1 0 26496 0 1 9828
box -48 -56 816 834
use sg13g2_nor3_1  _1756_
timestamp 1746816402
transform -1 0 25056 0 -1 11340
box -48 -56 528 834
use sg13g2_o21ai_1  _1757_
timestamp 1746816402
transform 1 0 25056 0 -1 11340
box -48 -56 538 834
use sg13g2_nor2b_1  _1758_
timestamp 1746816402
transform -1 0 26016 0 -1 11340
box -54 -56 528 834
use sg13g2_xnor2_1  _1759_
timestamp 1746816402
transform -1 0 25632 0 1 9828
box -48 -56 816 834
use sg13g2_o21ai_1  _1760_
timestamp 1746816402
transform -1 0 23136 0 -1 11340
box -48 -56 538 834
use sg13g2_nand3b_1  _1761_
timestamp 1746816402
transform -1 0 24576 0 1 9828
box -48 -56 720 834
use sg13g2_a21o_1  _1762_
timestamp 1746816402
transform 1 0 21984 0 -1 11340
box -48 -56 720 834
use sg13g2_a221oi_1  _1763_
timestamp 1746816402
transform 1 0 16032 0 1 11340
box -48 -56 816 834
use sg13g2_a22oi_1  _1764_
timestamp 1746816402
transform -1 0 15456 0 1 15876
box -48 -56 624 834
use sg13g2_o21ai_1  _1765_
timestamp 1746816402
transform 1 0 14784 0 1 17388
box -48 -56 538 834
use sg13g2_nand2_1  _1766_
timestamp 1746816402
transform 1 0 15264 0 -1 18900
box -48 -56 432 834
use sg13g2_o21ai_1  _1767_
timestamp 1746816402
transform 1 0 15168 0 1 18900
box -48 -56 538 834
use sg13g2_or3_1  _1768_
timestamp 1746816402
transform -1 0 16320 0 -1 18900
box -48 -56 720 834
use sg13g2_o21ai_1  _1769_
timestamp 1746816402
transform 1 0 14304 0 -1 18900
box -48 -56 538 834
use sg13g2_inv_1  _1770_
timestamp 1746816402
transform 1 0 14976 0 -1 21924
box -48 -56 336 834
use sg13g2_a21oi_1  _1771_
timestamp 1746816402
transform -1 0 15744 0 1 20412
box -48 -56 528 834
use sg13g2_o21ai_1  _1772_
timestamp 1746816402
transform 1 0 15264 0 -1 21924
box -48 -56 538 834
use sg13g2_a21oi_2  _1773_
timestamp 1746816402
transform -1 0 16512 0 -1 21924
box -48 -56 816 834
use sg13g2_xor2_1  _1774_
timestamp 1746816402
transform -1 0 23232 0 1 11340
box -48 -56 816 834
use sg13g2_a21oi_1  _1775_
timestamp 1746816402
transform 1 0 18528 0 1 11340
box -48 -56 528 834
use sg13g2_a21oi_1  _1776_
timestamp 1746816402
transform 1 0 27744 0 1 9828
box -48 -56 528 834
use sg13g2_xnor2_1  _1777_
timestamp 1746816402
transform -1 0 28512 0 1 11340
box -48 -56 816 834
use sg13g2_xnor2_1  _1778_
timestamp 1746816402
transform -1 0 27840 0 -1 11340
box -48 -56 816 834
use sg13g2_a21oi_1  _1779_
timestamp 1746816402
transform 1 0 24096 0 -1 11340
box -48 -56 528 834
use sg13g2_o21ai_1  _1780_
timestamp 1746816402
transform 1 0 23616 0 -1 11340
box -48 -56 538 834
use sg13g2_xor2_1  _1781_
timestamp 1746816402
transform -1 0 26976 0 1 11340
box -48 -56 816 834
use sg13g2_xnor2_1  _1782_
timestamp 1746816402
transform 1 0 26016 0 -1 11340
box -48 -56 816 834
use sg13g2_xnor2_1  _1783_
timestamp 1746816402
transform -1 0 27744 0 1 11340
box -48 -56 816 834
use sg13g2_a21oi_1  _1784_
timestamp 1746816402
transform 1 0 18528 0 -1 12852
box -48 -56 528 834
use sg13g2_o21ai_1  _1785_
timestamp 1746816402
transform 1 0 17856 0 -1 12852
box -48 -56 538 834
use sg13g2_and2_1  _1786_
timestamp 1746816402
transform -1 0 17664 0 1 15876
box -48 -56 528 834
use sg13g2_a221oi_1  _1787_
timestamp 1746816402
transform -1 0 17280 0 -1 17388
box -48 -56 816 834
use sg13g2_nor2b_1  _1788_
timestamp 1746816402
transform 1 0 16416 0 1 17388
box -54 -56 528 834
use sg13g2_a221oi_1  _1789_
timestamp 1746816402
transform 1 0 16896 0 1 17388
box -48 -56 816 834
use sg13g2_o21ai_1  _1790_
timestamp 1746816402
transform 1 0 18720 0 1 17388
box -48 -56 538 834
use sg13g2_a21oi_1  _1791_
timestamp 1746816402
transform -1 0 17472 0 -1 20412
box -48 -56 528 834
use sg13g2_a21oi_1  _1792_
timestamp 1746816402
transform -1 0 19008 0 -1 20412
box -48 -56 528 834
use sg13g2_o21ai_1  _1793_
timestamp 1746816402
transform 1 0 19104 0 1 20412
box -48 -56 538 834
use sg13g2_a21oi_2  _1794_
timestamp 1746816402
transform -1 0 19872 0 1 21924
box -48 -56 816 834
use sg13g2_a21o_1  _1795_
timestamp 1746816402
transform 1 0 6624 0 1 26460
box -48 -56 720 834
use sg13g2_nor3_1  _1796_
timestamp 1746816402
transform 1 0 26784 0 -1 18900
box -48 -56 528 834
use sg13g2_a21o_1  _1797_
timestamp 1746816402
transform -1 0 26784 0 -1 17388
box -48 -56 720 834
use sg13g2_nand2b_1  _1798_
timestamp 1746816402
transform -1 0 26304 0 -1 15876
box -48 -56 528 834
use sg13g2_nor4_1  _1799_
timestamp 1746816402
transform 1 0 24768 0 1 14364
box -48 -56 624 834
use sg13g2_nand3_1  _1800_
timestamp 1746816402
transform 1 0 25632 0 -1 17388
box -48 -56 528 834
use sg13g2_o21ai_1  _1801_
timestamp 1746816402
transform 1 0 26016 0 1 15876
box -48 -56 538 834
use sg13g2_nand3_1  _1802_
timestamp 1746816402
transform -1 0 27936 0 -1 17388
box -48 -56 528 834
use sg13g2_and3_2  _1803_
timestamp 1746816402
transform -1 0 27456 0 -1 17388
box -48 -56 720 834
use sg13g2_nor2_2  _1804_
timestamp 1746816402
transform 1 0 27456 0 1 18900
box -48 -56 624 834
use sg13g2_nand2_2  _1805_
timestamp 1746816402
transform -1 0 27168 0 1 15876
box -48 -56 624 834
use sg13g2_and2_1  _1806_
timestamp 1746816402
transform 1 0 29664 0 -1 17388
box -48 -56 528 834
use sg13g2_nor3_1  _1807_
timestamp 1746816402
transform -1 0 20448 0 1 17388
box -48 -56 528 834
use sg13g2_xnor2_1  _1808_
timestamp 1746816402
transform -1 0 24000 0 1 12852
box -48 -56 816 834
use sg13g2_nor2_1  _1809_
timestamp 1746816402
transform 1 0 23232 0 1 11340
box -48 -56 432 834
use sg13g2_nor2_1  _1810_
timestamp 1746816402
transform 1 0 21312 0 -1 15876
box -48 -56 432 834
use sg13g2_xnor2_1  _1811_
timestamp 1746816402
transform 1 0 21696 0 -1 15876
box -48 -56 816 834
use sg13g2_nor2_1  _1812_
timestamp 1746816402
transform -1 0 23232 0 1 15876
box -48 -56 432 834
use sg13g2_xor2_1  _1813_
timestamp 1746816402
transform 1 0 23328 0 -1 14364
box -48 -56 816 834
use sg13g2_nor2_1  _1814_
timestamp 1746816402
transform -1 0 26304 0 -1 12852
box -48 -56 432 834
use sg13g2_and3_1  _1815_
timestamp 1746816402
transform 1 0 23232 0 1 14364
box -48 -56 720 834
use sg13g2_a21oi_1  _1816_
timestamp 1746816402
transform -1 0 25728 0 1 12852
box -48 -56 528 834
use sg13g2_nor3_1  _1817_
timestamp 1746816402
transform -1 0 26208 0 1 12852
box -48 -56 528 834
use sg13g2_o21ai_1  _1818_
timestamp 1746816402
transform 1 0 26592 0 1 14364
box -48 -56 538 834
use sg13g2_a21oi_1  _1819_
timestamp 1746816402
transform 1 0 27072 0 1 14364
box -48 -56 528 834
use sg13g2_nor2b_1  _1820_
timestamp 1746816402
transform 1 0 27552 0 -1 14364
box -54 -56 528 834
use sg13g2_xnor2_1  _1821_
timestamp 1746816402
transform 1 0 26784 0 -1 14364
box -48 -56 816 834
use sg13g2_nor2_1  _1822_
timestamp 1746816402
transform -1 0 30240 0 -1 14364
box -48 -56 432 834
use sg13g2_nand3_1  _1823_
timestamp 1746816402
transform -1 0 24768 0 1 17388
box -48 -56 528 834
use sg13g2_nand3_1  _1824_
timestamp 1746816402
transform 1 0 26688 0 -1 15876
box -48 -56 528 834
use sg13g2_xor2_1  _1825_
timestamp 1746816402
transform -1 0 28032 0 -1 15876
box -48 -56 816 834
use sg13g2_nor2_1  _1826_
timestamp 1746816402
transform -1 0 27744 0 1 15876
box -48 -56 432 834
use sg13g2_nor2_1  _1827_
timestamp 1746816402
transform -1 0 27936 0 1 14364
box -48 -56 432 834
use sg13g2_xnor2_1  _1828_
timestamp 1746816402
transform -1 0 30528 0 -1 15876
box -48 -56 816 834
use sg13g2_nor2_1  _1829_
timestamp 1746816402
transform 1 0 29472 0 -1 14364
box -48 -56 432 834
use sg13g2_nand2_1  _1830_
timestamp 1746816402
transform 1 0 29664 0 1 11340
box -48 -56 432 834
use sg13g2_nor2_1  _1831_
timestamp 1746816402
transform 1 0 28896 0 1 11340
box -48 -56 432 834
use sg13g2_nor3_1  _1832_
timestamp 1746816402
transform 1 0 26016 0 1 20412
box -48 -56 528 834
use sg13g2_a21o_1  _1833_
timestamp 1746816402
transform 1 0 26688 0 -1 21924
box -48 -56 720 834
use sg13g2_nor3_1  _1834_
timestamp 1746816402
transform 1 0 25056 0 -1 21924
box -48 -56 528 834
use sg13g2_and2_1  _1835_
timestamp 1746816402
transform 1 0 30624 0 1 24948
box -48 -56 528 834
use sg13g2_nand3_1  _1836_
timestamp 1746816402
transform -1 0 26208 0 1 23436
box -48 -56 528 834
use sg13g2_o21ai_1  _1837_
timestamp 1746816402
transform 1 0 25344 0 1 21924
box -48 -56 538 834
use sg13g2_nand3_1  _1838_
timestamp 1746816402
transform 1 0 26304 0 1 21924
box -48 -56 528 834
use sg13g2_nor2_2  _1839_
timestamp 1746816402
transform -1 0 26592 0 -1 18900
box -48 -56 624 834
use sg13g2_and4_2  _1840_
timestamp 1746816402
transform -1 0 26688 0 -1 21924
box -48 -56 912 834
use sg13g2_o21ai_1  _1841_
timestamp 1746816402
transform 1 0 2496 0 1 24948
box -48 -56 538 834
use sg13g2_a21oi_1  _1842_
timestamp 1746816402
transform 1 0 3840 0 -1 23436
box -48 -56 528 834
use sg13g2_a21oi_1  _1843_
timestamp 1746816402
transform -1 0 3360 0 1 18900
box -48 -56 528 834
use sg13g2_and3_2  _1844_
timestamp 1746816402
transform 1 0 3168 0 1 17388
box -48 -56 720 834
use sg13g2_nor3_1  _1845_
timestamp 1746816402
transform 1 0 2208 0 1 17388
box -48 -56 528 834
use sg13g2_nor2_1  _1846_
timestamp 1746816402
transform 1 0 2592 0 -1 8316
box -48 -56 432 834
use sg13g2_and2_1  _1847_
timestamp 1746816402
transform 1 0 2976 0 -1 8316
box -48 -56 528 834
use sg13g2_nor3_1  _1848_
timestamp 1746816402
transform -1 0 4032 0 -1 9828
box -48 -56 528 834
use sg13g2_nor2b_1  _1849_
timestamp 1746816402
transform -1 0 3072 0 -1 9828
box -54 -56 528 834
use sg13g2_o21ai_1  _1850_
timestamp 1746816402
transform -1 0 2688 0 -1 6804
box -48 -56 538 834
use sg13g2_a21oi_1  _1851_
timestamp 1746816402
transform 1 0 2400 0 1 5292
box -48 -56 528 834
use sg13g2_a21oi_1  _1852_
timestamp 1746816402
transform -1 0 4320 0 1 5292
box -48 -56 528 834
use sg13g2_and3_1  _1853_
timestamp 1746816402
transform 1 0 4320 0 1 5292
box -48 -56 720 834
use sg13g2_nor3_1  _1854_
timestamp 1746816402
transform -1 0 6816 0 -1 6804
box -48 -56 528 834
use sg13g2_and3_1  _1855_
timestamp 1746816402
transform 1 0 5856 0 1 5292
box -48 -56 720 834
use sg13g2_o21ai_1  _1856_
timestamp 1746816402
transform -1 0 8448 0 1 3780
box -48 -56 538 834
use sg13g2_a21oi_1  _1857_
timestamp 1746816402
transform -1 0 7968 0 1 3780
box -48 -56 528 834
use sg13g2_and2_1  _1858_
timestamp 1746816402
transform 1 0 8448 0 1 5292
box -48 -56 528 834
use sg13g2_nor2_1  _1859_
timestamp 1746816402
transform -1 0 13536 0 1 3780
box -48 -56 432 834
use sg13g2_and2_1  _1860_
timestamp 1746816402
transform -1 0 14016 0 1 5292
box -48 -56 528 834
use sg13g2_nor3_1  _1861_
timestamp 1746816402
transform 1 0 12672 0 -1 5292
box -48 -56 528 834
use sg13g2_and2_1  _1862_
timestamp 1746816402
transform 1 0 13920 0 1 3780
box -48 -56 528 834
use sg13g2_o21ai_1  _1863_
timestamp 1746816402
transform -1 0 16512 0 1 5292
box -48 -56 538 834
use sg13g2_a21oi_1  _1864_
timestamp 1746816402
transform -1 0 16224 0 1 3780
box -48 -56 528 834
use sg13g2_nand2_1  _1865_
timestamp 1746816402
transform 1 0 20832 0 -1 5292
box -48 -56 432 834
use sg13g2_a21oi_1  _1866_
timestamp 1746816402
transform -1 0 22080 0 -1 5292
box -48 -56 528 834
use sg13g2_nor2_1  _1867_
timestamp 1746816402
transform 1 0 24192 0 -1 6804
box -48 -56 432 834
use sg13g2_nor3_1  _1868_
timestamp 1746816402
transform 1 0 21120 0 -1 6804
box -48 -56 528 834
use sg13g2_nor2_1  _1869_
timestamp 1746816402
transform -1 0 22464 0 -1 5292
box -48 -56 432 834
use sg13g2_o21ai_1  _1870_
timestamp 1746816402
transform -1 0 22080 0 1 6804
box -48 -56 538 834
use sg13g2_a21oi_1  _1871_
timestamp 1746816402
transform -1 0 21024 0 1 8316
box -48 -56 528 834
use sg13g2_nand2_1  _1872_
timestamp 1746816402
transform 1 0 25152 0 1 6804
box -48 -56 432 834
use sg13g2_o21ai_1  _1873_
timestamp 1746816402
transform 1 0 26112 0 1 6804
box -48 -56 538 834
use sg13g2_a21oi_1  _1874_
timestamp 1746816402
transform 1 0 26880 0 1 8316
box -48 -56 528 834
use sg13g2_nor2_1  _1875_
timestamp 1746816402
transform 1 0 26496 0 -1 9828
box -48 -56 432 834
use sg13g2_o21ai_1  _1876_
timestamp 1746816402
transform -1 0 27360 0 -1 9828
box -48 -56 538 834
use sg13g2_a21oi_1  _1877_
timestamp 1746816402
transform -1 0 27648 0 1 6804
box -48 -56 528 834
use sg13g2_xor2_1  _1878_
timestamp 1746816402
transform 1 0 13056 0 1 23436
box -48 -56 816 834
use sg13g2_xor2_1  _1879_
timestamp 1746816402
transform 1 0 5472 0 1 23436
box -48 -56 816 834
use sg13g2_xor2_1  _1880_
timestamp 1746816402
transform 1 0 6432 0 1 24948
box -48 -56 816 834
use sg13g2_nor3_1  _1881_
timestamp 1746816402
transform -1 0 11808 0 1 24948
box -48 -56 528 834
use sg13g2_nor3_1  _1882_
timestamp 1746816402
transform -1 0 13056 0 1 23436
box -48 -56 528 834
use sg13g2_nor2_1  _1883_
timestamp 1746816402
transform 1 0 10560 0 1 23436
box -48 -56 432 834
use sg13g2_nand2_2  _1884_
timestamp 1746816402
transform -1 0 17568 0 1 20412
box -48 -56 624 834
use sg13g2_and2_1  _1885_
timestamp 1746816402
transform 1 0 10272 0 1 26460
box -48 -56 528 834
use sg13g2_a221oi_1  _1886_
timestamp 1746816402
transform -1 0 13344 0 -1 26460
box -48 -56 816 834
use sg13g2_a21oi_1  _1887_
timestamp 1746816402
transform -1 0 12672 0 1 26460
box -48 -56 528 834
use sg13g2_and2_1  _1888_
timestamp 1746816402
transform 1 0 10752 0 1 26460
box -48 -56 528 834
use sg13g2_a221oi_1  _1889_
timestamp 1746816402
transform -1 0 12576 0 1 24948
box -48 -56 816 834
use sg13g2_a21oi_1  _1890_
timestamp 1746816402
transform 1 0 17472 0 -1 27972
box -48 -56 528 834
use sg13g2_nand3_1  _1891_
timestamp 1746816402
transform 1 0 11712 0 1 26460
box -48 -56 528 834
use sg13g2_a21oi_1  _1892_
timestamp 1746816402
transform -1 0 13824 0 -1 26460
box -48 -56 528 834
use sg13g2_a22oi_1  _1893_
timestamp 1746816402
transform -1 0 15072 0 1 24948
box -48 -56 624 834
use sg13g2_and2_1  _1894_
timestamp 1746816402
transform 1 0 11232 0 1 26460
box -48 -56 528 834
use sg13g2_a221oi_1  _1895_
timestamp 1746816402
transform 1 0 13152 0 -1 24948
box -48 -56 816 834
use sg13g2_a21oi_1  _1896_
timestamp 1746816402
transform 1 0 21024 0 1 24948
box -48 -56 528 834
use sg13g2_nand2_1  _1897_
timestamp 1746816402
transform 1 0 15936 0 1 24948
box -48 -56 432 834
use sg13g2_nand3_1  _1898_
timestamp 1746816402
transform 1 0 12672 0 1 24948
box -48 -56 528 834
use sg13g2_nand3_1  _1899_
timestamp 1746816402
transform 1 0 14592 0 -1 24948
box -48 -56 528 834
use sg13g2_a21oi_1  _1900_
timestamp 1746816402
transform 1 0 8352 0 1 26460
box -48 -56 528 834
use sg13g2_a21oi_1  _1901_
timestamp 1746816402
transform 1 0 9792 0 1 26460
box -48 -56 528 834
use sg13g2_mux2_1  _1902_
timestamp 1746816402
transform -1 0 20064 0 1 26460
box -48 -56 1008 834
use sg13g2_and2_1  _1903_
timestamp 1746816402
transform -1 0 13152 0 1 26460
box -48 -56 528 834
use sg13g2_a22oi_1  _1904_
timestamp 1746816402
transform 1 0 13152 0 1 26460
box -48 -56 624 834
use sg13g2_nand2_1  _1905_
timestamp 1746816402
transform 1 0 14784 0 -1 23436
box -48 -56 432 834
use sg13g2_o21ai_1  _1906_
timestamp 1746816402
transform 1 0 22752 0 -1 24948
box -48 -56 538 834
use sg13g2_and2_1  _1907_
timestamp 1746816402
transform -1 0 20544 0 1 26460
box -48 -56 528 834
use sg13g2_a22oi_1  _1908_
timestamp 1746816402
transform 1 0 17856 0 -1 26460
box -48 -56 624 834
use sg13g2_nand2_1  _1909_
timestamp 1746816402
transform 1 0 18432 0 1 14364
box -48 -56 432 834
use sg13g2_o21ai_1  _1910_
timestamp 1746816402
transform 1 0 21504 0 1 26460
box -48 -56 538 834
use sg13g2_nand3b_1  _1911_
timestamp 1746816402
transform 1 0 23424 0 -1 18900
box -48 -56 720 834
use sg13g2_nor3_1  _1912_
timestamp 1746816402
transform -1 0 25152 0 -1 18900
box -48 -56 528 834
use sg13g2_nand2b_1  _1913_
timestamp 1746816402
transform -1 0 25248 0 1 17388
box -48 -56 528 834
use sg13g2_nor4_1  _1914_
timestamp 1746816402
transform -1 0 24672 0 -1 18900
box -48 -56 624 834
use sg13g2_nor4_1  _1915_
timestamp 1746816402
transform -1 0 24384 0 1 18900
box -48 -56 624 834
use sg13g2_nor2_2  _1916_
timestamp 1746816402
transform -1 0 23808 0 -1 21924
box -48 -56 624 834
use sg13g2_nand4_1  _1917_
timestamp 1746816402
transform 1 0 23328 0 1 17388
box -48 -56 624 834
use sg13g2_nor4_1  _1918_
timestamp 1746816402
transform 1 0 22656 0 -1 18900
box -48 -56 624 834
use sg13g2_nor2b_1  _1919_
timestamp 1746816402
transform 1 0 22560 0 1 18900
box -54 -56 528 834
use sg13g2_or4_1  _1920_
timestamp 1746816402
transform -1 0 23328 0 1 17388
box -48 -56 816 834
use sg13g2_a21oi_1  _1921_
timestamp 1746816402
transform -1 0 22560 0 1 18900
box -48 -56 528 834
use sg13g2_nor3_1  _1922_
timestamp 1746816402
transform -1 0 23520 0 1 18900
box -48 -56 528 834
use sg13g2_mux2_1  _1923_
timestamp 1746816402
transform -1 0 24000 0 -1 20412
box -48 -56 1008 834
use sg13g2_nor2b_2  _1924_
timestamp 1746816402
transform 1 0 26208 0 1 18900
box -54 -56 720 834
use sg13g2_and2_1  _1925_
timestamp 1746816402
transform 1 0 30720 0 1 26460
box -48 -56 528 834
use sg13g2_o21ai_1  _1926_
timestamp 1746816402
transform -1 0 24000 0 1 23436
box -48 -56 538 834
use sg13g2_nor2_1  _1927_
timestamp 1746816402
transform 1 0 13728 0 -1 23436
box -48 -56 432 834
use sg13g2_o21ai_1  _1928_
timestamp 1746816402
transform -1 0 26304 0 -1 20412
box -48 -56 538 834
use sg13g2_nand2_1  _1929_
timestamp 1746816402
transform -1 0 29952 0 -1 11340
box -48 -56 432 834
use sg13g2_nor2b_1  _1930_
timestamp 1746816402
transform -1 0 30720 0 -1 18900
box -54 -56 528 834
use sg13g2_nand2b_1  _1931_
timestamp 1746816402
transform 1 0 27072 0 1 20412
box -48 -56 528 834
use sg13g2_xor2_1  _1932_
timestamp 1746816402
transform 1 0 27264 0 -1 26460
box -48 -56 816 834
use sg13g2_nor2_1  _1933_
timestamp 1746816402
transform -1 0 30336 0 -1 11340
box -48 -56 432 834
use sg13g2_nor2b_1  _1934_
timestamp 1746816402
transform 1 0 26880 0 1 23436
box -54 -56 528 834
use sg13g2_nand2_2  _1935_
timestamp 1746816402
transform -1 0 28128 0 1 20412
box -48 -56 624 834
use sg13g2_nor2_1  _1936_
timestamp 1746816402
transform -1 0 29664 0 1 11340
box -48 -56 432 834
use sg13g2_a21oi_1  _1937_
timestamp 1746816402
transform -1 0 26880 0 1 23436
box -48 -56 528 834
use sg13g2_a21oi_1  _1938_
timestamp 1746816402
transform -1 0 27936 0 1 24948
box -48 -56 528 834
use sg13g2_nor2_1  _1939_
timestamp 1746816402
transform 1 0 29184 0 -1 11340
box -48 -56 432 834
use sg13g2_a21oi_1  _1940_
timestamp 1746816402
transform -1 0 24480 0 1 23436
box -48 -56 528 834
use sg13g2_nand2_1  _1941_
timestamp 1746816402
transform 1 0 30336 0 1 12852
box -48 -56 432 834
use sg13g2_and3_1  _1942_
timestamp 1746816402
transform -1 0 28032 0 1 23436
box -48 -56 720 834
use sg13g2_nor3_1  _1943_
timestamp 1746816402
transform -1 0 30240 0 -1 18900
box -48 -56 528 834
use sg13g2_nand2_1  _1944_
timestamp 1746816402
transform -1 0 30912 0 1 11340
box -48 -56 432 834
use sg13g2_xnor2_1  _1945_
timestamp 1746816402
transform -1 0 28320 0 1 21924
box -48 -56 816 834
use sg13g2_o21ai_1  _1946_
timestamp 1746816402
transform 1 0 27168 0 -1 23436
box -48 -56 538 834
use sg13g2_a21oi_1  _1947_
timestamp 1746816402
transform -1 0 27072 0 1 20412
box -48 -56 528 834
use sg13g2_nor2_1  _1948_
timestamp 1746816402
transform -1 0 28896 0 1 11340
box -48 -56 432 834
use sg13g2_and2_1  _1949_
timestamp 1746816402
transform -1 0 31104 0 1 20412
box -48 -56 528 834
use sg13g2_nor3_1  _1950_
timestamp 1746816402
transform 1 0 27072 0 -1 24948
box -48 -56 528 834
use sg13g2_xnor2_1  _1951_
timestamp 1746816402
transform 1 0 28128 0 1 20412
box -48 -56 816 834
use sg13g2_nor2_1  _1952_
timestamp 1746816402
transform -1 0 30336 0 -1 12852
box -48 -56 432 834
use sg13g2_nand2_1  _1953_
timestamp 1746816402
transform -1 0 31008 0 1 15876
box -48 -56 432 834
use sg13g2_nor2b_1  _1954_
timestamp 1746816402
transform 1 0 27552 0 -1 20412
box -54 -56 528 834
use sg13g2_a21oi_1  _1955_
timestamp 1746816402
transform 1 0 27936 0 -1 21924
box -48 -56 528 834
use sg13g2_a21oi_1  _1956_
timestamp 1746816402
transform 1 0 27552 0 -1 24948
box -48 -56 528 834
use sg13g2_nor2_1  _1957_
timestamp 1746816402
transform 1 0 24576 0 1 18900
box -48 -56 432 834
use sg13g2_nand2_1  _1958_
timestamp 1746816402
transform -1 0 31392 0 1 15876
box -48 -56 432 834
use sg13g2_xnor2_1  _1959_
timestamp 1746816402
transform 1 0 26784 0 -1 20412
box -48 -56 816 834
use sg13g2_o21ai_1  _1960_
timestamp 1746816402
transform -1 0 27456 0 1 18900
box -48 -56 538 834
use sg13g2_nand3_1  _1961_
timestamp 1746816402
transform -1 0 26304 0 1 21924
box -48 -56 528 834
use sg13g2_nand2b_1  _1962_
timestamp 1746816402
transform -1 0 30720 0 -1 27972
box -48 -56 528 834
use sg13g2_nand4_1  _1963_
timestamp 1746816402
transform 1 0 24000 0 -1 24948
box -48 -56 624 834
use sg13g2_o21ai_1  _1964_
timestamp 1746816402
transform 1 0 24864 0 -1 24948
box -48 -56 538 834
use sg13g2_nand2b_1  _1965_
timestamp 1746816402
transform 1 0 26688 0 -1 26460
box -48 -56 528 834
use sg13g2_nor3_1  _1966_
timestamp 1746816402
transform 1 0 24480 0 -1 26460
box -48 -56 528 834
use sg13g2_a21oi_1  _1967_
timestamp 1746816402
transform 1 0 26304 0 -1 24948
box -48 -56 528 834
use sg13g2_nor3_1  _1968_
timestamp 1746816402
transform 1 0 26016 0 1 24948
box -48 -56 528 834
use sg13g2_a21oi_1  _1969_
timestamp 1746816402
transform -1 0 26976 0 1 24948
box -48 -56 528 834
use sg13g2_a22oi_1  _1970_
timestamp 1746816402
transform 1 0 24960 0 1 24948
box -48 -56 624 834
use sg13g2_nand2b_1  _1971_
timestamp 1746816402
transform -1 0 24960 0 1 23436
box -48 -56 528 834
use sg13g2_nand2_1  _1972_
timestamp 1746816402
transform 1 0 26112 0 -1 9828
box -48 -56 432 834
use sg13g2_o21ai_1  _1973_
timestamp 1746816402
transform 1 0 26976 0 1 24948
box -48 -56 538 834
use sg13g2_nor2_1  _1974_
timestamp 1746816402
transform 1 0 2400 0 1 26460
box -48 -56 432 834
use sg13g2_nor2_1  _1975_
timestamp 1746816402
transform 1 0 9504 0 1 20412
box -48 -56 432 834
use sg13g2_a21oi_1  _1976_
timestamp 1746816402
transform 1 0 9888 0 1 20412
box -48 -56 528 834
use sg13g2_o21ai_1  _1977_
timestamp 1746816402
transform -1 0 9600 0 -1 24948
box -48 -56 538 834
use sg13g2_nand2_1  _1978_
timestamp 1746816402
transform -1 0 11904 0 1 21924
box -48 -56 432 834
use sg13g2_o21ai_1  _1979_
timestamp 1746816402
transform 1 0 10080 0 1 23436
box -48 -56 538 834
use sg13g2_mux2_1  _1980_
timestamp 1746816402
transform 1 0 4128 0 -1 26460
box -48 -56 1008 834
use sg13g2_mux2_1  _1981_
timestamp 1746816402
transform -1 0 6432 0 1 24948
box -48 -56 1008 834
use sg13g2_mux2_1  _1982_
timestamp 1746816402
transform -1 0 5472 0 1 23436
box -48 -56 1008 834
use sg13g2_mux2_1  _1983_
timestamp 1746816402
transform 1 0 13824 0 1 23436
box -48 -56 1008 834
use sg13g2_a21o_1  _1984_
timestamp 1746816402
transform 1 0 21888 0 1 21924
box -48 -56 720 834
use sg13g2_dfrbp_1  _1985_
timestamp 1746816402
transform 1 0 9504 0 -1 27972
box -60 -56 2556 834
use sg13g2_tiehi  _1985__27
timestamp 1746816402
transform 1 0 5280 0 -1 24948
box -48 -56 432 834
use sg13g2_dfrbp_1  _1986_
timestamp 1746816402
transform 1 0 7008 0 -1 27972
box -60 -56 2556 834
use sg13g2_tiehi  _1986__18
timestamp 1746816402
transform 1 0 2112 0 1 24948
box -48 -56 432 834
use sg13g2_tiehi  _1987__59
timestamp 1746816402
transform 1 0 3264 0 -1 27972
box -48 -56 432 834
use sg13g2_dfrbp_1  _1987_
timestamp 1746816402
transform 1 0 8928 0 -1 26460
box -60 -56 2556 834
use sg13g2_dfrbp_1  _1988_
timestamp 1746816402
transform 1 0 4512 0 -1 27972
box -60 -56 2556 834
use sg13g2_tiehi  _1988__58
timestamp 1746816402
transform 1 0 960 0 -1 27972
box -48 -56 432 834
use sg13g2_dfrbp_1  _1989_
timestamp 1746816402
transform -1 0 14592 0 -1 27972
box -60 -56 2556 834
use sg13g2_tiehi  _1989__57
timestamp 1746816402
transform -1 0 14496 0 1 24948
box -48 -56 432 834
use sg13g2_dfrbp_1  _1990_
timestamp 1746816402
transform -1 0 30144 0 1 17388
box -60 -56 2556 834
use sg13g2_tiehi  _1990__56
timestamp 1746816402
transform -1 0 31296 0 -1 17388
box -48 -56 432 834
use sg13g2_tiehi  _1991__55
timestamp 1746816402
transform -1 0 21792 0 -1 17388
box -48 -56 432 834
use sg13g2_dfrbp_1  _1991_
timestamp 1746816402
transform 1 0 19872 0 1 15876
box -60 -56 2556 834
use sg13g2_dfrbp_1  _1992_
timestamp 1746816402
transform -1 0 22656 0 -1 12852
box -60 -56 2556 834
use sg13g2_tiehi  _1992__54
timestamp 1746816402
transform -1 0 22272 0 1 11340
box -48 -56 432 834
use sg13g2_dfrbp_1  _1993_
timestamp 1746816402
transform 1 0 22464 0 -1 15876
box -60 -56 2556 834
use sg13g2_tiehi  _1993__53
timestamp 1746816402
transform -1 0 24384 0 1 12852
box -48 -56 432 834
use sg13g2_tiehi  _1994__52
timestamp 1746816402
transform -1 0 29568 0 -1 12852
box -48 -56 432 834
use sg13g2_dfrbp_1  _1994_
timestamp 1746816402
transform -1 0 25920 0 -1 12852
box -60 -56 2556 834
use sg13g2_tiehi  _1995__51
timestamp 1746816402
transform -1 0 26688 0 -1 15876
box -48 -56 432 834
use sg13g2_dfrbp_1  _1995_
timestamp 1746816402
transform -1 0 26688 0 -1 14364
box -60 -56 2556 834
use sg13g2_tiehi  _1996__50
timestamp 1746816402
transform -1 0 29184 0 -1 12852
box -48 -56 432 834
use sg13g2_dfrbp_1  _1996_
timestamp 1746816402
transform 1 0 26304 0 -1 12852
box -60 -56 2556 834
use sg13g2_tiehi  _1997__49
timestamp 1746816402
transform -1 0 30624 0 -1 14364
box -48 -56 432 834
use sg13g2_dfrbp_1  _1997_
timestamp 1746816402
transform -1 0 29856 0 1 12852
box -60 -56 2556 834
use sg13g2_tiehi  _1998__48
timestamp 1746816402
transform -1 0 30912 0 -1 17388
box -48 -56 432 834
use sg13g2_dfrbp_1  _1998_
timestamp 1746816402
transform -1 0 30240 0 1 15876
box -60 -56 2556 834
use sg13g2_tiehi  _1999__47
timestamp 1746816402
transform -1 0 30624 0 1 15876
box -48 -56 432 834
use sg13g2_dfrbp_1  _1999_
timestamp 1746816402
transform -1 0 30528 0 1 14364
box -60 -56 2556 834
use sg13g2_tiehi  _2000__46
timestamp 1746816402
transform 1 0 1248 0 -1 26460
box -48 -56 432 834
use sg13g2_dfrbp_1  _2000_
timestamp 1746816402
transform -1 0 3072 0 1 23436
box -60 -56 2556 834
use sg13g2_dfrbp_1  _2001_
timestamp 1746816402
transform -1 0 3168 0 -1 18900
box -60 -56 2556 834
use sg13g2_tiehi  _2001__44
timestamp 1746816402
transform 1 0 1728 0 1 17388
box -48 -56 432 834
use sg13g2_dfrbp_1  _2002_
timestamp 1746816402
transform -1 0 3072 0 1 8316
box -60 -56 2556 834
use sg13g2_tiehi  _2002__42
timestamp 1746816402
transform 1 0 1728 0 -1 8316
box -48 -56 432 834
use sg13g2_tiehi  _2003__40
timestamp 1746816402
transform -1 0 4512 0 1 6804
box -48 -56 432 834
use sg13g2_dfrbp_1  _2003_
timestamp 1746816402
transform 1 0 2688 0 -1 6804
box -60 -56 2556 834
use sg13g2_dfrbp_1  _2004_
timestamp 1746816402
transform 1 0 4992 0 -1 5292
box -60 -56 2556 834
use sg13g2_tiehi  _2004__38
timestamp 1746816402
transform -1 0 6528 0 1 3780
box -48 -56 432 834
use sg13g2_tiehi  _2005__36
timestamp 1746816402
transform -1 0 9312 0 1 5292
box -48 -56 432 834
use sg13g2_dfrbp_1  _2005_
timestamp 1746816402
transform 1 0 7968 0 -1 5292
box -60 -56 2556 834
use sg13g2_dfrbp_1  _2006_
timestamp 1746816402
transform 1 0 13152 0 -1 5292
box -60 -56 2556 834
use sg13g2_tiehi  _2006__34
timestamp 1746816402
transform -1 0 14784 0 1 3780
box -48 -56 432 834
use sg13g2_dfrbp_1  _2007_
timestamp 1746816402
transform 1 0 16032 0 -1 5292
box -60 -56 2556 834
use sg13g2_tiehi  _2007__32
timestamp 1746816402
transform -1 0 17472 0 1 3780
box -48 -56 432 834
use sg13g2_tiehi  _2008__30
timestamp 1746816402
transform -1 0 24096 0 1 5292
box -48 -56 432 834
use sg13g2_dfrbp_1  _2008_
timestamp 1746816402
transform 1 0 21216 0 1 5292
box -60 -56 2556 834
use sg13g2_dfrbp_1  _2009_
timestamp 1746816402
transform 1 0 21024 0 1 8316
box -60 -56 2556 834
use sg13g2_tiehi  _2009__28
timestamp 1746816402
transform -1 0 23808 0 1 6804
box -48 -56 432 834
use sg13g2_tiehi  _2010__26
timestamp 1746816402
transform -1 0 28608 0 -1 8316
box -48 -56 432 834
use sg13g2_dfrbp_1  _2010_
timestamp 1746816402
transform 1 0 25728 0 -1 8316
box -60 -56 2556 834
use sg13g2_tiehi  _2011__24
timestamp 1746816402
transform 1 0 28224 0 1 9828
box -48 -56 432 834
use sg13g2_dfrbp_1  _2011_
timestamp 1746816402
transform -1 0 29856 0 -1 9828
box -60 -56 2556 834
use sg13g2_tiehi  _2012__22
timestamp 1746816402
transform 1 0 14592 0 -1 27972
box -48 -56 432 834
use sg13g2_dfrbp_1  _2012_
timestamp 1746816402
transform 1 0 13824 0 -1 26460
box -60 -56 2556 834
use sg13g2_dfrbp_1  _2013_
timestamp 1746816402
transform 1 0 16608 0 1 26460
box -60 -56 2556 834
use sg13g2_tiehi  _2013__21
timestamp 1746816402
transform -1 0 19008 0 -1 23436
box -48 -56 432 834
use sg13g2_dfrbp_1  _2014_
timestamp 1746816402
transform 1 0 16320 0 1 24948
box -60 -56 2556 834
use sg13g2_tiehi  _2014__20
timestamp 1746816402
transform -1 0 17856 0 -1 26460
box -48 -56 432 834
use sg13g2_dfrbp_1  _2015_
timestamp 1746816402
transform 1 0 21504 0 1 24948
box -60 -56 2556 834
use sg13g2_tiehi  _2015__19
timestamp 1746816402
transform 1 0 17472 0 1 21924
box -48 -56 432 834
use sg13g2_tiehi  _2016__17
timestamp 1746816402
transform -1 0 17952 0 -1 24948
box -48 -56 432 834
use sg13g2_dfrbp_1  _2016_
timestamp 1746816402
transform 1 0 15072 0 -1 24948
box -60 -56 2556 834
use sg13g2_dfrbp_1  _2017_
timestamp 1746816402
transform 1 0 19104 0 -1 27972
box -60 -56 2556 834
use sg13g2_tiehi  _2017__73
timestamp 1746816402
transform 1 0 17760 0 -1 21924
box -48 -56 432 834
use sg13g2_dfrbp_1  _2018_
timestamp 1746816402
transform 1 0 21888 0 -1 27972
box -60 -56 2556 834
use sg13g2_tiehi  _2018__72
timestamp 1746816402
transform 1 0 15552 0 -1 23436
box -48 -56 432 834
use sg13g2_dfrbp_1  _2019_
timestamp 1746816402
transform 1 0 21984 0 -1 26460
box -60 -56 2556 834
use sg13g2_tiehi  _2019__71
timestamp 1746816402
transform 1 0 18048 0 1 14364
box -48 -56 432 834
use sg13g2_tiehi  _2020__70
timestamp 1746816402
transform 1 0 21600 0 1 20412
box -48 -56 432 834
use sg13g2_dfrbp_1  _2020_
timestamp 1746816402
transform -1 0 23040 0 -1 20412
box -60 -56 2556 834
use sg13g2_dfrbp_1  _2021_
timestamp 1746816402
transform 1 0 26880 0 -1 27972
box -60 -56 2556 834
use sg13g2_tiehi  _2021__69
timestamp 1746816402
transform -1 0 31296 0 1 14364
box -48 -56 432 834
use sg13g2_dfrbp_1  _2022_
timestamp 1746816402
transform -1 0 30720 0 1 26460
box -60 -56 2556 834
use sg13g2_tiehi  _2022__67
timestamp 1746816402
transform -1 0 31200 0 -1 12852
box -48 -56 432 834
use sg13g2_dfrbp_1  _2023_
timestamp 1746816402
transform 1 0 28896 0 -1 26460
box -60 -56 2556 834
use sg13g2_tiehi  _2023__65
timestamp 1746816402
transform -1 0 30720 0 1 9828
box -48 -56 432 834
use sg13g2_dfrbp_1  _2024_
timestamp 1746816402
transform 1 0 28896 0 -1 24948
box -60 -56 2556 834
use sg13g2_tiehi  _2024__63
timestamp 1746816402
transform -1 0 31104 0 1 9828
box -48 -56 432 834
use sg13g2_dfrbp_1  _2025_
timestamp 1746816402
transform 1 0 28896 0 1 23436
box -60 -56 2556 834
use sg13g2_tiehi  _2025__61
timestamp 1746816402
transform -1 0 31104 0 -1 11340
box -48 -56 432 834
use sg13g2_dfrbp_1  _2026_
timestamp 1746816402
transform -1 0 31392 0 1 21924
box -60 -56 2556 834
use sg13g2_tiehi  _2026__45
timestamp 1746816402
transform -1 0 30720 0 -1 11340
box -48 -56 432 834
use sg13g2_dfrbp_1  _2027_
timestamp 1746816402
transform 1 0 28896 0 -1 21924
box -60 -56 2556 834
use sg13g2_tiehi  _2027__41
timestamp 1746816402
transform -1 0 31296 0 1 11340
box -48 -56 432 834
use sg13g2_dfrbp_1  _2028_
timestamp 1746816402
transform -1 0 31392 0 -1 20412
box -60 -56 2556 834
use sg13g2_tiehi  _2028__37
timestamp 1746816402
transform -1 0 30816 0 -1 12852
box -48 -56 432 834
use sg13g2_dfrbp_1  _2029_
timestamp 1746816402
transform 1 0 28896 0 1 18900
box -60 -56 2556 834
use sg13g2_tiehi  _2029__33
timestamp 1746816402
transform -1 0 31104 0 1 12852
box -48 -56 432 834
use sg13g2_dfrbp_1  _2030_
timestamp 1746816402
transform -1 0 29760 0 -1 18900
box -60 -56 2556 834
use sg13g2_tiehi  _2030__29
timestamp 1746816402
transform -1 0 31392 0 -1 15876
box -48 -56 432 834
use sg13g2_dfrbp_1  _2031_
timestamp 1746816402
transform -1 0 26880 0 -1 27972
box -60 -56 2556 834
use sg13g2_tiehi  _2031__25
timestamp 1746816402
transform -1 0 29184 0 -1 11340
box -48 -56 432 834
use sg13g2_dfrbp_1  _2032_
timestamp 1746816402
transform 1 0 14976 0 -1 27972
box -60 -56 2556 834
use sg13g2_tiehi  _2032__23
timestamp 1746816402
transform 1 0 15360 0 1 26460
box -48 -56 432 834
use sg13g2_tiehi  _2033__68
timestamp 1746816402
transform 1 0 2496 0 -1 27972
box -48 -56 432 834
use sg13g2_dfrbp_1  _2033_
timestamp 1746816402
transform 1 0 6432 0 -1 26460
box -60 -56 2556 834
use sg13g2_tiehi  _2034__66
timestamp 1746816402
transform -1 0 12192 0 -1 20412
box -48 -56 432 834
use sg13g2_dfrbp_1  _2034_
timestamp 1746816402
transform 1 0 9312 0 -1 20412
box -60 -56 2556 834
use sg13g2_dfrbp_1  _2035_
timestamp 1746816402
transform -1 0 8544 0 -1 24948
box -60 -56 2556 834
use sg13g2_tiehi  _2035__64
timestamp 1746816402
transform 1 0 5664 0 -1 24948
box -48 -56 432 834
use sg13g2_tiehi  _2036__62
timestamp 1746816402
transform 1 0 8928 0 1 24948
box -48 -56 432 834
use sg13g2_dfrbp_1  _2036_
timestamp 1746816402
transform 1 0 9792 0 -1 24948
box -60 -56 2556 834
use sg13g2_dfrbp_1  _2037_
timestamp 1746816402
transform -1 0 5280 0 1 26460
box -60 -56 2556 834
use sg13g2_tiehi  _2037__60
timestamp 1746816402
transform 1 0 1632 0 -1 26460
box -48 -56 432 834
use sg13g2_dfrbp_1  _2038_
timestamp 1746816402
transform 1 0 2976 0 1 24948
box -60 -56 2556 834
use sg13g2_tiehi  _2038__43
timestamp 1746816402
transform 1 0 1344 0 1 24948
box -48 -56 432 834
use sg13g2_dfrbp_1  _2039_
timestamp 1746816402
transform 1 0 1824 0 -1 24948
box -60 -56 2556 834
use sg13g2_tiehi  _2039__39
timestamp 1746816402
transform 1 0 672 0 -1 24948
box -48 -56 432 834
use sg13g2_dfrbp_1  _2040_
timestamp 1746816402
transform 1 0 14880 0 1 23436
box -60 -56 2556 834
use sg13g2_tiehi  _2040__35
timestamp 1746816402
transform -1 0 16320 0 -1 23436
box -48 -56 432 834
use sg13g2_dfrbp_1  _2041_
timestamp 1746816402
transform 1 0 22080 0 -1 23436
box -60 -56 2556 834
use sg13g2_tiehi  _2041__31
timestamp 1746816402
transform 1 0 17376 0 -1 21924
box -48 -56 432 834
use sg13g2_buf_2  clkbuf_0_clk
timestamp 1746816402
transform 1 0 15936 0 1 17388
box -48 -56 528 834
use sg13g2_buf_2  clkbuf_4_0_0_clk
timestamp 1746816402
transform -1 0 7968 0 1 14364
box -48 -56 528 834
use sg13g2_buf_2  clkbuf_4_1_0_clk
timestamp 1746816402
transform -1 0 8832 0 1 17388
box -48 -56 528 834
use sg13g2_buf_2  clkbuf_4_2_0_clk
timestamp 1746816402
transform 1 0 14880 0 -1 17388
box -48 -56 528 834
use sg13g2_buf_2  clkbuf_4_3_0_clk
timestamp 1746816402
transform 1 0 16320 0 -1 18900
box -48 -56 528 834
use sg13g2_buf_2  clkbuf_4_4_0_clk
timestamp 1746816402
transform 1 0 5952 0 -1 26460
box -48 -56 528 834
use sg13g2_buf_2  clkbuf_4_5_0_clk
timestamp 1746816402
transform 1 0 7968 0 1 24948
box -48 -56 528 834
use sg13g2_buf_2  clkbuf_4_6_0_clk
timestamp 1746816402
transform -1 0 11424 0 1 23436
box -48 -56 528 834
use sg13g2_buf_2  clkbuf_4_7_0_clk
timestamp 1746816402
transform -1 0 14592 0 -1 24948
box -48 -56 528 834
use sg13g2_buf_2  clkbuf_4_8_0_clk
timestamp 1746816402
transform -1 0 23616 0 -1 11340
box -48 -56 528 834
use sg13g2_buf_2  clkbuf_4_9_0_clk
timestamp 1746816402
transform 1 0 26208 0 1 12852
box -48 -56 528 834
use sg13g2_buf_2  clkbuf_4_10_0_clk
timestamp 1746816402
transform -1 0 29472 0 -1 14364
box -48 -56 528 834
use sg13g2_buf_2  clkbuf_4_11_0_clk
timestamp 1746816402
transform -1 0 31008 0 -1 15876
box -48 -56 528 834
use sg13g2_buf_2  clkbuf_4_12_0_clk
timestamp 1746816402
transform 1 0 23040 0 1 23436
box -48 -56 528 834
use sg13g2_buf_2  clkbuf_4_13_0_clk
timestamp 1746816402
transform 1 0 27648 0 -1 23436
box -48 -56 528 834
use sg13g2_buf_2  clkbuf_4_14_0_clk
timestamp 1746816402
transform -1 0 28896 0 -1 21924
box -48 -56 528 834
use sg13g2_buf_2  clkbuf_4_15_0_clk
timestamp 1746816402
transform 1 0 28320 0 1 21924
box -48 -56 528 834
use sg13g2_inv_1  clkload0
timestamp 1746816402
transform -1 0 17952 0 -1 18900
box -48 -56 336 834
use sg13g2_inv_1  clkload1
timestamp 1746816402
transform 1 0 7200 0 1 24948
box -48 -56 336 834
use sg13g2_inv_1  clkload2
timestamp 1746816402
transform -1 0 12576 0 -1 26460
box -48 -56 336 834
use sg13g2_inv_1  clkload3
timestamp 1746816402
transform 1 0 26304 0 1 14364
box -48 -56 336 834
use sg13g2_inv_1  clkload4
timestamp 1746816402
transform 1 0 31104 0 1 12852
box -48 -56 336 834
use sg13g2_inv_1  clkload5
timestamp 1746816402
transform -1 0 27552 0 1 21924
box -48 -56 336 834
use sg13g2_inv_1  clkload6
timestamp 1746816402
transform 1 0 31104 0 1 20412
box -48 -56 336 834
use sg13g2_tielo  controller_11
timestamp 1746816402
transform 1 0 1632 0 1 26460
box -48 -56 432 834
use sg13g2_tielo  controller_12
timestamp 1746816402
transform 1 0 2400 0 -1 26460
box -48 -56 432 834
use sg13g2_tielo  controller_13
timestamp 1746816402
transform 1 0 1344 0 -1 27972
box -48 -56 432 834
use sg13g2_tielo  controller_14
timestamp 1746816402
transform 1 0 1440 0 -1 24948
box -48 -56 432 834
use sg13g2_tielo  controller_15
timestamp 1746816402
transform 1 0 576 0 -1 27972
box -48 -56 432 834
use sg13g2_tielo  controller_16
timestamp 1746816402
transform 1 0 1248 0 1 26460
box -48 -56 432 834
use sg13g2_tiehi  controller_74
timestamp 1746816402
transform 1 0 864 0 1 26460
box -48 -56 432 834
use sg13g2_tiehi  controller_75
timestamp 1746816402
transform 1 0 1344 0 1 18900
box -48 -56 432 834
use sg13g2_buf_2  fanout315
timestamp 1746816402
transform -1 0 14112 0 1 24948
box -48 -56 528 834
use sg13g2_buf_2  fanout316
timestamp 1746816402
transform -1 0 13632 0 1 24948
box -48 -56 528 834
use sg13g2_buf_4  fanout317
timestamp 1746816402
transform 1 0 20160 0 -1 11340
box -48 -56 816 834
use sg13g2_buf_2  fanout318
timestamp 1746816402
transform 1 0 19776 0 1 11340
box -48 -56 528 834
use sg13g2_buf_4  fanout319
timestamp 1746816402
transform 1 0 21888 0 1 9828
box -48 -56 816 834
use sg13g2_buf_4  fanout320
timestamp 1746816402
transform -1 0 23712 0 1 20412
box -48 -56 816 834
use sg13g2_buf_4  fanout321
timestamp 1746816402
transform 1 0 19392 0 -1 11340
box -48 -56 816 834
use sg13g2_buf_2  fanout322
timestamp 1746816402
transform -1 0 21504 0 1 11340
box -48 -56 528 834
use sg13g2_buf_2  fanout323
timestamp 1746816402
transform 1 0 11136 0 -1 17388
box -48 -56 528 834
use sg13g2_buf_1  fanout324
timestamp 1746816402
transform 1 0 9888 0 1 17388
box -48 -56 432 834
use sg13g2_buf_2  fanout325
timestamp 1746816402
transform -1 0 10752 0 1 8316
box -48 -56 528 834
use sg13g2_buf_2  fanout326
timestamp 1746816402
transform 1 0 19200 0 1 17388
box -48 -56 528 834
use sg13g2_buf_2  fanout327
timestamp 1746816402
transform 1 0 13248 0 -1 18900
box -48 -56 528 834
use sg13g2_buf_2  fanout328
timestamp 1746816402
transform 1 0 9312 0 -1 18900
box -48 -56 528 834
use sg13g2_buf_2  fanout329
timestamp 1746816402
transform 1 0 17952 0 -1 18900
box -48 -56 528 834
use sg13g2_buf_2  fanout330
timestamp 1746816402
transform 1 0 13536 0 1 18900
box -48 -56 528 834
use sg13g2_buf_2  fanout331
timestamp 1746816402
transform -1 0 9216 0 1 11340
box -48 -56 528 834
use sg13g2_buf_1  fanout332
timestamp 1746816402
transform -1 0 6528 0 -1 14364
box -48 -56 432 834
use sg13g2_buf_2  fanout333
timestamp 1746816402
transform 1 0 19776 0 -1 23436
box -48 -56 528 834
use sg13g2_buf_2  fanout334
timestamp 1746816402
transform 1 0 3552 0 1 21924
box -48 -56 528 834
use sg13g2_buf_1  fanout335
timestamp 1746816402
transform 1 0 576 0 1 24948
box -48 -56 432 834
use sg13g2_buf_2  fanout336
timestamp 1746816402
transform -1 0 12000 0 -1 21924
box -48 -56 528 834
use sg13g2_buf_4  fanout337
timestamp 1746816402
transform -1 0 13248 0 -1 21924
box -48 -56 816 834
use sg13g2_buf_2  fanout338
timestamp 1746816402
transform -1 0 12960 0 1 15876
box -48 -56 528 834
use sg13g2_buf_2  fanout339
timestamp 1746816402
transform -1 0 13440 0 -1 17388
box -48 -56 528 834
use sg13g2_buf_2  fanout340
timestamp 1746816402
transform -1 0 11040 0 1 9828
box -48 -56 528 834
use sg13g2_buf_2  fanout341
timestamp 1746816402
transform -1 0 14112 0 1 9828
box -48 -56 528 834
use sg13g2_buf_4  fanout342
timestamp 1746816402
transform 1 0 11712 0 1 12852
box -48 -56 816 834
use sg13g2_buf_2  fanout343
timestamp 1746816402
transform 1 0 19008 0 1 11340
box -48 -56 528 834
use sg13g2_buf_2  fanout344
timestamp 1746816402
transform -1 0 10848 0 1 11340
box -48 -56 528 834
use sg13g2_buf_4  fanout345
timestamp 1746816402
transform 1 0 16224 0 1 20412
box -48 -56 816 834
use sg13g2_buf_2  fanout346
timestamp 1746816402
transform 1 0 16512 0 -1 12852
box -48 -56 528 834
use sg13g2_buf_2  fanout347
timestamp 1746816402
transform 1 0 10272 0 1 17388
box -48 -56 528 834
use sg13g2_buf_1  fanout348
timestamp 1746816402
transform -1 0 10560 0 1 18900
box -48 -56 432 834
use sg13g2_buf_2  fanout349
timestamp 1746816402
transform 1 0 11424 0 -1 18900
box -48 -56 528 834
use sg13g2_buf_2  fanout350
timestamp 1746816402
transform 1 0 16608 0 1 18900
box -48 -56 528 834
use sg13g2_buf_2  fanout351
timestamp 1746816402
transform -1 0 13056 0 -1 12852
box -48 -56 528 834
use sg13g2_buf_2  fanout352
timestamp 1746816402
transform -1 0 13056 0 -1 18900
box -48 -56 528 834
use sg13g2_buf_2  fanout353
timestamp 1746816402
transform 1 0 1152 0 1 12852
box -48 -56 528 834
use sg13g2_buf_2  fanout354
timestamp 1746816402
transform 1 0 9984 0 -1 18900
box -48 -56 528 834
use sg13g2_buf_2  fanout355
timestamp 1746816402
transform 1 0 10656 0 1 20412
box -48 -56 528 834
use sg13g2_buf_2  fanout356
timestamp 1746816402
transform 1 0 2688 0 1 20412
box -48 -56 528 834
use sg13g2_buf_1  fanout357
timestamp 1746816402
transform -1 0 7200 0 1 20412
box -48 -56 432 834
use sg13g2_buf_1  fanout358
timestamp 1746816402
transform -1 0 13344 0 -1 23436
box -48 -56 432 834
use sg13g2_buf_2  fanout359
timestamp 1746816402
transform -1 0 19968 0 -1 20412
box -48 -56 528 834
use sg13g2_buf_2  fanout360
timestamp 1746816402
transform -1 0 4416 0 -1 21924
box -48 -56 528 834
use sg13g2_buf_1  fanout361
timestamp 1746816402
transform 1 0 4896 0 -1 21924
box -48 -56 432 834
use sg13g2_buf_1  fanout362
timestamp 1746816402
transform -1 0 9408 0 1 20412
box -48 -56 432 834
use sg13g2_buf_2  fanout363
timestamp 1746816402
transform 1 0 13344 0 1 20412
box -48 -56 528 834
use sg13g2_buf_2  fanout364
timestamp 1746816402
transform 1 0 12000 0 -1 21924
box -48 -56 528 834
use sg13g2_buf_1  fanout365
timestamp 1746816402
transform 1 0 13152 0 1 18900
box -48 -56 432 834
use sg13g2_buf_2  fanout366
timestamp 1746816402
transform 1 0 10080 0 -1 15876
box -48 -56 528 834
use sg13g2_buf_2  fanout367
timestamp 1746816402
transform 1 0 13056 0 1 15876
box -48 -56 528 834
use sg13g2_buf_2  fanout368
timestamp 1746816402
transform -1 0 17184 0 1 15876
box -48 -56 528 834
use sg13g2_buf_1  fanout369
timestamp 1746816402
transform -1 0 15744 0 -1 15876
box -48 -56 432 834
use sg13g2_buf_4  fanout370
timestamp 1746816402
transform 1 0 3840 0 1 17388
box -48 -56 816 834
use sg13g2_buf_2  fanout371
timestamp 1746816402
transform -1 0 21024 0 1 24948
box -48 -56 528 834
use sg13g2_buf_2  fanout372
timestamp 1746816402
transform 1 0 15744 0 1 20412
box -48 -56 528 834
use sg13g2_buf_4  fanout373
timestamp 1746816402
transform -1 0 19200 0 1 15876
box -48 -56 816 834
use sg13g2_buf_4  fanout374
timestamp 1746816402
transform -1 0 19296 0 -1 14364
box -48 -56 816 834
use sg13g2_buf_2  fanout375
timestamp 1746816402
transform -1 0 8544 0 -1 20412
box -48 -56 528 834
use sg13g2_buf_2  fanout376
timestamp 1746816402
transform -1 0 9024 0 -1 20412
box -48 -56 528 834
use sg13g2_buf_2  fanout377
timestamp 1746816402
transform 1 0 11136 0 1 20412
box -48 -56 528 834
use sg13g2_buf_2  fanout378
timestamp 1746816402
transform -1 0 12096 0 1 18900
box -48 -56 528 834
use sg13g2_buf_2  fanout379
timestamp 1746816402
transform -1 0 27840 0 -1 21924
box -48 -56 528 834
use sg13g2_buf_2  fanout380
timestamp 1746816402
transform 1 0 23520 0 -1 24948
box -48 -56 528 834
use sg13g2_buf_2  fanout381
timestamp 1746816402
transform 1 0 26304 0 -1 20412
box -48 -56 528 834
use sg13g2_buf_2  fanout382
timestamp 1746816402
transform 1 0 17472 0 1 8316
box -48 -56 528 834
use sg13g2_buf_2  fanout383
timestamp 1746816402
transform -1 0 20544 0 -1 5292
box -48 -56 528 834
use sg13g2_buf_2  fanout384
timestamp 1746816402
transform 1 0 14976 0 1 3780
box -48 -56 528 834
use sg13g2_buf_2  fanout385
timestamp 1746816402
transform 1 0 9600 0 1 3780
box -48 -56 528 834
use sg13g2_buf_2  fanout386
timestamp 1746816402
transform -1 0 10848 0 1 3780
box -48 -56 528 834
use sg13g2_buf_2  fanout387
timestamp 1746816402
transform 1 0 6912 0 1 5292
box -48 -56 528 834
use sg13g2_buf_2  fanout388
timestamp 1746816402
transform -1 0 7968 0 -1 5292
box -48 -56 528 834
use sg13g2_buf_2  fanout389
timestamp 1746816402
transform 1 0 1920 0 1 6804
box -48 -56 528 834
use sg13g2_buf_2  fanout390
timestamp 1746816402
transform 1 0 5184 0 -1 6804
box -48 -56 528 834
use sg13g2_buf_2  fanout391
timestamp 1746816402
transform -1 0 1728 0 -1 8316
box -48 -56 528 834
use sg13g2_buf_2  fanout392
timestamp 1746816402
transform -1 0 27168 0 1 12852
box -48 -56 528 834
use sg13g2_buf_2  fanout393
timestamp 1746816402
transform -1 0 30336 0 1 12852
box -48 -56 528 834
use sg13g2_buf_2  fanout394
timestamp 1746816402
transform -1 0 26016 0 1 15876
box -48 -56 528 834
use sg13g2_buf_2  fanout395
timestamp 1746816402
transform 1 0 25632 0 -1 9828
box -48 -56 528 834
use sg13g2_buf_4  fanout396
timestamp 1746816402
transform 1 0 28032 0 -1 11340
box -48 -56 816 834
use sg13g2_buf_2  fanout397
timestamp 1746816402
transform -1 0 24480 0 1 6804
box -48 -56 528 834
use sg13g2_buf_4  fanout398
timestamp 1746816402
transform 1 0 24576 0 1 11340
box -48 -56 816 834
use sg13g2_buf_2  fanout399
timestamp 1746816402
transform 1 0 24672 0 1 6804
box -48 -56 528 834
use sg13g2_buf_4  fanout400
timestamp 1746816402
transform 1 0 25440 0 1 11340
box -48 -56 816 834
use sg13g2_buf_2  fanout401
timestamp 1746816402
transform 1 0 9888 0 -1 9828
box -48 -56 528 834
use sg13g2_buf_4  fanout402
timestamp 1746816402
transform 1 0 23904 0 1 14364
box -48 -56 816 834
use sg13g2_buf_2  fanout403
timestamp 1746816402
transform 1 0 8256 0 1 11340
box -48 -56 528 834
use sg13g2_buf_2  fanout404
timestamp 1746816402
transform 1 0 22656 0 -1 12852
box -48 -56 528 834
use sg13g2_buf_2  fanout405
timestamp 1746816402
transform 1 0 1344 0 -1 14364
box -48 -56 528 834
use sg13g2_buf_2  fanout406
timestamp 1746816402
transform 1 0 6528 0 -1 15876
box -48 -56 528 834
use sg13g2_buf_2  fanout407
timestamp 1746816402
transform -1 0 22848 0 1 15876
box -48 -56 528 834
use sg13g2_buf_4  fanout408
timestamp 1746816402
transform 1 0 26016 0 1 17388
box -48 -56 816 834
use sg13g2_buf_4  fanout409
timestamp 1746816402
transform 1 0 9792 0 1 24948
box -48 -56 816 834
use sg13g2_buf_1  fanout410
timestamp 1746816402
transform -1 0 7872 0 1 26460
box -48 -56 432 834
use sg13g2_buf_2  fanout411
timestamp 1746816402
transform -1 0 11328 0 1 24948
box -48 -56 528 834
use sg13g2_buf_4  fanout412
timestamp 1746816402
transform 1 0 18240 0 1 23436
box -48 -56 816 834
use sg13g2_buf_4  fanout413
timestamp 1746816402
transform 1 0 20352 0 1 20412
box -48 -56 816 834
use sg13g2_buf_2  fanout414
timestamp 1746816402
transform -1 0 19488 0 1 23436
box -48 -56 528 834
use sg13g2_buf_2  fanout415
timestamp 1746816402
transform -1 0 3264 0 -1 26460
box -48 -56 528 834
use sg13g2_buf_4  fanout416
timestamp 1746816402
transform -1 0 15360 0 1 26460
box -48 -56 816 834
use sg13g2_buf_4  fanout417
timestamp 1746816402
transform -1 0 21984 0 -1 26460
box -48 -56 816 834
use sg13g2_buf_2  fanout418
timestamp 1746816402
transform -1 0 18912 0 -1 24948
box -48 -56 528 834
use sg13g2_decap_8  FILLER_0_0
timestamp 1746816402
transform 1 0 576 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_7
timestamp 1746816402
transform 1 0 1248 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_14
timestamp 1746816402
transform 1 0 1920 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_21
timestamp 1746816402
transform 1 0 2592 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_28
timestamp 1746816402
transform 1 0 3264 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_35
timestamp 1746816402
transform 1 0 3936 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_42
timestamp 1746816402
transform 1 0 4608 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_49
timestamp 1746816402
transform 1 0 5280 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_56
timestamp 1746816402
transform 1 0 5952 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_63
timestamp 1746816402
transform 1 0 6624 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_70
timestamp 1746816402
transform 1 0 7296 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_77
timestamp 1746816402
transform 1 0 7968 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_84
timestamp 1746816402
transform 1 0 8640 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_91
timestamp 1746816402
transform 1 0 9312 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_98
timestamp 1746816402
transform 1 0 9984 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_105
timestamp 1746816402
transform 1 0 10656 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_112
timestamp 1746816402
transform 1 0 11328 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_119
timestamp 1746816402
transform 1 0 12000 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_126
timestamp 1746816402
transform 1 0 12672 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_133
timestamp 1746816402
transform 1 0 13344 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_140
timestamp 1746816402
transform 1 0 14016 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_147
timestamp 1746816402
transform 1 0 14688 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_154
timestamp 1746816402
transform 1 0 15360 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_161
timestamp 1746816402
transform 1 0 16032 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_168
timestamp 1746816402
transform 1 0 16704 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_175
timestamp 1746816402
transform 1 0 17376 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_182
timestamp 1746816402
transform 1 0 18048 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_189
timestamp 1746816402
transform 1 0 18720 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_196
timestamp 1746816402
transform 1 0 19392 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_203
timestamp 1746816402
transform 1 0 20064 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_210
timestamp 1746816402
transform 1 0 20736 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_217
timestamp 1746816402
transform 1 0 21408 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_224
timestamp 1746816402
transform 1 0 22080 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_231
timestamp 1746816402
transform 1 0 22752 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_238
timestamp 1746816402
transform 1 0 23424 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_245
timestamp 1746816402
transform 1 0 24096 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_252
timestamp 1746816402
transform 1 0 24768 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_259
timestamp 1746816402
transform 1 0 25440 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_266
timestamp 1746816402
transform 1 0 26112 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_273
timestamp 1746816402
transform 1 0 26784 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_280
timestamp 1746816402
transform 1 0 27456 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_287
timestamp 1746816402
transform 1 0 28128 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_294
timestamp 1746816402
transform 1 0 28800 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_301
timestamp 1746816402
transform 1 0 29472 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_308
timestamp 1746816402
transform 1 0 30144 0 1 756
box -48 -56 720 834
use sg13g2_decap_4  FILLER_0_315
timestamp 1746816402
transform 1 0 30816 0 1 756
box -48 -56 432 834
use sg13g2_fill_2  FILLER_0_319
timestamp 1746816402
transform 1 0 31200 0 1 756
box -48 -56 240 834
use sg13g2_decap_8  FILLER_1_0
timestamp 1746816402
transform 1 0 576 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_7
timestamp 1746816402
transform 1 0 1248 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_14
timestamp 1746816402
transform 1 0 1920 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_21
timestamp 1746816402
transform 1 0 2592 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_28
timestamp 1746816402
transform 1 0 3264 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_35
timestamp 1746816402
transform 1 0 3936 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_42
timestamp 1746816402
transform 1 0 4608 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_49
timestamp 1746816402
transform 1 0 5280 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_56
timestamp 1746816402
transform 1 0 5952 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_63
timestamp 1746816402
transform 1 0 6624 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_70
timestamp 1746816402
transform 1 0 7296 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_77
timestamp 1746816402
transform 1 0 7968 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_84
timestamp 1746816402
transform 1 0 8640 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_91
timestamp 1746816402
transform 1 0 9312 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_98
timestamp 1746816402
transform 1 0 9984 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_105
timestamp 1746816402
transform 1 0 10656 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_112
timestamp 1746816402
transform 1 0 11328 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_119
timestamp 1746816402
transform 1 0 12000 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_126
timestamp 1746816402
transform 1 0 12672 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_133
timestamp 1746816402
transform 1 0 13344 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_140
timestamp 1746816402
transform 1 0 14016 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_147
timestamp 1746816402
transform 1 0 14688 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_154
timestamp 1746816402
transform 1 0 15360 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_161
timestamp 1746816402
transform 1 0 16032 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_168
timestamp 1746816402
transform 1 0 16704 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_175
timestamp 1746816402
transform 1 0 17376 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_182
timestamp 1746816402
transform 1 0 18048 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_189
timestamp 1746816402
transform 1 0 18720 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_196
timestamp 1746816402
transform 1 0 19392 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_203
timestamp 1746816402
transform 1 0 20064 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_210
timestamp 1746816402
transform 1 0 20736 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_217
timestamp 1746816402
transform 1 0 21408 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_224
timestamp 1746816402
transform 1 0 22080 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_231
timestamp 1746816402
transform 1 0 22752 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_238
timestamp 1746816402
transform 1 0 23424 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_245
timestamp 1746816402
transform 1 0 24096 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_252
timestamp 1746816402
transform 1 0 24768 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_259
timestamp 1746816402
transform 1 0 25440 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_266
timestamp 1746816402
transform 1 0 26112 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_273
timestamp 1746816402
transform 1 0 26784 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_280
timestamp 1746816402
transform 1 0 27456 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_287
timestamp 1746816402
transform 1 0 28128 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_294
timestamp 1746816402
transform 1 0 28800 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_301
timestamp 1746816402
transform 1 0 29472 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_308
timestamp 1746816402
transform 1 0 30144 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_1_315
timestamp 1746816402
transform 1 0 30816 0 -1 2268
box -48 -56 432 834
use sg13g2_fill_2  FILLER_1_319
timestamp 1746816402
transform 1 0 31200 0 -1 2268
box -48 -56 240 834
use sg13g2_decap_8  FILLER_2_0
timestamp 1746816402
transform 1 0 576 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_7
timestamp 1746816402
transform 1 0 1248 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_14
timestamp 1746816402
transform 1 0 1920 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_21
timestamp 1746816402
transform 1 0 2592 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_28
timestamp 1746816402
transform 1 0 3264 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_35
timestamp 1746816402
transform 1 0 3936 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_42
timestamp 1746816402
transform 1 0 4608 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_49
timestamp 1746816402
transform 1 0 5280 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_56
timestamp 1746816402
transform 1 0 5952 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_63
timestamp 1746816402
transform 1 0 6624 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_70
timestamp 1746816402
transform 1 0 7296 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_77
timestamp 1746816402
transform 1 0 7968 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_84
timestamp 1746816402
transform 1 0 8640 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_91
timestamp 1746816402
transform 1 0 9312 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_98
timestamp 1746816402
transform 1 0 9984 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_105
timestamp 1746816402
transform 1 0 10656 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_112
timestamp 1746816402
transform 1 0 11328 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_119
timestamp 1746816402
transform 1 0 12000 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_126
timestamp 1746816402
transform 1 0 12672 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_133
timestamp 1746816402
transform 1 0 13344 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_140
timestamp 1746816402
transform 1 0 14016 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_147
timestamp 1746816402
transform 1 0 14688 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_154
timestamp 1746816402
transform 1 0 15360 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_161
timestamp 1746816402
transform 1 0 16032 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_168
timestamp 1746816402
transform 1 0 16704 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_175
timestamp 1746816402
transform 1 0 17376 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_182
timestamp 1746816402
transform 1 0 18048 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_189
timestamp 1746816402
transform 1 0 18720 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_196
timestamp 1746816402
transform 1 0 19392 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_203
timestamp 1746816402
transform 1 0 20064 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_210
timestamp 1746816402
transform 1 0 20736 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_217
timestamp 1746816402
transform 1 0 21408 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_224
timestamp 1746816402
transform 1 0 22080 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_231
timestamp 1746816402
transform 1 0 22752 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_238
timestamp 1746816402
transform 1 0 23424 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_245
timestamp 1746816402
transform 1 0 24096 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_252
timestamp 1746816402
transform 1 0 24768 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_259
timestamp 1746816402
transform 1 0 25440 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_266
timestamp 1746816402
transform 1 0 26112 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_273
timestamp 1746816402
transform 1 0 26784 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_280
timestamp 1746816402
transform 1 0 27456 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_287
timestamp 1746816402
transform 1 0 28128 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_294
timestamp 1746816402
transform 1 0 28800 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_301
timestamp 1746816402
transform 1 0 29472 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_308
timestamp 1746816402
transform 1 0 30144 0 1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_315
timestamp 1746816402
transform 1 0 30816 0 1 2268
box -48 -56 432 834
use sg13g2_fill_2  FILLER_2_319
timestamp 1746816402
transform 1 0 31200 0 1 2268
box -48 -56 240 834
use sg13g2_decap_8  FILLER_3_0
timestamp 1746816402
transform 1 0 576 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_7
timestamp 1746816402
transform 1 0 1248 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_14
timestamp 1746816402
transform 1 0 1920 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_21
timestamp 1746816402
transform 1 0 2592 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_28
timestamp 1746816402
transform 1 0 3264 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_35
timestamp 1746816402
transform 1 0 3936 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_42
timestamp 1746816402
transform 1 0 4608 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_49
timestamp 1746816402
transform 1 0 5280 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_56
timestamp 1746816402
transform 1 0 5952 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_63
timestamp 1746816402
transform 1 0 6624 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_70
timestamp 1746816402
transform 1 0 7296 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_77
timestamp 1746816402
transform 1 0 7968 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_84
timestamp 1746816402
transform 1 0 8640 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_91
timestamp 1746816402
transform 1 0 9312 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_98
timestamp 1746816402
transform 1 0 9984 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_105
timestamp 1746816402
transform 1 0 10656 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_112
timestamp 1746816402
transform 1 0 11328 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_119
timestamp 1746816402
transform 1 0 12000 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_126
timestamp 1746816402
transform 1 0 12672 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_133
timestamp 1746816402
transform 1 0 13344 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_140
timestamp 1746816402
transform 1 0 14016 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_147
timestamp 1746816402
transform 1 0 14688 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_154
timestamp 1746816402
transform 1 0 15360 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_161
timestamp 1746816402
transform 1 0 16032 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_168
timestamp 1746816402
transform 1 0 16704 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_175
timestamp 1746816402
transform 1 0 17376 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_182
timestamp 1746816402
transform 1 0 18048 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_189
timestamp 1746816402
transform 1 0 18720 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_196
timestamp 1746816402
transform 1 0 19392 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_203
timestamp 1746816402
transform 1 0 20064 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_210
timestamp 1746816402
transform 1 0 20736 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_217
timestamp 1746816402
transform 1 0 21408 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_224
timestamp 1746816402
transform 1 0 22080 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_231
timestamp 1746816402
transform 1 0 22752 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_238
timestamp 1746816402
transform 1 0 23424 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_245
timestamp 1746816402
transform 1 0 24096 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_252
timestamp 1746816402
transform 1 0 24768 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_259
timestamp 1746816402
transform 1 0 25440 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_266
timestamp 1746816402
transform 1 0 26112 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_273
timestamp 1746816402
transform 1 0 26784 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_280
timestamp 1746816402
transform 1 0 27456 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_287
timestamp 1746816402
transform 1 0 28128 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_294
timestamp 1746816402
transform 1 0 28800 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_301
timestamp 1746816402
transform 1 0 29472 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_308
timestamp 1746816402
transform 1 0 30144 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_315
timestamp 1746816402
transform 1 0 30816 0 -1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_3_319
timestamp 1746816402
transform 1 0 31200 0 -1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_4_0
timestamp 1746816402
transform 1 0 576 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_7
timestamp 1746816402
transform 1 0 1248 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_14
timestamp 1746816402
transform 1 0 1920 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_21
timestamp 1746816402
transform 1 0 2592 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_28
timestamp 1746816402
transform 1 0 3264 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_35
timestamp 1746816402
transform 1 0 3936 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_42
timestamp 1746816402
transform 1 0 4608 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_49
timestamp 1746816402
transform 1 0 5280 0 1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_4_56
timestamp 1746816402
transform 1 0 5952 0 1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_4_62
timestamp 1746816402
transform 1 0 6528 0 1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_4_69
timestamp 1746816402
transform 1 0 7200 0 1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_71
timestamp 1746816402
transform 1 0 7392 0 1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_85
timestamp 1746816402
transform 1 0 8736 0 1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_4_92
timestamp 1746816402
transform 1 0 9408 0 1 3780
box -48 -56 240 834
use sg13g2_fill_2  FILLER_4_99
timestamp 1746816402
transform 1 0 10080 0 1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_101
timestamp 1746816402
transform 1 0 10272 0 1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_107
timestamp 1746816402
transform 1 0 10848 0 1 3780
box -48 -56 720 834
use sg13g2_fill_1  FILLER_4_114
timestamp 1746816402
transform 1 0 11520 0 1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_119
timestamp 1746816402
transform 1 0 12000 0 1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_126
timestamp 1746816402
transform 1 0 12672 0 1 3780
box -48 -56 432 834
use sg13g2_fill_1  FILLER_4_130
timestamp 1746816402
transform 1 0 13056 0 1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_4_148
timestamp 1746816402
transform 1 0 14784 0 1 3780
box -48 -56 240 834
use sg13g2_fill_2  FILLER_4_155
timestamp 1746816402
transform 1 0 15456 0 1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_157
timestamp 1746816402
transform 1 0 15648 0 1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_163
timestamp 1746816402
transform 1 0 16224 0 1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_4_170
timestamp 1746816402
transform 1 0 16896 0 1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_4_176
timestamp 1746816402
transform 1 0 17472 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_183
timestamp 1746816402
transform 1 0 18144 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_190
timestamp 1746816402
transform 1 0 18816 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_197
timestamp 1746816402
transform 1 0 19488 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_204
timestamp 1746816402
transform 1 0 20160 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_211
timestamp 1746816402
transform 1 0 20832 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_218
timestamp 1746816402
transform 1 0 21504 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_225
timestamp 1746816402
transform 1 0 22176 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_232
timestamp 1746816402
transform 1 0 22848 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_239
timestamp 1746816402
transform 1 0 23520 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_246
timestamp 1746816402
transform 1 0 24192 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_253
timestamp 1746816402
transform 1 0 24864 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_260
timestamp 1746816402
transform 1 0 25536 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_267
timestamp 1746816402
transform 1 0 26208 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_274
timestamp 1746816402
transform 1 0 26880 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_281
timestamp 1746816402
transform 1 0 27552 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_288
timestamp 1746816402
transform 1 0 28224 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_295
timestamp 1746816402
transform 1 0 28896 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_302
timestamp 1746816402
transform 1 0 29568 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_309
timestamp 1746816402
transform 1 0 30240 0 1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_316
timestamp 1746816402
transform 1 0 30912 0 1 3780
box -48 -56 432 834
use sg13g2_fill_1  FILLER_4_320
timestamp 1746816402
transform 1 0 31296 0 1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_0
timestamp 1746816402
transform 1 0 576 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_7
timestamp 1746816402
transform 1 0 1248 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_14
timestamp 1746816402
transform 1 0 1920 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_21
timestamp 1746816402
transform 1 0 2592 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_28
timestamp 1746816402
transform 1 0 3264 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_35
timestamp 1746816402
transform 1 0 3936 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_42
timestamp 1746816402
transform 1 0 4608 0 -1 5292
box -48 -56 432 834
use sg13g2_fill_1  FILLER_5_120
timestamp 1746816402
transform 1 0 12096 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_4  FILLER_5_157
timestamp 1746816402
transform 1 0 15648 0 -1 5292
box -48 -56 432 834
use sg13g2_decap_8  FILLER_5_192
timestamp 1746816402
transform 1 0 19008 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_199
timestamp 1746816402
transform 1 0 19680 0 -1 5292
box -48 -56 432 834
use sg13g2_fill_2  FILLER_5_208
timestamp 1746816402
transform 1 0 20544 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_210
timestamp 1746816402
transform 1 0 20736 0 -1 5292
box -48 -56 144 834
use sg13g2_fill_1  FILLER_5_218
timestamp 1746816402
transform 1 0 21504 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_228
timestamp 1746816402
transform 1 0 22464 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_235
timestamp 1746816402
transform 1 0 23136 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_242
timestamp 1746816402
transform 1 0 23808 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_249
timestamp 1746816402
transform 1 0 24480 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_256
timestamp 1746816402
transform 1 0 25152 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_263
timestamp 1746816402
transform 1 0 25824 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_270
timestamp 1746816402
transform 1 0 26496 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_277
timestamp 1746816402
transform 1 0 27168 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_284
timestamp 1746816402
transform 1 0 27840 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_291
timestamp 1746816402
transform 1 0 28512 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_298
timestamp 1746816402
transform 1 0 29184 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_305
timestamp 1746816402
transform 1 0 29856 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_312
timestamp 1746816402
transform 1 0 30528 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_319
timestamp 1746816402
transform 1 0 31200 0 -1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_6_0
timestamp 1746816402
transform 1 0 576 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_7
timestamp 1746816402
transform 1 0 1248 0 1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_14
timestamp 1746816402
transform 1 0 1920 0 1 5292
box -48 -56 432 834
use sg13g2_fill_1  FILLER_6_18
timestamp 1746816402
transform 1 0 2304 0 1 5292
box -48 -56 144 834
use sg13g2_fill_1  FILLER_6_33
timestamp 1746816402
transform 1 0 3744 0 1 5292
box -48 -56 144 834
use sg13g2_fill_2  FILLER_6_80
timestamp 1746816402
transform 1 0 8256 0 1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_101
timestamp 1746816402
transform 1 0 10272 0 1 5292
box -48 -56 144 834
use sg13g2_fill_1  FILLER_6_166
timestamp 1746816402
transform 1 0 16512 0 1 5292
box -48 -56 144 834
use sg13g2_fill_1  FILLER_6_196
timestamp 1746816402
transform 1 0 19392 0 1 5292
box -48 -56 144 834
use sg13g2_fill_1  FILLER_6_214
timestamp 1746816402
transform 1 0 21120 0 1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_245
timestamp 1746816402
transform 1 0 24096 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_252
timestamp 1746816402
transform 1 0 24768 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_259
timestamp 1746816402
transform 1 0 25440 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_266
timestamp 1746816402
transform 1 0 26112 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_273
timestamp 1746816402
transform 1 0 26784 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_280
timestamp 1746816402
transform 1 0 27456 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_287
timestamp 1746816402
transform 1 0 28128 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_294
timestamp 1746816402
transform 1 0 28800 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_301
timestamp 1746816402
transform 1 0 29472 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_308
timestamp 1746816402
transform 1 0 30144 0 1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_315
timestamp 1746816402
transform 1 0 30816 0 1 5292
box -48 -56 432 834
use sg13g2_fill_2  FILLER_6_319
timestamp 1746816402
transform 1 0 31200 0 1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_7_0
timestamp 1746816402
transform 1 0 576 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_7
timestamp 1746816402
transform 1 0 1248 0 -1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_7_14
timestamp 1746816402
transform 1 0 1920 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_16
timestamp 1746816402
transform 1 0 2112 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_7_53
timestamp 1746816402
transform 1 0 5664 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_2  FILLER_7_65
timestamp 1746816402
transform 1 0 6816 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_109
timestamp 1746816402
transform 1 0 11040 0 -1 6804
box -48 -56 144 834
use sg13g2_decap_4  FILLER_7_123
timestamp 1746816402
transform 1 0 12384 0 -1 6804
box -48 -56 432 834
use sg13g2_decap_4  FILLER_7_145
timestamp 1746816402
transform 1 0 14496 0 -1 6804
box -48 -56 432 834
use sg13g2_fill_1  FILLER_7_149
timestamp 1746816402
transform 1 0 14880 0 -1 6804
box -48 -56 144 834
use sg13g2_decap_4  FILLER_7_176
timestamp 1746816402
transform 1 0 17472 0 -1 6804
box -48 -56 432 834
use sg13g2_decap_4  FILLER_7_188
timestamp 1746816402
transform 1 0 18624 0 -1 6804
box -48 -56 432 834
use sg13g2_fill_1  FILLER_7_192
timestamp 1746816402
transform 1 0 19008 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_7_219
timestamp 1746816402
transform 1 0 21600 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_7_230
timestamp 1746816402
transform 1 0 22656 0 -1 6804
box -48 -56 240 834
use sg13g2_decap_8  FILLER_7_250
timestamp 1746816402
transform 1 0 24576 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_257
timestamp 1746816402
transform 1 0 25248 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_264
timestamp 1746816402
transform 1 0 25920 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_271
timestamp 1746816402
transform 1 0 26592 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_278
timestamp 1746816402
transform 1 0 27264 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_285
timestamp 1746816402
transform 1 0 27936 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_292
timestamp 1746816402
transform 1 0 28608 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_299
timestamp 1746816402
transform 1 0 29280 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_306
timestamp 1746816402
transform 1 0 29952 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_313
timestamp 1746816402
transform 1 0 30624 0 -1 6804
box -48 -56 720 834
use sg13g2_fill_1  FILLER_7_320
timestamp 1746816402
transform 1 0 31296 0 -1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_0
timestamp 1746816402
transform 1 0 576 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_7
timestamp 1746816402
transform 1 0 1248 0 1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_8_70
timestamp 1746816402
transform 1 0 7296 0 1 6804
box -48 -56 240 834
use sg13g2_fill_2  FILLER_8_85
timestamp 1746816402
transform 1 0 8736 0 1 6804
box -48 -56 240 834
use sg13g2_fill_2  FILLER_8_107
timestamp 1746816402
transform 1 0 10848 0 1 6804
box -48 -56 240 834
use sg13g2_decap_4  FILLER_8_117
timestamp 1746816402
transform 1 0 11808 0 1 6804
box -48 -56 432 834
use sg13g2_decap_4  FILLER_8_137
timestamp 1746816402
transform 1 0 13728 0 1 6804
box -48 -56 432 834
use sg13g2_decap_4  FILLER_8_168
timestamp 1746816402
transform 1 0 16704 0 1 6804
box -48 -56 432 834
use sg13g2_fill_1  FILLER_8_172
timestamp 1746816402
transform 1 0 17088 0 1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_8_205
timestamp 1746816402
transform 1 0 20256 0 1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_8_229
timestamp 1746816402
transform 1 0 22560 0 1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_8_242
timestamp 1746816402
transform 1 0 23808 0 1 6804
box -48 -56 240 834
use sg13g2_fill_2  FILLER_8_249
timestamp 1746816402
transform 1 0 24480 0 1 6804
box -48 -56 240 834
use sg13g2_decap_4  FILLER_8_260
timestamp 1746816402
transform 1 0 25536 0 1 6804
box -48 -56 432 834
use sg13g2_fill_2  FILLER_8_264
timestamp 1746816402
transform 1 0 25920 0 1 6804
box -48 -56 240 834
use sg13g2_decap_4  FILLER_8_271
timestamp 1746816402
transform 1 0 26592 0 1 6804
box -48 -56 432 834
use sg13g2_fill_2  FILLER_8_275
timestamp 1746816402
transform 1 0 26976 0 1 6804
box -48 -56 240 834
use sg13g2_decap_8  FILLER_8_282
timestamp 1746816402
transform 1 0 27648 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_289
timestamp 1746816402
transform 1 0 28320 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_296
timestamp 1746816402
transform 1 0 28992 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_303
timestamp 1746816402
transform 1 0 29664 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_310
timestamp 1746816402
transform 1 0 30336 0 1 6804
box -48 -56 720 834
use sg13g2_decap_4  FILLER_8_317
timestamp 1746816402
transform 1 0 31008 0 1 6804
box -48 -56 432 834
use sg13g2_decap_8  FILLER_9_0
timestamp 1746816402
transform 1 0 576 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_4  FILLER_9_16
timestamp 1746816402
transform 1 0 2112 0 -1 8316
box -48 -56 432 834
use sg13g2_fill_1  FILLER_9_20
timestamp 1746816402
transform 1 0 2496 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_9_30
timestamp 1746816402
transform 1 0 3456 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_32
timestamp 1746816402
transform 1 0 3648 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_9_41
timestamp 1746816402
transform 1 0 4512 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_43
timestamp 1746816402
transform 1 0 4704 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_4  FILLER_9_50
timestamp 1746816402
transform 1 0 5376 0 -1 8316
box -48 -56 432 834
use sg13g2_fill_2  FILLER_9_64
timestamp 1746816402
transform 1 0 6720 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_66
timestamp 1746816402
transform 1 0 6912 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_4  FILLER_9_108
timestamp 1746816402
transform 1 0 10944 0 -1 8316
box -48 -56 432 834
use sg13g2_decap_4  FILLER_9_122
timestamp 1746816402
transform 1 0 12288 0 -1 8316
box -48 -56 432 834
use sg13g2_fill_1  FILLER_9_131
timestamp 1746816402
transform 1 0 13152 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_9_138
timestamp 1746816402
transform 1 0 13824 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_140
timestamp 1746816402
transform 1 0 14016 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_4  FILLER_9_169
timestamp 1746816402
transform 1 0 16800 0 -1 8316
box -48 -56 432 834
use sg13g2_decap_4  FILLER_9_188
timestamp 1746816402
transform 1 0 18624 0 -1 8316
box -48 -56 432 834
use sg13g2_fill_2  FILLER_9_210
timestamp 1746816402
transform 1 0 20736 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_212
timestamp 1746816402
transform 1 0 20928 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_9_222
timestamp 1746816402
transform 1 0 21888 0 -1 8316
box -48 -56 240 834
use sg13g2_decap_8  FILLER_9_292
timestamp 1746816402
transform 1 0 28608 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_299
timestamp 1746816402
transform 1 0 29280 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_306
timestamp 1746816402
transform 1 0 29952 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_313
timestamp 1746816402
transform 1 0 30624 0 -1 8316
box -48 -56 720 834
use sg13g2_fill_1  FILLER_9_320
timestamp 1746816402
transform 1 0 31296 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_10_26
timestamp 1746816402
transform 1 0 3072 0 1 8316
box -48 -56 240 834
use sg13g2_fill_2  FILLER_10_75
timestamp 1746816402
transform 1 0 7776 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_77
timestamp 1746816402
transform 1 0 7968 0 1 8316
box -48 -56 144 834
use sg13g2_decap_4  FILLER_10_83
timestamp 1746816402
transform 1 0 8544 0 1 8316
box -48 -56 432 834
use sg13g2_fill_2  FILLER_10_87
timestamp 1746816402
transform 1 0 8928 0 1 8316
box -48 -56 240 834
use sg13g2_fill_2  FILLER_10_99
timestamp 1746816402
transform 1 0 10080 0 1 8316
box -48 -56 240 834
use sg13g2_decap_4  FILLER_10_111
timestamp 1746816402
transform 1 0 11232 0 1 8316
box -48 -56 432 834
use sg13g2_decap_4  FILLER_10_145
timestamp 1746816402
transform 1 0 14496 0 1 8316
box -48 -56 432 834
use sg13g2_fill_1  FILLER_10_149
timestamp 1746816402
transform 1 0 14880 0 1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_10_160
timestamp 1746816402
transform 1 0 15936 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_175
timestamp 1746816402
transform 1 0 17376 0 1 8316
box -48 -56 144 834
use sg13g2_decap_4  FILLER_10_181
timestamp 1746816402
transform 1 0 17952 0 1 8316
box -48 -56 432 834
use sg13g2_fill_1  FILLER_10_185
timestamp 1746816402
transform 1 0 18336 0 1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_10_191
timestamp 1746816402
transform 1 0 18912 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_193
timestamp 1746816402
transform 1 0 19104 0 1 8316
box -48 -56 144 834
use sg13g2_fill_1  FILLER_10_207
timestamp 1746816402
transform 1 0 20448 0 1 8316
box -48 -56 144 834
use sg13g2_decap_4  FILLER_10_239
timestamp 1746816402
transform 1 0 23520 0 1 8316
box -48 -56 432 834
use sg13g2_fill_2  FILLER_10_243
timestamp 1746816402
transform 1 0 23904 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_261
timestamp 1746816402
transform 1 0 25632 0 1 8316
box -48 -56 144 834
use sg13g2_fill_1  FILLER_10_279
timestamp 1746816402
transform 1 0 27360 0 1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_298
timestamp 1746816402
transform 1 0 29184 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_305
timestamp 1746816402
transform 1 0 29856 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_312
timestamp 1746816402
transform 1 0 30528 0 1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_10_319
timestamp 1746816402
transform 1 0 31200 0 1 8316
box -48 -56 240 834
use sg13g2_fill_2  FILLER_11_0
timestamp 1746816402
transform 1 0 576 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_2
timestamp 1746816402
transform 1 0 768 0 -1 9828
box -48 -56 144 834
use sg13g2_fill_2  FILLER_11_15
timestamp 1746816402
transform 1 0 2016 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_2  FILLER_11_45
timestamp 1746816402
transform 1 0 4896 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_57
timestamp 1746816402
transform 1 0 6048 0 -1 9828
box -48 -56 144 834
use sg13g2_fill_2  FILLER_11_62
timestamp 1746816402
transform 1 0 6528 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_2  FILLER_11_115
timestamp 1746816402
transform 1 0 11616 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_117
timestamp 1746816402
transform 1 0 11808 0 -1 9828
box -48 -56 144 834
use sg13g2_fill_2  FILLER_11_128
timestamp 1746816402
transform 1 0 12864 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_130
timestamp 1746816402
transform 1 0 13056 0 -1 9828
box -48 -56 144 834
use sg13g2_fill_1  FILLER_11_135
timestamp 1746816402
transform 1 0 13536 0 -1 9828
box -48 -56 144 834
use sg13g2_decap_4  FILLER_11_166
timestamp 1746816402
transform 1 0 16512 0 -1 9828
box -48 -56 432 834
use sg13g2_fill_1  FILLER_11_170
timestamp 1746816402
transform 1 0 16896 0 -1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_305
timestamp 1746816402
transform 1 0 29856 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_312
timestamp 1746816402
transform 1 0 30528 0 -1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_11_319
timestamp 1746816402
transform 1 0 31200 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_2  FILLER_12_72
timestamp 1746816402
transform 1 0 7488 0 1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_12_74
timestamp 1746816402
transform 1 0 7680 0 1 9828
box -48 -56 144 834
use sg13g2_fill_1  FILLER_12_80
timestamp 1746816402
transform 1 0 8256 0 1 9828
box -48 -56 144 834
use sg13g2_fill_2  FILLER_12_94
timestamp 1746816402
transform 1 0 9600 0 1 9828
box -48 -56 240 834
use sg13g2_fill_2  FILLER_12_101
timestamp 1746816402
transform 1 0 10272 0 1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_12_103
timestamp 1746816402
transform 1 0 10464 0 1 9828
box -48 -56 144 834
use sg13g2_fill_2  FILLER_12_109
timestamp 1746816402
transform 1 0 11040 0 1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_12_135
timestamp 1746816402
transform 1 0 13536 0 1 9828
box -48 -56 144 834
use sg13g2_fill_2  FILLER_12_157
timestamp 1746816402
transform 1 0 15648 0 1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_12_159
timestamp 1746816402
transform 1 0 15840 0 1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_12_186
timestamp 1746816402
transform 1 0 18432 0 1 9828
box -48 -56 720 834
use sg13g2_fill_1  FILLER_12_197
timestamp 1746816402
transform 1 0 19488 0 1 9828
box -48 -56 144 834
use sg13g2_decap_4  FILLER_12_203
timestamp 1746816402
transform 1 0 20064 0 1 9828
box -48 -56 432 834
use sg13g2_fill_2  FILLER_12_207
timestamp 1746816402
transform 1 0 20448 0 1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_12_217
timestamp 1746816402
transform 1 0 21408 0 1 9828
box -48 -56 144 834
use sg13g2_fill_2  FILLER_12_250
timestamp 1746816402
transform 1 0 24576 0 1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_12_252
timestamp 1746816402
transform 1 0 24768 0 1 9828
box -48 -56 144 834
use sg13g2_fill_1  FILLER_12_261
timestamp 1746816402
transform 1 0 25632 0 1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_12_301
timestamp 1746816402
transform 1 0 29472 0 1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_12_308
timestamp 1746816402
transform 1 0 30144 0 1 9828
box -48 -56 240 834
use sg13g2_fill_2  FILLER_12_318
timestamp 1746816402
transform 1 0 31104 0 1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_12_320
timestamp 1746816402
transform 1 0 31296 0 1 9828
box -48 -56 144 834
use sg13g2_fill_2  FILLER_13_0
timestamp 1746816402
transform 1 0 576 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_2  FILLER_13_14
timestamp 1746816402
transform 1 0 1920 0 -1 11340
box -48 -56 240 834
use sg13g2_decap_4  FILLER_13_38
timestamp 1746816402
transform 1 0 4224 0 -1 11340
box -48 -56 432 834
use sg13g2_fill_2  FILLER_13_42
timestamp 1746816402
transform 1 0 4608 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_2  FILLER_13_49
timestamp 1746816402
transform 1 0 5280 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_13_51
timestamp 1746816402
transform 1 0 5472 0 -1 11340
box -48 -56 144 834
use sg13g2_decap_4  FILLER_13_57
timestamp 1746816402
transform 1 0 6048 0 -1 11340
box -48 -56 432 834
use sg13g2_fill_2  FILLER_13_61
timestamp 1746816402
transform 1 0 6432 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_2  FILLER_13_78
timestamp 1746816402
transform 1 0 8064 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_13_80
timestamp 1746816402
transform 1 0 8256 0 -1 11340
box -48 -56 144 834
use sg13g2_decap_4  FILLER_13_86
timestamp 1746816402
transform 1 0 8832 0 -1 11340
box -48 -56 432 834
use sg13g2_fill_2  FILLER_13_90
timestamp 1746816402
transform 1 0 9216 0 -1 11340
box -48 -56 240 834
use sg13g2_decap_4  FILLER_13_107
timestamp 1746816402
transform 1 0 10848 0 -1 11340
box -48 -56 432 834
use sg13g2_fill_2  FILLER_13_123
timestamp 1746816402
transform 1 0 12384 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_13_125
timestamp 1746816402
transform 1 0 12576 0 -1 11340
box -48 -56 144 834
use sg13g2_decap_4  FILLER_13_161
timestamp 1746816402
transform 1 0 16032 0 -1 11340
box -48 -56 432 834
use sg13g2_fill_1  FILLER_13_165
timestamp 1746816402
transform 1 0 16416 0 -1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_13_194
timestamp 1746816402
transform 1 0 19200 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_2  FILLER_13_220
timestamp 1746816402
transform 1 0 21696 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_13_222
timestamp 1746816402
transform 1 0 21888 0 -1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_13_273
timestamp 1746816402
transform 1 0 26784 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_13_275
timestamp 1746816402
transform 1 0 26976 0 -1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_13_284
timestamp 1746816402
transform 1 0 27840 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_2  FILLER_13_318
timestamp 1746816402
transform 1 0 31104 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_13_320
timestamp 1746816402
transform 1 0 31296 0 -1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_14_0
timestamp 1746816402
transform 1 0 576 0 1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_14_2
timestamp 1746816402
transform 1 0 768 0 1 11340
box -48 -56 144 834
use sg13g2_fill_1  FILLER_14_107
timestamp 1746816402
transform 1 0 10848 0 1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_14_139
timestamp 1746816402
transform 1 0 13920 0 1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_14_141
timestamp 1746816402
transform 1 0 14112 0 1 11340
box -48 -56 144 834
use sg13g2_fill_1  FILLER_14_155
timestamp 1746816402
transform 1 0 15456 0 1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_14_180
timestamp 1746816402
transform 1 0 17856 0 1 11340
box -48 -56 240 834
use sg13g2_fill_2  FILLER_14_197
timestamp 1746816402
transform 1 0 19488 0 1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_14_199
timestamp 1746816402
transform 1 0 19680 0 1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_14_226
timestamp 1746816402
transform 1 0 22272 0 1 11340
box -48 -56 240 834
use sg13g2_fill_2  FILLER_14_240
timestamp 1746816402
transform 1 0 23616 0 1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_14_242
timestamp 1746816402
transform 1 0 23808 0 1 11340
box -48 -56 144 834
use sg13g2_fill_1  FILLER_14_249
timestamp 1746816402
transform 1 0 24480 0 1 11340
box -48 -56 144 834
use sg13g2_fill_1  FILLER_14_258
timestamp 1746816402
transform 1 0 25344 0 1 11340
box -48 -56 144 834
use sg13g2_fill_1  FILLER_14_307
timestamp 1746816402
transform 1 0 30048 0 1 11340
box -48 -56 144 834
use sg13g2_fill_1  FILLER_14_320
timestamp 1746816402
transform 1 0 31296 0 1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_15_26
timestamp 1746816402
transform 1 0 3072 0 -1 12852
box -48 -56 720 834
use sg13g2_fill_2  FILLER_15_33
timestamp 1746816402
transform 1 0 3744 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_2  FILLER_15_52
timestamp 1746816402
transform 1 0 5568 0 -1 12852
box -48 -56 240 834
use sg13g2_decap_4  FILLER_15_62
timestamp 1746816402
transform 1 0 6528 0 -1 12852
box -48 -56 432 834
use sg13g2_fill_1  FILLER_15_66
timestamp 1746816402
transform 1 0 6912 0 -1 12852
box -48 -56 144 834
use sg13g2_fill_1  FILLER_15_75
timestamp 1746816402
transform 1 0 7776 0 -1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_15_90
timestamp 1746816402
transform 1 0 9216 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_15_92
timestamp 1746816402
transform 1 0 9408 0 -1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_15_106
timestamp 1746816402
transform 1 0 10752 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_2  FILLER_15_122
timestamp 1746816402
transform 1 0 12288 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_15_124
timestamp 1746816402
transform 1 0 12480 0 -1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_15_141
timestamp 1746816402
transform 1 0 14112 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_15_143
timestamp 1746816402
transform 1 0 14304 0 -1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_15_163
timestamp 1746816402
transform 1 0 16224 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_15_165
timestamp 1746816402
transform 1 0 16416 0 -1 12852
box -48 -56 144 834
use sg13g2_decap_4  FILLER_15_174
timestamp 1746816402
transform 1 0 17280 0 -1 12852
box -48 -56 432 834
use sg13g2_fill_2  FILLER_15_178
timestamp 1746816402
transform 1 0 17664 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_2  FILLER_15_185
timestamp 1746816402
transform 1 0 18336 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_2  FILLER_15_192
timestamp 1746816402
transform 1 0 19008 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_15_194
timestamp 1746816402
transform 1 0 19200 0 -1 12852
box -48 -56 144 834
use sg13g2_fill_1  FILLER_15_203
timestamp 1746816402
transform 1 0 20064 0 -1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_15_235
timestamp 1746816402
transform 1 0 23136 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_15_237
timestamp 1746816402
transform 1 0 23328 0 -1 12852
box -48 -56 144 834
use sg13g2_fill_1  FILLER_15_310
timestamp 1746816402
transform 1 0 30336 0 -1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_15_319
timestamp 1746816402
transform 1 0 31200 0 -1 12852
box -48 -56 240 834
use sg13g2_decap_4  FILLER_16_0
timestamp 1746816402
transform 1 0 576 0 1 12852
box -48 -56 432 834
use sg13g2_fill_2  FILLER_16_4
timestamp 1746816402
transform 1 0 960 0 1 12852
box -48 -56 240 834
use sg13g2_fill_2  FILLER_16_11
timestamp 1746816402
transform 1 0 1632 0 1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_16_13
timestamp 1746816402
transform 1 0 1824 0 1 12852
box -48 -56 144 834
use sg13g2_decap_4  FILLER_16_19
timestamp 1746816402
transform 1 0 2400 0 1 12852
box -48 -56 432 834
use sg13g2_decap_4  FILLER_16_31
timestamp 1746816402
transform 1 0 3552 0 1 12852
box -48 -56 432 834
use sg13g2_fill_2  FILLER_16_51
timestamp 1746816402
transform 1 0 5472 0 1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_16_62
timestamp 1746816402
transform 1 0 6528 0 1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_16_90
timestamp 1746816402
transform 1 0 9216 0 1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_16_92
timestamp 1746816402
transform 1 0 9408 0 1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_16_98
timestamp 1746816402
transform 1 0 9984 0 1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_16_100
timestamp 1746816402
transform 1 0 10176 0 1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_16_108
timestamp 1746816402
transform 1 0 10944 0 1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_16_110
timestamp 1746816402
transform 1 0 11136 0 1 12852
box -48 -56 144 834
use sg13g2_fill_1  FILLER_16_124
timestamp 1746816402
transform 1 0 12480 0 1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_16_140
timestamp 1746816402
transform 1 0 14016 0 1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_16_157
timestamp 1746816402
transform 1 0 15648 0 1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_16_189
timestamp 1746816402
transform 1 0 18720 0 1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_16_191
timestamp 1746816402
transform 1 0 18912 0 1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_16_277
timestamp 1746816402
transform 1 0 27168 0 1 12852
box -48 -56 240 834
use sg13g2_decap_4  FILLER_17_0
timestamp 1746816402
transform 1 0 576 0 -1 14364
box -48 -56 432 834
use sg13g2_fill_1  FILLER_17_34
timestamp 1746816402
transform 1 0 3840 0 -1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_17_43
timestamp 1746816402
transform 1 0 4704 0 -1 14364
box -48 -56 240 834
use sg13g2_fill_2  FILLER_17_62
timestamp 1746816402
transform 1 0 6528 0 -1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_17_64
timestamp 1746816402
transform 1 0 6720 0 -1 14364
box -48 -56 144 834
use sg13g2_decap_4  FILLER_17_81
timestamp 1746816402
transform 1 0 8352 0 -1 14364
box -48 -56 432 834
use sg13g2_fill_2  FILLER_17_100
timestamp 1746816402
transform 1 0 10176 0 -1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_17_102
timestamp 1746816402
transform 1 0 10368 0 -1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_17_112
timestamp 1746816402
transform 1 0 11328 0 -1 14364
box -48 -56 240 834
use sg13g2_fill_2  FILLER_17_120
timestamp 1746816402
transform 1 0 12096 0 -1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_17_130
timestamp 1746816402
transform 1 0 13056 0 -1 14364
box -48 -56 144 834
use sg13g2_fill_1  FILLER_17_141
timestamp 1746816402
transform 1 0 14112 0 -1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_17_152
timestamp 1746816402
transform 1 0 15168 0 -1 14364
box -48 -56 240 834
use sg13g2_fill_2  FILLER_17_163
timestamp 1746816402
transform 1 0 16224 0 -1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_17_165
timestamp 1746816402
transform 1 0 16416 0 -1 14364
box -48 -56 144 834
use sg13g2_fill_1  FILLER_17_195
timestamp 1746816402
transform 1 0 19296 0 -1 14364
box -48 -56 144 834
use sg13g2_fill_1  FILLER_17_245
timestamp 1746816402
transform 1 0 24096 0 -1 14364
box -48 -56 144 834
use sg13g2_fill_1  FILLER_17_272
timestamp 1746816402
transform 1 0 26688 0 -1 14364
box -48 -56 144 834
use sg13g2_fill_1  FILLER_17_286
timestamp 1746816402
transform 1 0 28032 0 -1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_17_313
timestamp 1746816402
transform 1 0 30624 0 -1 14364
box -48 -56 240 834
use sg13g2_fill_2  FILLER_17_319
timestamp 1746816402
transform 1 0 31200 0 -1 14364
box -48 -56 240 834
use sg13g2_decap_8  FILLER_18_0
timestamp 1746816402
transform 1 0 576 0 1 14364
box -48 -56 720 834
use sg13g2_decap_4  FILLER_18_19
timestamp 1746816402
transform 1 0 2400 0 1 14364
box -48 -56 432 834
use sg13g2_fill_2  FILLER_18_23
timestamp 1746816402
transform 1 0 2784 0 1 14364
box -48 -56 240 834
use sg13g2_decap_4  FILLER_18_30
timestamp 1746816402
transform 1 0 3456 0 1 14364
box -48 -56 432 834
use sg13g2_fill_1  FILLER_18_39
timestamp 1746816402
transform 1 0 4320 0 1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_18_53
timestamp 1746816402
transform 1 0 5664 0 1 14364
box -48 -56 240 834
use sg13g2_decap_4  FILLER_18_63
timestamp 1746816402
transform 1 0 6624 0 1 14364
box -48 -56 432 834
use sg13g2_fill_2  FILLER_18_88
timestamp 1746816402
transform 1 0 9024 0 1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_18_90
timestamp 1746816402
transform 1 0 9216 0 1 14364
box -48 -56 144 834
use sg13g2_decap_4  FILLER_18_109
timestamp 1746816402
transform 1 0 11040 0 1 14364
box -48 -56 432 834
use sg13g2_fill_1  FILLER_18_113
timestamp 1746816402
transform 1 0 11424 0 1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_18_136
timestamp 1746816402
transform 1 0 13632 0 1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_18_146
timestamp 1746816402
transform 1 0 14592 0 1 14364
box -48 -56 144 834
use sg13g2_decap_4  FILLER_18_156
timestamp 1746816402
transform 1 0 15552 0 1 14364
box -48 -56 432 834
use sg13g2_decap_8  FILLER_18_173
timestamp 1746816402
transform 1 0 17184 0 1 14364
box -48 -56 720 834
use sg13g2_fill_2  FILLER_18_180
timestamp 1746816402
transform 1 0 17856 0 1 14364
box -48 -56 240 834
use sg13g2_fill_2  FILLER_18_210
timestamp 1746816402
transform 1 0 20736 0 1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_18_212
timestamp 1746816402
transform 1 0 20928 0 1 14364
box -48 -56 144 834
use sg13g2_fill_1  FILLER_18_226
timestamp 1746816402
transform 1 0 22272 0 1 14364
box -48 -56 144 834
use sg13g2_fill_1  FILLER_18_251
timestamp 1746816402
transform 1 0 24672 0 1 14364
box -48 -56 144 834
use sg13g2_fill_1  FILLER_18_285
timestamp 1746816402
transform 1 0 27936 0 1 14364
box -48 -56 144 834
use sg13g2_fill_1  FILLER_18_320
timestamp 1746816402
transform 1 0 31296 0 1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_19_0
timestamp 1746816402
transform 1 0 576 0 -1 15876
box -48 -56 720 834
use sg13g2_fill_1  FILLER_19_7
timestamp 1746816402
transform 1 0 1248 0 -1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_19_16
timestamp 1746816402
transform 1 0 2112 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_19_25
timestamp 1746816402
transform 1 0 2976 0 -1 15876
box -48 -56 144 834
use sg13g2_decap_4  FILLER_19_55
timestamp 1746816402
transform 1 0 5856 0 -1 15876
box -48 -56 432 834
use sg13g2_fill_1  FILLER_19_72
timestamp 1746816402
transform 1 0 7488 0 -1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_19_79
timestamp 1746816402
transform 1 0 8160 0 -1 15876
box -48 -56 144 834
use sg13g2_decap_4  FILLER_19_84
timestamp 1746816402
transform 1 0 8640 0 -1 15876
box -48 -56 432 834
use sg13g2_fill_2  FILLER_19_92
timestamp 1746816402
transform 1 0 9408 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_19_104
timestamp 1746816402
transform 1 0 10560 0 -1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_19_119
timestamp 1746816402
transform 1 0 12000 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_2  FILLER_19_126
timestamp 1746816402
transform 1 0 12672 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_2  FILLER_19_209
timestamp 1746816402
transform 1 0 20640 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_2  FILLER_19_254
timestamp 1746816402
transform 1 0 24960 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_19_277
timestamp 1746816402
transform 1 0 27168 0 -1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_20_0
timestamp 1746816402
transform 1 0 576 0 1 15876
box -48 -56 720 834
use sg13g2_fill_1  FILLER_20_7
timestamp 1746816402
transform 1 0 1248 0 1 15876
box -48 -56 144 834
use sg13g2_decap_4  FILLER_20_43
timestamp 1746816402
transform 1 0 4704 0 1 15876
box -48 -56 432 834
use sg13g2_fill_1  FILLER_20_47
timestamp 1746816402
transform 1 0 5088 0 1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_20_61
timestamp 1746816402
transform 1 0 6432 0 1 15876
box -48 -56 240 834
use sg13g2_fill_2  FILLER_20_107
timestamp 1746816402
transform 1 0 10848 0 1 15876
box -48 -56 240 834
use sg13g2_decap_4  FILLER_20_118
timestamp 1746816402
transform 1 0 11904 0 1 15876
box -48 -56 432 834
use sg13g2_fill_2  FILLER_20_122
timestamp 1746816402
transform 1 0 12288 0 1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_20_129
timestamp 1746816402
transform 1 0 12960 0 1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_20_140
timestamp 1746816402
transform 1 0 14016 0 1 15876
box -48 -56 240 834
use sg13g2_fill_2  FILLER_20_147
timestamp 1746816402
transform 1 0 14688 0 1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_20_161
timestamp 1746816402
transform 1 0 16032 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_178
timestamp 1746816402
transform 1 0 17664 0 1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_20_184
timestamp 1746816402
transform 1 0 18240 0 1 15876
box -48 -56 240 834
use sg13g2_fill_2  FILLER_20_199
timestamp 1746816402
transform 1 0 19680 0 1 15876
box -48 -56 240 834
use sg13g2_fill_2  FILLER_20_236
timestamp 1746816402
transform 1 0 23232 0 1 15876
box -48 -56 240 834
use sg13g2_fill_2  FILLER_20_248
timestamp 1746816402
transform 1 0 24384 0 1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_20_250
timestamp 1746816402
transform 1 0 24576 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_270
timestamp 1746816402
transform 1 0 26496 0 1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_20_277
timestamp 1746816402
transform 1 0 27168 0 1 15876
box -48 -56 240 834
use sg13g2_decap_8  FILLER_21_0
timestamp 1746816402
transform 1 0 576 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_7
timestamp 1746816402
transform 1 0 1248 0 -1 17388
box -48 -56 720 834
use sg13g2_fill_2  FILLER_21_14
timestamp 1746816402
transform 1 0 1920 0 -1 17388
box -48 -56 240 834
use sg13g2_decap_4  FILLER_21_21
timestamp 1746816402
transform 1 0 2592 0 -1 17388
box -48 -56 432 834
use sg13g2_fill_1  FILLER_21_66
timestamp 1746816402
transform 1 0 6912 0 -1 17388
box -48 -56 144 834
use sg13g2_fill_1  FILLER_21_75
timestamp 1746816402
transform 1 0 7776 0 -1 17388
box -48 -56 144 834
use sg13g2_fill_1  FILLER_21_92
timestamp 1746816402
transform 1 0 9408 0 -1 17388
box -48 -56 144 834
use sg13g2_fill_2  FILLER_21_99
timestamp 1746816402
transform 1 0 10080 0 -1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_21_101
timestamp 1746816402
transform 1 0 10272 0 -1 17388
box -48 -56 144 834
use sg13g2_fill_2  FILLER_21_146
timestamp 1746816402
transform 1 0 14592 0 -1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_21_148
timestamp 1746816402
transform 1 0 14784 0 -1 17388
box -48 -56 144 834
use sg13g2_fill_2  FILLER_21_201
timestamp 1746816402
transform 1 0 19872 0 -1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_21_203
timestamp 1746816402
transform 1 0 20064 0 -1 17388
box -48 -56 144 834
use sg13g2_fill_2  FILLER_21_226
timestamp 1746816402
transform 1 0 22272 0 -1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_21_260
timestamp 1746816402
transform 1 0 25536 0 -1 17388
box -48 -56 144 834
use sg13g2_fill_1  FILLER_21_320
timestamp 1746816402
transform 1 0 31296 0 -1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_22_0
timestamp 1746816402
transform 1 0 576 0 1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_22_7
timestamp 1746816402
transform 1 0 1248 0 1 17388
box -48 -56 432 834
use sg13g2_fill_1  FILLER_22_11
timestamp 1746816402
transform 1 0 1632 0 1 17388
box -48 -56 144 834
use sg13g2_fill_1  FILLER_22_16
timestamp 1746816402
transform 1 0 2112 0 1 17388
box -48 -56 144 834
use sg13g2_fill_2  FILLER_22_61
timestamp 1746816402
transform 1 0 6432 0 1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_22_63
timestamp 1746816402
transform 1 0 6624 0 1 17388
box -48 -56 144 834
use sg13g2_fill_1  FILLER_22_80
timestamp 1746816402
transform 1 0 8256 0 1 17388
box -48 -56 144 834
use sg13g2_fill_2  FILLER_22_111
timestamp 1746816402
transform 1 0 11232 0 1 17388
box -48 -56 240 834
use sg13g2_fill_2  FILLER_22_153
timestamp 1746816402
transform 1 0 15264 0 1 17388
box -48 -56 240 834
use sg13g2_fill_2  FILLER_22_199
timestamp 1746816402
transform 1 0 19680 0 1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_22_201
timestamp 1746816402
transform 1 0 19872 0 1 17388
box -48 -56 144 834
use sg13g2_fill_2  FILLER_22_227
timestamp 1746816402
transform 1 0 22368 0 1 17388
box -48 -56 240 834
use sg13g2_fill_2  FILLER_22_257
timestamp 1746816402
transform 1 0 25248 0 1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_22_259
timestamp 1746816402
transform 1 0 25440 0 1 17388
box -48 -56 144 834
use sg13g2_fill_2  FILLER_22_318
timestamp 1746816402
transform 1 0 31104 0 1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_22_320
timestamp 1746816402
transform 1 0 31296 0 1 17388
box -48 -56 144 834
use sg13g2_fill_1  FILLER_23_0
timestamp 1746816402
transform 1 0 576 0 -1 18900
box -48 -56 144 834
use sg13g2_fill_1  FILLER_23_41
timestamp 1746816402
transform 1 0 4512 0 -1 18900
box -48 -56 144 834
use sg13g2_fill_2  FILLER_23_50
timestamp 1746816402
transform 1 0 5376 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_23_52
timestamp 1746816402
transform 1 0 5568 0 -1 18900
box -48 -56 144 834
use sg13g2_fill_1  FILLER_23_85
timestamp 1746816402
transform 1 0 8736 0 -1 18900
box -48 -56 144 834
use sg13g2_fill_2  FILLER_23_96
timestamp 1746816402
transform 1 0 9792 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_2  FILLER_23_118
timestamp 1746816402
transform 1 0 11904 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_2  FILLER_23_130
timestamp 1746816402
transform 1 0 13056 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_23_142
timestamp 1746816402
transform 1 0 14208 0 -1 18900
box -48 -56 144 834
use sg13g2_fill_2  FILLER_23_217
timestamp 1746816402
transform 1 0 21408 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_23_219
timestamp 1746816402
transform 1 0 21600 0 -1 18900
box -48 -56 144 834
use sg13g2_fill_2  FILLER_23_236
timestamp 1746816402
transform 1 0 23232 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_2  FILLER_23_271
timestamp 1746816402
transform 1 0 26592 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_2  FILLER_23_319
timestamp 1746816402
transform 1 0 31200 0 -1 18900
box -48 -56 240 834
use sg13g2_decap_4  FILLER_24_4
timestamp 1746816402
transform 1 0 960 0 1 18900
box -48 -56 432 834
use sg13g2_fill_2  FILLER_24_21
timestamp 1746816402
transform 1 0 2592 0 1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_24_23
timestamp 1746816402
transform 1 0 2784 0 1 18900
box -48 -56 144 834
use sg13g2_fill_2  FILLER_24_44
timestamp 1746816402
transform 1 0 4800 0 1 18900
box -48 -56 240 834
use sg13g2_decap_4  FILLER_24_70
timestamp 1746816402
transform 1 0 7296 0 1 18900
box -48 -56 432 834
use sg13g2_decap_4  FILLER_24_79
timestamp 1746816402
transform 1 0 8160 0 1 18900
box -48 -56 432 834
use sg13g2_fill_1  FILLER_24_83
timestamp 1746816402
transform 1 0 8544 0 1 18900
box -48 -56 144 834
use sg13g2_decap_4  FILLER_24_104
timestamp 1746816402
transform 1 0 10560 0 1 18900
box -48 -56 432 834
use sg13g2_fill_2  FILLER_24_113
timestamp 1746816402
transform 1 0 11424 0 1 18900
box -48 -56 240 834
use sg13g2_decap_4  FILLER_24_120
timestamp 1746816402
transform 1 0 12096 0 1 18900
box -48 -56 432 834
use sg13g2_fill_1  FILLER_24_124
timestamp 1746816402
transform 1 0 12480 0 1 18900
box -48 -56 144 834
use sg13g2_fill_2  FILLER_24_177
timestamp 1746816402
transform 1 0 17568 0 1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_24_179
timestamp 1746816402
transform 1 0 17760 0 1 18900
box -48 -56 144 834
use sg13g2_fill_2  FILLER_24_191
timestamp 1746816402
transform 1 0 18912 0 1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_24_193
timestamp 1746816402
transform 1 0 19104 0 1 18900
box -48 -56 144 834
use sg13g2_fill_2  FILLER_24_203
timestamp 1746816402
transform 1 0 20064 0 1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_24_205
timestamp 1746816402
transform 1 0 20256 0 1 18900
box -48 -56 144 834
use sg13g2_fill_1  FILLER_24_219
timestamp 1746816402
transform 1 0 21600 0 1 18900
box -48 -56 144 834
use sg13g2_fill_2  FILLER_24_239
timestamp 1746816402
transform 1 0 23520 0 1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_24_241
timestamp 1746816402
transform 1 0 23712 0 1 18900
box -48 -56 144 834
use sg13g2_fill_2  FILLER_24_248
timestamp 1746816402
transform 1 0 24384 0 1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_24_274
timestamp 1746816402
transform 1 0 26880 0 1 18900
box -48 -56 144 834
use sg13g2_fill_2  FILLER_25_13
timestamp 1746816402
transform 1 0 1824 0 -1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_25_15
timestamp 1746816402
transform 1 0 2016 0 -1 20412
box -48 -56 144 834
use sg13g2_fill_1  FILLER_25_26
timestamp 1746816402
transform 1 0 3072 0 -1 20412
box -48 -56 144 834
use sg13g2_fill_2  FILLER_25_40
timestamp 1746816402
transform 1 0 4416 0 -1 20412
box -48 -56 240 834
use sg13g2_fill_2  FILLER_25_72
timestamp 1746816402
transform 1 0 7488 0 -1 20412
box -48 -56 240 834
use sg13g2_fill_2  FILLER_25_88
timestamp 1746816402
transform 1 0 9024 0 -1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_25_90
timestamp 1746816402
transform 1 0 9216 0 -1 20412
box -48 -56 144 834
use sg13g2_fill_1  FILLER_25_146
timestamp 1746816402
transform 1 0 14592 0 -1 20412
box -48 -56 144 834
use sg13g2_fill_1  FILLER_25_152
timestamp 1746816402
transform 1 0 15168 0 -1 20412
box -48 -56 144 834
use sg13g2_fill_1  FILLER_25_165
timestamp 1746816402
transform 1 0 16416 0 -1 20412
box -48 -56 144 834
use sg13g2_fill_1  FILLER_25_181
timestamp 1746816402
transform 1 0 17952 0 -1 20412
box -48 -56 144 834
use sg13g2_fill_1  FILLER_25_196
timestamp 1746816402
transform 1 0 19392 0 -1 20412
box -48 -56 144 834
use sg13g2_fill_1  FILLER_25_207
timestamp 1746816402
transform 1 0 20448 0 -1 20412
box -48 -56 144 834
use sg13g2_fill_2  FILLER_25_244
timestamp 1746816402
transform 1 0 24000 0 -1 20412
box -48 -56 240 834
use sg13g2_fill_2  FILLER_25_261
timestamp 1746816402
transform 1 0 25632 0 -1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_26_4
timestamp 1746816402
transform 1 0 960 0 1 20412
box -48 -56 144 834
use sg13g2_fill_2  FILLER_26_41
timestamp 1746816402
transform 1 0 4512 0 1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_26_64
timestamp 1746816402
transform 1 0 6720 0 1 20412
box -48 -56 144 834
use sg13g2_fill_1  FILLER_26_92
timestamp 1746816402
transform 1 0 9408 0 1 20412
box -48 -56 144 834
use sg13g2_fill_2  FILLER_26_102
timestamp 1746816402
transform 1 0 10368 0 1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_26_104
timestamp 1746816402
transform 1 0 10560 0 1 20412
box -48 -56 144 834
use sg13g2_fill_1  FILLER_26_177
timestamp 1746816402
transform 1 0 17568 0 1 20412
box -48 -56 144 834
use sg13g2_fill_2  FILLER_26_203
timestamp 1746816402
transform 1 0 20064 0 1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_26_205
timestamp 1746816402
transform 1 0 20256 0 1 20412
box -48 -56 144 834
use sg13g2_fill_1  FILLER_26_214
timestamp 1746816402
transform 1 0 21120 0 1 20412
box -48 -56 144 834
use sg13g2_fill_1  FILLER_26_223
timestamp 1746816402
transform 1 0 21984 0 1 20412
box -48 -56 144 834
use sg13g2_fill_2  FILLER_26_241
timestamp 1746816402
transform 1 0 23712 0 1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_26_270
timestamp 1746816402
transform 1 0 26496 0 1 20412
box -48 -56 144 834
use sg13g2_fill_1  FILLER_27_4
timestamp 1746816402
transform 1 0 960 0 -1 21924
box -48 -56 144 834
use sg13g2_fill_2  FILLER_27_33
timestamp 1746816402
transform 1 0 3744 0 -1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_27_69
timestamp 1746816402
transform 1 0 7200 0 -1 21924
box -48 -56 144 834
use sg13g2_fill_2  FILLER_27_88
timestamp 1746816402
transform 1 0 9024 0 -1 21924
box -48 -56 240 834
use sg13g2_fill_2  FILLER_27_195
timestamp 1746816402
transform 1 0 19296 0 -1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_27_197
timestamp 1746816402
transform 1 0 19488 0 -1 21924
box -48 -56 144 834
use sg13g2_fill_1  FILLER_27_227
timestamp 1746816402
transform 1 0 22368 0 -1 21924
box -48 -56 144 834
use sg13g2_fill_1  FILLER_27_242
timestamp 1746816402
transform 1 0 23808 0 -1 21924
box -48 -56 144 834
use sg13g2_fill_1  FILLER_27_284
timestamp 1746816402
transform 1 0 27840 0 -1 21924
box -48 -56 144 834
use sg13g2_fill_2  FILLER_28_23
timestamp 1746816402
transform 1 0 2784 0 1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_28_25
timestamp 1746816402
transform 1 0 2976 0 1 21924
box -48 -56 144 834
use sg13g2_fill_2  FILLER_28_41
timestamp 1746816402
transform 1 0 4512 0 1 21924
box -48 -56 240 834
use sg13g2_fill_2  FILLER_28_66
timestamp 1746816402
transform 1 0 6912 0 1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_28_68
timestamp 1746816402
transform 1 0 7104 0 1 21924
box -48 -56 144 834
use sg13g2_fill_2  FILLER_28_160
timestamp 1746816402
transform 1 0 15936 0 1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_28_175
timestamp 1746816402
transform 1 0 17376 0 1 21924
box -48 -56 144 834
use sg13g2_fill_2  FILLER_28_201
timestamp 1746816402
transform 1 0 19872 0 1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_28_211
timestamp 1746816402
transform 1 0 20832 0 1 21924
box -48 -56 144 834
use sg13g2_fill_2  FILLER_28_220
timestamp 1746816402
transform 1 0 21696 0 1 21924
box -48 -56 240 834
use sg13g2_fill_2  FILLER_28_255
timestamp 1746816402
transform 1 0 25056 0 1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_28_257
timestamp 1746816402
transform 1 0 25248 0 1 21924
box -48 -56 144 834
use sg13g2_fill_1  FILLER_28_294
timestamp 1746816402
transform 1 0 28800 0 1 21924
box -48 -56 144 834
use sg13g2_fill_2  FILLER_29_0
timestamp 1746816402
transform 1 0 576 0 -1 23436
box -48 -56 240 834
use sg13g2_fill_2  FILLER_29_39
timestamp 1746816402
transform 1 0 4320 0 -1 23436
box -48 -56 240 834
use sg13g2_fill_2  FILLER_29_69
timestamp 1746816402
transform 1 0 7200 0 -1 23436
box -48 -56 240 834
use sg13g2_fill_2  FILLER_29_97
timestamp 1746816402
transform 1 0 9888 0 -1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_29_99
timestamp 1746816402
transform 1 0 10080 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_29_115
timestamp 1746816402
transform 1 0 11616 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_29_121
timestamp 1746816402
transform 1 0 12192 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_29_146
timestamp 1746816402
transform 1 0 14592 0 -1 23436
box -48 -56 240 834
use sg13g2_fill_2  FILLER_29_164
timestamp 1746816402
transform 1 0 16320 0 -1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_29_192
timestamp 1746816402
transform 1 0 19008 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_29_197
timestamp 1746816402
transform 1 0 19488 0 -1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_29_199
timestamp 1746816402
transform 1 0 19680 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_29_258
timestamp 1746816402
transform 1 0 25344 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_29_267
timestamp 1746816402
transform 1 0 26208 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_29_319
timestamp 1746816402
transform 1 0 31200 0 -1 23436
box -48 -56 240 834
use sg13g2_fill_2  FILLER_30_26
timestamp 1746816402
transform 1 0 3072 0 1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_30_28
timestamp 1746816402
transform 1 0 3264 0 1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_30_64
timestamp 1746816402
transform 1 0 6720 0 1 23436
box -48 -56 240 834
use sg13g2_fill_2  FILLER_30_71
timestamp 1746816402
transform 1 0 7392 0 1 23436
box -48 -56 240 834
use sg13g2_fill_2  FILLER_30_113
timestamp 1746816402
transform 1 0 11424 0 1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_30_124
timestamp 1746816402
transform 1 0 12480 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_148
timestamp 1746816402
transform 1 0 14784 0 1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_30_216
timestamp 1746816402
transform 1 0 21312 0 1 23436
box -48 -56 240 834
use sg13g2_fill_2  FILLER_30_267
timestamp 1746816402
transform 1 0 26208 0 1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_31_0
timestamp 1746816402
transform 1 0 576 0 -1 24948
box -48 -56 144 834
use sg13g2_fill_1  FILLER_31_48
timestamp 1746816402
transform 1 0 5184 0 -1 24948
box -48 -56 144 834
use sg13g2_fill_1  FILLER_31_83
timestamp 1746816402
transform 1 0 8544 0 -1 24948
box -48 -56 144 834
use sg13g2_fill_2  FILLER_31_94
timestamp 1746816402
transform 1 0 9600 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_2  FILLER_31_139
timestamp 1746816402
transform 1 0 13920 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_31_181
timestamp 1746816402
transform 1 0 17952 0 -1 24948
box -48 -56 144 834
use sg13g2_fill_2  FILLER_31_191
timestamp 1746816402
transform 1 0 18912 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_31_198
timestamp 1746816402
transform 1 0 19584 0 -1 24948
box -48 -56 144 834
use sg13g2_fill_1  FILLER_32_82
timestamp 1746816402
transform 1 0 8448 0 1 24948
box -48 -56 144 834
use sg13g2_fill_1  FILLER_32_95
timestamp 1746816402
transform 1 0 9696 0 1 24948
box -48 -56 144 834
use sg13g2_fill_1  FILLER_32_125
timestamp 1746816402
transform 1 0 12576 0 1 24948
box -48 -56 144 834
use sg13g2_fill_1  FILLER_32_190
timestamp 1746816402
transform 1 0 18816 0 1 24948
box -48 -56 144 834
use sg13g2_fill_1  FILLER_32_253
timestamp 1746816402
transform 1 0 24864 0 1 24948
box -48 -56 144 834
use sg13g2_fill_1  FILLER_32_285
timestamp 1746816402
transform 1 0 27936 0 1 24948
box -48 -56 144 834
use sg13g2_fill_2  FILLER_32_318
timestamp 1746816402
transform 1 0 31104 0 1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_32_320
timestamp 1746816402
transform 1 0 31296 0 1 24948
box -48 -56 144 834
use sg13g2_fill_2  FILLER_33_4
timestamp 1746816402
transform 1 0 960 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_33_6
timestamp 1746816402
transform 1 0 1152 0 -1 26460
box -48 -56 144 834
use sg13g2_fill_1  FILLER_33_277
timestamp 1746816402
transform 1 0 27168 0 -1 26460
box -48 -56 144 834
use sg13g2_fill_2  FILLER_34_0
timestamp 1746816402
transform 1 0 576 0 1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_34_2
timestamp 1746816402
transform 1 0 768 0 1 26460
box -48 -56 144 834
use sg13g2_fill_2  FILLER_34_70
timestamp 1746816402
transform 1 0 7296 0 1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_34_95
timestamp 1746816402
transform 1 0 9696 0 1 26460
box -48 -56 144 834
use sg13g2_fill_1  FILLER_34_217
timestamp 1746816402
transform 1 0 21408 0 1 26460
box -48 -56 144 834
use sg13g2_fill_2  FILLER_34_286
timestamp 1746816402
transform 1 0 28032 0 1 26460
box -48 -56 240 834
use sg13g2_fill_2  FILLER_34_319
timestamp 1746816402
transform 1 0 31200 0 1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_35_119
timestamp 1746816402
transform 1 0 12000 0 -1 27972
box -48 -56 144 834
use sg13g2_fill_2  FILLER_35_219
timestamp 1746816402
transform 1 0 21600 0 -1 27972
box -48 -56 240 834
use sg13g2_fill_1  FILLER_35_221
timestamp 1746816402
transform 1 0 21792 0 -1 27972
box -48 -56 144 834
use sg13g2_fill_2  FILLER_35_319
timestamp 1746816402
transform 1 0 31200 0 -1 27972
box -48 -56 240 834
use sg13g2_dlygate4sd3_1  hold1
timestamp 1746816402
transform 1 0 22080 0 1 20412
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold2
timestamp 1746816402
transform -1 0 26304 0 1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold3
timestamp 1746816402
transform -1 0 27168 0 1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold4
timestamp 1746816402
transform -1 0 4512 0 -1 27972
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold5
timestamp 1746816402
transform 1 0 8832 0 1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold6
timestamp 1746816402
transform 1 0 11424 0 -1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold7
timestamp 1746816402
transform -1 0 15936 0 1 24948
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold8
timestamp 1746816402
transform -1 0 19680 0 -1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold9
timestamp 1746816402
transform 1 0 15744 0 1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold10
timestamp 1746816402
transform 1 0 18912 0 1 24948
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold11
timestamp 1746816402
transform -1 0 17472 0 -1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold12
timestamp 1746816402
transform 1 0 13728 0 1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold13
timestamp 1746816402
transform -1 0 25440 0 1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold14
timestamp 1746816402
transform -1 0 23712 0 1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold15
timestamp 1746816402
transform -1 0 24576 0 1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold16
timestamp 1746816402
transform -1 0 22848 0 1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold17
timestamp 1746816402
transform 1 0 28800 0 -1 17388
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold18
timestamp 1746816402
transform -1 0 29472 0 -1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold19
timestamp 1746816402
transform 1 0 29472 0 -1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold20
timestamp 1746816402
transform -1 0 29472 0 1 9828
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold21
timestamp 1746816402
transform 1 0 27456 0 1 8316
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold22
timestamp 1746816402
transform -1 0 29184 0 1 8316
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold23
timestamp 1746816402
transform -1 0 26880 0 1 8316
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold24
timestamp 1746816402
transform 1 0 2496 0 -1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold25
timestamp 1746816402
transform -1 0 4224 0 1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold26
timestamp 1746816402
transform -1 0 24864 0 1 24948
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold27
timestamp 1746816402
transform 1 0 21408 0 -1 24948
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold28
timestamp 1746816402
transform -1 0 12480 0 1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold29
timestamp 1746816402
transform 1 0 28032 0 1 18900
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold30
timestamp 1746816402
transform 1 0 28032 0 -1 20412
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold31
timestamp 1746816402
transform -1 0 22944 0 -1 8316
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold32
timestamp 1746816402
transform -1 0 21888 0 -1 8316
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold33
timestamp 1746816402
transform 1 0 12288 0 -1 24948
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold34
timestamp 1746816402
transform 1 0 5760 0 1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold35
timestamp 1746816402
transform 1 0 7584 0 1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold36
timestamp 1746816402
transform -1 0 28896 0 -1 15876
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold37
timestamp 1746816402
transform 1 0 28896 0 -1 15876
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold38
timestamp 1746816402
transform -1 0 21408 0 1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold39
timestamp 1746816402
transform 1 0 18240 0 -1 27972
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold40
timestamp 1746816402
transform -1 0 31200 0 -1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold41
timestamp 1746816402
transform -1 0 28896 0 1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold42
timestamp 1746816402
transform 1 0 1920 0 -1 21924
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold43
timestamp 1746816402
transform -1 0 4032 0 -1 18900
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold44
timestamp 1746816402
transform -1 0 29760 0 1 20412
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold45
timestamp 1746816402
transform -1 0 28992 0 -1 14364
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold46
timestamp 1746816402
transform -1 0 23712 0 -1 6804
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold47
timestamp 1746816402
transform -1 0 30624 0 1 20412
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold48
timestamp 1746816402
transform -1 0 18240 0 1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold49
timestamp 1746816402
transform -1 0 25248 0 1 12852
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold50
timestamp 1746816402
transform 1 0 5088 0 -1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold51
timestamp 1746816402
transform 1 0 4320 0 -1 24948
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold52
timestamp 1746816402
transform 1 0 3264 0 -1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold53
timestamp 1746816402
transform -1 0 29760 0 1 24948
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold54
timestamp 1746816402
transform 1 0 28032 0 -1 24948
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold55
timestamp 1746816402
transform 1 0 20448 0 -1 14364
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold56
timestamp 1746816402
transform 1 0 22368 0 1 14364
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold57
timestamp 1746816402
transform -1 0 30240 0 -1 27972
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold58
timestamp 1746816402
transform -1 0 11328 0 -1 5292
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold59
timestamp 1746816402
transform -1 0 8256 0 1 5292
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold60
timestamp 1746816402
transform 1 0 4992 0 1 5292
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold61
timestamp 1746816402
transform -1 0 12480 0 1 20412
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold62
timestamp 1746816402
transform -1 0 28800 0 -1 17388
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold63
timestamp 1746816402
transform 1 0 4992 0 1 6804
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold64
timestamp 1746816402
transform -1 0 3744 0 1 5292
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold65
timestamp 1746816402
transform -1 0 28896 0 1 24948
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold66
timestamp 1746816402
transform -1 0 30624 0 1 24948
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold67
timestamp 1746816402
transform 1 0 22368 0 1 12852
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold68
timestamp 1746816402
transform -1 0 28896 0 -1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold69
timestamp 1746816402
transform -1 0 28032 0 1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold70
timestamp 1746816402
transform -1 0 27648 0 1 17388
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold71
timestamp 1746816402
transform -1 0 21792 0 1 17388
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold72
timestamp 1746816402
transform 1 0 7392 0 -1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold73
timestamp 1746816402
transform 1 0 19488 0 1 5292
box -48 -56 912 834
use sg13g2_buf_1  input1
timestamp 1746816402
transform -1 0 31200 0 -1 14364
box -48 -56 432 834
use sg13g2_buf_1  input2
timestamp 1746816402
transform 1 0 8544 0 1 24948
box -48 -56 432 834
use sg13g2_buf_2  input3
timestamp 1746816402
transform -1 0 31104 0 1 17388
box -48 -56 528 834
use sg13g2_buf_2  input4
timestamp 1746816402
transform -1 0 30624 0 1 17388
box -48 -56 528 834
use sg13g2_buf_2  input5
timestamp 1746816402
transform -1 0 31200 0 -1 18900
box -48 -56 528 834
use sg13g2_buf_2  input6
timestamp 1746816402
transform 1 0 20928 0 -1 24948
box -48 -56 528 834
use sg13g2_buf_2  input7
timestamp 1746816402
transform -1 0 31200 0 -1 27972
box -48 -56 528 834
use sg13g2_buf_2  input8
timestamp 1746816402
transform -1 0 25824 0 -1 24948
box -48 -56 528 834
use sg13g2_buf_2  input9
timestamp 1746816402
transform -1 0 26688 0 -1 26460
box -48 -56 528 834
use sg13g2_buf_2  input10
timestamp 1746816402
transform -1 0 25440 0 -1 26460
box -48 -56 528 834
use sg13g2_buf_8  rgb_buffers\[0\]
timestamp 1746816402
transform -1 0 9888 0 -1 23436
box -48 -56 1296 834
use sg13g2_buf_8  rgb_buffers\[1\]
timestamp 1746816402
transform -1 0 7200 0 -1 23436
box -48 -56 1296 834
use sg13g2_buf_8  rgb_buffers\[2\]
timestamp 1746816402
transform -1 0 1824 0 -1 20412
box -48 -56 1296 834
use sg13g2_buf_8  rgb_buffers\[3\]
timestamp 1746816402
transform -1 0 1824 0 1 21924
box -48 -56 1296 834
use sg13g2_buf_2  rgb_buffers\[4\]
timestamp 1746816402
transform 1 0 3360 0 -1 23436
box -48 -56 528 834
use sg13g2_buf_1  rgb_buffers\[5\]
timestamp 1746816402
transform -1 0 4032 0 -1 20412
box -48 -56 432 834
use sg13g2_buf_2  rgb_buffers\[6\]
timestamp 1746816402
transform 1 0 11904 0 1 21924
box -48 -56 528 834
use sg13g2_buf_2  rgb_buffers\[7\]
timestamp 1746816402
transform 1 0 16512 0 -1 21924
box -48 -56 528 834
use sg13g2_buf_8  rgb_buffers\[8\]
timestamp 1746816402
transform -1 0 9888 0 1 21924
box -48 -56 1296 834
use sg13g2_buf_2  rgb_buffers\[9\]
timestamp 1746816402
transform 1 0 6240 0 1 23436
box -48 -56 528 834
use sg13g2_buf_1  rgb_buffers\[10\]
timestamp 1746816402
transform -1 0 960 0 1 18900
box -48 -56 432 834
use sg13g2_buf_1  rgb_buffers\[11\]
timestamp 1746816402
transform -1 0 960 0 -1 26460
box -48 -56 432 834
use sg13g2_buf_1  rgb_buffers\[12\]
timestamp 1746816402
transform -1 0 1344 0 1 24948
box -48 -56 432 834
use sg13g2_buf_1  rgb_buffers\[13\]
timestamp 1746816402
transform -1 0 4032 0 1 20412
box -48 -56 432 834
use sg13g2_buf_8  rgb_buffers\[14\]
timestamp 1746816402
transform -1 0 13632 0 1 21924
box -48 -56 1296 834
use sg13g2_buf_8  rgb_buffers\[15\]
timestamp 1746816402
transform -1 0 17376 0 1 21924
box -48 -56 1296 834
use sg13g2_buf_1  rgb_buffers\[16\]
timestamp 1746816402
transform -1 0 9696 0 1 24948
box -48 -56 432 834
use sg13g2_buf_1  rgb_buffers\[17\]
timestamp 1746816402
transform -1 0 5472 0 1 21924
box -48 -56 432 834
use sg13g2_buf_1  rgb_buffers\[18\]
timestamp 1746816402
transform -1 0 960 0 1 20412
box -48 -56 432 834
use sg13g2_buf_1  rgb_buffers\[19\]
timestamp 1746816402
transform -1 0 960 0 -1 21924
box -48 -56 432 834
use sg13g2_buf_1  rgb_buffers\[20\]
timestamp 1746816402
transform -1 0 1440 0 -1 24948
box -48 -56 432 834
use sg13g2_buf_1  rgb_buffers\[21\]
timestamp 1746816402
transform -1 0 4416 0 -1 20412
box -48 -56 432 834
use sg13g2_buf_8  rgb_buffers\[22\]
timestamp 1746816402
transform -1 0 15456 0 1 21924
box -48 -56 1296 834
use sg13g2_buf_8  rgb_buffers\[23\]
timestamp 1746816402
transform -1 0 17760 0 -1 23436
box -48 -56 1296 834
<< labels >>
flabel metal5 s 27638 712 28078 28016 0 FreeSans 3200 90 0 0 VGND
port 1 nsew
flabel metal5 s 19864 712 20304 28016 0 FreeSans 3200 90 0 0 VGND
port 1 nsew
flabel metal5 s 12090 712 12530 28016 0 FreeSans 3200 90 0 0 VGND
port 1 nsew
flabel metal5 s 4316 712 4756 28016 0 FreeSans 3200 90 0 0 VGND
port 1 nsew
flabel metal5 s 26398 712 26838 28016 0 FreeSans 3200 90 0 0 VPWR
port 2 nsew
flabel metal5 s 18624 712 19064 28016 0 FreeSans 3200 90 0 0 VPWR
port 2 nsew
flabel metal5 s 10850 712 11290 28016 0 FreeSans 3200 90 0 0 VPWR
port 2 nsew
flabel metal5 s 3076 712 3516 28016 0 FreeSans 3200 90 0 0 VPWR
port 2 nsew
flabel metal3 s 11576 28600 11656 29000 0 FreeSans 400 90 0 0 b6
port 3 nsew
flabel metal3 s 14648 28600 14728 29000 0 FreeSans 400 90 0 0 b7
port 4 nsew
flabel metal3 s 30008 28600 30088 29000 0 FreeSans 400 90 0 0 clk
port 5 nsew
flabel metal2 s 0 8864 400 8944 0 FreeSans 400 0 0 0 db[0]
port 6 nsew
flabel metal2 s 0 8444 400 8524 0 FreeSans 400 0 0 0 db[1]
port 7 nsew
flabel metal2 s 0 8024 400 8104 0 FreeSans 400 0 0 0 db[2]
port 8 nsew
flabel metal2 s 0 7604 400 7684 0 FreeSans 400 0 0 0 db[3]
port 9 nsew
flabel metal2 s 0 7184 400 7264 0 FreeSans 400 0 0 0 db[4]
port 10 nsew
flabel metal2 s 0 6764 400 6844 0 FreeSans 400 0 0 0 db[5]
port 11 nsew
flabel metal2 s 0 6344 400 6424 0 FreeSans 400 0 0 0 db[6]
port 12 nsew
flabel metal2 s 0 5924 400 6004 0 FreeSans 400 0 0 0 db[7]
port 13 nsew
flabel metal2 s 0 15584 400 15664 0 FreeSans 400 0 0 0 dg[0]
port 14 nsew
flabel metal2 s 0 15164 400 15244 0 FreeSans 400 0 0 0 dg[1]
port 15 nsew
flabel metal2 s 0 14744 400 14824 0 FreeSans 400 0 0 0 dg[2]
port 16 nsew
flabel metal2 s 0 14324 400 14404 0 FreeSans 400 0 0 0 dg[3]
port 17 nsew
flabel metal2 s 0 13904 400 13984 0 FreeSans 400 0 0 0 dg[4]
port 18 nsew
flabel metal2 s 0 13484 400 13564 0 FreeSans 400 0 0 0 dg[5]
port 19 nsew
flabel metal2 s 0 13064 400 13144 0 FreeSans 400 0 0 0 dg[6]
port 20 nsew
flabel metal2 s 0 12644 400 12724 0 FreeSans 400 0 0 0 dg[7]
port 21 nsew
flabel metal2 s 0 22304 400 22384 0 FreeSans 400 0 0 0 dr[0]
port 22 nsew
flabel metal2 s 0 21884 400 21964 0 FreeSans 400 0 0 0 dr[1]
port 23 nsew
flabel metal2 s 0 21464 400 21544 0 FreeSans 400 0 0 0 dr[2]
port 24 nsew
flabel metal2 s 0 21044 400 21124 0 FreeSans 400 0 0 0 dr[3]
port 25 nsew
flabel metal2 s 0 20624 400 20704 0 FreeSans 400 0 0 0 dr[4]
port 26 nsew
flabel metal2 s 0 20204 400 20284 0 FreeSans 400 0 0 0 dr[5]
port 27 nsew
flabel metal2 s 0 19784 400 19864 0 FreeSans 400 0 0 0 dr[6]
port 28 nsew
flabel metal2 s 0 19364 400 19444 0 FreeSans 400 0 0 0 dr[7]
port 29 nsew
flabel metal3 s 30776 28600 30856 29000 0 FreeSans 400 90 0 0 ena
port 30 nsew
flabel metal3 s 12344 28600 12424 29000 0 FreeSans 400 90 0 0 g6
port 31 nsew
flabel metal3 s 15416 28600 15496 29000 0 FreeSans 400 90 0 0 g7
port 32 nsew
flabel metal3 s 9272 28600 9352 29000 0 FreeSans 400 90 0 0 hblank
port 33 nsew
flabel metal3 s 10808 28600 10888 29000 0 FreeSans 400 90 0 0 hsync
port 34 nsew
flabel metal3 s 13112 28600 13192 29000 0 FreeSans 400 90 0 0 r6
port 35 nsew
flabel metal3 s 16184 28600 16264 29000 0 FreeSans 400 90 0 0 r7
port 36 nsew
flabel metal3 s 29240 28600 29320 29000 0 FreeSans 400 90 0 0 rst_n
port 37 nsew
flabel metal3 s 28472 28600 28552 29000 0 FreeSans 400 90 0 0 ui_in[0]
port 38 nsew
flabel metal3 s 27704 28600 27784 29000 0 FreeSans 400 90 0 0 ui_in[1]
port 39 nsew
flabel metal3 s 26936 28600 27016 29000 0 FreeSans 400 90 0 0 ui_in[2]
port 40 nsew
flabel metal3 s 26168 28600 26248 29000 0 FreeSans 400 90 0 0 ui_in[3]
port 41 nsew
flabel metal3 s 25400 28600 25480 29000 0 FreeSans 400 90 0 0 ui_in[4]
port 42 nsew
flabel metal3 s 24632 28600 24712 29000 0 FreeSans 400 90 0 0 ui_in[5]
port 43 nsew
flabel metal3 s 23864 28600 23944 29000 0 FreeSans 400 90 0 0 ui_in[6]
port 44 nsew
flabel metal3 s 23096 28600 23176 29000 0 FreeSans 400 90 0 0 ui_in[7]
port 45 nsew
flabel metal3 s 3896 28600 3976 29000 0 FreeSans 400 90 0 0 uio_oe[0]
port 46 nsew
flabel metal3 s 3128 28600 3208 29000 0 FreeSans 400 90 0 0 uio_oe[1]
port 47 nsew
flabel metal3 s 8504 28600 8584 29000 0 FreeSans 400 90 0 0 uio_out2
port 48 nsew
flabel metal3 s 7736 28600 7816 29000 0 FreeSans 400 90 0 0 uio_out3
port 49 nsew
flabel metal3 s 6968 28600 7048 29000 0 FreeSans 400 90 0 0 uio_out4
port 50 nsew
flabel metal3 s 6200 28600 6280 29000 0 FreeSans 400 90 0 0 uio_out5
port 51 nsew
flabel metal3 s 5432 28600 5512 29000 0 FreeSans 400 90 0 0 uio_out6
port 52 nsew
flabel metal3 s 4664 28600 4744 29000 0 FreeSans 400 90 0 0 uio_out7
port 53 nsew
flabel metal3 s 10040 28600 10120 29000 0 FreeSans 400 90 0 0 vblank
port 54 nsew
flabel metal3 s 13880 28600 13960 29000 0 FreeSans 400 90 0 0 vsync
port 55 nsew
<< properties >>
string FIXED_BBOX 0 0 32000 29000
string GDS_END 2284076
string GDS_FILE ../gds/controller.gds
string GDS_START 257850
<< end >>
