magic
tech ihp-sg13g2
timestamp 1747537721
<< nwell >>
rect -24 175 408 417
<< pwell >>
rect 11 28 373 157
rect -13 -28 397 28
<< nmos >>
rect 58 70 71 144
rect 109 70 122 144
rect 160 70 173 144
rect 262 70 275 144
rect 313 70 326 144
<< pmos >>
rect 58 206 71 318
rect 109 206 122 318
rect 160 206 173 318
rect 262 206 275 318
rect 313 206 326 318
<< ndiff >>
rect 24 137 58 144
rect 24 121 31 137
rect 47 121 58 137
rect 24 93 58 121
rect 24 77 31 93
rect 47 77 58 93
rect 24 70 58 77
rect 71 93 109 144
rect 71 77 82 93
rect 98 77 109 93
rect 71 70 109 77
rect 122 70 160 144
rect 173 93 207 144
rect 173 77 184 93
rect 200 77 207 93
rect 173 70 207 77
rect 228 93 262 144
rect 228 77 235 93
rect 251 77 262 93
rect 228 70 262 77
rect 275 70 313 144
rect 326 93 360 144
rect 326 77 337 93
rect 353 77 360 93
rect 326 70 360 77
<< pdiff >>
rect 24 311 58 318
rect 24 295 31 311
rect 47 295 58 311
rect 24 271 58 295
rect 24 255 31 271
rect 47 255 58 271
rect 24 229 58 255
rect 24 213 31 229
rect 47 213 58 229
rect 24 206 58 213
rect 71 311 109 318
rect 71 295 82 311
rect 98 295 109 311
rect 71 271 109 295
rect 71 255 82 271
rect 98 255 109 271
rect 71 206 109 255
rect 122 271 160 318
rect 122 255 133 271
rect 149 255 160 271
rect 122 206 160 255
rect 173 311 207 318
rect 173 295 184 311
rect 200 295 207 311
rect 173 206 207 295
rect 228 311 262 318
rect 228 295 235 311
rect 251 295 262 311
rect 228 206 262 295
rect 275 311 313 318
rect 275 295 286 311
rect 302 295 313 311
rect 275 271 313 295
rect 275 255 286 271
rect 302 255 313 271
rect 275 206 313 255
rect 326 311 360 318
rect 326 295 337 311
rect 353 295 360 311
rect 326 271 360 295
rect 326 255 337 271
rect 353 255 360 271
rect 326 206 360 255
<< ndiffc >>
rect 31 121 47 137
rect 31 77 47 93
rect 82 77 98 93
rect 184 77 200 93
rect 235 77 251 93
rect 337 77 353 93
<< pdiffc >>
rect 31 295 47 311
rect 31 255 47 271
rect 31 213 47 229
rect 82 295 98 311
rect 82 255 98 271
rect 133 255 149 271
rect 184 295 200 311
rect 235 295 251 311
rect 286 295 302 311
rect 286 255 302 271
rect 337 295 353 311
rect 337 255 353 271
<< psubdiff >>
rect 0 8 384 15
rect 0 -8 16 8
rect 32 -8 64 8
rect 80 -8 112 8
rect 128 -8 160 8
rect 176 -8 208 8
rect 224 -8 256 8
rect 272 -8 304 8
rect 320 -8 352 8
rect 368 -8 384 8
rect 0 -15 384 -8
<< nsubdiff >>
rect 0 386 384 393
rect 0 370 16 386
rect 32 370 64 386
rect 80 370 112 386
rect 128 370 160 386
rect 176 370 208 386
rect 224 370 256 386
rect 272 370 304 386
rect 320 370 352 386
rect 368 370 384 386
rect 0 363 384 370
<< psubdiffcont >>
rect 16 -8 32 8
rect 64 -8 80 8
rect 112 -8 128 8
rect 160 -8 176 8
rect 208 -8 224 8
rect 256 -8 272 8
rect 304 -8 320 8
rect 352 -8 368 8
<< nsubdiffcont >>
rect 16 370 32 386
rect 64 370 80 386
rect 112 370 128 386
rect 160 370 176 386
rect 208 370 224 386
rect 256 370 272 386
rect 304 370 320 386
rect 352 370 368 386
<< poly >>
rect 58 318 71 336
rect 109 318 122 336
rect 160 318 173 336
rect 262 318 275 336
rect 313 318 326 336
rect 58 190 71 206
rect 109 190 122 206
rect 160 190 173 206
rect 262 190 275 206
rect 313 190 326 206
rect 26 183 71 190
rect 26 167 37 183
rect 53 167 71 183
rect 26 160 71 167
rect 100 183 130 190
rect 100 167 107 183
rect 123 167 130 183
rect 100 160 130 167
rect 160 183 205 190
rect 160 167 177 183
rect 193 167 205 183
rect 160 160 205 167
rect 230 183 275 190
rect 230 167 241 183
rect 257 167 275 183
rect 230 160 275 167
rect 304 183 334 190
rect 304 167 311 183
rect 327 167 334 183
rect 304 160 334 167
rect 58 144 71 160
rect 109 144 122 160
rect 160 144 173 160
rect 262 144 275 160
rect 313 144 326 160
rect 58 52 71 70
rect 109 52 122 70
rect 160 52 173 70
rect 262 52 275 70
rect 313 52 326 70
<< polycont >>
rect 37 167 53 183
rect 107 167 123 183
rect 177 167 193 183
rect 241 167 257 183
rect 311 167 327 183
<< metal1 >>
rect 0 386 384 400
rect 0 370 16 386
rect 32 370 64 386
rect 80 370 112 386
rect 128 370 160 386
rect 176 370 208 386
rect 224 370 256 386
rect 272 370 304 386
rect 320 370 352 386
rect 368 370 384 386
rect 0 356 384 370
rect 26 311 52 316
rect 26 295 31 311
rect 47 295 52 311
rect 26 271 52 295
rect 26 255 31 271
rect 47 255 52 271
rect 26 229 52 255
rect 77 311 205 316
rect 77 295 82 311
rect 98 295 184 311
rect 200 295 205 311
rect 77 271 103 295
rect 179 290 205 295
rect 230 311 256 356
rect 230 295 235 311
rect 251 295 256 311
rect 230 290 256 295
rect 281 311 307 316
rect 281 295 286 311
rect 302 295 307 311
rect 77 255 82 271
rect 98 255 103 271
rect 77 250 103 255
rect 128 271 154 276
rect 281 271 307 295
rect 128 255 133 271
rect 149 255 286 271
rect 302 255 307 271
rect 128 250 307 255
rect 332 311 358 356
rect 332 295 337 311
rect 353 295 358 311
rect 332 271 358 295
rect 332 255 337 271
rect 353 255 358 271
rect 332 250 358 255
rect 26 213 31 229
rect 47 213 374 229
rect 26 208 374 213
rect 25 183 64 190
rect 25 167 37 183
rect 53 167 64 183
rect 25 157 64 167
rect 88 183 136 190
rect 88 167 107 183
rect 123 167 136 183
rect 88 157 136 167
rect 154 183 200 190
rect 154 167 177 183
rect 193 167 200 183
rect 154 157 200 167
rect 26 121 31 137
rect 47 121 154 137
rect 26 116 154 121
rect 172 116 200 157
rect 218 183 270 190
rect 218 167 241 183
rect 257 167 270 183
rect 218 157 270 167
rect 288 183 338 190
rect 288 167 311 183
rect 327 167 338 183
rect 288 157 338 167
rect 218 116 248 157
rect 356 137 374 208
rect 281 116 374 137
rect 26 93 52 116
rect 128 98 154 116
rect 281 98 307 116
rect 26 77 31 93
rect 47 77 52 93
rect 26 72 52 77
rect 77 93 103 98
rect 77 77 82 93
rect 98 77 103 93
rect 77 22 103 77
rect 128 93 307 98
rect 128 77 184 93
rect 200 77 235 93
rect 251 77 307 93
rect 128 72 307 77
rect 332 93 358 98
rect 332 77 337 93
rect 353 77 358 93
rect 332 22 358 77
rect 0 8 384 22
rect 0 -8 16 8
rect 32 -8 64 8
rect 80 -8 112 8
rect 128 -8 160 8
rect 176 -8 208 8
rect 224 -8 256 8
rect 272 -8 304 8
rect 320 -8 352 8
rect 368 -8 384 8
rect 0 -22 384 -8
<< labels >>
flabel metal1 s 0 -22 384 22 0 FreeSans 200 0 0 0 VSS
port 3 nsew
flabel metal1 s 0 356 384 400 0 FreeSans 200 0 0 0 VDD
port 5 nsew
flabel metal1 s 25 157 64 190 0 FreeSans 200 0 0 0 C1
port 6 nsew
flabel metal1 s 356 116 374 229 0 FreeSans 200 0 0 0 Y
port 7 nsew
flabel metal1 s 88 157 136 190 0 FreeSans 200 0 0 0 B2
port 8 nsew
flabel metal1 s 172 116 200 190 0 FreeSans 200 0 0 0 B1
port 9 nsew
flabel metal1 s 288 157 338 190 0 FreeSans 200 0 0 0 A2
port 10 nsew
flabel metal1 s 218 116 248 190 0 FreeSans 200 0 0 0 A1
port 11 nsew
<< properties >>
string FIXED_BBOX 0 0 384 378
string GDS_END 144844
string GDS_FILE ../gds/controller.gds
string GDS_START 139132
<< end >>
