magic
tech ihp-sg13g2
magscale 1 2
timestamp 1747056179
<< metal1 >>
rect 576 27992 31392 28016
rect 576 27952 4352 27992
rect 4720 27952 12126 27992
rect 12494 27952 19900 27992
rect 20268 27952 27674 27992
rect 28042 27952 31392 27992
rect 576 27928 31392 27952
rect 2091 27824 2133 27833
rect 2091 27784 2092 27824
rect 2132 27784 2133 27824
rect 2091 27775 2133 27784
rect 2475 27824 2517 27833
rect 2475 27784 2476 27824
rect 2516 27784 2517 27824
rect 2475 27775 2517 27784
rect 2938 27824 2996 27825
rect 2938 27784 2947 27824
rect 2987 27784 2996 27824
rect 2938 27783 2996 27784
rect 4090 27824 4148 27825
rect 4090 27784 4099 27824
rect 4139 27784 4148 27824
rect 4090 27783 4148 27784
rect 5163 27824 5205 27833
rect 5163 27784 5164 27824
rect 5204 27784 5205 27824
rect 5163 27775 5205 27784
rect 13035 27824 13077 27833
rect 13035 27784 13036 27824
rect 13076 27784 13077 27824
rect 13035 27775 13077 27784
rect 13515 27824 13557 27833
rect 13515 27784 13516 27824
rect 13556 27784 13557 27824
rect 13515 27775 13557 27784
rect 19467 27824 19509 27833
rect 19467 27784 19468 27824
rect 19508 27784 19509 27824
rect 19467 27775 19509 27784
rect 19738 27824 19796 27825
rect 19738 27784 19747 27824
rect 19787 27784 19796 27824
rect 19738 27783 19796 27784
rect 22443 27824 22485 27833
rect 22443 27784 22444 27824
rect 22484 27784 22485 27824
rect 22443 27775 22485 27784
rect 27867 27824 27909 27833
rect 27867 27784 27868 27824
rect 27908 27784 27909 27824
rect 27867 27775 27909 27784
rect 6058 27740 6116 27741
rect 6058 27700 6067 27740
rect 6107 27700 6116 27740
rect 6058 27699 6116 27700
rect 6603 27740 6645 27749
rect 6603 27700 6604 27740
rect 6644 27700 6645 27740
rect 6603 27691 6645 27700
rect 6874 27740 6932 27741
rect 6874 27700 6883 27740
rect 6923 27700 6932 27740
rect 6874 27699 6932 27700
rect 9946 27740 10004 27741
rect 9946 27700 9955 27740
rect 9995 27700 10004 27740
rect 9946 27699 10004 27700
rect 12250 27740 12308 27741
rect 12250 27700 12259 27740
rect 12299 27700 12308 27740
rect 12250 27699 12308 27700
rect 13786 27740 13844 27741
rect 13786 27700 13795 27740
rect 13835 27700 13844 27740
rect 13786 27699 13844 27700
rect 13899 27740 13941 27749
rect 13899 27700 13900 27740
rect 13940 27700 13941 27740
rect 13899 27691 13941 27700
rect 19930 27740 19988 27741
rect 19930 27700 19939 27740
rect 19979 27700 19988 27740
rect 19930 27699 19988 27700
rect 4294 27675 4336 27684
rect 843 27656 885 27665
rect 843 27616 844 27656
rect 884 27616 885 27656
rect 843 27607 885 27616
rect 1035 27656 1077 27665
rect 1035 27616 1036 27656
rect 1076 27616 1077 27656
rect 1035 27607 1077 27616
rect 1611 27656 1653 27665
rect 1611 27616 1612 27656
rect 1652 27616 1653 27656
rect 1611 27607 1653 27616
rect 1801 27656 1843 27665
rect 1801 27616 1802 27656
rect 1842 27616 1843 27656
rect 1801 27607 1843 27616
rect 2002 27656 2044 27665
rect 2002 27616 2003 27656
rect 2043 27616 2044 27656
rect 2002 27607 2044 27616
rect 2170 27656 2228 27657
rect 2170 27616 2179 27656
rect 2219 27616 2228 27656
rect 2170 27615 2228 27616
rect 2374 27656 2416 27665
rect 2374 27616 2375 27656
rect 2415 27616 2416 27656
rect 2374 27607 2416 27616
rect 2565 27656 2607 27665
rect 2565 27616 2566 27656
rect 2606 27616 2607 27656
rect 2565 27607 2607 27616
rect 2763 27656 2805 27665
rect 2763 27616 2764 27656
rect 2804 27616 2805 27656
rect 2763 27607 2805 27616
rect 2954 27656 2996 27665
rect 2954 27616 2955 27656
rect 2995 27616 2996 27656
rect 2954 27607 2996 27616
rect 3154 27656 3196 27665
rect 3154 27616 3155 27656
rect 3195 27616 3196 27656
rect 3154 27607 3196 27616
rect 3322 27656 3380 27657
rect 3322 27616 3331 27656
rect 3371 27616 3380 27656
rect 3322 27615 3380 27616
rect 3915 27656 3957 27665
rect 3915 27616 3916 27656
rect 3956 27616 3957 27656
rect 3915 27607 3957 27616
rect 4111 27651 4153 27660
rect 4111 27611 4112 27651
rect 4152 27611 4153 27651
rect 4294 27635 4295 27675
rect 4335 27635 4336 27675
rect 4294 27626 4336 27635
rect 4491 27656 4533 27665
rect 4111 27602 4153 27611
rect 4491 27616 4492 27656
rect 4532 27616 4533 27656
rect 4491 27607 4533 27616
rect 5067 27656 5109 27665
rect 5067 27616 5068 27656
rect 5108 27616 5109 27656
rect 5067 27607 5109 27616
rect 5242 27656 5300 27657
rect 5242 27616 5251 27656
rect 5291 27616 5300 27656
rect 5242 27615 5300 27616
rect 5743 27656 5801 27657
rect 5743 27616 5752 27656
rect 5792 27616 5801 27656
rect 5743 27615 5801 27616
rect 6223 27656 6281 27657
rect 6223 27616 6232 27656
rect 6272 27616 6281 27656
rect 6223 27615 6281 27616
rect 6400 27656 6442 27665
rect 7258 27656 7316 27657
rect 6400 27616 6401 27656
rect 6441 27616 6442 27656
rect 6400 27607 6442 27616
rect 6699 27647 6741 27656
rect 6699 27607 6700 27647
rect 6740 27607 6741 27647
rect 7258 27616 7267 27656
rect 7307 27616 7316 27656
rect 7258 27615 7316 27616
rect 9679 27656 9737 27657
rect 9679 27616 9688 27656
rect 9728 27616 9737 27656
rect 9679 27615 9737 27616
rect 11866 27656 11924 27657
rect 11866 27616 11875 27656
rect 11915 27616 11924 27656
rect 11866 27615 11924 27616
rect 12634 27656 12692 27657
rect 12634 27616 12643 27656
rect 12683 27616 12692 27656
rect 12634 27615 12692 27616
rect 12747 27656 12789 27665
rect 12747 27616 12748 27656
rect 12788 27616 12789 27656
rect 12747 27607 12789 27616
rect 13227 27656 13269 27665
rect 13227 27616 13228 27656
rect 13268 27616 13269 27656
rect 13693 27656 13735 27665
rect 16282 27656 16340 27657
rect 13227 27607 13269 27616
rect 13361 27624 13419 27625
rect 6699 27598 6741 27607
rect 13361 27584 13370 27624
rect 13410 27584 13419 27624
rect 13693 27616 13694 27656
rect 13734 27616 13735 27656
rect 13693 27607 13735 27616
rect 13995 27647 14037 27656
rect 13995 27607 13996 27647
rect 14036 27607 14037 27647
rect 16282 27616 16291 27656
rect 16331 27616 16340 27656
rect 16282 27615 16340 27616
rect 16666 27656 16724 27657
rect 16666 27616 16675 27656
rect 16715 27616 16724 27656
rect 16666 27615 16724 27616
rect 17242 27656 17300 27657
rect 17242 27616 17251 27656
rect 17291 27616 17300 27656
rect 17242 27615 17300 27616
rect 19659 27656 19701 27665
rect 19659 27616 19660 27656
rect 19700 27616 19701 27656
rect 19659 27607 19701 27616
rect 21850 27656 21908 27657
rect 21850 27616 21859 27656
rect 21899 27616 21908 27656
rect 21850 27615 21908 27616
rect 24346 27656 24404 27657
rect 24346 27616 24355 27656
rect 24395 27616 24404 27656
rect 24346 27615 24404 27616
rect 24939 27656 24981 27665
rect 24939 27616 24940 27656
rect 24980 27616 24981 27656
rect 24939 27607 24981 27616
rect 25789 27656 25831 27665
rect 25789 27616 25790 27656
rect 25830 27616 25831 27656
rect 25789 27607 25831 27616
rect 25899 27656 25941 27665
rect 25899 27616 25900 27656
rect 25940 27616 25941 27656
rect 25899 27607 25941 27616
rect 26091 27656 26133 27665
rect 26091 27616 26092 27656
rect 26132 27616 26133 27656
rect 26091 27607 26133 27616
rect 26274 27647 26320 27656
rect 26274 27607 26275 27647
rect 26315 27607 26320 27647
rect 13995 27598 14037 27607
rect 26274 27598 26320 27607
rect 26754 27647 26800 27656
rect 26754 27607 26755 27647
rect 26795 27607 26800 27647
rect 26754 27598 26800 27607
rect 27234 27647 27280 27656
rect 27234 27607 27235 27647
rect 27275 27607 27280 27647
rect 27234 27598 27280 27607
rect 27714 27647 27760 27656
rect 27714 27607 27715 27647
rect 27755 27607 27760 27647
rect 27714 27598 27760 27607
rect 28194 27647 28240 27656
rect 28194 27607 28195 27647
rect 28235 27607 28240 27647
rect 28194 27598 28240 27607
rect 28674 27647 28720 27656
rect 28674 27607 28675 27647
rect 28715 27607 28720 27647
rect 28674 27598 28720 27607
rect 29154 27647 29200 27656
rect 29154 27607 29155 27647
rect 29195 27607 29200 27647
rect 29154 27598 29200 27607
rect 30882 27647 30928 27656
rect 30882 27607 30883 27647
rect 30923 27607 30928 27647
rect 30882 27598 30928 27607
rect 13361 27583 13419 27584
rect 5578 27572 5636 27573
rect 5578 27532 5587 27572
rect 5627 27532 5636 27572
rect 5578 27531 5636 27532
rect 9514 27572 9572 27573
rect 9514 27532 9523 27572
rect 9563 27532 9572 27572
rect 9514 27531 9572 27532
rect 16875 27572 16917 27581
rect 16875 27532 16876 27572
rect 16916 27532 16917 27572
rect 16875 27523 16917 27532
rect 22234 27572 22292 27573
rect 22234 27532 22243 27572
rect 22283 27532 22292 27572
rect 22234 27531 22292 27532
rect 24730 27572 24788 27573
rect 24730 27532 24739 27572
rect 24779 27532 24788 27572
rect 24730 27531 24788 27532
rect 26427 27572 26469 27581
rect 26427 27532 26428 27572
rect 26468 27532 26469 27572
rect 26427 27523 26469 27532
rect 26907 27572 26949 27581
rect 26907 27532 26908 27572
rect 26948 27532 26949 27572
rect 26907 27523 26949 27532
rect 27387 27572 27429 27581
rect 27387 27532 27388 27572
rect 27428 27532 27429 27572
rect 27387 27523 27429 27532
rect 28347 27572 28389 27581
rect 28347 27532 28348 27572
rect 28388 27532 28389 27572
rect 28347 27523 28389 27532
rect 28827 27572 28869 27581
rect 28827 27532 28828 27572
rect 28868 27532 28869 27572
rect 28827 27523 28869 27532
rect 29307 27572 29349 27581
rect 29307 27532 29308 27572
rect 29348 27532 29349 27572
rect 29307 27523 29349 27532
rect 31035 27572 31077 27581
rect 31035 27532 31036 27572
rect 31076 27532 31077 27572
rect 31035 27523 31077 27532
rect 1419 27488 1461 27497
rect 1419 27448 1420 27488
rect 1460 27448 1461 27488
rect 1419 27439 1461 27448
rect 1611 27488 1653 27497
rect 1611 27448 1612 27488
rect 1652 27448 1653 27488
rect 1611 27439 1653 27448
rect 3723 27488 3765 27497
rect 3723 27448 3724 27488
rect 3764 27448 3765 27488
rect 3723 27439 3765 27448
rect 4395 27488 4437 27497
rect 4395 27448 4396 27488
rect 4436 27448 4437 27488
rect 4395 27439 4437 27448
rect 4875 27488 4917 27497
rect 4875 27448 4876 27488
rect 4916 27448 4917 27488
rect 4875 27439 4917 27448
rect 19179 27488 19221 27497
rect 19179 27448 19180 27488
rect 19220 27448 19221 27488
rect 19179 27439 19221 27448
rect 25611 27488 25653 27497
rect 25611 27448 25612 27488
rect 25652 27448 25653 27488
rect 25611 27439 25653 27448
rect 29643 27488 29685 27497
rect 29643 27448 29644 27488
rect 29684 27448 29685 27488
rect 29643 27439 29685 27448
rect 30027 27488 30069 27497
rect 30027 27448 30028 27488
rect 30068 27448 30069 27488
rect 30027 27439 30069 27448
rect 30411 27488 30453 27497
rect 30411 27448 30412 27488
rect 30452 27448 30453 27488
rect 30411 27439 30453 27448
rect 843 27404 885 27413
rect 843 27364 844 27404
rect 884 27364 885 27404
rect 843 27355 885 27364
rect 3322 27404 3380 27405
rect 3322 27364 3331 27404
rect 3371 27364 3380 27404
rect 3322 27363 3380 27364
rect 6394 27404 6452 27405
rect 6394 27364 6403 27404
rect 6443 27364 6452 27404
rect 6394 27363 6452 27364
rect 9195 27404 9237 27413
rect 9195 27364 9196 27404
rect 9236 27364 9237 27404
rect 9195 27355 9237 27364
rect 14379 27404 14421 27413
rect 14379 27364 14380 27404
rect 14420 27364 14421 27404
rect 14379 27355 14421 27364
rect 19467 27404 19509 27413
rect 19467 27364 19468 27404
rect 19508 27364 19509 27404
rect 19467 27355 19509 27364
rect 22827 27404 22869 27413
rect 22827 27364 22828 27404
rect 22868 27364 22869 27404
rect 22827 27355 22869 27364
rect 25803 27404 25845 27413
rect 25803 27364 25804 27404
rect 25844 27364 25845 27404
rect 25803 27355 25845 27364
rect 576 27236 31392 27260
rect 576 27196 3112 27236
rect 3480 27196 10886 27236
rect 11254 27196 18660 27236
rect 19028 27196 26434 27236
rect 26802 27196 31392 27236
rect 576 27172 31392 27196
rect 891 27068 933 27077
rect 891 27028 892 27068
rect 932 27028 933 27068
rect 891 27019 933 27028
rect 1978 27068 2036 27069
rect 1978 27028 1987 27068
rect 2027 27028 2036 27068
rect 1978 27027 2036 27028
rect 2362 27068 2420 27069
rect 2362 27028 2371 27068
rect 2411 27028 2420 27068
rect 2362 27027 2420 27028
rect 9675 27068 9717 27077
rect 9675 27028 9676 27068
rect 9716 27028 9717 27068
rect 9675 27019 9717 27028
rect 12171 27068 12213 27077
rect 12171 27028 12172 27068
rect 12212 27028 12213 27068
rect 12171 27019 12213 27028
rect 17355 27068 17397 27077
rect 17355 27028 17356 27068
rect 17396 27028 17397 27068
rect 17355 27019 17397 27028
rect 20523 27068 20565 27077
rect 20523 27028 20524 27068
rect 20564 27028 20565 27068
rect 20523 27019 20565 27028
rect 21675 27068 21717 27077
rect 21675 27028 21676 27068
rect 21716 27028 21717 27068
rect 21675 27019 21717 27028
rect 23499 27068 23541 27077
rect 23499 27028 23500 27068
rect 23540 27028 23541 27068
rect 23499 27019 23541 27028
rect 29115 27068 29157 27077
rect 29115 27028 29116 27068
rect 29156 27028 29157 27068
rect 29115 27019 29157 27028
rect 29643 27068 29685 27077
rect 29643 27028 29644 27068
rect 29684 27028 29685 27068
rect 29643 27019 29685 27028
rect 3531 26984 3573 26993
rect 3531 26944 3532 26984
rect 3572 26944 3573 26984
rect 3531 26935 3573 26944
rect 3915 26984 3957 26993
rect 3915 26944 3916 26984
rect 3956 26944 3957 26984
rect 3915 26935 3957 26944
rect 15435 26984 15477 26993
rect 15435 26944 15436 26984
rect 15476 26944 15477 26984
rect 15435 26935 15477 26944
rect 19371 26984 19413 26993
rect 19371 26944 19372 26984
rect 19412 26944 19413 26984
rect 19371 26935 19413 26944
rect 21483 26984 21525 26993
rect 21483 26944 21484 26984
rect 21524 26944 21525 26984
rect 21483 26935 21525 26944
rect 27147 26984 27189 26993
rect 27147 26944 27148 26984
rect 27188 26944 27189 26984
rect 27147 26935 27189 26944
rect 27723 26984 27765 26993
rect 27723 26944 27724 26984
rect 27764 26944 27765 26984
rect 27723 26935 27765 26944
rect 28779 26984 28821 26993
rect 28779 26944 28780 26984
rect 28820 26944 28821 26984
rect 28779 26935 28821 26944
rect 31083 26984 31125 26993
rect 31083 26944 31084 26984
rect 31124 26944 31125 26984
rect 31083 26935 31125 26944
rect 651 26900 693 26909
rect 651 26860 652 26900
rect 692 26860 693 26900
rect 651 26851 693 26860
rect 1419 26900 1461 26909
rect 1419 26860 1420 26900
rect 1460 26860 1461 26900
rect 1419 26851 1461 26860
rect 1659 26900 1701 26909
rect 1659 26860 1660 26900
rect 1700 26860 1701 26900
rect 1659 26851 1701 26860
rect 13227 26900 13269 26909
rect 29355 26900 29397 26909
rect 13227 26860 13228 26900
rect 13268 26860 13269 26900
rect 13227 26851 13269 26860
rect 13458 26891 13504 26900
rect 13458 26851 13459 26891
rect 13499 26851 13504 26891
rect 29355 26860 29356 26900
rect 29396 26860 29397 26900
rect 17373 26858 17431 26859
rect 13458 26842 13504 26851
rect 14040 26849 14082 26858
rect 1035 26816 1077 26825
rect 1035 26776 1036 26816
rect 1076 26776 1077 26816
rect 1035 26767 1077 26776
rect 1210 26816 1268 26817
rect 1210 26776 1219 26816
rect 1259 26776 1268 26816
rect 1210 26775 1268 26776
rect 1803 26816 1845 26825
rect 1803 26776 1804 26816
rect 1844 26776 1845 26816
rect 1803 26767 1845 26776
rect 1978 26816 2036 26817
rect 1978 26776 1987 26816
rect 2027 26776 2036 26816
rect 1978 26775 2036 26776
rect 2194 26816 2236 26825
rect 2194 26776 2195 26816
rect 2235 26776 2236 26816
rect 2194 26767 2236 26776
rect 2362 26816 2420 26817
rect 2362 26776 2371 26816
rect 2411 26776 2420 26816
rect 2362 26775 2420 26776
rect 2571 26816 2613 26825
rect 2571 26776 2572 26816
rect 2612 26776 2613 26816
rect 2571 26767 2613 26776
rect 2763 26816 2805 26825
rect 2763 26776 2764 26816
rect 2804 26776 2805 26816
rect 2763 26767 2805 26776
rect 2955 26816 2997 26825
rect 2955 26776 2956 26816
rect 2996 26776 2997 26816
rect 2955 26767 2997 26776
rect 3147 26816 3189 26825
rect 3147 26776 3148 26816
rect 3188 26776 3189 26816
rect 3147 26767 3189 26776
rect 4779 26816 4821 26825
rect 4779 26776 4780 26816
rect 4820 26776 4821 26816
rect 4779 26767 4821 26776
rect 5338 26816 5396 26817
rect 5338 26776 5347 26816
rect 5387 26776 5396 26816
rect 5338 26775 5396 26776
rect 7467 26816 7509 26825
rect 7467 26776 7468 26816
rect 7508 26776 7509 26816
rect 7467 26767 7509 26776
rect 8523 26816 8565 26825
rect 8523 26776 8524 26816
rect 8564 26776 8565 26816
rect 8523 26767 8565 26776
rect 8667 26816 8709 26825
rect 8667 26776 8668 26816
rect 8708 26776 8709 26816
rect 8667 26767 8709 26776
rect 9003 26816 9045 26825
rect 9003 26776 9004 26816
rect 9044 26776 9045 26816
rect 9003 26767 9045 26776
rect 9867 26816 9909 26825
rect 9867 26776 9868 26816
rect 9908 26776 9909 26816
rect 9867 26767 9909 26776
rect 10234 26816 10292 26817
rect 10234 26776 10243 26816
rect 10283 26776 10292 26816
rect 10234 26775 10292 26776
rect 13035 26816 13077 26825
rect 13035 26776 13036 26816
rect 13076 26776 13077 26816
rect 13035 26767 13077 26776
rect 13323 26816 13365 26825
rect 13323 26776 13324 26816
rect 13364 26776 13365 26816
rect 13323 26767 13365 26776
rect 13552 26816 13610 26817
rect 13552 26776 13561 26816
rect 13601 26776 13610 26816
rect 13552 26775 13610 26776
rect 13707 26816 13749 26825
rect 13707 26776 13708 26816
rect 13748 26776 13749 26816
rect 13707 26767 13749 26776
rect 13821 26816 13879 26817
rect 13821 26776 13830 26816
rect 13870 26776 13879 26816
rect 13821 26775 13879 26776
rect 13944 26816 13986 26825
rect 13944 26776 13945 26816
rect 13985 26776 13986 26816
rect 14040 26809 14041 26849
rect 14081 26809 14082 26849
rect 14040 26800 14082 26809
rect 14314 26816 14372 26817
rect 13944 26767 13986 26776
rect 14314 26776 14323 26816
rect 14363 26776 14372 26816
rect 14314 26775 14372 26776
rect 14571 26816 14613 26825
rect 14571 26776 14572 26816
rect 14612 26776 14613 26816
rect 14571 26767 14613 26776
rect 14762 26816 14804 26825
rect 14762 26776 14763 26816
rect 14803 26776 14804 26816
rect 14762 26767 14804 26776
rect 15099 26816 15141 26825
rect 15099 26776 15100 26816
rect 15140 26776 15141 26816
rect 15099 26767 15141 26776
rect 15234 26816 15292 26817
rect 15234 26776 15243 26816
rect 15283 26776 15292 26816
rect 15234 26775 15292 26776
rect 15723 26816 15765 26825
rect 15723 26776 15724 26816
rect 15764 26776 15765 26816
rect 15723 26767 15765 26776
rect 15915 26816 15957 26825
rect 15915 26776 15916 26816
rect 15956 26776 15957 26816
rect 15915 26767 15957 26776
rect 16875 26816 16917 26825
rect 16875 26776 16876 26816
rect 16916 26776 16917 26816
rect 16875 26767 16917 26776
rect 17259 26816 17301 26825
rect 17373 26818 17382 26858
rect 17422 26818 17431 26858
rect 18456 26849 18498 26858
rect 29355 26851 29397 26860
rect 30411 26900 30453 26909
rect 30411 26860 30412 26900
rect 30452 26860 30453 26900
rect 30411 26851 30453 26860
rect 30891 26900 30933 26909
rect 30891 26860 30892 26900
rect 30932 26860 30933 26900
rect 30891 26851 30933 26860
rect 17373 26817 17431 26818
rect 17259 26776 17260 26816
rect 17300 26776 17301 26816
rect 17259 26767 17301 26776
rect 17500 26816 17558 26817
rect 17500 26776 17509 26816
rect 17549 26776 17558 26816
rect 17500 26775 17558 26776
rect 18031 26816 18089 26817
rect 18031 26776 18040 26816
rect 18080 26776 18089 26816
rect 18031 26775 18089 26776
rect 18216 26816 18258 26825
rect 18216 26776 18217 26816
rect 18257 26776 18258 26816
rect 18216 26767 18258 26776
rect 18333 26816 18391 26817
rect 18333 26776 18342 26816
rect 18382 26776 18391 26816
rect 18456 26809 18457 26849
rect 18497 26809 18498 26849
rect 18456 26800 18498 26809
rect 18555 26816 18597 26825
rect 18333 26775 18391 26776
rect 18555 26776 18556 26816
rect 18596 26776 18597 26816
rect 18555 26767 18597 26776
rect 18796 26816 18854 26817
rect 18796 26776 18805 26816
rect 18845 26776 18854 26816
rect 18796 26775 18854 26776
rect 18931 26816 18989 26817
rect 18931 26776 18940 26816
rect 18980 26776 18989 26816
rect 18931 26775 18989 26776
rect 19066 26816 19124 26817
rect 19066 26776 19075 26816
rect 19115 26776 19124 26816
rect 19066 26775 19124 26776
rect 19171 26816 19229 26817
rect 19171 26776 19180 26816
rect 19220 26776 19229 26816
rect 19171 26775 19229 26776
rect 19563 26816 19605 26825
rect 19563 26776 19564 26816
rect 19604 26776 19605 26816
rect 19563 26767 19605 26776
rect 20427 26816 20469 26825
rect 20427 26776 20428 26816
rect 20468 26776 20469 26816
rect 20427 26767 20469 26776
rect 20619 26816 20661 26825
rect 20619 26776 20620 26816
rect 20660 26776 20661 26816
rect 20619 26767 20661 26776
rect 20811 26816 20853 26825
rect 20811 26776 20812 26816
rect 20852 26776 20853 26816
rect 20811 26767 20853 26776
rect 22299 26816 22341 26825
rect 22299 26776 22300 26816
rect 22340 26776 22341 26816
rect 22299 26767 22341 26776
rect 23307 26816 23349 26825
rect 23307 26776 23308 26816
rect 23348 26776 23349 26816
rect 23307 26767 23349 26776
rect 24171 26816 24213 26825
rect 24171 26776 24172 26816
rect 24212 26776 24213 26816
rect 24171 26767 24213 26776
rect 26362 26816 26420 26817
rect 26362 26776 26371 26816
rect 26411 26776 26420 26816
rect 26362 26775 26420 26776
rect 26941 26816 26983 26825
rect 26941 26776 26942 26816
rect 26982 26776 26983 26816
rect 26941 26767 26983 26776
rect 27051 26816 27093 26825
rect 27051 26776 27052 26816
rect 27092 26776 27093 26816
rect 27051 26767 27093 26776
rect 27253 26816 27295 26825
rect 27253 26776 27254 26816
rect 27294 26776 27295 26816
rect 27253 26767 27295 26776
rect 27418 26816 27476 26817
rect 27418 26776 27427 26816
rect 27467 26776 27476 26816
rect 27418 26775 27476 26776
rect 27723 26816 27765 26825
rect 27723 26776 27724 26816
rect 27764 26776 27765 26816
rect 27723 26767 27765 26776
rect 27895 26816 27953 26817
rect 27895 26776 27904 26816
rect 27944 26776 27953 26816
rect 27895 26775 27953 26776
rect 28384 26816 28426 26825
rect 28384 26776 28385 26816
rect 28425 26776 28426 26816
rect 28384 26767 28426 26776
rect 28587 26816 28629 26825
rect 28587 26776 28588 26816
rect 28628 26776 28629 26816
rect 28587 26767 28629 26776
rect 29547 26816 29589 26825
rect 29547 26776 29548 26816
rect 29588 26776 29589 26816
rect 29547 26767 29589 26776
rect 29732 26813 29774 26822
rect 29732 26773 29733 26813
rect 29773 26773 29774 26813
rect 29732 26764 29774 26773
rect 29920 26816 29962 26825
rect 29920 26776 29921 26816
rect 29961 26776 29962 26816
rect 29920 26767 29962 26776
rect 30123 26816 30165 26825
rect 30123 26776 30124 26816
rect 30164 26776 30165 26816
rect 30123 26767 30165 26776
rect 30315 26816 30357 26825
rect 30315 26776 30316 26816
rect 30356 26776 30357 26816
rect 30315 26767 30357 26776
rect 30507 26816 30549 26825
rect 30507 26776 30508 26816
rect 30548 26776 30549 26816
rect 30507 26767 30549 26776
rect 4954 26732 5012 26733
rect 4954 26692 4963 26732
rect 5003 26692 5012 26732
rect 4954 26691 5012 26692
rect 8314 26732 8372 26733
rect 8314 26692 8323 26732
rect 8363 26692 8372 26732
rect 8314 26691 8372 26692
rect 15579 26732 15621 26741
rect 15579 26692 15580 26732
rect 15620 26692 15621 26732
rect 15579 26683 15621 26692
rect 24442 26732 24500 26733
rect 24442 26692 24451 26732
rect 24491 26692 24500 26732
rect 24442 26691 24500 26692
rect 26746 26732 26804 26733
rect 26746 26692 26755 26732
rect 26795 26692 26804 26732
rect 26746 26691 26804 26692
rect 28059 26732 28101 26741
rect 28059 26692 28060 26732
rect 28100 26692 28101 26732
rect 28059 26683 28101 26692
rect 1131 26648 1173 26657
rect 1131 26608 1132 26648
rect 1172 26608 1173 26648
rect 1131 26599 1173 26608
rect 2746 26648 2804 26649
rect 2746 26608 2755 26648
rect 2795 26608 2804 26648
rect 2746 26607 2804 26608
rect 3130 26648 3188 26649
rect 3130 26608 3139 26648
rect 3179 26608 3188 26648
rect 3130 26607 3188 26608
rect 4107 26648 4149 26657
rect 4107 26608 4108 26648
rect 4148 26608 4149 26648
rect 4107 26599 4149 26608
rect 7275 26648 7317 26657
rect 7275 26608 7276 26648
rect 7316 26608 7317 26648
rect 7275 26599 7317 26608
rect 8139 26648 8181 26657
rect 8139 26608 8140 26648
rect 8180 26608 8181 26648
rect 8139 26599 8181 26608
rect 8619 26648 8661 26657
rect 8619 26608 8620 26648
rect 8660 26608 8661 26648
rect 8619 26599 8661 26608
rect 12363 26648 12405 26657
rect 12363 26608 12364 26648
rect 12404 26608 12405 26648
rect 12363 26599 12405 26608
rect 13227 26648 13269 26657
rect 13227 26608 13228 26648
rect 13268 26608 13269 26648
rect 13227 26599 13269 26608
rect 14091 26648 14133 26657
rect 14091 26608 14092 26648
rect 14132 26608 14133 26648
rect 14091 26599 14133 26608
rect 14667 26648 14709 26657
rect 14667 26608 14668 26648
rect 14708 26608 14709 26648
rect 14667 26599 14709 26608
rect 15147 26648 15189 26657
rect 15147 26608 15148 26648
rect 15188 26608 15189 26648
rect 15147 26599 15189 26608
rect 16587 26648 16629 26657
rect 16587 26608 16588 26648
rect 16628 26608 16629 26648
rect 16587 26599 16629 26608
rect 16762 26648 16820 26649
rect 16762 26608 16771 26648
rect 16811 26608 16820 26648
rect 16762 26607 16820 26608
rect 17067 26648 17109 26657
rect 17067 26608 17068 26648
rect 17108 26608 17109 26648
rect 17067 26599 17109 26608
rect 17866 26648 17924 26649
rect 17866 26608 17875 26648
rect 17915 26608 17924 26648
rect 17866 26607 17924 26608
rect 18603 26648 18645 26657
rect 18603 26608 18604 26648
rect 18644 26608 18645 26648
rect 18603 26599 18645 26608
rect 20235 26648 20277 26657
rect 20235 26608 20236 26648
rect 20276 26608 20277 26648
rect 20235 26599 20277 26608
rect 22635 26648 22677 26657
rect 22635 26608 22636 26648
rect 22676 26608 22677 26648
rect 22635 26599 22677 26608
rect 28395 26648 28437 26657
rect 28395 26608 28396 26648
rect 28436 26608 28437 26648
rect 28395 26599 28437 26608
rect 29931 26648 29973 26657
rect 29931 26608 29932 26648
rect 29972 26608 29973 26648
rect 29931 26599 29973 26608
rect 30651 26648 30693 26657
rect 30651 26608 30652 26648
rect 30692 26608 30693 26648
rect 30651 26599 30693 26608
rect 576 26480 31392 26504
rect 576 26440 4352 26480
rect 4720 26440 12126 26480
rect 12494 26440 19900 26480
rect 20268 26440 27674 26480
rect 28042 26440 31392 26480
rect 576 26416 31392 26440
rect 5163 26312 5205 26321
rect 5163 26272 5164 26312
rect 5204 26272 5205 26312
rect 5163 26263 5205 26272
rect 11211 26312 11253 26321
rect 11211 26272 11212 26312
rect 11252 26272 11253 26312
rect 11211 26263 11253 26272
rect 11770 26312 11828 26313
rect 11770 26272 11779 26312
rect 11819 26272 11828 26312
rect 11770 26271 11828 26272
rect 12154 26312 12212 26313
rect 12154 26272 12163 26312
rect 12203 26272 12212 26312
rect 12154 26271 12212 26272
rect 14938 26312 14996 26313
rect 14938 26272 14947 26312
rect 14987 26272 14996 26312
rect 14938 26271 14996 26272
rect 15988 26312 16046 26313
rect 15988 26272 15997 26312
rect 16037 26272 16046 26312
rect 15988 26271 16046 26272
rect 17530 26312 17588 26313
rect 17530 26272 17539 26312
rect 17579 26272 17588 26312
rect 17530 26271 17588 26272
rect 19275 26312 19317 26321
rect 19275 26272 19276 26312
rect 19316 26272 19317 26312
rect 19275 26263 19317 26272
rect 21099 26312 21141 26321
rect 21099 26272 21100 26312
rect 21140 26272 21141 26312
rect 21099 26263 21141 26272
rect 24651 26312 24693 26321
rect 24651 26272 24652 26312
rect 24692 26272 24693 26312
rect 24651 26263 24693 26272
rect 30315 26312 30357 26321
rect 30315 26272 30316 26312
rect 30356 26272 30357 26312
rect 30315 26263 30357 26272
rect 30603 26312 30645 26321
rect 30603 26272 30604 26312
rect 30644 26272 30645 26312
rect 30603 26263 30645 26272
rect 30987 26312 31029 26321
rect 30987 26272 30988 26312
rect 31028 26272 31029 26312
rect 30987 26263 31029 26272
rect 2187 26228 2229 26237
rect 2187 26188 2188 26228
rect 2228 26188 2229 26228
rect 2187 26179 2229 26188
rect 12778 26228 12836 26229
rect 12778 26188 12787 26228
rect 12827 26188 12836 26228
rect 12778 26187 12836 26188
rect 15161 26228 15203 26237
rect 15161 26188 15162 26228
rect 15202 26188 15203 26228
rect 15161 26179 15203 26188
rect 17163 26228 17205 26237
rect 17163 26188 17164 26228
rect 17204 26188 17205 26228
rect 17163 26179 17205 26188
rect 23002 26228 23060 26229
rect 23002 26188 23011 26228
rect 23051 26188 23060 26228
rect 23002 26187 23060 26188
rect 27805 26228 27847 26237
rect 27805 26188 27806 26228
rect 27846 26188 27847 26228
rect 27805 26179 27847 26188
rect 28011 26228 28053 26237
rect 28011 26188 28012 26228
rect 28052 26188 28053 26228
rect 28011 26179 28053 26188
rect 651 26144 693 26153
rect 651 26104 652 26144
rect 692 26104 693 26144
rect 651 26095 693 26104
rect 826 26144 884 26145
rect 826 26104 835 26144
rect 875 26104 884 26144
rect 826 26103 884 26104
rect 1357 26144 1415 26145
rect 1357 26104 1366 26144
rect 1406 26104 1415 26144
rect 1357 26103 1415 26104
rect 1978 26144 2036 26145
rect 1978 26104 1987 26144
rect 2027 26104 2036 26144
rect 1978 26103 2036 26104
rect 2283 26144 2325 26153
rect 2283 26104 2284 26144
rect 2324 26104 2325 26144
rect 2283 26095 2325 26104
rect 2470 26144 2512 26153
rect 2470 26104 2471 26144
rect 2511 26104 2512 26144
rect 2470 26095 2512 26104
rect 2666 26144 2708 26153
rect 2666 26104 2667 26144
rect 2707 26104 2708 26144
rect 2666 26095 2708 26104
rect 3226 26144 3284 26145
rect 3226 26104 3235 26144
rect 3275 26104 3284 26144
rect 3226 26103 3284 26104
rect 5773 26144 5831 26145
rect 5773 26104 5782 26144
rect 5822 26104 5831 26144
rect 5773 26103 5831 26104
rect 5931 26144 5973 26153
rect 5931 26104 5932 26144
rect 5972 26104 5973 26144
rect 5931 26095 5973 26104
rect 6106 26144 6164 26145
rect 6106 26104 6115 26144
rect 6155 26104 6164 26144
rect 6106 26103 6164 26104
rect 6219 26144 6261 26153
rect 6219 26104 6220 26144
rect 6260 26104 6261 26144
rect 6219 26095 6261 26104
rect 7083 26144 7125 26153
rect 7083 26104 7084 26144
rect 7124 26104 7125 26144
rect 7083 26095 7125 26104
rect 7947 26144 7989 26153
rect 7947 26104 7948 26144
rect 7988 26104 7989 26144
rect 7947 26095 7989 26104
rect 8283 26144 8325 26153
rect 8283 26104 8284 26144
rect 8324 26104 8325 26144
rect 8283 26095 8325 26104
rect 8427 26144 8469 26153
rect 8427 26104 8428 26144
rect 8468 26104 8469 26144
rect 8427 26095 8469 26104
rect 9387 26144 9429 26153
rect 9387 26104 9388 26144
rect 9428 26104 9429 26144
rect 9387 26095 9429 26104
rect 9850 26144 9908 26145
rect 9850 26104 9859 26144
rect 9899 26104 9908 26144
rect 9850 26103 9908 26104
rect 10539 26144 10581 26153
rect 10539 26104 10540 26144
rect 10580 26104 10581 26144
rect 10539 26095 10581 26104
rect 11053 26144 11111 26145
rect 11053 26104 11062 26144
rect 11102 26104 11111 26144
rect 11053 26103 11111 26104
rect 11307 26144 11349 26153
rect 11307 26104 11308 26144
rect 11348 26104 11349 26144
rect 11307 26095 11349 26104
rect 11536 26144 11594 26145
rect 11536 26104 11545 26144
rect 11585 26104 11594 26144
rect 11536 26103 11594 26104
rect 11674 26144 11732 26145
rect 11674 26104 11683 26144
rect 11723 26104 11732 26144
rect 11674 26103 11732 26104
rect 11993 26144 12035 26153
rect 11993 26104 11994 26144
rect 12034 26104 12035 26144
rect 11993 26095 12035 26104
rect 12267 26144 12309 26153
rect 12267 26104 12268 26144
rect 12308 26104 12309 26144
rect 12267 26095 12309 26104
rect 12943 26144 13001 26145
rect 12943 26104 12952 26144
rect 12992 26104 13001 26144
rect 13398 26144 13440 26153
rect 12943 26103 13001 26104
rect 13083 26102 13125 26111
rect 1162 26060 1220 26061
rect 1162 26020 1171 26060
rect 1211 26020 1220 26060
rect 1162 26019 1220 26020
rect 2859 26060 2901 26069
rect 2859 26020 2860 26060
rect 2900 26020 2901 26060
rect 2859 26011 2901 26020
rect 5578 26060 5636 26061
rect 5578 26020 5587 26060
rect 5627 26020 5636 26060
rect 5578 26019 5636 26020
rect 9297 26060 9339 26069
rect 13083 26062 13084 26102
rect 13124 26062 13125 26102
rect 13398 26104 13399 26144
rect 13439 26104 13440 26144
rect 13398 26095 13440 26104
rect 13546 26144 13604 26145
rect 13956 26144 14014 26145
rect 13546 26104 13555 26144
rect 13595 26104 13604 26144
rect 13546 26103 13604 26104
rect 13851 26135 13893 26144
rect 13851 26095 13852 26135
rect 13892 26095 13893 26135
rect 13956 26104 13965 26144
rect 14005 26104 14014 26144
rect 13956 26103 14014 26104
rect 14187 26144 14229 26153
rect 14187 26104 14188 26144
rect 14228 26104 14229 26144
rect 14187 26095 14229 26104
rect 14371 26144 14429 26145
rect 14371 26104 14380 26144
rect 14420 26104 14429 26144
rect 14371 26103 14429 26104
rect 14620 26144 14678 26145
rect 14620 26104 14629 26144
rect 14669 26104 14678 26144
rect 14620 26103 14678 26104
rect 14842 26144 14900 26145
rect 14842 26104 14851 26144
rect 14891 26104 14900 26144
rect 14842 26103 14900 26104
rect 15339 26144 15381 26153
rect 15339 26104 15340 26144
rect 15380 26104 15381 26144
rect 14510 26102 14568 26103
rect 13851 26086 13893 26095
rect 9297 26020 9298 26060
rect 9338 26020 9339 26060
rect 9297 26011 9339 26020
rect 10858 26060 10916 26061
rect 10858 26020 10867 26060
rect 10907 26020 10916 26060
rect 10858 26019 10916 26020
rect 11442 26051 11488 26060
rect 13083 26053 13125 26062
rect 13227 26060 13269 26069
rect 14510 26062 14519 26102
rect 14559 26062 14568 26102
rect 15339 26095 15381 26104
rect 15531 26144 15573 26153
rect 15531 26104 15532 26144
rect 15572 26104 15573 26144
rect 15531 26095 15573 26104
rect 15754 26144 15812 26145
rect 15754 26104 15763 26144
rect 15803 26104 15812 26144
rect 15754 26103 15812 26104
rect 16090 26144 16148 26145
rect 16858 26144 16916 26145
rect 16090 26104 16099 26144
rect 16139 26104 16148 26144
rect 16090 26103 16148 26104
rect 16203 26135 16245 26144
rect 16203 26095 16204 26135
rect 16244 26095 16245 26135
rect 16858 26104 16867 26144
rect 16907 26104 16916 26144
rect 17648 26144 17690 26153
rect 16858 26103 16916 26104
rect 17467 26133 17509 26142
rect 16203 26086 16245 26095
rect 17467 26093 17468 26133
rect 17508 26093 17509 26133
rect 17648 26104 17649 26144
rect 17689 26104 17690 26144
rect 17648 26095 17690 26104
rect 17751 26144 17793 26153
rect 18010 26144 18068 26145
rect 17751 26104 17752 26144
rect 17792 26104 17793 26144
rect 17751 26095 17793 26104
rect 17883 26135 17925 26144
rect 17883 26095 17884 26135
rect 17924 26095 17925 26135
rect 18010 26104 18019 26144
rect 18059 26104 18068 26144
rect 18010 26103 18068 26104
rect 18411 26144 18453 26153
rect 18411 26104 18412 26144
rect 18452 26104 18453 26144
rect 18411 26095 18453 26104
rect 18538 26144 18596 26145
rect 18538 26104 18547 26144
rect 18587 26104 18596 26144
rect 18538 26103 18596 26104
rect 18652 26144 18710 26145
rect 18652 26104 18661 26144
rect 18701 26104 18710 26144
rect 18652 26103 18710 26104
rect 18987 26144 19029 26153
rect 18987 26104 18988 26144
rect 19028 26104 19029 26144
rect 18987 26095 19029 26104
rect 19301 26144 19359 26145
rect 19301 26104 19310 26144
rect 19350 26104 19359 26144
rect 19301 26103 19359 26104
rect 20139 26144 20181 26153
rect 20139 26104 20140 26144
rect 20180 26104 20181 26144
rect 20139 26095 20181 26104
rect 20427 26144 20469 26153
rect 20427 26104 20428 26144
rect 20468 26104 20469 26144
rect 20427 26095 20469 26104
rect 21250 26144 21308 26145
rect 21250 26104 21259 26144
rect 21299 26104 21308 26144
rect 21250 26103 21308 26104
rect 21698 26144 21740 26153
rect 21698 26104 21699 26144
rect 21739 26104 21740 26144
rect 22245 26146 22303 26147
rect 22245 26106 22254 26146
rect 22294 26106 22303 26146
rect 22245 26105 22303 26106
rect 22378 26144 22436 26145
rect 21562 26102 21620 26103
rect 17467 26084 17509 26093
rect 17883 26086 17925 26095
rect 14510 26061 14568 26062
rect 11442 26011 11443 26051
rect 11483 26011 11488 26051
rect 13227 26020 13228 26060
rect 13268 26020 13269 26060
rect 13227 26011 13269 26020
rect 16683 26060 16725 26069
rect 16683 26020 16684 26060
rect 16724 26020 16725 26060
rect 16683 26011 16725 26020
rect 17259 26060 17301 26069
rect 21387 26060 21429 26069
rect 21562 26062 21571 26102
rect 21611 26062 21620 26102
rect 21698 26095 21740 26104
rect 22378 26104 22387 26144
rect 22427 26104 22436 26144
rect 22924 26144 22966 26153
rect 22378 26103 22436 26104
rect 22683 26102 22725 26111
rect 21562 26061 21620 26062
rect 22683 26062 22684 26102
rect 22724 26062 22725 26102
rect 22924 26104 22925 26144
rect 22965 26104 22966 26144
rect 22924 26095 22966 26104
rect 23386 26144 23444 26145
rect 23386 26104 23395 26144
rect 23435 26104 23444 26144
rect 23386 26103 23444 26104
rect 23499 26144 23541 26153
rect 23499 26104 23500 26144
rect 23540 26104 23541 26144
rect 23499 26095 23541 26104
rect 23979 26144 24021 26153
rect 23979 26104 23980 26144
rect 24020 26104 24021 26144
rect 23979 26095 24021 26104
rect 26746 26144 26804 26145
rect 26746 26104 26755 26144
rect 26795 26104 26804 26144
rect 26746 26103 26804 26104
rect 27303 26144 27345 26153
rect 27303 26104 27304 26144
rect 27344 26104 27345 26144
rect 27303 26095 27345 26104
rect 27418 26144 27476 26145
rect 27418 26104 27427 26144
rect 27467 26104 27476 26144
rect 27418 26103 27476 26104
rect 27531 26144 27573 26153
rect 28299 26144 28341 26153
rect 27531 26104 27532 26144
rect 27572 26104 27573 26144
rect 27531 26095 27573 26104
rect 28107 26135 28149 26144
rect 28107 26095 28108 26135
rect 28148 26095 28149 26135
rect 28299 26104 28300 26144
rect 28340 26104 28341 26144
rect 28299 26095 28341 26104
rect 28491 26144 28533 26153
rect 28491 26104 28492 26144
rect 28532 26104 28533 26144
rect 28491 26095 28533 26104
rect 28683 26144 28725 26153
rect 28683 26104 28684 26144
rect 28724 26104 28725 26144
rect 28683 26095 28725 26104
rect 28875 26144 28917 26153
rect 28875 26104 28876 26144
rect 28916 26104 28917 26144
rect 28875 26095 28917 26104
rect 29068 26144 29110 26153
rect 29068 26104 29069 26144
rect 29109 26104 29110 26144
rect 29068 26095 29110 26104
rect 29259 26144 29301 26153
rect 29259 26104 29260 26144
rect 29300 26104 29301 26144
rect 29259 26095 29301 26104
rect 29451 26144 29493 26153
rect 29451 26104 29452 26144
rect 29492 26104 29493 26144
rect 29451 26095 29493 26104
rect 29641 26144 29683 26153
rect 29641 26104 29642 26144
rect 29682 26104 29683 26144
rect 29641 26095 29683 26104
rect 30219 26144 30261 26153
rect 30219 26104 30220 26144
rect 30260 26104 30261 26144
rect 30219 26095 30261 26104
rect 30411 26144 30453 26153
rect 30411 26104 30412 26144
rect 30452 26104 30453 26144
rect 30411 26095 30453 26104
rect 28107 26086 28149 26095
rect 17259 26020 17260 26060
rect 17300 26020 17301 26060
rect 17259 26011 17301 26020
rect 19218 26051 19264 26060
rect 19218 26011 19219 26051
rect 19259 26011 19264 26051
rect 21387 26020 21388 26060
rect 21428 26020 21429 26060
rect 22683 26053 22725 26062
rect 22810 26060 22868 26061
rect 21387 26011 21429 26020
rect 22810 26020 22819 26060
rect 22859 26020 22868 26060
rect 22810 26019 22868 26020
rect 24826 26060 24884 26061
rect 24826 26020 24835 26060
rect 24875 26020 24884 26060
rect 24826 26019 24884 26020
rect 27130 26060 27188 26061
rect 27130 26020 27139 26060
rect 27179 26020 27188 26060
rect 27130 26019 27188 26020
rect 27627 26060 27669 26069
rect 27627 26020 27628 26060
rect 27668 26020 27669 26060
rect 27627 26011 27669 26020
rect 30027 26060 30069 26069
rect 30027 26020 30028 26060
rect 30068 26020 30069 26060
rect 30027 26011 30069 26020
rect 11442 26002 11488 26011
rect 19218 26002 19264 26011
rect 826 25976 884 25977
rect 826 25936 835 25976
rect 875 25936 884 25976
rect 826 25935 884 25936
rect 1803 25976 1845 25985
rect 1803 25936 1804 25976
rect 1844 25936 1845 25976
rect 1803 25927 1845 25936
rect 2650 25976 2708 25977
rect 2650 25936 2659 25976
rect 2699 25936 2708 25976
rect 2650 25935 2708 25936
rect 12459 25976 12501 25985
rect 12459 25936 12460 25976
rect 12500 25936 12501 25976
rect 12459 25927 12501 25936
rect 13323 25976 13365 25985
rect 13323 25936 13324 25976
rect 13364 25936 13365 25976
rect 13323 25927 13365 25936
rect 16491 25976 16533 25985
rect 16491 25936 16492 25976
rect 16532 25936 16533 25976
rect 16491 25927 16533 25936
rect 19083 25976 19125 25985
rect 19083 25936 19084 25976
rect 19124 25936 19125 25976
rect 19083 25927 19125 25936
rect 21483 25976 21525 25985
rect 21483 25936 21484 25976
rect 21524 25936 21525 25976
rect 21483 25927 21525 25936
rect 23674 25976 23732 25977
rect 23674 25936 23683 25976
rect 23723 25936 23732 25976
rect 23674 25935 23732 25936
rect 28299 25976 28341 25985
rect 28299 25936 28300 25976
rect 28340 25936 28341 25976
rect 28299 25927 28341 25936
rect 29787 25976 29829 25985
rect 29787 25936 29788 25976
rect 29828 25936 29829 25976
rect 29787 25927 29829 25936
rect 6219 25892 6261 25901
rect 6219 25852 6220 25892
rect 6260 25852 6261 25892
rect 6219 25843 6261 25852
rect 6411 25892 6453 25901
rect 6411 25852 6412 25892
rect 6452 25852 6453 25892
rect 6411 25843 6453 25852
rect 7275 25892 7317 25901
rect 7275 25852 7276 25892
rect 7316 25852 7317 25892
rect 7275 25843 7317 25852
rect 8314 25892 8372 25893
rect 8314 25852 8323 25892
rect 8363 25852 8372 25892
rect 8314 25851 8372 25852
rect 9195 25892 9237 25901
rect 9195 25852 9196 25892
rect 9236 25852 9237 25892
rect 9195 25843 9237 25852
rect 11979 25892 12021 25901
rect 11979 25852 11980 25892
rect 12020 25852 12021 25892
rect 11979 25843 12021 25852
rect 13803 25892 13845 25901
rect 13803 25852 13804 25892
rect 13844 25852 13845 25892
rect 13803 25843 13845 25852
rect 14091 25892 14133 25901
rect 14091 25852 14092 25892
rect 14132 25852 14133 25892
rect 14091 25843 14133 25852
rect 14475 25892 14517 25901
rect 14475 25852 14476 25892
rect 14516 25852 14517 25892
rect 14475 25843 14517 25852
rect 15147 25892 15189 25901
rect 15147 25852 15148 25892
rect 15188 25852 15189 25892
rect 15147 25843 15189 25852
rect 15435 25892 15477 25901
rect 15435 25852 15436 25892
rect 15476 25852 15477 25892
rect 15435 25843 15477 25852
rect 15867 25892 15909 25901
rect 15867 25852 15868 25892
rect 15908 25852 15909 25892
rect 15867 25843 15909 25852
rect 18507 25892 18549 25901
rect 18507 25852 18508 25892
rect 18548 25852 18549 25892
rect 18507 25843 18549 25852
rect 19738 25892 19796 25893
rect 19738 25852 19747 25892
rect 19787 25852 19796 25892
rect 19738 25851 19796 25852
rect 22426 25892 22484 25893
rect 22426 25852 22435 25892
rect 22475 25852 22484 25892
rect 22426 25851 22484 25852
rect 27802 25892 27860 25893
rect 27802 25852 27811 25892
rect 27851 25852 27860 25892
rect 27802 25851 27860 25852
rect 28683 25892 28725 25901
rect 28683 25852 28684 25892
rect 28724 25852 28725 25892
rect 28683 25843 28725 25852
rect 29163 25892 29205 25901
rect 29163 25852 29164 25892
rect 29204 25852 29205 25892
rect 29163 25843 29205 25852
rect 29451 25892 29493 25901
rect 29451 25852 29452 25892
rect 29492 25852 29493 25892
rect 29451 25843 29493 25852
rect 576 25724 31392 25748
rect 576 25684 3112 25724
rect 3480 25684 10886 25724
rect 11254 25684 18660 25724
rect 19028 25684 26434 25724
rect 26802 25684 31392 25724
rect 576 25660 31392 25684
rect 2475 25556 2517 25565
rect 2475 25516 2476 25556
rect 2516 25516 2517 25556
rect 2475 25507 2517 25516
rect 3435 25556 3477 25565
rect 3435 25516 3436 25556
rect 3476 25516 3477 25556
rect 3435 25507 3477 25516
rect 4683 25556 4725 25565
rect 4683 25516 4684 25556
rect 4724 25516 4725 25556
rect 4683 25507 4725 25516
rect 9099 25556 9141 25565
rect 9099 25516 9100 25556
rect 9140 25516 9141 25556
rect 9099 25507 9141 25516
rect 10923 25556 10965 25565
rect 10923 25516 10924 25556
rect 10964 25516 10965 25556
rect 10923 25507 10965 25516
rect 13306 25556 13364 25557
rect 13306 25516 13315 25556
rect 13355 25516 13364 25556
rect 13306 25515 13364 25516
rect 14091 25556 14133 25565
rect 14091 25516 14092 25556
rect 14132 25516 14133 25556
rect 14091 25507 14133 25516
rect 14571 25556 14613 25565
rect 14571 25516 14572 25556
rect 14612 25516 14613 25556
rect 14571 25507 14613 25516
rect 20986 25556 21044 25557
rect 20986 25516 20995 25556
rect 21035 25516 21044 25556
rect 20986 25515 21044 25516
rect 23019 25556 23061 25565
rect 23019 25516 23020 25556
rect 23060 25516 23061 25556
rect 23019 25507 23061 25516
rect 24747 25556 24789 25565
rect 24747 25516 24748 25556
rect 24788 25516 24789 25556
rect 24747 25507 24789 25516
rect 29739 25556 29781 25565
rect 29739 25516 29740 25556
rect 29780 25516 29781 25556
rect 29739 25507 29781 25516
rect 4875 25472 4917 25481
rect 4875 25432 4876 25472
rect 4916 25432 4917 25472
rect 4875 25423 4917 25432
rect 12939 25472 12981 25481
rect 12939 25432 12940 25472
rect 12980 25432 12981 25472
rect 12939 25423 12981 25432
rect 15898 25472 15956 25473
rect 15898 25432 15907 25472
rect 15947 25432 15956 25472
rect 15898 25431 15956 25432
rect 19851 25472 19893 25481
rect 19851 25432 19852 25472
rect 19892 25432 19893 25472
rect 19851 25423 19893 25432
rect 21291 25472 21333 25481
rect 21291 25432 21292 25472
rect 21332 25432 21333 25472
rect 21291 25423 21333 25432
rect 30027 25472 30069 25481
rect 30027 25432 30028 25472
rect 30068 25432 30069 25472
rect 30027 25423 30069 25432
rect 30411 25472 30453 25481
rect 30411 25432 30412 25472
rect 30452 25432 30453 25472
rect 30411 25423 30453 25432
rect 30795 25472 30837 25481
rect 30795 25432 30796 25472
rect 30836 25432 30837 25472
rect 30795 25423 30837 25432
rect 9850 25388 9908 25389
rect 9850 25348 9859 25388
rect 9899 25348 9908 25388
rect 9850 25347 9908 25348
rect 10395 25388 10437 25397
rect 10395 25348 10396 25388
rect 10436 25348 10437 25388
rect 10395 25339 10437 25348
rect 13035 25388 13077 25397
rect 13035 25348 13036 25388
rect 13076 25348 13077 25388
rect 13035 25339 13077 25348
rect 16875 25388 16917 25397
rect 16875 25348 16876 25388
rect 16916 25348 16917 25388
rect 14523 25337 14565 25346
rect 16875 25339 16917 25348
rect 17338 25388 17396 25389
rect 17338 25348 17347 25388
rect 17387 25348 17396 25388
rect 17338 25347 17396 25348
rect 19354 25388 19412 25389
rect 19354 25348 19363 25388
rect 19403 25348 19412 25388
rect 19354 25347 19412 25348
rect 25402 25388 25460 25389
rect 25402 25348 25411 25388
rect 25451 25348 25460 25388
rect 25402 25347 25460 25348
rect 29259 25346 29301 25355
rect 843 25304 885 25313
rect 843 25264 844 25304
rect 884 25264 885 25304
rect 843 25255 885 25264
rect 1018 25304 1076 25305
rect 1018 25264 1027 25304
rect 1067 25264 1076 25304
rect 1018 25263 1076 25264
rect 1131 25304 1173 25313
rect 1131 25264 1132 25304
rect 1172 25264 1173 25304
rect 1131 25255 1173 25264
rect 1995 25304 2037 25313
rect 1995 25264 1996 25304
rect 2036 25264 2037 25304
rect 1995 25255 2037 25264
rect 2187 25304 2229 25313
rect 3147 25304 3189 25313
rect 2187 25264 2188 25304
rect 2228 25264 2229 25304
rect 2187 25255 2229 25264
rect 2859 25295 2901 25304
rect 2859 25255 2860 25295
rect 2900 25255 2901 25295
rect 3147 25264 3148 25304
rect 3188 25264 3189 25304
rect 3147 25255 3189 25264
rect 4107 25304 4149 25313
rect 4107 25264 4108 25304
rect 4148 25264 4149 25304
rect 4107 25255 4149 25264
rect 4378 25304 4436 25305
rect 4378 25264 4387 25304
rect 4427 25264 4436 25304
rect 4378 25263 4436 25264
rect 4491 25304 4533 25313
rect 4491 25264 4492 25304
rect 4532 25264 4533 25304
rect 4491 25255 4533 25264
rect 6778 25304 6836 25305
rect 6778 25264 6787 25304
rect 6827 25264 6836 25304
rect 6778 25263 6836 25264
rect 7371 25304 7413 25313
rect 7371 25264 7372 25304
rect 7412 25264 7413 25304
rect 7371 25255 7413 25264
rect 7755 25304 7797 25313
rect 7755 25264 7756 25304
rect 7796 25264 7797 25304
rect 7755 25255 7797 25264
rect 8811 25304 8853 25313
rect 8811 25264 8812 25304
rect 8852 25264 8853 25304
rect 8811 25255 8853 25264
rect 9147 25304 9189 25313
rect 9147 25264 9148 25304
rect 9188 25264 9189 25304
rect 9147 25255 9189 25264
rect 9291 25304 9333 25313
rect 9291 25264 9292 25304
rect 9332 25264 9333 25304
rect 9291 25255 9333 25264
rect 9718 25304 9760 25313
rect 9718 25264 9719 25304
rect 9759 25264 9760 25304
rect 9718 25255 9760 25264
rect 9963 25304 10005 25313
rect 9963 25264 9964 25304
rect 10004 25264 10005 25304
rect 9963 25255 10005 25264
rect 10186 25304 10244 25305
rect 10186 25264 10195 25304
rect 10235 25264 10244 25304
rect 10186 25263 10244 25264
rect 10827 25304 10869 25313
rect 10827 25264 10828 25304
rect 10868 25264 10869 25304
rect 10827 25255 10869 25264
rect 11020 25304 11078 25305
rect 11020 25264 11029 25304
rect 11069 25264 11078 25304
rect 11020 25263 11078 25264
rect 11403 25304 11445 25313
rect 11403 25264 11404 25304
rect 11444 25264 11445 25304
rect 11403 25255 11445 25264
rect 11787 25304 11829 25313
rect 11787 25264 11788 25304
rect 11828 25264 11829 25304
rect 11787 25255 11829 25264
rect 12154 25304 12212 25305
rect 12154 25264 12163 25304
rect 12203 25264 12212 25304
rect 12154 25263 12212 25264
rect 12267 25304 12309 25313
rect 12267 25264 12268 25304
rect 12308 25264 12309 25304
rect 12267 25255 12309 25264
rect 12708 25304 12766 25305
rect 12708 25264 12717 25304
rect 12757 25264 12766 25304
rect 12708 25263 12766 25264
rect 12878 25304 12920 25313
rect 12878 25264 12879 25304
rect 12919 25264 12920 25304
rect 12878 25255 12920 25264
rect 13156 25304 13198 25313
rect 13156 25264 13157 25304
rect 13197 25264 13198 25304
rect 13156 25255 13198 25264
rect 13309 25304 13351 25313
rect 13309 25264 13310 25304
rect 13350 25264 13351 25304
rect 13309 25255 13351 25264
rect 13603 25304 13661 25305
rect 13603 25264 13612 25304
rect 13652 25264 13661 25304
rect 13603 25263 13661 25264
rect 13803 25304 13845 25313
rect 13803 25264 13804 25304
rect 13844 25264 13845 25304
rect 13803 25255 13845 25264
rect 13978 25304 14036 25305
rect 13978 25264 13987 25304
rect 14027 25264 14036 25304
rect 13978 25263 14036 25264
rect 14091 25304 14133 25313
rect 14091 25264 14092 25304
rect 14132 25264 14133 25304
rect 14091 25255 14133 25264
rect 14283 25304 14325 25313
rect 14283 25264 14284 25304
rect 14324 25264 14325 25304
rect 14283 25255 14325 25264
rect 14397 25304 14455 25305
rect 14397 25264 14406 25304
rect 14446 25264 14455 25304
rect 14523 25297 14524 25337
rect 14564 25297 14565 25337
rect 19755 25337 19797 25346
rect 14523 25288 14565 25297
rect 14746 25304 14804 25305
rect 14397 25263 14455 25264
rect 14746 25264 14755 25304
rect 14795 25264 14804 25304
rect 14746 25263 14804 25264
rect 15062 25304 15104 25313
rect 15062 25264 15063 25304
rect 15103 25264 15104 25304
rect 15062 25255 15104 25264
rect 15610 25304 15668 25305
rect 15610 25264 15619 25304
rect 15659 25264 15668 25304
rect 15610 25263 15668 25264
rect 15723 25304 15765 25313
rect 15723 25264 15724 25304
rect 15764 25264 15765 25304
rect 15723 25255 15765 25264
rect 16395 25304 16437 25313
rect 16395 25264 16396 25304
rect 16436 25264 16437 25304
rect 16395 25255 16437 25264
rect 16483 25304 16541 25305
rect 16483 25264 16492 25304
rect 16532 25264 16541 25304
rect 16483 25263 16541 25264
rect 16779 25304 16821 25313
rect 16779 25264 16780 25304
rect 16820 25264 16821 25304
rect 16779 25255 16821 25264
rect 17082 25304 17124 25313
rect 17082 25264 17083 25304
rect 17123 25264 17124 25304
rect 17082 25255 17124 25264
rect 17218 25304 17276 25305
rect 17218 25264 17227 25304
rect 17267 25264 17276 25304
rect 17218 25263 17276 25264
rect 17451 25304 17493 25313
rect 17451 25264 17452 25304
rect 17492 25264 17493 25304
rect 17451 25255 17493 25264
rect 17962 25304 18020 25305
rect 17962 25264 17971 25304
rect 18011 25264 18020 25304
rect 17962 25263 18020 25264
rect 18202 25304 18260 25305
rect 18202 25264 18211 25304
rect 18251 25264 18260 25304
rect 18202 25263 18260 25264
rect 18616 25304 18674 25305
rect 18616 25264 18625 25304
rect 18665 25264 18674 25304
rect 18616 25263 18674 25264
rect 18891 25304 18933 25313
rect 18891 25264 18892 25304
rect 18932 25264 18933 25304
rect 18891 25255 18933 25264
rect 19222 25304 19264 25313
rect 19222 25264 19223 25304
rect 19263 25264 19264 25304
rect 19222 25255 19264 25264
rect 19465 25304 19507 25313
rect 19465 25264 19466 25304
rect 19506 25264 19507 25304
rect 19755 25297 19756 25337
rect 19796 25297 19797 25337
rect 20012 25337 20054 25346
rect 19755 25288 19797 25297
rect 19882 25304 19940 25305
rect 19465 25255 19507 25264
rect 19882 25264 19891 25304
rect 19931 25264 19940 25304
rect 20012 25297 20013 25337
rect 20053 25297 20054 25337
rect 20012 25288 20054 25297
rect 20331 25304 20373 25313
rect 19882 25263 19940 25264
rect 20331 25264 20332 25304
rect 20372 25264 20373 25304
rect 20331 25255 20373 25264
rect 20698 25304 20756 25305
rect 20698 25264 20707 25304
rect 20747 25264 20756 25304
rect 20698 25263 20756 25264
rect 20811 25304 20853 25313
rect 20811 25264 20812 25304
rect 20852 25264 20853 25304
rect 20811 25255 20853 25264
rect 21291 25304 21333 25313
rect 21291 25264 21292 25304
rect 21332 25264 21333 25304
rect 21291 25255 21333 25264
rect 21483 25304 21525 25313
rect 21483 25264 21484 25304
rect 21524 25264 21525 25304
rect 21483 25255 21525 25264
rect 22347 25304 22389 25313
rect 22347 25264 22348 25304
rect 22388 25264 22389 25304
rect 22347 25255 22389 25264
rect 22714 25304 22772 25305
rect 22714 25264 22723 25304
rect 22763 25264 22772 25304
rect 22714 25263 22772 25264
rect 22818 25304 22876 25305
rect 22818 25264 22827 25304
rect 22867 25264 22876 25304
rect 22818 25263 22876 25264
rect 23211 25304 23253 25313
rect 23211 25264 23212 25304
rect 23252 25264 23253 25304
rect 23211 25255 23253 25264
rect 24075 25304 24117 25313
rect 24075 25264 24076 25304
rect 24116 25264 24117 25304
rect 24075 25255 24117 25264
rect 24939 25304 24981 25313
rect 24939 25264 24940 25304
rect 24980 25264 24981 25304
rect 24939 25255 24981 25264
rect 25227 25304 25269 25313
rect 25227 25264 25228 25304
rect 25268 25264 25269 25304
rect 25227 25255 25269 25264
rect 27322 25304 27380 25305
rect 27322 25264 27331 25304
rect 27371 25264 27380 25304
rect 27322 25263 27380 25264
rect 28587 25304 28629 25313
rect 29259 25306 29260 25346
rect 29300 25306 29301 25346
rect 28587 25264 28588 25304
rect 28628 25264 28629 25304
rect 28587 25255 28629 25264
rect 29061 25304 29119 25305
rect 29061 25264 29070 25304
rect 29110 25264 29119 25304
rect 29259 25297 29301 25306
rect 29451 25304 29493 25313
rect 29061 25263 29119 25264
rect 29451 25264 29452 25304
rect 29492 25264 29493 25304
rect 29451 25255 29493 25264
rect 29644 25304 29686 25313
rect 29644 25264 29645 25304
rect 29685 25264 29686 25304
rect 29644 25255 29686 25264
rect 29835 25304 29877 25313
rect 29835 25264 29836 25304
rect 29876 25264 29877 25304
rect 29835 25255 29877 25264
rect 2859 25246 2901 25255
rect 922 25220 980 25221
rect 922 25180 931 25220
rect 971 25180 980 25220
rect 922 25179 980 25180
rect 2763 25220 2805 25229
rect 2763 25180 2764 25220
rect 2804 25180 2805 25220
rect 2763 25171 2805 25180
rect 4697 25220 4739 25229
rect 4697 25180 4698 25220
rect 4738 25180 4739 25220
rect 4697 25171 4739 25180
rect 7162 25220 7220 25221
rect 7162 25180 7171 25220
rect 7211 25180 7220 25220
rect 7162 25179 7220 25180
rect 8122 25220 8180 25221
rect 8122 25180 8131 25220
rect 8171 25180 8180 25220
rect 8122 25179 8180 25180
rect 16192 25220 16234 25229
rect 16192 25180 16193 25220
rect 16233 25180 16234 25220
rect 16192 25171 16234 25180
rect 19546 25220 19604 25221
rect 19546 25180 19555 25220
rect 19595 25180 19604 25220
rect 19546 25179 19604 25180
rect 23883 25220 23925 25229
rect 23883 25180 23884 25220
rect 23924 25180 23925 25220
rect 23883 25171 23925 25180
rect 27706 25220 27764 25221
rect 27706 25180 27715 25220
rect 27755 25180 27764 25220
rect 27706 25179 27764 25180
rect 27898 25220 27956 25221
rect 27898 25180 27907 25220
rect 27947 25180 27956 25220
rect 27898 25179 27956 25180
rect 28765 25220 28807 25229
rect 28765 25180 28766 25220
rect 28806 25180 28807 25220
rect 28765 25171 28807 25180
rect 28858 25220 28916 25221
rect 28858 25180 28867 25220
rect 28907 25180 28916 25220
rect 28858 25179 28916 25180
rect 1323 25136 1365 25145
rect 1323 25096 1324 25136
rect 1364 25096 1365 25136
rect 1323 25087 1365 25096
rect 2331 25136 2373 25145
rect 2331 25096 2332 25136
rect 2372 25096 2373 25136
rect 2331 25087 2373 25096
rect 7851 25136 7893 25145
rect 7851 25096 7852 25136
rect 7892 25096 7893 25136
rect 7851 25087 7893 25096
rect 10042 25136 10100 25137
rect 10042 25096 10051 25136
rect 10091 25096 10100 25136
rect 10042 25095 10100 25096
rect 10827 25136 10869 25145
rect 10827 25096 10828 25136
rect 10868 25096 10869 25136
rect 10827 25087 10869 25096
rect 11290 25136 11348 25137
rect 11290 25096 11299 25136
rect 11339 25096 11348 25136
rect 11290 25095 11348 25096
rect 12555 25136 12597 25145
rect 12555 25096 12556 25136
rect 12596 25096 12597 25136
rect 12555 25087 12597 25096
rect 13515 25136 13557 25145
rect 13515 25096 13516 25136
rect 13556 25096 13557 25136
rect 13515 25087 13557 25096
rect 14842 25136 14900 25137
rect 14842 25096 14851 25136
rect 14891 25096 14900 25136
rect 14842 25095 14900 25096
rect 14955 25136 14997 25145
rect 14955 25096 14956 25136
rect 14996 25096 14997 25136
rect 14955 25087 14997 25096
rect 16282 25136 16340 25137
rect 16282 25096 16291 25136
rect 16331 25096 16340 25136
rect 16282 25095 16340 25096
rect 17530 25136 17588 25137
rect 17530 25096 17539 25136
rect 17579 25096 17588 25136
rect 17530 25095 17588 25096
rect 18010 25136 18068 25137
rect 18010 25096 18019 25136
rect 18059 25096 18068 25136
rect 18010 25095 18068 25096
rect 18778 25136 18836 25137
rect 18778 25096 18787 25136
rect 18827 25096 18836 25136
rect 18778 25095 18836 25096
rect 19083 25136 19125 25145
rect 19083 25096 19084 25136
rect 19124 25096 19125 25136
rect 19083 25087 19125 25096
rect 20187 25136 20229 25145
rect 20187 25096 20188 25136
rect 20228 25096 20229 25136
rect 20187 25087 20229 25096
rect 21675 25136 21717 25145
rect 21675 25096 21676 25136
rect 21716 25096 21717 25136
rect 21675 25087 21717 25096
rect 22731 25136 22773 25145
rect 22731 25096 22732 25136
rect 22772 25096 22773 25136
rect 22731 25087 22773 25096
rect 25018 25136 25076 25137
rect 25018 25096 25027 25136
rect 25067 25096 25076 25136
rect 25018 25095 25076 25096
rect 28971 25136 29013 25145
rect 28971 25096 28972 25136
rect 29012 25096 29013 25136
rect 28971 25087 29013 25096
rect 29355 25136 29397 25145
rect 29355 25096 29356 25136
rect 29396 25096 29397 25136
rect 29355 25087 29397 25096
rect 576 24968 31392 24992
rect 576 24928 4352 24968
rect 4720 24928 12126 24968
rect 12494 24928 19900 24968
rect 20268 24928 27674 24968
rect 28042 24928 31392 24968
rect 576 24904 31392 24928
rect 2955 24800 2997 24809
rect 2955 24760 2956 24800
rect 2996 24760 2997 24800
rect 2955 24751 2997 24760
rect 4491 24800 4533 24809
rect 4491 24760 4492 24800
rect 4532 24760 4533 24800
rect 4491 24751 4533 24760
rect 7467 24800 7509 24809
rect 7467 24760 7468 24800
rect 7508 24760 7509 24800
rect 7467 24751 7509 24760
rect 8139 24800 8181 24809
rect 8139 24760 8140 24800
rect 8180 24760 8181 24800
rect 8139 24751 8181 24760
rect 8523 24800 8565 24809
rect 8523 24760 8524 24800
rect 8564 24760 8565 24800
rect 8523 24751 8565 24760
rect 8890 24800 8948 24801
rect 8890 24760 8899 24800
rect 8939 24760 8948 24800
rect 8890 24759 8948 24760
rect 13402 24800 13460 24801
rect 13402 24760 13411 24800
rect 13451 24760 13460 24800
rect 13402 24759 13460 24760
rect 14763 24800 14805 24809
rect 14763 24760 14764 24800
rect 14804 24760 14805 24800
rect 14763 24751 14805 24760
rect 15178 24800 15236 24801
rect 15178 24760 15187 24800
rect 15227 24760 15236 24800
rect 15178 24759 15236 24760
rect 17539 24800 17597 24801
rect 17539 24760 17548 24800
rect 17588 24760 17597 24800
rect 17539 24759 17597 24760
rect 18778 24800 18836 24801
rect 18778 24760 18787 24800
rect 18827 24760 18836 24800
rect 18778 24759 18836 24760
rect 22587 24800 22629 24809
rect 22587 24760 22588 24800
rect 22628 24760 22629 24800
rect 22587 24751 22629 24760
rect 23002 24800 23060 24801
rect 23002 24760 23011 24800
rect 23051 24760 23060 24800
rect 23002 24759 23060 24760
rect 634 24716 692 24717
rect 634 24676 643 24716
rect 683 24676 692 24716
rect 634 24675 692 24676
rect 4875 24716 4917 24725
rect 4875 24676 4876 24716
rect 4916 24676 4917 24716
rect 4875 24667 4917 24676
rect 5146 24716 5204 24717
rect 5146 24676 5155 24716
rect 5195 24676 5204 24716
rect 5146 24675 5204 24676
rect 8800 24716 8842 24725
rect 8800 24676 8801 24716
rect 8841 24676 8842 24716
rect 8800 24667 8842 24676
rect 17818 24716 17876 24717
rect 17818 24676 17827 24716
rect 17867 24676 17876 24716
rect 17818 24675 17876 24676
rect 18219 24716 18261 24725
rect 18219 24676 18220 24716
rect 18260 24676 18261 24716
rect 18219 24667 18261 24676
rect 19930 24716 19988 24717
rect 19930 24676 19939 24716
rect 19979 24676 19988 24716
rect 19930 24675 19988 24676
rect 22234 24716 22292 24717
rect 22234 24676 22243 24716
rect 22283 24676 22292 24716
rect 22234 24675 22292 24676
rect 25498 24716 25556 24717
rect 25498 24676 25507 24716
rect 25547 24676 25556 24716
rect 25498 24675 25556 24676
rect 26074 24716 26132 24717
rect 26074 24676 26083 24716
rect 26123 24676 26132 24716
rect 26074 24675 26132 24676
rect 1018 24632 1076 24633
rect 1018 24592 1027 24632
rect 1067 24592 1076 24632
rect 1018 24591 1076 24592
rect 3819 24632 3861 24641
rect 3819 24592 3820 24632
rect 3860 24592 3861 24632
rect 3819 24583 3861 24592
rect 4011 24632 4053 24641
rect 4011 24592 4012 24632
rect 4052 24592 4053 24632
rect 4011 24583 4053 24592
rect 4395 24632 4437 24641
rect 4395 24592 4396 24632
rect 4436 24592 4437 24632
rect 4395 24583 4437 24592
rect 4971 24632 5013 24641
rect 4971 24592 4972 24632
rect 5012 24592 5013 24632
rect 4971 24583 5013 24592
rect 5530 24632 5588 24633
rect 5530 24592 5539 24632
rect 5579 24592 5588 24632
rect 5530 24591 5588 24592
rect 7659 24632 7701 24641
rect 7659 24592 7660 24632
rect 7700 24592 7701 24632
rect 7659 24583 7701 24592
rect 8043 24632 8085 24641
rect 8043 24592 8044 24632
rect 8084 24592 8085 24632
rect 8043 24583 8085 24592
rect 8427 24632 8469 24641
rect 8427 24592 8428 24632
rect 8468 24592 8469 24632
rect 8427 24583 8469 24592
rect 9003 24632 9045 24641
rect 11386 24632 11444 24633
rect 9003 24592 9004 24632
rect 9044 24592 9045 24632
rect 8602 24590 8660 24591
rect 8602 24550 8611 24590
rect 8651 24550 8660 24590
rect 9003 24583 9045 24592
rect 9099 24623 9141 24632
rect 9099 24583 9100 24623
rect 9140 24583 9141 24623
rect 11386 24592 11395 24632
rect 11435 24592 11444 24632
rect 11386 24591 11444 24592
rect 11979 24632 12021 24641
rect 11979 24592 11980 24632
rect 12020 24592 12021 24632
rect 11979 24583 12021 24592
rect 12843 24632 12885 24641
rect 12843 24592 12844 24632
rect 12884 24592 12885 24632
rect 12843 24583 12885 24592
rect 12958 24632 13000 24641
rect 12958 24592 12959 24632
rect 12999 24592 13000 24632
rect 12958 24583 13000 24592
rect 13131 24632 13173 24641
rect 13131 24592 13132 24632
rect 13172 24592 13173 24632
rect 13131 24583 13173 24592
rect 13515 24632 13557 24641
rect 13515 24592 13516 24632
rect 13556 24592 13557 24632
rect 13515 24583 13557 24592
rect 13899 24632 13941 24641
rect 13899 24592 13900 24632
rect 13940 24592 13941 24632
rect 13899 24583 13941 24592
rect 14091 24632 14133 24641
rect 14091 24592 14092 24632
rect 14132 24592 14133 24632
rect 14091 24583 14133 24592
rect 15373 24632 15431 24633
rect 15373 24592 15382 24632
rect 15422 24592 15431 24632
rect 15373 24591 15431 24592
rect 16395 24632 16437 24641
rect 17146 24632 17204 24633
rect 16395 24592 16396 24632
rect 16436 24592 16437 24632
rect 16395 24583 16437 24592
rect 16578 24623 16624 24632
rect 16578 24583 16579 24623
rect 16619 24583 16624 24623
rect 17146 24592 17155 24632
rect 17195 24592 17204 24632
rect 17146 24591 17204 24592
rect 17739 24632 17781 24641
rect 17739 24592 17740 24632
rect 17780 24592 17781 24632
rect 17739 24583 17781 24592
rect 17914 24632 17972 24633
rect 17914 24592 17923 24632
rect 17963 24592 17972 24632
rect 17914 24591 17972 24592
rect 18027 24632 18069 24641
rect 18027 24592 18028 24632
rect 18068 24592 18069 24632
rect 18027 24583 18069 24592
rect 18394 24632 18452 24633
rect 18394 24592 18403 24632
rect 18443 24592 18452 24632
rect 18394 24591 18452 24592
rect 18730 24632 18788 24633
rect 18730 24592 18739 24632
rect 18779 24592 18788 24632
rect 18730 24591 18788 24592
rect 19018 24632 19076 24633
rect 19018 24592 19027 24632
rect 19067 24592 19076 24632
rect 19018 24591 19076 24592
rect 19258 24632 19316 24633
rect 19258 24592 19267 24632
rect 19307 24592 19316 24632
rect 19258 24591 19316 24592
rect 19450 24632 19508 24633
rect 19450 24592 19459 24632
rect 19499 24592 19508 24632
rect 19450 24591 19508 24592
rect 21850 24632 21908 24633
rect 21850 24592 21859 24632
rect 21899 24592 21908 24632
rect 21850 24591 21908 24592
rect 22443 24632 22485 24641
rect 22443 24592 22444 24632
rect 22484 24592 22485 24632
rect 22443 24583 22485 24592
rect 22923 24632 22965 24641
rect 22923 24592 22924 24632
rect 22964 24592 22965 24632
rect 22923 24583 22965 24592
rect 25114 24632 25172 24633
rect 25114 24592 25123 24632
rect 25163 24592 25172 24632
rect 25114 24591 25172 24592
rect 25707 24632 25749 24641
rect 25707 24592 25708 24632
rect 25748 24592 25749 24632
rect 25707 24583 25749 24592
rect 25899 24632 25941 24641
rect 25899 24592 25900 24632
rect 25940 24592 25941 24632
rect 25899 24583 25941 24592
rect 26458 24632 26516 24633
rect 26458 24592 26467 24632
rect 26507 24592 26516 24632
rect 26458 24591 26516 24592
rect 28909 24632 28967 24633
rect 28909 24592 28918 24632
rect 28958 24592 28967 24632
rect 28909 24591 28967 24592
rect 29067 24632 29109 24641
rect 29067 24592 29068 24632
rect 29108 24592 29109 24632
rect 29067 24583 29109 24592
rect 29259 24632 29301 24641
rect 29259 24592 29260 24632
rect 29300 24592 29301 24632
rect 29259 24583 29301 24592
rect 29835 24632 29877 24641
rect 29835 24592 29836 24632
rect 29876 24592 29877 24632
rect 29835 24583 29877 24592
rect 30027 24632 30069 24641
rect 30027 24592 30028 24632
rect 30068 24592 30069 24632
rect 30027 24583 30069 24592
rect 9099 24574 9141 24583
rect 16578 24574 16624 24583
rect 8602 24549 8660 24550
rect 9466 24548 9524 24549
rect 9466 24508 9475 24548
rect 9515 24508 9524 24548
rect 9466 24507 9524 24508
rect 11770 24548 11828 24549
rect 11770 24508 11779 24548
rect 11819 24508 11828 24548
rect 11770 24507 11828 24508
rect 16731 24548 16773 24557
rect 16731 24508 16732 24548
rect 16772 24508 16773 24548
rect 16731 24499 16773 24508
rect 28714 24548 28772 24549
rect 28714 24508 28723 24548
rect 28763 24508 28772 24548
rect 28714 24507 28772 24508
rect 2571 24464 2613 24473
rect 2571 24424 2572 24464
rect 2612 24424 2613 24464
rect 2571 24415 2613 24424
rect 12843 24464 12885 24473
rect 12843 24424 12844 24464
rect 12884 24424 12885 24464
rect 12843 24415 12885 24424
rect 17242 24464 17300 24465
rect 17242 24424 17251 24464
rect 17291 24424 17300 24464
rect 17242 24423 17300 24424
rect 18447 24464 18489 24473
rect 18447 24424 18448 24464
rect 18488 24424 18489 24464
rect 18447 24415 18489 24424
rect 23211 24464 23253 24473
rect 23211 24424 23212 24464
rect 23252 24424 23253 24464
rect 23211 24415 23253 24424
rect 29451 24464 29493 24473
rect 29451 24424 29452 24464
rect 29492 24424 29493 24464
rect 29451 24415 29493 24424
rect 30219 24464 30261 24473
rect 30219 24424 30220 24464
rect 30260 24424 30261 24464
rect 30219 24415 30261 24424
rect 30603 24464 30645 24473
rect 30603 24424 30604 24464
rect 30644 24424 30645 24464
rect 30603 24415 30645 24424
rect 30987 24464 31029 24473
rect 30987 24424 30988 24464
rect 31028 24424 31029 24464
rect 30987 24415 31029 24424
rect 3147 24380 3189 24389
rect 3147 24340 3148 24380
rect 3188 24340 3189 24380
rect 3147 24331 3189 24340
rect 12651 24380 12693 24389
rect 12651 24340 12652 24380
rect 12692 24340 12693 24380
rect 12651 24331 12693 24340
rect 15723 24380 15765 24389
rect 15723 24340 15724 24380
rect 15764 24340 15765 24380
rect 15723 24331 15765 24340
rect 20331 24380 20373 24389
rect 20331 24340 20332 24380
rect 20372 24340 20373 24380
rect 20331 24331 20373 24340
rect 22731 24380 22773 24389
rect 22731 24340 22732 24380
rect 22772 24340 22773 24380
rect 22731 24331 22773 24340
rect 25707 24380 25749 24389
rect 25707 24340 25708 24380
rect 25748 24340 25749 24380
rect 25707 24331 25749 24340
rect 28395 24380 28437 24389
rect 28395 24340 28396 24380
rect 28436 24340 28437 24380
rect 28395 24331 28437 24340
rect 29163 24380 29205 24389
rect 29163 24340 29164 24380
rect 29204 24340 29205 24380
rect 29163 24331 29205 24340
rect 29835 24380 29877 24389
rect 29835 24340 29836 24380
rect 29876 24340 29877 24380
rect 29835 24331 29877 24340
rect 576 24212 31392 24236
rect 576 24172 3112 24212
rect 3480 24172 10886 24212
rect 11254 24172 18660 24212
rect 19028 24172 26434 24212
rect 26802 24172 31392 24212
rect 576 24148 31392 24172
rect 1114 24044 1172 24045
rect 1114 24004 1123 24044
rect 1163 24004 1172 24044
rect 1114 24003 1172 24004
rect 6778 24044 6836 24045
rect 6778 24004 6787 24044
rect 6827 24004 6836 24044
rect 6778 24003 6836 24004
rect 12699 24044 12741 24053
rect 12699 24004 12700 24044
rect 12740 24004 12741 24044
rect 12699 23995 12741 24004
rect 16587 24044 16629 24053
rect 16587 24004 16588 24044
rect 16628 24004 16629 24044
rect 16587 23995 16629 24004
rect 19258 24044 19316 24045
rect 19258 24004 19267 24044
rect 19307 24004 19316 24044
rect 19258 24003 19316 24004
rect 21946 24044 22004 24045
rect 21946 24004 21955 24044
rect 21995 24004 22004 24044
rect 21946 24003 22004 24004
rect 23787 24044 23829 24053
rect 23787 24004 23788 24044
rect 23828 24004 23829 24044
rect 23787 23995 23829 24004
rect 25882 24044 25940 24045
rect 25882 24004 25891 24044
rect 25931 24004 25940 24044
rect 25882 24003 25940 24004
rect 27435 24044 27477 24053
rect 27435 24004 27436 24044
rect 27476 24004 27477 24044
rect 27435 23995 27477 24004
rect 28587 24044 28629 24053
rect 28587 24004 28588 24044
rect 28628 24004 28629 24044
rect 28587 23995 28629 24004
rect 29835 24044 29877 24053
rect 29835 24004 29836 24044
rect 29876 24004 29877 24044
rect 29835 23995 29877 24004
rect 651 23960 693 23969
rect 651 23920 652 23960
rect 692 23920 693 23960
rect 651 23911 693 23920
rect 3339 23960 3381 23969
rect 3339 23920 3340 23960
rect 3380 23920 3381 23960
rect 3339 23911 3381 23920
rect 12843 23960 12885 23969
rect 12843 23920 12844 23960
rect 12884 23920 12885 23960
rect 12843 23911 12885 23920
rect 15627 23960 15669 23969
rect 15627 23920 15628 23960
rect 15668 23920 15669 23960
rect 15627 23911 15669 23920
rect 20331 23960 20373 23969
rect 20331 23920 20332 23960
rect 20372 23920 20373 23960
rect 20331 23911 20373 23920
rect 30298 23960 30356 23961
rect 30298 23920 30307 23960
rect 30347 23920 30356 23960
rect 30298 23919 30356 23920
rect 20554 23904 20612 23905
rect 3531 23876 3573 23885
rect 3531 23836 3532 23876
rect 3572 23836 3573 23876
rect 8241 23876 8283 23885
rect 3531 23827 3573 23836
rect 6429 23834 6471 23843
rect 651 23792 693 23801
rect 651 23752 652 23792
rect 692 23752 693 23792
rect 651 23743 693 23752
rect 768 23792 826 23793
rect 768 23752 777 23792
rect 817 23752 826 23792
rect 768 23751 826 23752
rect 939 23792 981 23801
rect 939 23752 940 23792
rect 980 23752 981 23792
rect 939 23743 981 23752
rect 1411 23792 1469 23793
rect 1411 23752 1420 23792
rect 1460 23752 1469 23792
rect 1411 23751 1469 23752
rect 2283 23792 2325 23801
rect 2283 23752 2284 23792
rect 2324 23752 2325 23792
rect 2283 23743 2325 23752
rect 2667 23792 2709 23801
rect 2667 23752 2668 23792
rect 2708 23752 2709 23792
rect 2667 23743 2709 23752
rect 2938 23792 2996 23793
rect 2938 23752 2947 23792
rect 2987 23752 2996 23792
rect 2938 23751 2996 23752
rect 3898 23792 3956 23793
rect 3898 23752 3907 23792
rect 3947 23752 3956 23792
rect 3898 23751 3956 23752
rect 6123 23792 6165 23801
rect 6123 23752 6124 23792
rect 6164 23752 6165 23792
rect 6429 23794 6430 23834
rect 6470 23794 6471 23834
rect 8241 23836 8242 23876
rect 8282 23836 8283 23876
rect 8241 23827 8283 23836
rect 9771 23876 9813 23885
rect 9771 23836 9772 23876
rect 9812 23836 9813 23876
rect 9771 23827 9813 23836
rect 15130 23876 15188 23877
rect 15130 23836 15139 23876
rect 15179 23836 15188 23876
rect 15130 23835 15188 23836
rect 15723 23876 15765 23885
rect 15723 23836 15724 23876
rect 15764 23836 15765 23876
rect 20554 23864 20563 23904
rect 20603 23864 20612 23904
rect 20554 23863 20612 23864
rect 21291 23876 21333 23885
rect 21969 23876 22011 23885
rect 15723 23827 15765 23836
rect 21291 23836 21292 23876
rect 21332 23836 21333 23876
rect 21291 23827 21333 23836
rect 21522 23867 21568 23876
rect 21522 23827 21523 23867
rect 21563 23827 21568 23867
rect 21969 23836 21970 23876
rect 22010 23836 22011 23876
rect 21969 23827 22011 23836
rect 22618 23876 22676 23877
rect 22618 23836 22627 23876
rect 22667 23836 22676 23876
rect 22618 23835 22676 23836
rect 28923 23876 28965 23885
rect 28923 23836 28924 23876
rect 28964 23836 28965 23876
rect 28923 23827 28965 23836
rect 30507 23834 30549 23843
rect 21522 23818 21568 23827
rect 6429 23785 6471 23794
rect 6781 23792 6823 23801
rect 6123 23743 6165 23752
rect 6781 23752 6782 23792
rect 6822 23752 6823 23792
rect 6781 23743 6823 23752
rect 7075 23792 7133 23793
rect 7075 23752 7084 23792
rect 7124 23752 7133 23792
rect 7075 23751 7133 23752
rect 7786 23792 7844 23793
rect 7786 23752 7795 23792
rect 7835 23752 7844 23792
rect 7786 23751 7844 23752
rect 8331 23792 8373 23801
rect 8331 23752 8332 23792
rect 8372 23752 8373 23792
rect 8331 23743 8373 23752
rect 9003 23792 9045 23801
rect 9003 23752 9004 23792
rect 9044 23752 9045 23792
rect 9003 23743 9045 23752
rect 9195 23792 9237 23801
rect 9195 23752 9196 23792
rect 9236 23752 9237 23792
rect 9195 23743 9237 23752
rect 9850 23792 9908 23793
rect 9850 23752 9859 23792
rect 9899 23752 9908 23792
rect 9850 23751 9908 23752
rect 10522 23792 10580 23793
rect 10522 23752 10531 23792
rect 10571 23752 10580 23792
rect 10522 23751 10580 23752
rect 11163 23792 11205 23801
rect 11163 23752 11164 23792
rect 11204 23752 11205 23792
rect 11163 23743 11205 23752
rect 11307 23792 11349 23801
rect 11307 23752 11308 23792
rect 11348 23752 11349 23792
rect 11307 23743 11349 23752
rect 12267 23792 12309 23801
rect 12267 23752 12268 23792
rect 12308 23752 12309 23792
rect 12267 23743 12309 23752
rect 12555 23792 12597 23801
rect 12555 23752 12556 23792
rect 12596 23752 12597 23792
rect 12555 23743 12597 23752
rect 14746 23792 14804 23793
rect 14746 23752 14755 23792
rect 14795 23752 14804 23792
rect 14746 23751 14804 23752
rect 15387 23792 15429 23801
rect 15387 23752 15388 23792
rect 15428 23752 15429 23792
rect 15387 23743 15429 23752
rect 15566 23792 15608 23801
rect 15566 23752 15567 23792
rect 15607 23752 15608 23792
rect 15566 23743 15608 23752
rect 15850 23792 15908 23793
rect 15850 23752 15859 23792
rect 15899 23752 15908 23792
rect 15850 23751 15908 23752
rect 16070 23792 16128 23793
rect 16070 23752 16079 23792
rect 16119 23752 16128 23792
rect 16070 23751 16128 23752
rect 16208 23792 16250 23801
rect 16208 23752 16209 23792
rect 16249 23752 16250 23792
rect 16208 23743 16250 23752
rect 16311 23792 16353 23801
rect 16311 23752 16312 23792
rect 16352 23752 16353 23792
rect 16311 23743 16353 23752
rect 16435 23792 16493 23793
rect 16435 23752 16444 23792
rect 16484 23752 16493 23792
rect 16435 23751 16493 23752
rect 16570 23792 16628 23793
rect 16570 23752 16579 23792
rect 16619 23752 16628 23792
rect 16570 23751 16628 23752
rect 16875 23792 16917 23801
rect 16875 23752 16876 23792
rect 16916 23752 16917 23792
rect 16875 23743 16917 23752
rect 17242 23792 17300 23793
rect 17242 23752 17251 23792
rect 17291 23752 17300 23792
rect 17242 23751 17300 23752
rect 17643 23792 17685 23801
rect 17643 23752 17644 23792
rect 17684 23752 17685 23792
rect 17643 23743 17685 23752
rect 18202 23792 18260 23793
rect 18202 23752 18211 23792
rect 18251 23752 18260 23792
rect 18202 23751 18260 23752
rect 18315 23792 18357 23801
rect 18315 23752 18316 23792
rect 18356 23752 18357 23792
rect 18315 23743 18357 23752
rect 18970 23792 19028 23793
rect 18970 23752 18979 23792
rect 19019 23752 19028 23792
rect 18970 23751 19028 23752
rect 19083 23792 19125 23801
rect 19083 23752 19084 23792
rect 19124 23752 19125 23792
rect 19083 23743 19125 23752
rect 19740 23792 19782 23801
rect 19740 23752 19741 23792
rect 19781 23752 19782 23792
rect 19740 23743 19782 23752
rect 19851 23792 19893 23801
rect 19851 23752 19852 23792
rect 19892 23752 19893 23792
rect 19851 23743 19893 23752
rect 20506 23792 20564 23793
rect 20506 23752 20515 23792
rect 20555 23752 20564 23792
rect 20506 23751 20564 23752
rect 21003 23792 21045 23801
rect 21003 23752 21004 23792
rect 21044 23752 21045 23792
rect 21003 23743 21045 23752
rect 21387 23792 21429 23801
rect 21387 23752 21388 23792
rect 21428 23752 21429 23792
rect 21387 23743 21429 23752
rect 21616 23792 21674 23793
rect 21616 23752 21625 23792
rect 21665 23752 21674 23792
rect 21616 23751 21674 23752
rect 22059 23792 22101 23801
rect 22059 23752 22060 23792
rect 22100 23752 22101 23792
rect 22059 23743 22101 23752
rect 22498 23792 22556 23793
rect 22498 23752 22507 23792
rect 22547 23752 22556 23792
rect 22498 23751 22556 23752
rect 22731 23792 22773 23801
rect 22731 23752 22732 23792
rect 22772 23752 22773 23792
rect 22731 23743 22773 23752
rect 23115 23792 23157 23801
rect 23115 23752 23116 23792
rect 23156 23752 23157 23792
rect 23115 23743 23157 23752
rect 23979 23792 24021 23801
rect 23979 23752 23980 23792
rect 24020 23752 24021 23792
rect 23979 23743 24021 23752
rect 24939 23792 24981 23801
rect 24939 23752 24940 23792
rect 24980 23752 24981 23792
rect 24939 23743 24981 23752
rect 25147 23792 25205 23793
rect 25147 23752 25156 23792
rect 25196 23752 25205 23792
rect 25147 23751 25205 23752
rect 25306 23792 25364 23793
rect 25306 23752 25315 23792
rect 25355 23752 25364 23792
rect 25306 23751 25364 23752
rect 25450 23792 25508 23793
rect 25450 23752 25459 23792
rect 25499 23752 25508 23792
rect 25450 23751 25508 23752
rect 25594 23792 25652 23793
rect 25594 23752 25603 23792
rect 25643 23752 25652 23792
rect 25594 23751 25652 23752
rect 25716 23792 25774 23793
rect 25716 23752 25725 23792
rect 25765 23752 25774 23792
rect 25716 23751 25774 23752
rect 25888 23792 25930 23801
rect 25888 23752 25889 23792
rect 25929 23752 25930 23792
rect 25888 23743 25930 23752
rect 26179 23792 26237 23793
rect 26179 23752 26188 23792
rect 26228 23752 26237 23792
rect 26179 23751 26237 23752
rect 27243 23792 27285 23801
rect 27243 23752 27244 23792
rect 27284 23752 27285 23792
rect 27243 23743 27285 23752
rect 28107 23792 28149 23801
rect 28107 23752 28108 23792
rect 28148 23752 28149 23792
rect 28107 23743 28149 23752
rect 28395 23792 28437 23801
rect 28395 23752 28396 23792
rect 28436 23752 28437 23792
rect 28395 23743 28437 23752
rect 28759 23792 28817 23793
rect 28759 23752 28768 23792
rect 28808 23752 28817 23792
rect 28759 23751 28817 23752
rect 29355 23792 29397 23801
rect 29355 23752 29356 23792
rect 29396 23752 29397 23792
rect 29355 23743 29397 23752
rect 29739 23792 29781 23801
rect 29739 23752 29740 23792
rect 29780 23752 29781 23792
rect 29739 23743 29781 23752
rect 29931 23792 29973 23801
rect 29931 23752 29932 23792
rect 29972 23752 29973 23792
rect 29931 23743 29973 23752
rect 30123 23792 30165 23801
rect 30123 23752 30124 23792
rect 30164 23752 30165 23792
rect 30123 23743 30165 23752
rect 30314 23792 30356 23801
rect 30314 23752 30315 23792
rect 30355 23752 30356 23792
rect 30507 23794 30508 23834
rect 30548 23794 30549 23834
rect 30507 23785 30549 23794
rect 30692 23792 30734 23801
rect 30314 23743 30356 23752
rect 30692 23752 30693 23792
rect 30733 23752 30734 23792
rect 30692 23743 30734 23752
rect 30891 23792 30933 23801
rect 30891 23752 30892 23792
rect 30932 23752 30933 23792
rect 30891 23743 30933 23752
rect 31083 23792 31125 23801
rect 31083 23752 31084 23792
rect 31124 23752 31125 23792
rect 31083 23743 31125 23752
rect 1120 23708 1162 23717
rect 1120 23668 1121 23708
rect 1161 23668 1162 23708
rect 1120 23659 1162 23668
rect 3051 23708 3093 23717
rect 3051 23668 3052 23708
rect 3092 23668 3093 23708
rect 3051 23659 3093 23668
rect 6219 23708 6261 23717
rect 6219 23668 6220 23708
rect 6260 23668 6261 23708
rect 6219 23659 6261 23668
rect 6987 23708 7029 23717
rect 6987 23668 6988 23708
rect 7028 23668 7029 23708
rect 6987 23659 7029 23668
rect 10347 23708 10389 23717
rect 10347 23668 10348 23708
rect 10388 23668 10389 23708
rect 10347 23659 10389 23668
rect 11866 23708 11924 23709
rect 11866 23668 11875 23708
rect 11915 23668 11924 23708
rect 11866 23667 11924 23668
rect 17163 23708 17205 23717
rect 17163 23668 17164 23708
rect 17204 23668 17205 23708
rect 17163 23659 17205 23668
rect 24250 23708 24308 23709
rect 24250 23668 24259 23708
rect 24299 23668 24308 23708
rect 24250 23667 24308 23668
rect 30603 23708 30645 23717
rect 30603 23668 30604 23708
rect 30644 23668 30645 23708
rect 30603 23659 30645 23668
rect 1323 23624 1365 23633
rect 1323 23584 1324 23624
rect 1364 23584 1365 23624
rect 1323 23575 1365 23584
rect 1611 23624 1653 23633
rect 1611 23584 1612 23624
rect 1652 23584 1653 23624
rect 1611 23575 1653 23584
rect 5835 23624 5877 23633
rect 5835 23584 5836 23624
rect 5876 23584 5877 23624
rect 5835 23575 5877 23584
rect 6315 23624 6357 23633
rect 6315 23584 6316 23624
rect 6356 23584 6357 23624
rect 6315 23575 6357 23584
rect 6603 23624 6645 23633
rect 6603 23584 6604 23624
rect 6644 23584 6645 23624
rect 6603 23575 6645 23584
rect 7563 23624 7605 23633
rect 7563 23584 7564 23624
rect 7604 23584 7605 23624
rect 7563 23575 7605 23584
rect 8026 23624 8084 23625
rect 8026 23584 8035 23624
rect 8075 23584 8084 23624
rect 8026 23583 8084 23584
rect 9195 23624 9237 23633
rect 9195 23584 9196 23624
rect 9236 23584 9237 23624
rect 9195 23575 9237 23584
rect 9466 23624 9524 23625
rect 9466 23584 9475 23624
rect 9515 23584 9524 23624
rect 9466 23583 9524 23584
rect 10138 23624 10196 23625
rect 10138 23584 10147 23624
rect 10187 23584 10196 23624
rect 10138 23583 10196 23584
rect 11002 23624 11060 23625
rect 11002 23584 11011 23624
rect 11051 23584 11060 23624
rect 11002 23583 11060 23584
rect 16731 23624 16773 23633
rect 16731 23584 16732 23624
rect 16772 23584 16773 23624
rect 16731 23575 16773 23584
rect 18603 23624 18645 23633
rect 18603 23584 18604 23624
rect 18644 23584 18645 23624
rect 18603 23575 18645 23584
rect 19546 23624 19604 23625
rect 19546 23584 19555 23624
rect 19595 23584 19604 23624
rect 19546 23583 19604 23584
rect 20811 23624 20853 23633
rect 20811 23584 20812 23624
rect 20852 23584 20853 23624
rect 20811 23575 20853 23584
rect 21082 23624 21140 23625
rect 21082 23584 21091 23624
rect 21131 23584 21140 23624
rect 21082 23583 21140 23584
rect 22810 23624 22868 23625
rect 22810 23584 22819 23624
rect 22859 23584 22868 23624
rect 22810 23583 22868 23584
rect 25498 23624 25556 23625
rect 25498 23584 25507 23624
rect 25547 23584 25556 23624
rect 25498 23583 25556 23584
rect 26091 23624 26133 23633
rect 26091 23584 26092 23624
rect 26132 23584 26133 23624
rect 26091 23575 26133 23584
rect 26571 23624 26613 23633
rect 26571 23584 26572 23624
rect 26612 23584 26613 23624
rect 26571 23575 26613 23584
rect 28282 23624 28340 23625
rect 28282 23584 28291 23624
rect 28331 23584 28340 23624
rect 28282 23583 28340 23584
rect 29242 23624 29300 23625
rect 29242 23584 29251 23624
rect 29291 23584 29300 23624
rect 29242 23583 29300 23584
rect 29547 23624 29589 23633
rect 29547 23584 29548 23624
rect 29588 23584 29589 23624
rect 29547 23575 29589 23584
rect 30987 23624 31029 23633
rect 30987 23584 30988 23624
rect 31028 23584 31029 23624
rect 30987 23575 31029 23584
rect 576 23456 31392 23480
rect 576 23416 4352 23456
rect 4720 23416 12126 23456
rect 12494 23416 19900 23456
rect 20268 23416 27674 23456
rect 28042 23416 31392 23456
rect 576 23392 31392 23416
rect 2955 23288 2997 23297
rect 2955 23248 2956 23288
rect 2996 23248 2997 23288
rect 2955 23239 2997 23248
rect 3915 23288 3957 23297
rect 3915 23248 3916 23288
rect 3956 23248 3957 23288
rect 3915 23239 3957 23248
rect 4491 23288 4533 23297
rect 4491 23248 4492 23288
rect 4532 23248 4533 23288
rect 4491 23239 4533 23248
rect 5434 23288 5492 23289
rect 5434 23248 5443 23288
rect 5483 23248 5492 23288
rect 5434 23247 5492 23248
rect 6795 23288 6837 23297
rect 6795 23248 6796 23288
rect 6836 23248 6837 23288
rect 6795 23239 6837 23248
rect 7258 23288 7316 23289
rect 7258 23248 7267 23288
rect 7307 23248 7316 23288
rect 7258 23247 7316 23248
rect 7899 23288 7941 23297
rect 7899 23248 7900 23288
rect 7940 23248 7941 23288
rect 7899 23239 7941 23248
rect 11787 23288 11829 23297
rect 11787 23248 11788 23288
rect 11828 23248 11829 23288
rect 11787 23239 11829 23248
rect 13882 23288 13940 23289
rect 13882 23248 13891 23288
rect 13931 23248 13940 23288
rect 13882 23247 13940 23248
rect 15243 23288 15285 23297
rect 15243 23248 15244 23288
rect 15284 23248 15285 23288
rect 15243 23239 15285 23248
rect 16443 23288 16485 23297
rect 16443 23248 16444 23288
rect 16484 23248 16485 23288
rect 16443 23239 16485 23248
rect 19738 23288 19796 23289
rect 19738 23248 19747 23288
rect 19787 23248 19796 23288
rect 19738 23247 19796 23248
rect 20698 23288 20756 23289
rect 20698 23248 20707 23288
rect 20747 23248 20756 23288
rect 20698 23247 20756 23248
rect 26763 23288 26805 23297
rect 26763 23248 26764 23288
rect 26804 23248 26805 23288
rect 26763 23239 26805 23248
rect 30027 23288 30069 23297
rect 30027 23248 30028 23288
rect 30068 23248 30069 23288
rect 30027 23239 30069 23248
rect 634 23204 692 23205
rect 634 23164 643 23204
rect 683 23164 692 23204
rect 634 23163 692 23164
rect 6267 23204 6309 23213
rect 6267 23164 6268 23204
rect 6308 23164 6309 23204
rect 6267 23155 6309 23164
rect 7738 23204 7796 23205
rect 7738 23164 7747 23204
rect 7787 23164 7796 23204
rect 7738 23163 7796 23164
rect 16971 23204 17013 23213
rect 16971 23164 16972 23204
rect 17012 23164 17013 23204
rect 16971 23155 17013 23164
rect 20091 23204 20133 23213
rect 20091 23164 20092 23204
rect 20132 23164 20133 23204
rect 20091 23155 20133 23164
rect 20605 23204 20647 23213
rect 20605 23164 20606 23204
rect 20646 23164 20647 23204
rect 20605 23155 20647 23164
rect 20811 23204 20853 23213
rect 20811 23164 20812 23204
rect 20852 23164 20853 23204
rect 20811 23155 20853 23164
rect 24250 23204 24308 23205
rect 24250 23164 24259 23204
rect 24299 23164 24308 23204
rect 24250 23163 24308 23164
rect 1018 23120 1076 23121
rect 1018 23080 1027 23120
rect 1067 23080 1076 23120
rect 1018 23079 1076 23080
rect 3435 23120 3477 23129
rect 3435 23080 3436 23120
rect 3476 23080 3477 23120
rect 3435 23071 3477 23080
rect 3819 23120 3861 23129
rect 3819 23080 3820 23120
rect 3860 23080 3861 23120
rect 3819 23071 3861 23080
rect 4299 23120 4341 23129
rect 4299 23080 4300 23120
rect 4340 23080 4341 23120
rect 4299 23071 4341 23080
rect 5163 23120 5205 23129
rect 5163 23080 5164 23120
rect 5204 23080 5205 23120
rect 5163 23071 5205 23080
rect 5722 23120 5780 23121
rect 6891 23120 6933 23129
rect 5722 23080 5731 23120
rect 5771 23080 5780 23120
rect 5722 23079 5780 23080
rect 6114 23111 6160 23120
rect 6114 23071 6115 23111
rect 6155 23071 6160 23111
rect 6891 23080 6892 23120
rect 6932 23080 6933 23120
rect 6891 23071 6933 23080
rect 7083 23120 7125 23129
rect 7083 23080 7084 23120
rect 7124 23080 7125 23120
rect 7083 23071 7125 23080
rect 7279 23115 7321 23124
rect 7279 23075 7280 23115
rect 7320 23075 7321 23115
rect 7659 23120 7701 23129
rect 6114 23062 6160 23071
rect 7279 23066 7321 23075
rect 7419 23078 7461 23087
rect 7419 23038 7420 23078
rect 7460 23038 7461 23078
rect 7659 23080 7660 23120
rect 7700 23080 7701 23120
rect 7659 23071 7701 23080
rect 8091 23120 8133 23129
rect 8091 23080 8092 23120
rect 8132 23080 8133 23120
rect 8091 23071 8133 23080
rect 8235 23120 8277 23129
rect 8235 23080 8236 23120
rect 8276 23080 8277 23120
rect 8235 23071 8277 23080
rect 8410 23120 8468 23121
rect 8410 23080 8419 23120
rect 8459 23080 8468 23120
rect 8410 23079 8468 23080
rect 8950 23120 8992 23129
rect 8950 23080 8951 23120
rect 8991 23080 8992 23120
rect 8950 23071 8992 23080
rect 9195 23120 9237 23129
rect 9195 23080 9196 23120
rect 9236 23080 9237 23120
rect 9195 23071 9237 23080
rect 9850 23120 9908 23121
rect 9850 23080 9859 23120
rect 9899 23080 9908 23120
rect 9850 23079 9908 23080
rect 11979 23120 12021 23129
rect 11979 23080 11980 23120
rect 12020 23080 12021 23120
rect 11979 23071 12021 23080
rect 12651 23120 12693 23129
rect 12651 23080 12652 23120
rect 12692 23080 12693 23120
rect 12651 23071 12693 23080
rect 13323 23120 13365 23129
rect 13323 23080 13324 23120
rect 13364 23080 13365 23120
rect 14000 23120 14042 23129
rect 13323 23071 13365 23080
rect 13819 23109 13861 23118
rect 13819 23069 13820 23109
rect 13860 23069 13861 23109
rect 14000 23080 14001 23120
rect 14041 23080 14042 23120
rect 14000 23071 14042 23080
rect 14103 23120 14145 23129
rect 14103 23080 14104 23120
rect 14144 23080 14145 23120
rect 14103 23071 14145 23080
rect 14234 23120 14292 23121
rect 14234 23080 14243 23120
rect 14283 23080 14292 23120
rect 14234 23079 14292 23080
rect 14362 23120 14420 23121
rect 14362 23080 14371 23120
rect 14411 23080 14420 23120
rect 14362 23079 14420 23080
rect 14571 23120 14613 23129
rect 14571 23080 14572 23120
rect 14612 23080 14613 23120
rect 14571 23071 14613 23080
rect 15547 23120 15605 23121
rect 15547 23080 15556 23120
rect 15596 23080 15605 23120
rect 15547 23079 15605 23080
rect 15706 23120 15764 23121
rect 15706 23080 15715 23120
rect 15755 23080 15764 23120
rect 15706 23079 15764 23080
rect 15831 23120 15873 23129
rect 15831 23080 15832 23120
rect 15872 23080 15873 23120
rect 15831 23071 15873 23080
rect 15994 23120 16052 23121
rect 15994 23080 16003 23120
rect 16043 23080 16052 23120
rect 15994 23079 16052 23080
rect 16096 23120 16154 23121
rect 16096 23080 16105 23120
rect 16145 23080 16154 23120
rect 16096 23079 16154 23080
rect 16234 23120 16292 23121
rect 16234 23080 16243 23120
rect 16283 23080 16292 23120
rect 16234 23079 16292 23080
rect 17067 23120 17109 23129
rect 17067 23080 17068 23120
rect 17108 23080 17109 23120
rect 17067 23071 17109 23080
rect 17296 23120 17354 23121
rect 17296 23080 17305 23120
rect 17345 23080 17354 23120
rect 17296 23079 17354 23080
rect 17451 23120 17493 23129
rect 17451 23080 17452 23120
rect 17492 23080 17493 23120
rect 17451 23071 17493 23080
rect 17626 23120 17684 23121
rect 17626 23080 17635 23120
rect 17675 23080 17684 23120
rect 17626 23079 17684 23080
rect 17931 23120 17973 23129
rect 17931 23080 17932 23120
rect 17972 23080 17973 23120
rect 17931 23071 17973 23080
rect 18123 23120 18165 23129
rect 18123 23080 18124 23120
rect 18164 23080 18165 23120
rect 18123 23071 18165 23080
rect 18307 23120 18365 23121
rect 18307 23080 18316 23120
rect 18356 23080 18365 23120
rect 18307 23079 18365 23080
rect 18556 23120 18614 23121
rect 18556 23080 18565 23120
rect 18605 23080 18614 23120
rect 18556 23079 18614 23080
rect 19467 23120 19509 23129
rect 19467 23080 19468 23120
rect 19508 23080 19509 23120
rect 18430 23078 18488 23079
rect 13819 23060 13861 23069
rect 5338 23036 5396 23037
rect 5338 22996 5347 23036
rect 5387 22996 5396 23036
rect 5338 22995 5396 22996
rect 5914 23036 5972 23037
rect 5914 22996 5923 23036
rect 5963 22996 5972 23036
rect 7419 23029 7461 23038
rect 7546 23036 7604 23037
rect 5914 22995 5972 22996
rect 7546 22996 7555 23036
rect 7595 22996 7604 23036
rect 7546 22995 7604 22996
rect 9082 23036 9140 23037
rect 9082 22996 9091 23036
rect 9131 22996 9140 23036
rect 9082 22995 9140 22996
rect 9291 23036 9333 23045
rect 9291 22996 9292 23036
rect 9332 22996 9333 23036
rect 9291 22987 9333 22996
rect 9483 23036 9525 23045
rect 9483 22996 9484 23036
rect 9524 22996 9525 23036
rect 9483 22987 9525 22996
rect 17186 23036 17228 23045
rect 18430 23038 18439 23078
rect 18479 23038 18488 23078
rect 19467 23071 19509 23080
rect 19642 23120 19700 23121
rect 19642 23080 19651 23120
rect 19691 23080 19700 23120
rect 19642 23079 19700 23080
rect 19961 23120 20003 23129
rect 21082 23120 21140 23121
rect 19961 23080 19962 23120
rect 20002 23080 20003 23120
rect 19961 23071 20003 23080
rect 20907 23111 20949 23120
rect 20907 23071 20908 23111
rect 20948 23071 20949 23111
rect 21082 23080 21091 23120
rect 21131 23080 21140 23120
rect 21082 23079 21140 23080
rect 21771 23120 21813 23129
rect 21771 23080 21772 23120
rect 21812 23080 21813 23120
rect 21771 23071 21813 23080
rect 22731 23120 22773 23129
rect 22731 23080 22732 23120
rect 22772 23080 22773 23120
rect 22731 23071 22773 23080
rect 23595 23120 23637 23129
rect 23595 23080 23596 23120
rect 23636 23080 23637 23120
rect 23595 23071 23637 23080
rect 23830 23120 23872 23129
rect 24075 23120 24117 23129
rect 23830 23080 23831 23120
rect 23871 23080 23872 23120
rect 23830 23071 23872 23080
rect 23970 23111 24016 23120
rect 23970 23071 23971 23111
rect 24011 23071 24016 23111
rect 24075 23080 24076 23120
rect 24116 23080 24117 23120
rect 24075 23071 24117 23080
rect 26170 23120 26228 23121
rect 26170 23080 26179 23120
rect 26219 23080 26228 23120
rect 26170 23079 26228 23080
rect 28666 23120 28724 23121
rect 28666 23080 28675 23120
rect 28715 23080 28724 23120
rect 28666 23079 28724 23080
rect 29050 23120 29108 23121
rect 29050 23080 29059 23120
rect 29099 23080 29108 23120
rect 29050 23079 29108 23080
rect 30027 23120 30069 23129
rect 30027 23080 30028 23120
rect 30068 23080 30069 23120
rect 30027 23071 30069 23080
rect 30219 23120 30261 23129
rect 30219 23080 30220 23120
rect 30260 23080 30261 23120
rect 30219 23071 30261 23080
rect 31179 23120 31221 23129
rect 31179 23080 31180 23120
rect 31220 23080 31221 23120
rect 31179 23071 31221 23080
rect 20907 23062 20949 23071
rect 23970 23062 24016 23071
rect 18430 23037 18488 23038
rect 17186 22996 17187 23036
rect 17227 22996 17228 23036
rect 17186 22987 17228 22996
rect 20331 23036 20373 23045
rect 20331 22996 20332 23036
rect 20372 22996 20373 23036
rect 20331 22987 20373 22996
rect 26554 23036 26612 23037
rect 26554 22996 26563 23036
rect 26603 22996 26612 23036
rect 26554 22995 26612 22996
rect 8811 22952 8853 22961
rect 8811 22912 8812 22952
rect 8852 22912 8853 22952
rect 8811 22903 8853 22912
rect 11403 22952 11445 22961
rect 11403 22912 11404 22952
rect 11444 22912 11445 22952
rect 11403 22903 11445 22912
rect 18027 22952 18069 22961
rect 18027 22912 18028 22952
rect 18068 22912 18069 22952
rect 18027 22903 18069 22912
rect 18603 22952 18645 22961
rect 18603 22912 18604 22952
rect 18644 22912 18645 22952
rect 18603 22903 18645 22912
rect 22923 22952 22965 22961
rect 22923 22912 22924 22952
rect 22964 22912 22965 22952
rect 22923 22903 22965 22912
rect 23787 22952 23829 22961
rect 23787 22912 23788 22952
rect 23828 22912 23829 22952
rect 23787 22903 23829 22912
rect 29259 22952 29301 22961
rect 29259 22912 29260 22952
rect 29300 22912 29301 22952
rect 29259 22903 29301 22912
rect 29643 22952 29685 22961
rect 29643 22912 29644 22952
rect 29684 22912 29685 22952
rect 29643 22903 29685 22912
rect 30411 22952 30453 22961
rect 30411 22912 30412 22952
rect 30452 22912 30453 22952
rect 30411 22903 30453 22912
rect 30795 22952 30837 22961
rect 30795 22912 30796 22952
rect 30836 22912 30837 22952
rect 30795 22903 30837 22912
rect 2571 22868 2613 22877
rect 2571 22828 2572 22868
rect 2612 22828 2613 22868
rect 2571 22819 2613 22828
rect 8410 22868 8468 22869
rect 8410 22828 8419 22868
rect 8459 22828 8468 22868
rect 8410 22827 8468 22828
rect 12922 22868 12980 22869
rect 12922 22828 12931 22868
rect 12971 22828 12980 22868
rect 12922 22827 12980 22828
rect 16107 22868 16149 22877
rect 16107 22828 16108 22868
rect 16148 22828 16149 22868
rect 16107 22819 16149 22828
rect 17626 22868 17684 22869
rect 17626 22828 17635 22868
rect 17675 22828 17684 22868
rect 17626 22827 17684 22828
rect 18795 22868 18837 22877
rect 18795 22828 18796 22868
rect 18836 22828 18837 22868
rect 18795 22819 18837 22828
rect 19947 22868 19989 22877
rect 19947 22828 19948 22868
rect 19988 22828 19989 22868
rect 19947 22819 19989 22828
rect 22059 22868 22101 22877
rect 22059 22828 22060 22868
rect 22100 22828 22101 22868
rect 22059 22819 22101 22828
rect 576 22700 31392 22724
rect 576 22660 3112 22700
rect 3480 22660 10886 22700
rect 11254 22660 18660 22700
rect 19028 22660 26434 22700
rect 26802 22660 31392 22700
rect 576 22636 31392 22660
rect 6394 22532 6452 22533
rect 6394 22492 6403 22532
rect 6443 22492 6452 22532
rect 6394 22491 6452 22492
rect 10731 22532 10773 22541
rect 10731 22492 10732 22532
rect 10772 22492 10773 22532
rect 10731 22483 10773 22492
rect 16299 22532 16341 22541
rect 16299 22492 16300 22532
rect 16340 22492 16341 22532
rect 16299 22483 16341 22492
rect 21099 22532 21141 22541
rect 21099 22492 21100 22532
rect 21140 22492 21141 22532
rect 21099 22483 21141 22492
rect 21723 22532 21765 22541
rect 21723 22492 21724 22532
rect 21764 22492 21765 22532
rect 21723 22483 21765 22492
rect 24363 22532 24405 22541
rect 24363 22492 24364 22532
rect 24404 22492 24405 22532
rect 24363 22483 24405 22492
rect 25210 22532 25268 22533
rect 25210 22492 25219 22532
rect 25259 22492 25268 22532
rect 25210 22491 25268 22492
rect 26571 22532 26613 22541
rect 26571 22492 26572 22532
rect 26612 22492 26613 22532
rect 26571 22483 26613 22492
rect 27051 22532 27093 22541
rect 27051 22492 27052 22532
rect 27092 22492 27093 22532
rect 27051 22483 27093 22492
rect 8218 22448 8276 22449
rect 8218 22408 8227 22448
rect 8267 22408 8276 22448
rect 8218 22407 8276 22408
rect 10347 22448 10389 22457
rect 10347 22408 10348 22448
rect 10388 22408 10389 22448
rect 10347 22399 10389 22408
rect 12843 22448 12885 22457
rect 12843 22408 12844 22448
rect 12884 22408 12885 22448
rect 12843 22399 12885 22408
rect 17451 22448 17493 22457
rect 17451 22408 17452 22448
rect 17492 22408 17493 22448
rect 17451 22399 17493 22408
rect 30603 22448 30645 22457
rect 30603 22408 30604 22448
rect 30644 22408 30645 22448
rect 30603 22399 30645 22408
rect 30987 22448 31029 22457
rect 30987 22408 30988 22448
rect 31028 22408 31029 22448
rect 30987 22399 31029 22408
rect 747 22364 789 22373
rect 747 22324 748 22364
rect 788 22324 789 22364
rect 747 22315 789 22324
rect 4570 22364 4628 22365
rect 4570 22324 4579 22364
rect 4619 22324 4628 22364
rect 4570 22323 4628 22324
rect 5146 22364 5204 22365
rect 5146 22324 5155 22364
rect 5195 22324 5204 22364
rect 5146 22323 5204 22324
rect 5355 22364 5397 22373
rect 5355 22324 5356 22364
rect 5396 22324 5397 22364
rect 1450 22322 1508 22323
rect 1450 22282 1459 22322
rect 1499 22282 1508 22322
rect 5355 22315 5397 22324
rect 5570 22364 5612 22373
rect 5570 22324 5571 22364
rect 5611 22324 5612 22364
rect 5570 22315 5612 22324
rect 5835 22364 5877 22373
rect 7179 22364 7221 22373
rect 5835 22324 5836 22364
rect 5876 22324 5877 22364
rect 5835 22315 5877 22324
rect 6066 22355 6112 22364
rect 6066 22315 6067 22355
rect 6107 22315 6112 22355
rect 7179 22324 7180 22364
rect 7220 22324 7221 22364
rect 7179 22315 7221 22324
rect 7371 22364 7413 22373
rect 7371 22324 7372 22364
rect 7412 22324 7413 22364
rect 7371 22315 7413 22324
rect 7947 22364 7989 22373
rect 7947 22324 7948 22364
rect 7988 22324 7989 22364
rect 7947 22315 7989 22324
rect 8122 22364 8180 22365
rect 8122 22324 8131 22364
rect 8171 22324 8180 22364
rect 8122 22323 8180 22324
rect 8698 22364 8756 22365
rect 8698 22324 8707 22364
rect 8747 22324 8756 22364
rect 8698 22323 8756 22324
rect 12634 22364 12692 22365
rect 12634 22324 12643 22364
rect 12683 22324 12692 22364
rect 12634 22323 12692 22324
rect 14907 22364 14949 22373
rect 14907 22324 14908 22364
rect 14948 22324 14949 22364
rect 14907 22315 14949 22324
rect 16570 22364 16628 22365
rect 16570 22324 16579 22364
rect 16619 22324 16628 22364
rect 16570 22323 16628 22324
rect 16971 22364 17013 22373
rect 16971 22324 16972 22364
rect 17012 22324 17013 22364
rect 16971 22315 17013 22324
rect 17547 22364 17589 22373
rect 17547 22324 17548 22364
rect 17588 22324 17589 22364
rect 17547 22315 17589 22324
rect 21370 22364 21428 22365
rect 21370 22324 21379 22364
rect 21419 22324 21428 22364
rect 21370 22323 21428 22324
rect 22059 22364 22101 22373
rect 22059 22324 22060 22364
rect 22100 22324 22101 22364
rect 22059 22315 22101 22324
rect 6066 22306 6112 22315
rect 6689 22313 6747 22314
rect 1450 22281 1508 22282
rect 1803 22280 1845 22289
rect 1803 22240 1804 22280
rect 1844 22240 1845 22280
rect 1803 22231 1845 22240
rect 1947 22280 1989 22289
rect 1947 22240 1948 22280
rect 1988 22240 1989 22280
rect 1947 22231 1989 22240
rect 2571 22280 2613 22289
rect 2571 22240 2572 22280
rect 2612 22240 2613 22280
rect 2571 22231 2613 22240
rect 2955 22280 2997 22289
rect 2955 22240 2956 22280
rect 2996 22240 2997 22280
rect 2955 22231 2997 22240
rect 3514 22280 3572 22281
rect 3514 22240 3523 22280
rect 3563 22240 3572 22280
rect 3514 22239 3572 22240
rect 3627 22280 3669 22289
rect 3627 22240 3628 22280
rect 3668 22240 3669 22280
rect 3627 22231 3669 22240
rect 4054 22280 4096 22289
rect 4054 22240 4055 22280
rect 4095 22240 4096 22280
rect 4054 22231 4096 22240
rect 4186 22280 4244 22281
rect 4186 22240 4195 22280
rect 4235 22240 4244 22280
rect 4186 22239 4244 22240
rect 4299 22280 4341 22289
rect 4299 22240 4300 22280
rect 4340 22240 4341 22280
rect 4299 22231 4341 22240
rect 4954 22280 5012 22281
rect 4954 22240 4963 22280
rect 5003 22240 5012 22280
rect 4954 22239 5012 22240
rect 5451 22280 5493 22289
rect 5451 22240 5452 22280
rect 5492 22240 5493 22280
rect 5451 22231 5493 22240
rect 5668 22280 5710 22289
rect 5668 22240 5669 22280
rect 5709 22240 5710 22280
rect 5668 22231 5710 22240
rect 5931 22280 5973 22289
rect 5931 22240 5932 22280
rect 5972 22240 5973 22280
rect 5931 22231 5973 22240
rect 6160 22280 6218 22281
rect 6160 22240 6169 22280
rect 6209 22240 6218 22280
rect 6160 22239 6218 22240
rect 6400 22280 6442 22289
rect 6400 22240 6401 22280
rect 6441 22240 6442 22280
rect 6689 22273 6698 22313
rect 6738 22273 6747 22313
rect 25503 22313 25545 22322
rect 6689 22272 6747 22273
rect 6838 22280 6880 22289
rect 6400 22231 6442 22240
rect 6838 22240 6839 22280
rect 6879 22240 6880 22280
rect 6838 22231 6880 22240
rect 6970 22280 7028 22281
rect 6970 22240 6979 22280
rect 7019 22240 7028 22280
rect 6970 22239 7028 22240
rect 7083 22280 7125 22289
rect 7083 22240 7084 22280
rect 7124 22240 7125 22280
rect 7083 22231 7125 22240
rect 7546 22280 7604 22281
rect 7546 22240 7555 22280
rect 7595 22240 7604 22280
rect 7546 22239 7604 22240
rect 8506 22280 8564 22281
rect 8506 22240 8515 22280
rect 8555 22240 8564 22280
rect 8506 22239 8564 22240
rect 8938 22280 8996 22281
rect 8938 22240 8947 22280
rect 8987 22240 8996 22280
rect 8938 22239 8996 22240
rect 9867 22280 9909 22289
rect 9867 22240 9868 22280
rect 9908 22240 9909 22280
rect 9867 22231 9909 22240
rect 12250 22280 12308 22281
rect 12250 22240 12259 22280
rect 12299 22240 12308 22280
rect 12250 22239 12308 22240
rect 13233 22280 13291 22281
rect 13233 22240 13242 22280
rect 13282 22240 13291 22280
rect 13233 22239 13291 22240
rect 13515 22280 13557 22289
rect 13515 22240 13516 22280
rect 13556 22240 13557 22280
rect 13515 22231 13557 22240
rect 13978 22280 14036 22281
rect 13978 22240 13987 22280
rect 14027 22240 14036 22280
rect 13978 22239 14036 22240
rect 14698 22280 14756 22281
rect 14698 22240 14707 22280
rect 14747 22240 14756 22280
rect 14698 22239 14756 22240
rect 15243 22280 15285 22289
rect 15243 22240 15244 22280
rect 15284 22240 15285 22280
rect 15243 22231 15285 22240
rect 15387 22280 15429 22289
rect 15387 22240 15388 22280
rect 15428 22240 15429 22280
rect 15387 22231 15429 22240
rect 15531 22280 15573 22289
rect 15531 22240 15532 22280
rect 15572 22240 15573 22280
rect 15531 22231 15573 22240
rect 15706 22280 15764 22281
rect 15706 22240 15715 22280
rect 15755 22240 15764 22280
rect 15706 22239 15764 22240
rect 15819 22280 15861 22289
rect 15819 22240 15820 22280
rect 15860 22240 15861 22280
rect 15819 22231 15861 22240
rect 16011 22280 16053 22289
rect 16011 22240 16012 22280
rect 16052 22240 16053 22280
rect 16011 22231 16053 22240
rect 16142 22280 16200 22281
rect 16142 22240 16151 22280
rect 16191 22240 16200 22280
rect 16142 22239 16200 22240
rect 16252 22280 16310 22281
rect 16252 22240 16261 22280
rect 16301 22240 16310 22280
rect 16252 22239 16310 22240
rect 16450 22280 16508 22281
rect 16450 22240 16459 22280
rect 16499 22240 16508 22280
rect 16450 22239 16508 22240
rect 16683 22280 16725 22289
rect 16683 22240 16684 22280
rect 16724 22240 16725 22280
rect 16683 22231 16725 22240
rect 17146 22280 17204 22281
rect 17146 22240 17155 22280
rect 17195 22240 17204 22280
rect 17146 22239 17204 22240
rect 18027 22280 18069 22289
rect 18027 22240 18028 22280
rect 18068 22240 18069 22280
rect 18027 22231 18069 22240
rect 18607 22280 18665 22281
rect 18607 22240 18616 22280
rect 18656 22240 18665 22280
rect 18607 22239 18665 22240
rect 19162 22280 19220 22281
rect 19162 22240 19171 22280
rect 19211 22240 19220 22280
rect 19162 22239 19220 22240
rect 21238 22280 21280 22289
rect 21238 22240 21239 22280
rect 21279 22240 21280 22280
rect 21238 22231 21280 22240
rect 21483 22280 21525 22289
rect 21483 22240 21484 22280
rect 21524 22240 21525 22280
rect 21483 22231 21525 22240
rect 21867 22280 21909 22289
rect 21867 22240 21868 22280
rect 21908 22240 21909 22280
rect 21867 22231 21909 22240
rect 22426 22280 22484 22281
rect 22426 22240 22435 22280
rect 22475 22240 22484 22280
rect 22426 22239 22484 22240
rect 24939 22280 24981 22289
rect 24939 22240 24940 22280
rect 24980 22240 24981 22280
rect 25503 22273 25504 22313
rect 25544 22273 25545 22313
rect 25503 22264 25545 22273
rect 25594 22280 25652 22281
rect 24939 22231 24981 22240
rect 25594 22240 25603 22280
rect 25643 22240 25652 22280
rect 25594 22239 25652 22240
rect 25899 22280 25941 22289
rect 25899 22240 25900 22280
rect 25940 22240 25941 22280
rect 25899 22231 25941 22240
rect 26763 22280 26805 22289
rect 26763 22240 26764 22280
rect 26804 22240 26805 22280
rect 26763 22231 26805 22240
rect 26890 22280 26948 22281
rect 26890 22240 26899 22280
rect 26939 22240 26948 22280
rect 26890 22239 26948 22240
rect 26995 22280 27053 22281
rect 26995 22240 27004 22280
rect 27044 22240 27053 22280
rect 26995 22239 27053 22240
rect 29146 22280 29204 22281
rect 29146 22240 29155 22280
rect 29195 22240 29204 22280
rect 29146 22239 29204 22240
rect 29725 22280 29767 22289
rect 29725 22240 29726 22280
rect 29766 22240 29767 22280
rect 29725 22231 29767 22240
rect 30019 22280 30077 22281
rect 30019 22240 30028 22280
rect 30068 22240 30077 22280
rect 30019 22239 30077 22240
rect 30219 22280 30261 22289
rect 30219 22240 30220 22280
rect 30260 22240 30261 22280
rect 30219 22231 30261 22240
rect 30394 22280 30452 22281
rect 30394 22240 30403 22280
rect 30443 22240 30452 22280
rect 30394 22239 30452 22240
rect 1594 22196 1652 22197
rect 1594 22156 1603 22196
rect 1643 22156 1652 22196
rect 1594 22155 1652 22156
rect 4378 22196 4436 22197
rect 4378 22156 4387 22196
rect 4427 22156 4436 22196
rect 4378 22155 4436 22156
rect 7851 22196 7893 22205
rect 7851 22156 7852 22196
rect 7892 22156 7893 22196
rect 7851 22147 7893 22156
rect 13131 22196 13173 22205
rect 13131 22156 13132 22196
rect 13172 22156 13173 22196
rect 13131 22147 13173 22156
rect 14379 22196 14421 22205
rect 14379 22156 14380 22196
rect 14420 22156 14421 22196
rect 14379 22147 14421 22156
rect 15610 22196 15668 22197
rect 15610 22156 15619 22196
rect 15659 22156 15668 22196
rect 15610 22155 15668 22156
rect 18778 22196 18836 22197
rect 18778 22156 18787 22196
rect 18827 22156 18836 22196
rect 18778 22155 18836 22156
rect 27226 22196 27284 22197
rect 27226 22156 27235 22196
rect 27275 22156 27284 22196
rect 27226 22155 27284 22156
rect 29530 22196 29588 22197
rect 29530 22156 29539 22196
rect 29579 22156 29588 22196
rect 29530 22155 29588 22156
rect 987 22112 1029 22121
rect 987 22072 988 22112
rect 1028 22072 1029 22112
rect 987 22063 1029 22072
rect 1258 22112 1316 22113
rect 1258 22072 1267 22112
rect 1307 22072 1316 22112
rect 1258 22071 1316 22072
rect 1899 22112 1941 22121
rect 1899 22072 1900 22112
rect 1940 22072 1941 22112
rect 1899 22063 1941 22072
rect 3051 22112 3093 22121
rect 3051 22072 3052 22112
rect 3092 22072 3093 22112
rect 3051 22063 3093 22072
rect 3915 22112 3957 22121
rect 3915 22072 3916 22112
rect 3956 22072 3957 22112
rect 3915 22063 3957 22072
rect 4666 22112 4724 22113
rect 4666 22072 4675 22112
rect 4715 22072 4724 22112
rect 4666 22071 4724 22072
rect 6603 22112 6645 22121
rect 6603 22072 6604 22112
rect 6644 22072 6645 22112
rect 6603 22063 6645 22072
rect 9147 22112 9189 22121
rect 9147 22072 9148 22112
rect 9188 22072 9189 22112
rect 9147 22063 9189 22072
rect 9675 22112 9717 22121
rect 9675 22072 9676 22112
rect 9716 22072 9717 22112
rect 9675 22063 9717 22072
rect 9946 22112 10004 22113
rect 9946 22072 9955 22112
rect 9995 22072 10004 22112
rect 9946 22071 10004 22072
rect 16762 22112 16820 22113
rect 16762 22072 16771 22112
rect 16811 22072 16820 22112
rect 16762 22071 16820 22072
rect 17835 22112 17877 22121
rect 17835 22072 17836 22112
rect 17876 22072 17877 22112
rect 17835 22063 17877 22072
rect 18106 22112 18164 22113
rect 18106 22072 18115 22112
rect 18155 22072 18164 22112
rect 18106 22071 18164 22072
rect 18442 22112 18500 22113
rect 18442 22072 18451 22112
rect 18491 22072 18500 22112
rect 18442 22071 18500 22072
rect 21562 22112 21620 22113
rect 21562 22072 21571 22112
rect 21611 22072 21620 22112
rect 21562 22071 21620 22072
rect 24747 22112 24789 22121
rect 24747 22072 24748 22112
rect 24788 22072 24789 22112
rect 24747 22063 24789 22072
rect 25018 22112 25076 22113
rect 25018 22072 25027 22112
rect 25067 22072 25076 22112
rect 25018 22071 25076 22072
rect 25738 22112 25796 22113
rect 25738 22072 25747 22112
rect 25787 22072 25796 22112
rect 25738 22071 25796 22072
rect 29818 22112 29876 22113
rect 29818 22072 29827 22112
rect 29867 22072 29876 22112
rect 29818 22071 29876 22072
rect 29931 22112 29973 22121
rect 29931 22072 29932 22112
rect 29972 22072 29973 22112
rect 29931 22063 29973 22072
rect 30315 22112 30357 22121
rect 30315 22072 30316 22112
rect 30356 22072 30357 22112
rect 30315 22063 30357 22072
rect 576 21944 31392 21968
rect 576 21904 4352 21944
rect 4720 21904 12126 21944
rect 12494 21904 19900 21944
rect 20268 21904 27674 21944
rect 28042 21904 31392 21944
rect 576 21880 31392 21904
rect 874 21776 932 21777
rect 874 21736 883 21776
rect 923 21736 932 21776
rect 874 21735 932 21736
rect 5434 21776 5492 21777
rect 5434 21736 5443 21776
rect 5483 21736 5492 21776
rect 5434 21735 5492 21736
rect 5547 21776 5589 21785
rect 5547 21736 5548 21776
rect 5588 21736 5589 21776
rect 5547 21727 5589 21736
rect 6106 21776 6164 21777
rect 6106 21736 6115 21776
rect 6155 21736 6164 21776
rect 6106 21735 6164 21736
rect 6586 21776 6644 21777
rect 6586 21736 6595 21776
rect 6635 21736 6644 21776
rect 6586 21735 6644 21736
rect 6987 21776 7029 21785
rect 6987 21736 6988 21776
rect 7028 21736 7029 21776
rect 6987 21727 7029 21736
rect 7659 21776 7701 21785
rect 7659 21736 7660 21776
rect 7700 21736 7701 21776
rect 7659 21727 7701 21736
rect 9531 21776 9573 21785
rect 9531 21736 9532 21776
rect 9572 21736 9573 21776
rect 9531 21727 9573 21736
rect 11434 21776 11492 21777
rect 11434 21736 11443 21776
rect 11483 21736 11492 21776
rect 11434 21735 11492 21736
rect 13323 21776 13365 21785
rect 13323 21736 13324 21776
rect 13364 21736 13365 21776
rect 13323 21727 13365 21736
rect 15034 21776 15092 21777
rect 15034 21736 15043 21776
rect 15083 21736 15092 21776
rect 15034 21735 15092 21736
rect 18075 21776 18117 21785
rect 18075 21736 18076 21776
rect 18116 21736 18117 21776
rect 18075 21727 18117 21736
rect 18778 21776 18836 21777
rect 18778 21736 18787 21776
rect 18827 21736 18836 21776
rect 18778 21735 18836 21736
rect 24699 21776 24741 21785
rect 24699 21736 24700 21776
rect 24740 21736 24741 21776
rect 24699 21727 24741 21736
rect 25515 21776 25557 21785
rect 25515 21736 25516 21776
rect 25556 21736 25557 21776
rect 25515 21727 25557 21736
rect 28011 21776 28053 21785
rect 28011 21736 28012 21776
rect 28052 21736 28053 21776
rect 28011 21727 28053 21736
rect 5175 21692 5217 21701
rect 5175 21652 5176 21692
rect 5216 21652 5217 21692
rect 5175 21643 5217 21652
rect 5655 21692 5697 21701
rect 5655 21652 5656 21692
rect 5696 21652 5697 21692
rect 5655 21643 5697 21652
rect 6806 21692 6848 21701
rect 6806 21652 6807 21692
rect 6847 21652 6848 21692
rect 6806 21643 6848 21652
rect 8218 21692 8276 21693
rect 8218 21652 8227 21692
rect 8267 21652 8276 21692
rect 8218 21651 8276 21652
rect 9034 21692 9092 21693
rect 9034 21652 9043 21692
rect 9083 21652 9092 21692
rect 9034 21651 9092 21652
rect 10954 21692 11012 21693
rect 10954 21652 10963 21692
rect 11003 21652 11012 21692
rect 10954 21651 11012 21652
rect 16203 21692 16245 21701
rect 16203 21652 16204 21692
rect 16244 21652 16245 21692
rect 16203 21643 16245 21652
rect 16971 21692 17013 21701
rect 16971 21652 16972 21692
rect 17012 21652 17013 21692
rect 16971 21643 17013 21652
rect 17722 21692 17780 21693
rect 17722 21652 17731 21692
rect 17771 21652 17780 21692
rect 17722 21651 17780 21652
rect 20619 21692 20661 21701
rect 20619 21652 20620 21692
rect 20660 21652 20661 21692
rect 20619 21643 20661 21652
rect 25323 21692 25365 21701
rect 25323 21652 25324 21692
rect 25364 21652 25365 21692
rect 23962 21650 24020 21651
rect 1066 21608 1124 21609
rect 1066 21568 1075 21608
rect 1115 21568 1124 21608
rect 1306 21608 1364 21609
rect 1066 21567 1124 21568
rect 1179 21566 1221 21575
rect 1306 21568 1315 21608
rect 1355 21568 1364 21608
rect 1306 21567 1364 21568
rect 1419 21608 1461 21617
rect 1419 21568 1420 21608
rect 1460 21568 1461 21608
rect 1179 21526 1180 21566
rect 1220 21526 1221 21566
rect 1419 21559 1461 21568
rect 1786 21608 1844 21609
rect 1786 21568 1795 21608
rect 1835 21568 1844 21608
rect 1786 21567 1844 21568
rect 2571 21608 2613 21617
rect 2571 21568 2572 21608
rect 2612 21568 2613 21608
rect 2571 21559 2613 21568
rect 2800 21608 2858 21609
rect 2800 21568 2809 21608
rect 2849 21568 2858 21608
rect 2800 21567 2858 21568
rect 2955 21608 2997 21617
rect 2955 21568 2956 21608
rect 2996 21568 2997 21608
rect 2955 21559 2997 21568
rect 3130 21608 3188 21609
rect 3130 21568 3139 21608
rect 3179 21568 3188 21608
rect 3130 21567 3188 21568
rect 3514 21608 3572 21609
rect 3514 21568 3523 21608
rect 3563 21568 3572 21608
rect 3514 21567 3572 21568
rect 3637 21608 3679 21617
rect 3637 21568 3638 21608
rect 3678 21568 3679 21608
rect 3637 21559 3679 21568
rect 4354 21608 4412 21609
rect 4354 21568 4363 21608
rect 4403 21568 4412 21608
rect 4354 21567 4412 21568
rect 4587 21608 4629 21617
rect 4587 21568 4588 21608
rect 4628 21568 4629 21608
rect 4587 21559 4629 21568
rect 4856 21608 4914 21609
rect 4856 21568 4865 21608
rect 4905 21568 4914 21608
rect 4856 21567 4914 21568
rect 4971 21608 5013 21617
rect 4971 21568 4972 21608
rect 5012 21568 5013 21608
rect 4971 21559 5013 21568
rect 5338 21608 5396 21609
rect 5338 21568 5347 21608
rect 5387 21568 5396 21608
rect 5338 21567 5396 21568
rect 5794 21608 5852 21609
rect 5794 21568 5803 21608
rect 5843 21568 5852 21608
rect 6490 21608 6548 21609
rect 5794 21567 5852 21568
rect 6027 21566 6069 21575
rect 6490 21568 6499 21608
rect 6539 21568 6548 21608
rect 6490 21567 6548 21568
rect 7083 21608 7125 21617
rect 7083 21568 7084 21608
rect 7124 21568 7125 21608
rect 1179 21517 1221 21526
rect 1515 21524 1557 21533
rect 1515 21484 1516 21524
rect 1556 21484 1557 21524
rect 1515 21475 1557 21484
rect 2475 21524 2517 21533
rect 2475 21484 2476 21524
rect 2516 21484 2517 21524
rect 2475 21475 2517 21484
rect 2690 21524 2732 21533
rect 2690 21484 2691 21524
rect 2731 21484 2732 21524
rect 2690 21475 2732 21484
rect 4474 21524 4532 21525
rect 4474 21484 4483 21524
rect 4523 21484 4532 21524
rect 4474 21483 4532 21484
rect 4683 21524 4725 21533
rect 4683 21484 4684 21524
rect 4724 21484 4725 21524
rect 4683 21475 4725 21484
rect 5908 21524 5950 21533
rect 5908 21484 5909 21524
rect 5949 21484 5950 21524
rect 6027 21526 6028 21566
rect 6068 21526 6069 21566
rect 7083 21559 7125 21568
rect 7300 21608 7342 21617
rect 7300 21568 7301 21608
rect 7341 21568 7342 21608
rect 7300 21559 7342 21568
rect 7453 21608 7495 21617
rect 8139 21608 8181 21617
rect 7453 21568 7454 21608
rect 7494 21568 7495 21608
rect 7453 21559 7495 21568
rect 7755 21599 7797 21608
rect 7755 21559 7756 21599
rect 7796 21559 7797 21599
rect 7755 21550 7797 21559
rect 7899 21566 7941 21575
rect 6027 21517 6069 21526
rect 7202 21524 7244 21533
rect 5908 21475 5950 21484
rect 7202 21484 7203 21524
rect 7243 21484 7244 21524
rect 7899 21526 7900 21566
rect 7940 21526 7941 21566
rect 8139 21568 8140 21608
rect 8180 21568 8181 21608
rect 8139 21559 8181 21568
rect 8719 21608 8777 21609
rect 8719 21568 8728 21608
rect 8768 21568 8777 21608
rect 8719 21567 8777 21568
rect 9229 21608 9287 21609
rect 11119 21608 11177 21609
rect 9229 21568 9238 21608
rect 9278 21568 9287 21608
rect 9229 21567 9287 21568
rect 9378 21599 9424 21608
rect 9378 21559 9379 21599
rect 9419 21559 9424 21599
rect 9378 21550 9424 21559
rect 9858 21599 9904 21608
rect 9858 21559 9859 21599
rect 9899 21559 9904 21599
rect 9858 21550 9904 21559
rect 10338 21599 10384 21608
rect 10338 21559 10339 21599
rect 10379 21559 10384 21599
rect 11119 21568 11128 21608
rect 11168 21568 11177 21608
rect 11119 21567 11177 21568
rect 11599 21608 11657 21609
rect 11599 21568 11608 21608
rect 11648 21568 11657 21608
rect 11599 21567 11657 21568
rect 11787 21608 11829 21617
rect 11787 21568 11788 21608
rect 11828 21568 11829 21608
rect 11787 21559 11829 21568
rect 12843 21608 12885 21617
rect 12843 21568 12844 21608
rect 12884 21568 12885 21608
rect 12843 21559 12885 21568
rect 13227 21608 13269 21617
rect 13227 21568 13228 21608
rect 13268 21568 13269 21608
rect 13227 21559 13269 21568
rect 13654 21608 13696 21617
rect 13654 21568 13655 21608
rect 13695 21568 13696 21608
rect 13654 21559 13696 21568
rect 13899 21608 13941 21617
rect 13899 21568 13900 21608
rect 13940 21568 13941 21608
rect 13899 21559 13941 21568
rect 14362 21608 14420 21609
rect 14362 21568 14371 21608
rect 14411 21568 14420 21608
rect 14362 21567 14420 21568
rect 15322 21608 15380 21609
rect 15322 21568 15331 21608
rect 15371 21568 15380 21608
rect 15322 21567 15380 21568
rect 15723 21608 15765 21617
rect 15723 21568 15724 21608
rect 15764 21568 15765 21608
rect 15723 21559 15765 21568
rect 15915 21608 15957 21617
rect 15915 21568 15916 21608
rect 15956 21568 15957 21608
rect 15915 21559 15957 21568
rect 16107 21608 16149 21617
rect 16107 21568 16108 21608
rect 16148 21568 16149 21608
rect 16107 21559 16149 21568
rect 16299 21608 16341 21617
rect 16299 21568 16300 21608
rect 16340 21568 16341 21608
rect 16299 21559 16341 21568
rect 16587 21608 16629 21617
rect 16587 21568 16588 21608
rect 16628 21568 16629 21608
rect 16587 21559 16629 21568
rect 16779 21608 16821 21617
rect 16779 21568 16780 21608
rect 16820 21568 16821 21608
rect 16779 21559 16821 21568
rect 17067 21608 17109 21617
rect 17067 21568 17068 21608
rect 17108 21568 17109 21608
rect 17067 21559 17109 21568
rect 17296 21608 17354 21609
rect 17296 21568 17305 21608
rect 17345 21568 17354 21608
rect 17296 21567 17354 21568
rect 17410 21608 17468 21609
rect 17410 21568 17419 21608
rect 17459 21568 17468 21608
rect 17410 21567 17468 21568
rect 17643 21608 17685 21617
rect 18891 21608 18933 21617
rect 17643 21568 17644 21608
rect 17684 21568 17685 21608
rect 17643 21559 17685 21568
rect 17922 21599 17968 21608
rect 17922 21559 17923 21599
rect 17963 21559 17968 21599
rect 18891 21568 18892 21608
rect 18932 21568 18933 21608
rect 18891 21559 18933 21568
rect 19851 21608 19893 21617
rect 19851 21568 19852 21608
rect 19892 21568 19893 21608
rect 19851 21559 19893 21568
rect 20235 21608 20277 21617
rect 20235 21568 20236 21608
rect 20276 21568 20277 21608
rect 20235 21559 20277 21568
rect 20506 21608 20564 21609
rect 20506 21568 20515 21608
rect 20555 21568 20564 21608
rect 20506 21567 20564 21568
rect 21099 21608 21141 21617
rect 21099 21568 21100 21608
rect 21140 21568 21141 21608
rect 21099 21559 21141 21568
rect 21466 21608 21524 21609
rect 21466 21568 21475 21608
rect 21515 21568 21524 21608
rect 21466 21567 21524 21568
rect 23595 21608 23637 21617
rect 23962 21610 23971 21650
rect 24011 21610 24020 21650
rect 25323 21643 25365 21652
rect 23962 21609 24020 21610
rect 23595 21568 23596 21608
rect 23636 21568 23637 21608
rect 23595 21559 23637 21568
rect 23770 21608 23828 21609
rect 23770 21568 23779 21608
rect 23819 21568 23828 21608
rect 23770 21567 23828 21568
rect 24096 21608 24138 21617
rect 24096 21568 24097 21608
rect 24137 21568 24138 21608
rect 24096 21559 24138 21568
rect 24394 21608 24452 21609
rect 25114 21608 25172 21609
rect 24394 21568 24403 21608
rect 24443 21568 24452 21608
rect 24394 21567 24452 21568
rect 24546 21599 24592 21608
rect 24546 21559 24547 21599
rect 24587 21559 24592 21599
rect 25114 21568 25123 21608
rect 25163 21568 25172 21608
rect 25114 21567 25172 21568
rect 27418 21608 27476 21609
rect 27418 21568 27427 21608
rect 27467 21568 27476 21608
rect 27418 21567 27476 21568
rect 27802 21608 27860 21609
rect 27802 21568 27811 21608
rect 27851 21568 27860 21608
rect 27802 21567 27860 21568
rect 29914 21608 29972 21609
rect 29914 21568 29923 21608
rect 29963 21568 29972 21608
rect 29914 21567 29972 21568
rect 30298 21608 30356 21609
rect 30298 21568 30307 21608
rect 30347 21568 30356 21608
rect 30298 21567 30356 21568
rect 10338 21550 10384 21559
rect 17922 21550 17968 21559
rect 24546 21550 24592 21559
rect 7899 21517 7941 21526
rect 8026 21524 8084 21525
rect 7202 21475 7244 21484
rect 8026 21484 8035 21524
rect 8075 21484 8084 21524
rect 8026 21483 8084 21484
rect 8554 21524 8612 21525
rect 8554 21484 8563 21524
rect 8603 21484 8612 21524
rect 8554 21483 8612 21484
rect 10011 21524 10053 21533
rect 10011 21484 10012 21524
rect 10052 21484 10053 21524
rect 10011 21475 10053 21484
rect 10491 21524 10533 21533
rect 10491 21484 10492 21524
rect 10532 21484 10533 21524
rect 10491 21475 10533 21484
rect 13786 21524 13844 21525
rect 13786 21484 13795 21524
rect 13835 21484 13844 21524
rect 13786 21483 13844 21484
rect 13995 21524 14037 21533
rect 13995 21484 13996 21524
rect 14036 21484 14037 21524
rect 13995 21475 14037 21484
rect 14187 21524 14229 21533
rect 14187 21484 14188 21524
rect 14228 21484 14229 21524
rect 14187 21475 14229 21484
rect 14763 21524 14805 21533
rect 14763 21484 14764 21524
rect 14804 21484 14805 21524
rect 14763 21475 14805 21484
rect 14938 21524 14996 21525
rect 14938 21484 14947 21524
rect 14987 21484 14996 21524
rect 14938 21483 14996 21484
rect 15514 21524 15572 21525
rect 15514 21484 15523 21524
rect 15563 21484 15572 21524
rect 15514 21483 15572 21484
rect 17186 21524 17228 21533
rect 17186 21484 17187 21524
rect 17227 21484 17228 21524
rect 17186 21475 17228 21484
rect 17530 21524 17588 21525
rect 17530 21484 17539 21524
rect 17579 21484 17588 21524
rect 17530 21483 17588 21484
rect 18603 21524 18645 21533
rect 18603 21484 18604 21524
rect 18644 21484 18645 21524
rect 18603 21475 18645 21484
rect 19450 21524 19508 21525
rect 19450 21484 19459 21524
rect 19499 21484 19508 21524
rect 19450 21483 19508 21484
rect 24267 21524 24309 21533
rect 24267 21484 24268 21524
rect 24308 21484 24309 21524
rect 24267 21475 24309 21484
rect 14667 21440 14709 21449
rect 14667 21400 14668 21440
rect 14708 21400 14709 21440
rect 14667 21391 14709 21400
rect 23403 21440 23445 21449
rect 23403 21400 23404 21440
rect 23444 21400 23445 21440
rect 23403 21391 23445 21400
rect 24171 21440 24213 21449
rect 24171 21400 24172 21440
rect 24212 21400 24213 21440
rect 24171 21391 24213 21400
rect 25094 21440 25136 21449
rect 25094 21400 25095 21440
rect 25135 21400 25136 21440
rect 25094 21391 25136 21400
rect 30507 21440 30549 21449
rect 30507 21400 30508 21440
rect 30548 21400 30549 21440
rect 30507 21391 30549 21400
rect 30891 21440 30933 21449
rect 30891 21400 30892 21440
rect 30932 21400 30933 21440
rect 30891 21391 30933 21400
rect 2187 21356 2229 21365
rect 2187 21316 2188 21356
rect 2228 21316 2229 21356
rect 2187 21307 2229 21316
rect 3130 21356 3188 21357
rect 3130 21316 3139 21356
rect 3179 21316 3188 21356
rect 3130 21315 3188 21316
rect 3802 21356 3860 21357
rect 3802 21316 3811 21356
rect 3851 21316 3860 21356
rect 3802 21315 3860 21316
rect 5163 21356 5205 21365
rect 5163 21316 5164 21356
rect 5204 21316 5205 21356
rect 5163 21307 5205 21316
rect 6795 21356 6837 21365
rect 6795 21316 6796 21356
rect 6836 21316 6837 21356
rect 6795 21307 6837 21316
rect 7450 21356 7508 21357
rect 7450 21316 7459 21356
rect 7499 21316 7508 21356
rect 7450 21315 7508 21316
rect 12459 21356 12501 21365
rect 12459 21316 12460 21356
rect 12500 21316 12501 21356
rect 12459 21307 12501 21316
rect 15723 21356 15765 21365
rect 15723 21316 15724 21356
rect 15764 21316 15765 21356
rect 15723 21307 15765 21316
rect 16587 21356 16629 21365
rect 16587 21316 16588 21356
rect 16628 21316 16629 21356
rect 16587 21307 16629 21316
rect 18363 21356 18405 21365
rect 18363 21316 18364 21356
rect 18404 21316 18405 21356
rect 18363 21307 18405 21316
rect 19083 21356 19125 21365
rect 19083 21316 19084 21356
rect 19124 21316 19125 21356
rect 19083 21307 19125 21316
rect 20907 21356 20949 21365
rect 20907 21316 20908 21356
rect 20948 21316 20949 21356
rect 20907 21307 20949 21316
rect 23770 21356 23828 21357
rect 23770 21316 23779 21356
rect 23819 21316 23828 21356
rect 23770 21315 23828 21316
rect 576 21188 31392 21212
rect 576 21148 3112 21188
rect 3480 21148 10886 21188
rect 11254 21148 18660 21188
rect 19028 21148 26434 21188
rect 26802 21148 31392 21188
rect 576 21124 31392 21148
rect 6315 21020 6357 21029
rect 6315 20980 6316 21020
rect 6356 20980 6357 21020
rect 6315 20971 6357 20980
rect 7930 21020 7988 21021
rect 7930 20980 7939 21020
rect 7979 20980 7988 21020
rect 7930 20979 7988 20980
rect 9003 21020 9045 21029
rect 9003 20980 9004 21020
rect 9044 20980 9045 21020
rect 9003 20971 9045 20980
rect 10347 21020 10389 21029
rect 10347 20980 10348 21020
rect 10388 20980 10389 21020
rect 10347 20971 10389 20980
rect 24555 21020 24597 21029
rect 24555 20980 24556 21020
rect 24596 20980 24597 21020
rect 24555 20971 24597 20980
rect 25227 21020 25269 21029
rect 25227 20980 25228 21020
rect 25268 20980 25269 21020
rect 25227 20971 25269 20980
rect 29739 21020 29781 21029
rect 29739 20980 29740 21020
rect 29780 20980 29781 21020
rect 29739 20971 29781 20980
rect 30075 21020 30117 21029
rect 30075 20980 30076 21020
rect 30116 20980 30117 21020
rect 30075 20971 30117 20980
rect 30507 21020 30549 21029
rect 30507 20980 30508 21020
rect 30548 20980 30549 21020
rect 30507 20971 30549 20980
rect 1803 20936 1845 20945
rect 1803 20896 1804 20936
rect 1844 20896 1845 20936
rect 1803 20887 1845 20896
rect 2170 20936 2228 20937
rect 2170 20896 2179 20936
rect 2219 20896 2228 20936
rect 2170 20895 2228 20896
rect 5067 20936 5109 20945
rect 5067 20896 5068 20936
rect 5108 20896 5109 20936
rect 5067 20887 5109 20896
rect 9771 20936 9813 20945
rect 9771 20896 9772 20936
rect 9812 20896 9813 20936
rect 9771 20887 9813 20896
rect 14763 20936 14805 20945
rect 14763 20896 14764 20936
rect 14804 20896 14805 20936
rect 14763 20887 14805 20896
rect 20794 20936 20852 20937
rect 20794 20896 20803 20936
rect 20843 20896 20852 20936
rect 20794 20895 20852 20896
rect 27243 20936 27285 20945
rect 27243 20896 27244 20936
rect 27284 20896 27285 20936
rect 27243 20887 27285 20896
rect 30891 20936 30933 20945
rect 30891 20896 30892 20936
rect 30932 20896 30933 20936
rect 30891 20887 30933 20896
rect 843 20852 885 20861
rect 1323 20852 1365 20861
rect 843 20812 844 20852
rect 884 20812 885 20852
rect 843 20803 885 20812
rect 1074 20843 1120 20852
rect 1074 20803 1075 20843
rect 1115 20803 1120 20843
rect 1323 20812 1324 20852
rect 1364 20812 1365 20852
rect 1323 20803 1365 20812
rect 1899 20852 1941 20861
rect 1899 20812 1900 20852
rect 1940 20812 1941 20852
rect 1899 20803 1941 20812
rect 2074 20852 2132 20853
rect 2074 20812 2083 20852
rect 2123 20812 2132 20852
rect 2074 20811 2132 20812
rect 2650 20852 2708 20853
rect 5386 20852 5444 20853
rect 2650 20812 2659 20852
rect 2699 20812 2708 20852
rect 2650 20811 2708 20812
rect 3666 20843 3712 20852
rect 3666 20803 3667 20843
rect 3707 20803 3712 20843
rect 5386 20812 5395 20852
rect 5435 20812 5444 20852
rect 5386 20811 5444 20812
rect 7275 20852 7317 20861
rect 7275 20812 7276 20852
rect 7316 20812 7317 20852
rect 7275 20803 7317 20812
rect 9387 20852 9429 20861
rect 9387 20812 9388 20852
rect 9428 20812 9429 20852
rect 13396 20852 13438 20861
rect 9387 20803 9429 20812
rect 12795 20810 12837 20819
rect 1074 20794 1120 20803
rect 3666 20794 3712 20803
rect 8043 20779 8085 20788
rect 939 20768 981 20777
rect 939 20728 940 20768
rect 980 20728 981 20768
rect 939 20719 981 20728
rect 1168 20768 1226 20769
rect 1168 20728 1177 20768
rect 1217 20728 1226 20768
rect 1168 20727 1226 20728
rect 1498 20768 1556 20769
rect 1498 20728 1507 20768
rect 1547 20728 1556 20768
rect 1498 20727 1556 20728
rect 2458 20768 2516 20769
rect 2458 20728 2467 20768
rect 2507 20728 2516 20768
rect 2458 20727 2516 20728
rect 3181 20768 3239 20769
rect 3181 20728 3190 20768
rect 3230 20728 3239 20768
rect 3181 20727 3239 20728
rect 3531 20768 3573 20777
rect 3531 20728 3532 20768
rect 3572 20728 3573 20768
rect 3531 20719 3573 20728
rect 3760 20768 3818 20769
rect 3760 20728 3769 20768
rect 3809 20728 3818 20768
rect 3760 20727 3818 20728
rect 4090 20768 4148 20769
rect 4090 20728 4099 20768
rect 4139 20728 4148 20768
rect 4090 20727 4148 20728
rect 4203 20768 4245 20777
rect 4203 20728 4204 20768
rect 4244 20728 4245 20768
rect 4203 20719 4245 20728
rect 5581 20768 5639 20769
rect 5581 20728 5590 20768
rect 5630 20728 5639 20768
rect 5581 20727 5639 20728
rect 5835 20768 5877 20777
rect 5835 20728 5836 20768
rect 5876 20728 5877 20768
rect 5835 20719 5877 20728
rect 6010 20768 6068 20769
rect 6010 20728 6019 20768
rect 6059 20728 6068 20768
rect 6010 20727 6068 20728
rect 6210 20768 6268 20769
rect 6210 20728 6219 20768
rect 6259 20728 6268 20768
rect 6210 20727 6268 20728
rect 6411 20768 6453 20777
rect 6411 20728 6412 20768
rect 6452 20728 6453 20768
rect 6411 20719 6453 20728
rect 6603 20768 6645 20777
rect 6603 20728 6604 20768
rect 6644 20728 6645 20768
rect 6603 20719 6645 20728
rect 6778 20768 6836 20769
rect 6778 20728 6787 20768
rect 6827 20728 6836 20768
rect 6778 20727 6836 20728
rect 6946 20768 7004 20769
rect 6946 20728 6955 20768
rect 6995 20728 7004 20768
rect 6946 20727 7004 20728
rect 7066 20768 7124 20769
rect 7066 20728 7075 20768
rect 7115 20728 7124 20768
rect 7066 20727 7124 20728
rect 7179 20768 7221 20777
rect 7179 20728 7180 20768
rect 7220 20728 7221 20768
rect 7179 20719 7221 20728
rect 7611 20768 7653 20777
rect 7611 20728 7612 20768
rect 7652 20728 7653 20768
rect 7611 20719 7653 20728
rect 7755 20768 7797 20777
rect 7755 20728 7756 20768
rect 7796 20728 7797 20768
rect 7755 20719 7797 20728
rect 7930 20768 7988 20769
rect 7930 20728 7939 20768
rect 7979 20728 7988 20768
rect 8043 20739 8044 20779
rect 8084 20739 8085 20779
rect 8043 20730 8085 20739
rect 8180 20768 8238 20769
rect 7930 20727 7988 20728
rect 8180 20728 8189 20768
rect 8229 20728 8238 20768
rect 8180 20727 8238 20728
rect 8314 20768 8372 20769
rect 8314 20728 8323 20768
rect 8363 20728 8372 20768
rect 8314 20727 8372 20728
rect 8491 20768 8549 20769
rect 8491 20728 8500 20768
rect 8540 20728 8549 20768
rect 8491 20727 8549 20728
rect 8698 20768 8756 20769
rect 8698 20728 8707 20768
rect 8747 20728 8756 20768
rect 8698 20727 8756 20728
rect 9675 20768 9717 20777
rect 9675 20728 9676 20768
rect 9716 20728 9717 20768
rect 9675 20719 9717 20728
rect 9867 20768 9909 20777
rect 9867 20728 9868 20768
rect 9908 20728 9909 20768
rect 9867 20719 9909 20728
rect 10155 20768 10197 20777
rect 10155 20728 10156 20768
rect 10196 20728 10197 20768
rect 10155 20719 10197 20728
rect 11019 20768 11061 20777
rect 12795 20770 12796 20810
rect 12836 20770 12837 20810
rect 13396 20812 13397 20852
rect 13437 20812 13438 20852
rect 13396 20803 13438 20812
rect 14091 20852 14133 20861
rect 14091 20812 14092 20852
rect 14132 20812 14133 20852
rect 14091 20803 14133 20812
rect 14283 20852 14325 20861
rect 14283 20812 14284 20852
rect 14324 20812 14325 20852
rect 14283 20803 14325 20812
rect 14859 20852 14901 20861
rect 14859 20812 14860 20852
rect 14900 20812 14901 20852
rect 14859 20803 14901 20812
rect 15130 20852 15188 20853
rect 15130 20812 15139 20852
rect 15179 20812 15188 20852
rect 15130 20811 15188 20812
rect 15339 20852 15381 20861
rect 15339 20812 15340 20852
rect 15380 20812 15381 20852
rect 15339 20803 15381 20812
rect 17067 20852 17109 20861
rect 17067 20812 17068 20852
rect 17108 20812 17109 20852
rect 17067 20803 17109 20812
rect 17242 20852 17300 20853
rect 17242 20812 17251 20852
rect 17291 20812 17300 20852
rect 17242 20811 17300 20812
rect 17818 20852 17876 20853
rect 17818 20812 17827 20852
rect 17867 20812 17876 20852
rect 17818 20811 17876 20812
rect 18010 20852 18068 20853
rect 18010 20812 18019 20852
rect 18059 20812 18068 20852
rect 18010 20811 18068 20812
rect 18586 20852 18644 20853
rect 18586 20812 18595 20852
rect 18635 20812 18644 20852
rect 18586 20811 18644 20812
rect 23194 20852 23252 20853
rect 23194 20812 23203 20852
rect 23243 20812 23252 20852
rect 23194 20811 23252 20812
rect 30315 20852 30357 20861
rect 30315 20812 30316 20852
rect 30356 20812 30357 20852
rect 19266 20801 19312 20810
rect 11019 20728 11020 20768
rect 11060 20728 11061 20768
rect 11019 20719 11061 20728
rect 11695 20768 11753 20769
rect 11695 20728 11704 20768
rect 11744 20728 11753 20768
rect 11695 20727 11753 20728
rect 11863 20768 11921 20769
rect 11863 20728 11872 20768
rect 11912 20728 11921 20768
rect 11863 20727 11921 20728
rect 12313 20768 12371 20769
rect 12313 20728 12322 20768
rect 12362 20728 12371 20768
rect 12795 20761 12837 20770
rect 12922 20768 12980 20769
rect 12313 20727 12371 20728
rect 12922 20728 12931 20768
rect 12971 20728 12980 20768
rect 12922 20727 12980 20728
rect 13035 20768 13077 20777
rect 13035 20728 13036 20768
rect 13076 20728 13077 20768
rect 13035 20719 13077 20728
rect 13282 20768 13340 20769
rect 13282 20728 13291 20768
rect 13331 20728 13340 20768
rect 13282 20727 13340 20728
rect 13513 20768 13555 20777
rect 13513 20728 13514 20768
rect 13554 20728 13555 20768
rect 13513 20719 13555 20728
rect 13750 20768 13792 20777
rect 13750 20728 13751 20768
rect 13791 20728 13792 20768
rect 13750 20719 13792 20728
rect 13882 20768 13940 20769
rect 13882 20728 13891 20768
rect 13931 20728 13940 20768
rect 13882 20727 13940 20728
rect 13995 20768 14037 20777
rect 13995 20728 13996 20768
rect 14036 20728 14037 20768
rect 13995 20719 14037 20728
rect 14458 20768 14516 20769
rect 14458 20728 14467 20768
rect 14507 20728 14516 20768
rect 14458 20727 14516 20728
rect 14998 20768 15040 20777
rect 14998 20728 14999 20768
rect 15039 20728 15040 20768
rect 14998 20719 15040 20728
rect 15243 20768 15285 20777
rect 15243 20728 15244 20768
rect 15284 20728 15285 20768
rect 15243 20719 15285 20728
rect 16111 20768 16169 20769
rect 16111 20728 16120 20768
rect 16160 20728 16169 20768
rect 16111 20727 16169 20728
rect 16294 20768 16336 20777
rect 16294 20728 16295 20768
rect 16335 20728 16336 20768
rect 16294 20719 16336 20728
rect 16474 20768 16532 20769
rect 16474 20728 16483 20768
rect 16523 20728 16532 20768
rect 16474 20727 16532 20728
rect 16726 20768 16768 20777
rect 16726 20728 16727 20768
rect 16767 20728 16768 20768
rect 16726 20719 16768 20728
rect 16858 20768 16916 20769
rect 16858 20728 16867 20768
rect 16907 20728 16916 20768
rect 16858 20727 16916 20728
rect 16971 20768 17013 20777
rect 16971 20728 16972 20768
rect 17012 20728 17013 20768
rect 16971 20719 17013 20728
rect 17626 20768 17684 20769
rect 17626 20728 17635 20768
rect 17675 20728 17684 20768
rect 17626 20727 17684 20728
rect 18394 20768 18452 20769
rect 18394 20728 18403 20768
rect 18443 20728 18452 20768
rect 18394 20727 18452 20728
rect 18730 20768 18788 20769
rect 18730 20728 18739 20768
rect 18779 20728 18788 20768
rect 19266 20761 19267 20801
rect 19307 20761 19312 20801
rect 21087 20801 21129 20810
rect 30315 20803 30357 20812
rect 19266 20752 19312 20761
rect 20032 20768 20074 20777
rect 18730 20727 18788 20728
rect 20032 20728 20033 20768
rect 20073 20728 20074 20768
rect 20032 20719 20074 20728
rect 20323 20768 20381 20769
rect 20323 20728 20332 20768
rect 20372 20728 20381 20768
rect 20323 20727 20381 20728
rect 20619 20768 20661 20777
rect 20619 20728 20620 20768
rect 20660 20728 20661 20768
rect 21087 20761 21088 20801
rect 21128 20761 21129 20801
rect 21087 20752 21129 20761
rect 21178 20768 21236 20769
rect 20619 20719 20661 20728
rect 21178 20728 21187 20768
rect 21227 20728 21236 20768
rect 21178 20727 21236 20728
rect 21660 20768 21702 20777
rect 21660 20728 21661 20768
rect 21701 20728 21702 20768
rect 21660 20719 21702 20728
rect 21771 20768 21813 20777
rect 21771 20728 21772 20768
rect 21812 20728 21813 20768
rect 21771 20719 21813 20728
rect 22347 20768 22389 20777
rect 22347 20728 22348 20768
rect 22388 20728 22389 20768
rect 22347 20719 22389 20728
rect 22466 20768 22508 20777
rect 22466 20728 22467 20768
rect 22507 20728 22508 20768
rect 22466 20719 22508 20728
rect 22576 20768 22634 20769
rect 22576 20728 22585 20768
rect 22625 20728 22634 20768
rect 22576 20727 22634 20728
rect 23403 20768 23445 20777
rect 23403 20728 23404 20768
rect 23444 20728 23445 20768
rect 23403 20719 23445 20728
rect 23626 20768 23684 20769
rect 23626 20728 23635 20768
rect 23675 20728 23684 20768
rect 23626 20727 23684 20728
rect 23835 20768 23877 20777
rect 23835 20728 23836 20768
rect 23876 20728 23877 20768
rect 23835 20719 23877 20728
rect 24250 20768 24308 20769
rect 24250 20728 24259 20768
rect 24299 20728 24308 20768
rect 24250 20727 24308 20728
rect 24922 20768 24980 20769
rect 24922 20728 24931 20768
rect 24971 20728 24980 20768
rect 24922 20727 24980 20728
rect 25241 20768 25283 20777
rect 25241 20728 25242 20768
rect 25282 20728 25283 20768
rect 25241 20719 25283 20728
rect 26091 20768 26133 20777
rect 26091 20728 26092 20768
rect 26132 20728 26133 20768
rect 26091 20719 26133 20728
rect 26379 20768 26421 20777
rect 26379 20728 26380 20768
rect 26420 20728 26421 20768
rect 26379 20719 26421 20728
rect 29146 20768 29204 20769
rect 29146 20728 29155 20768
rect 29195 20728 29204 20768
rect 29146 20727 29204 20728
rect 29739 20768 29781 20777
rect 29739 20728 29740 20768
rect 29780 20728 29781 20768
rect 29739 20719 29781 20728
rect 29931 20768 29973 20777
rect 29931 20728 29932 20768
rect 29972 20728 29973 20768
rect 29931 20719 29973 20728
rect 30507 20768 30549 20777
rect 30507 20728 30508 20768
rect 30548 20728 30549 20768
rect 30507 20719 30549 20728
rect 30699 20768 30741 20777
rect 30699 20728 30700 20768
rect 30740 20728 30741 20768
rect 30699 20719 30741 20728
rect 9014 20684 9056 20693
rect 9014 20644 9015 20684
rect 9055 20644 9056 20684
rect 9014 20635 9056 20644
rect 13114 20684 13172 20685
rect 13114 20644 13123 20684
rect 13163 20644 13172 20684
rect 13114 20643 13172 20644
rect 15946 20684 16004 20685
rect 15946 20644 15955 20684
rect 15995 20644 16004 20684
rect 15946 20643 16004 20644
rect 19419 20684 19461 20693
rect 19419 20644 19420 20684
rect 19460 20644 19461 20684
rect 19419 20635 19461 20644
rect 24363 20684 24405 20693
rect 24363 20644 24364 20684
rect 24404 20644 24405 20684
rect 24363 20635 24405 20644
rect 24569 20684 24611 20693
rect 24569 20644 24570 20684
rect 24610 20644 24611 20684
rect 24569 20635 24611 20644
rect 27051 20684 27093 20693
rect 27051 20644 27052 20684
rect 27092 20644 27093 20684
rect 27051 20635 27093 20644
rect 29530 20684 29588 20685
rect 29530 20644 29539 20684
rect 29579 20644 29588 20684
rect 29530 20643 29588 20644
rect 2986 20600 3044 20601
rect 2986 20560 2995 20600
rect 3035 20560 3044 20600
rect 2986 20559 3044 20560
rect 3435 20600 3477 20609
rect 3435 20560 3436 20600
rect 3476 20560 3477 20600
rect 3435 20551 3477 20560
rect 4491 20600 4533 20609
rect 4491 20560 4492 20600
rect 4532 20560 4533 20600
rect 4491 20551 4533 20560
rect 5931 20600 5973 20609
rect 5931 20560 5932 20600
rect 5972 20560 5973 20600
rect 5931 20551 5973 20560
rect 6699 20600 6741 20609
rect 6699 20560 6700 20600
rect 6740 20560 6741 20600
rect 6699 20551 6741 20560
rect 7450 20600 7508 20601
rect 7450 20560 7459 20600
rect 7499 20560 7508 20600
rect 7450 20559 7508 20560
rect 8794 20600 8852 20601
rect 8794 20560 8803 20600
rect 8843 20560 8852 20600
rect 8794 20559 8852 20560
rect 9147 20600 9189 20609
rect 9147 20560 9148 20600
rect 9188 20560 9189 20600
rect 9147 20551 9189 20560
rect 9994 20600 10052 20601
rect 9994 20560 10003 20600
rect 10043 20560 10052 20600
rect 9994 20559 10052 20560
rect 10906 20600 10964 20601
rect 10906 20560 10915 20600
rect 10955 20560 10964 20600
rect 10906 20559 10964 20560
rect 11211 20600 11253 20609
rect 11211 20560 11212 20600
rect 11252 20560 11253 20600
rect 11211 20551 11253 20560
rect 11530 20600 11588 20601
rect 11530 20560 11539 20600
rect 11579 20560 11588 20600
rect 11530 20559 11588 20560
rect 12027 20600 12069 20609
rect 12027 20560 12028 20600
rect 12068 20560 12069 20600
rect 12027 20551 12069 20560
rect 12507 20600 12549 20609
rect 12507 20560 12508 20600
rect 12548 20560 12549 20600
rect 12507 20551 12549 20560
rect 13594 20600 13652 20601
rect 13594 20560 13603 20600
rect 13643 20560 13652 20600
rect 13594 20559 13652 20560
rect 16395 20600 16437 20609
rect 16395 20560 16396 20600
rect 16436 20560 16437 20600
rect 16395 20551 16437 20560
rect 17338 20600 17396 20601
rect 17338 20560 17347 20600
rect 17387 20560 17396 20600
rect 17338 20559 17396 20560
rect 18106 20600 18164 20601
rect 18106 20560 18115 20600
rect 18155 20560 18164 20600
rect 18106 20559 18164 20560
rect 18939 20600 18981 20609
rect 18939 20560 18940 20600
rect 18980 20560 18981 20600
rect 18939 20551 18981 20560
rect 20122 20600 20180 20601
rect 20122 20560 20131 20600
rect 20171 20560 20180 20600
rect 20122 20559 20180 20560
rect 20235 20600 20277 20609
rect 20235 20560 20236 20600
rect 20276 20560 20277 20600
rect 20235 20551 20277 20560
rect 20475 20600 20517 20609
rect 20475 20560 20476 20600
rect 20516 20560 20517 20600
rect 20475 20551 20517 20560
rect 21298 20600 21356 20601
rect 21298 20560 21307 20600
rect 21347 20560 21356 20600
rect 21298 20559 21356 20560
rect 21466 20600 21524 20601
rect 21466 20560 21475 20600
rect 21515 20560 21524 20600
rect 21466 20559 21524 20560
rect 22251 20600 22293 20609
rect 22251 20560 22252 20600
rect 22292 20560 22293 20600
rect 22251 20551 22293 20560
rect 25018 20600 25076 20601
rect 25018 20560 25027 20600
rect 25067 20560 25076 20600
rect 25018 20559 25076 20560
rect 25419 20600 25461 20609
rect 25419 20560 25420 20600
rect 25460 20560 25461 20600
rect 25419 20551 25461 20560
rect 576 20432 31392 20456
rect 576 20392 4352 20432
rect 4720 20392 12126 20432
rect 12494 20392 19900 20432
rect 20268 20392 27674 20432
rect 28042 20392 31392 20432
rect 576 20368 31392 20392
rect 1131 20264 1173 20273
rect 1131 20224 1132 20264
rect 1172 20224 1173 20264
rect 1131 20215 1173 20224
rect 2362 20264 2420 20265
rect 2362 20224 2371 20264
rect 2411 20224 2420 20264
rect 2362 20223 2420 20224
rect 3627 20264 3669 20273
rect 3627 20224 3628 20264
rect 3668 20224 3669 20264
rect 3627 20215 3669 20224
rect 4059 20264 4101 20273
rect 4059 20224 4060 20264
rect 4100 20224 4101 20264
rect 4059 20215 4101 20224
rect 5434 20264 5492 20265
rect 5434 20224 5443 20264
rect 5483 20224 5492 20264
rect 9562 20264 9620 20265
rect 5434 20223 5492 20224
rect 6615 20222 6657 20231
rect 9562 20224 9571 20264
rect 9611 20224 9620 20264
rect 9562 20223 9620 20224
rect 10443 20264 10485 20273
rect 10443 20224 10444 20264
rect 10484 20224 10485 20264
rect 1594 20180 1652 20181
rect 1594 20140 1603 20180
rect 1643 20140 1652 20180
rect 1594 20139 1652 20140
rect 3424 20180 3466 20189
rect 3424 20140 3425 20180
rect 3465 20140 3466 20180
rect 6615 20182 6616 20222
rect 6656 20182 6657 20222
rect 10443 20215 10485 20224
rect 13803 20264 13845 20273
rect 13803 20224 13804 20264
rect 13844 20224 13845 20264
rect 13803 20215 13845 20224
rect 14074 20264 14132 20265
rect 14074 20224 14083 20264
rect 14123 20224 14132 20264
rect 14074 20223 14132 20224
rect 14554 20264 14612 20265
rect 14554 20224 14563 20264
rect 14603 20224 14612 20264
rect 14554 20223 14612 20224
rect 16474 20264 16532 20265
rect 16474 20224 16483 20264
rect 16523 20224 16532 20264
rect 16474 20223 16532 20224
rect 18682 20264 18740 20265
rect 18682 20224 18691 20264
rect 18731 20224 18740 20264
rect 18682 20223 18740 20224
rect 19851 20264 19893 20273
rect 19851 20224 19852 20264
rect 19892 20224 19893 20264
rect 19851 20215 19893 20224
rect 21579 20264 21621 20273
rect 21579 20224 21580 20264
rect 21620 20224 21621 20264
rect 21579 20215 21621 20224
rect 23979 20264 24021 20273
rect 23979 20224 23980 20264
rect 24020 20224 24021 20264
rect 23979 20215 24021 20224
rect 28875 20264 28917 20273
rect 28875 20224 28876 20264
rect 28916 20224 28917 20264
rect 28875 20215 28917 20224
rect 6615 20173 6657 20182
rect 7258 20180 7316 20181
rect 3424 20131 3466 20140
rect 7258 20140 7267 20180
rect 7307 20140 7316 20180
rect 7258 20139 7316 20140
rect 8043 20180 8085 20189
rect 8043 20140 8044 20180
rect 8084 20140 8085 20180
rect 5818 20138 5876 20139
rect 843 20096 885 20105
rect 843 20056 844 20096
rect 884 20056 885 20096
rect 1282 20096 1340 20097
rect 843 20047 885 20056
rect 977 20093 1035 20094
rect 977 20053 986 20093
rect 1026 20053 1035 20093
rect 1282 20056 1291 20096
rect 1331 20056 1340 20096
rect 1282 20055 1340 20056
rect 1516 20096 1558 20105
rect 1516 20056 1517 20096
rect 1557 20056 1558 20096
rect 977 20052 1035 20053
rect 1516 20047 1558 20056
rect 1762 20096 1820 20097
rect 1762 20056 1771 20096
rect 1811 20056 1820 20096
rect 1762 20055 1820 20056
rect 1995 20096 2037 20105
rect 1995 20056 1996 20096
rect 2036 20056 2037 20096
rect 1995 20047 2037 20056
rect 2266 20096 2324 20097
rect 2266 20056 2275 20096
rect 2315 20056 2324 20096
rect 2266 20055 2324 20056
rect 2582 20096 2624 20105
rect 2582 20056 2583 20096
rect 2623 20056 2624 20096
rect 2582 20047 2624 20056
rect 3051 20096 3093 20105
rect 3051 20056 3052 20096
rect 3092 20056 3093 20096
rect 3051 20047 3093 20056
rect 3280 20096 3338 20097
rect 3915 20096 3957 20105
rect 3280 20056 3289 20096
rect 3329 20056 3338 20096
rect 3280 20055 3338 20056
rect 3723 20087 3765 20096
rect 3723 20047 3724 20087
rect 3764 20047 3765 20087
rect 3915 20056 3916 20096
rect 3956 20056 3957 20096
rect 3915 20047 3957 20056
rect 4203 20096 4245 20105
rect 4203 20056 4204 20096
rect 4244 20056 4245 20096
rect 4203 20047 4245 20056
rect 4378 20096 4436 20097
rect 4378 20056 4387 20096
rect 4427 20056 4436 20096
rect 4378 20055 4436 20056
rect 4534 20096 4576 20105
rect 4534 20056 4535 20096
rect 4575 20056 4576 20096
rect 4534 20047 4576 20056
rect 4779 20096 4821 20105
rect 4779 20056 4780 20096
rect 4820 20056 4821 20096
rect 4779 20047 4821 20056
rect 5083 20096 5141 20097
rect 5083 20056 5092 20096
rect 5132 20056 5141 20096
rect 5083 20055 5141 20056
rect 5242 20096 5300 20097
rect 5242 20056 5251 20096
rect 5291 20056 5300 20096
rect 5242 20055 5300 20056
rect 5367 20096 5409 20105
rect 5818 20098 5827 20138
rect 5867 20098 5876 20138
rect 5818 20097 5876 20098
rect 6394 20138 6452 20139
rect 6394 20098 6403 20138
rect 6443 20098 6452 20138
rect 6394 20097 6452 20098
rect 6826 20138 6884 20139
rect 6826 20098 6835 20138
rect 6875 20098 6884 20138
rect 8043 20131 8085 20140
rect 9147 20180 9189 20189
rect 9147 20140 9148 20180
rect 9188 20140 9189 20180
rect 9147 20131 9189 20140
rect 9782 20180 9824 20189
rect 9782 20140 9783 20180
rect 9823 20140 9824 20180
rect 9782 20131 9824 20140
rect 10923 20180 10965 20189
rect 10923 20140 10924 20180
rect 10964 20140 10965 20180
rect 10923 20131 10965 20140
rect 12459 20180 12501 20189
rect 12459 20140 12460 20180
rect 12500 20140 12501 20180
rect 12459 20131 12501 20140
rect 12970 20180 13028 20181
rect 12970 20140 12979 20180
rect 13019 20140 13028 20180
rect 12970 20139 13028 20140
rect 14187 20180 14229 20189
rect 14187 20140 14188 20180
rect 14228 20140 14229 20180
rect 14187 20131 14229 20140
rect 15133 20180 15175 20189
rect 15133 20140 15134 20180
rect 15174 20140 15175 20180
rect 15133 20131 15175 20140
rect 16971 20180 17013 20189
rect 16971 20140 16972 20180
rect 17012 20140 17013 20180
rect 16971 20131 17013 20140
rect 19546 20180 19604 20181
rect 19546 20140 19555 20180
rect 19595 20140 19604 20180
rect 19546 20139 19604 20140
rect 22138 20180 22196 20181
rect 22138 20140 22147 20180
rect 22187 20140 22196 20180
rect 22138 20139 22196 20140
rect 25131 20180 25173 20189
rect 25131 20140 25132 20180
rect 25172 20140 25173 20180
rect 25131 20131 25173 20140
rect 29211 20180 29253 20189
rect 29211 20140 29212 20180
rect 29252 20140 29253 20180
rect 29211 20131 29253 20140
rect 30267 20180 30309 20189
rect 30267 20140 30268 20180
rect 30308 20140 30309 20180
rect 30267 20131 30309 20140
rect 6826 20097 6884 20098
rect 5367 20056 5368 20096
rect 5408 20056 5409 20096
rect 5367 20047 5409 20056
rect 5530 20096 5588 20097
rect 5530 20056 5539 20096
rect 5579 20056 5588 20096
rect 5530 20055 5588 20056
rect 5652 20096 5710 20097
rect 5652 20056 5661 20096
rect 5701 20056 5710 20096
rect 6939 20096 6981 20105
rect 5652 20055 5710 20056
rect 5931 20054 5973 20063
rect 3723 20038 3765 20047
rect 1402 20012 1460 20013
rect 1402 19972 1411 20012
rect 1451 19972 1460 20012
rect 1402 19971 1460 19972
rect 1882 20012 1940 20013
rect 1882 19972 1891 20012
rect 1931 19972 1940 20012
rect 1882 19971 1940 19972
rect 2091 20012 2133 20021
rect 2091 19972 2092 20012
rect 2132 19972 2133 20012
rect 2091 19963 2133 19972
rect 2955 20012 2997 20021
rect 4666 20012 4724 20013
rect 2955 19972 2956 20012
rect 2996 19972 2997 20012
rect 2955 19963 2997 19972
rect 3186 20003 3232 20012
rect 3186 19963 3187 20003
rect 3227 19963 3232 20003
rect 4666 19972 4675 20012
rect 4715 19972 4724 20012
rect 4666 19971 4724 19972
rect 4875 20012 4917 20021
rect 4875 19972 4876 20012
rect 4916 19972 4917 20012
rect 5931 20014 5932 20054
rect 5972 20014 5973 20054
rect 6250 20054 6308 20055
rect 5931 20005 5973 20014
rect 6123 20012 6165 20021
rect 6250 20014 6259 20054
rect 6299 20014 6308 20054
rect 6250 20013 6308 20014
rect 6535 20054 6577 20063
rect 6535 20014 6536 20054
rect 6576 20014 6577 20054
rect 6939 20056 6940 20096
rect 6980 20056 6981 20096
rect 6939 20047 6981 20056
rect 7179 20096 7221 20105
rect 7179 20056 7180 20096
rect 7220 20056 7221 20096
rect 7179 20047 7221 20056
rect 7563 20096 7605 20105
rect 7563 20056 7564 20096
rect 7604 20056 7605 20096
rect 7563 20047 7605 20056
rect 7682 20096 7724 20105
rect 7682 20056 7683 20096
rect 7723 20056 7724 20096
rect 7682 20047 7724 20056
rect 7792 20096 7850 20097
rect 7792 20056 7801 20096
rect 7841 20056 7850 20096
rect 7792 20055 7850 20056
rect 7947 20096 7989 20105
rect 7947 20056 7948 20096
rect 7988 20056 7989 20096
rect 7947 20047 7989 20056
rect 8139 20096 8181 20105
rect 8139 20056 8140 20096
rect 8180 20056 8181 20096
rect 8139 20047 8181 20056
rect 8278 20096 8320 20105
rect 8278 20056 8279 20096
rect 8319 20056 8320 20096
rect 8278 20047 8320 20056
rect 8523 20096 8565 20105
rect 8523 20056 8524 20096
rect 8564 20056 8565 20096
rect 8523 20047 8565 20056
rect 8811 20096 8853 20105
rect 8811 20056 8812 20096
rect 8852 20056 8853 20096
rect 8811 20047 8853 20056
rect 9003 20096 9045 20105
rect 9003 20056 9004 20096
rect 9044 20056 9045 20096
rect 9003 20047 9045 20056
rect 9291 20096 9333 20105
rect 9291 20056 9292 20096
rect 9332 20056 9333 20096
rect 9291 20047 9333 20056
rect 9466 20096 9524 20097
rect 9466 20056 9475 20096
rect 9515 20056 9524 20096
rect 10155 20096 10197 20105
rect 9466 20055 9524 20056
rect 9915 20054 9957 20063
rect 4875 19963 4917 19972
rect 6123 19972 6124 20012
rect 6164 19972 6165 20012
rect 6535 20005 6577 20014
rect 6692 20012 6734 20021
rect 6123 19963 6165 19972
rect 6692 19972 6693 20012
rect 6733 19972 6734 20012
rect 6692 19963 6734 19972
rect 7066 20012 7124 20013
rect 7066 19972 7075 20012
rect 7115 19972 7124 20012
rect 7066 19971 7124 19972
rect 7467 20012 7509 20021
rect 7467 19972 7468 20012
rect 7508 19972 7509 20012
rect 7467 19963 7509 19972
rect 8410 20012 8468 20013
rect 8410 19972 8419 20012
rect 8459 19972 8468 20012
rect 8410 19971 8468 19972
rect 8619 20012 8661 20021
rect 8619 19972 8620 20012
rect 8660 19972 8661 20012
rect 9915 20014 9916 20054
rect 9956 20014 9957 20054
rect 10155 20056 10156 20096
rect 10196 20056 10197 20096
rect 10155 20047 10197 20056
rect 10538 20096 10580 20105
rect 10538 20056 10539 20096
rect 10579 20056 10580 20096
rect 10538 20047 10580 20056
rect 10658 20096 10700 20105
rect 10658 20056 10659 20096
rect 10699 20056 10700 20096
rect 10658 20047 10700 20056
rect 10768 20096 10826 20097
rect 10768 20056 10777 20096
rect 10817 20056 10826 20096
rect 10768 20055 10826 20056
rect 11019 20096 11061 20105
rect 11019 20056 11020 20096
rect 11060 20056 11061 20096
rect 11019 20047 11061 20056
rect 11138 20096 11180 20105
rect 11138 20056 11139 20096
rect 11179 20056 11180 20096
rect 11138 20047 11180 20056
rect 11248 20096 11306 20097
rect 11248 20056 11257 20096
rect 11297 20056 11306 20096
rect 11248 20055 11306 20056
rect 11979 20096 12021 20105
rect 11979 20056 11980 20096
rect 12020 20056 12021 20096
rect 11979 20047 12021 20056
rect 12346 20096 12404 20097
rect 12346 20056 12355 20096
rect 12395 20056 12404 20096
rect 12346 20055 12404 20056
rect 12665 20096 12707 20105
rect 12665 20056 12666 20096
rect 12706 20056 12707 20096
rect 12665 20047 12707 20056
rect 13165 20096 13223 20097
rect 13165 20056 13174 20096
rect 13214 20056 13223 20096
rect 13165 20055 13223 20056
rect 13371 20096 13413 20105
rect 13371 20056 13372 20096
rect 13412 20056 13413 20096
rect 13371 20047 13413 20056
rect 13492 20096 13534 20105
rect 13492 20056 13493 20096
rect 13533 20056 13534 20096
rect 13492 20047 13534 20056
rect 13611 20096 13653 20105
rect 13611 20056 13612 20096
rect 13652 20056 13653 20096
rect 13611 20047 13653 20056
rect 13981 20096 14023 20105
rect 14464 20096 14506 20105
rect 13981 20056 13982 20096
rect 14022 20056 14023 20096
rect 13981 20047 14023 20056
rect 14283 20087 14325 20096
rect 14283 20047 14284 20087
rect 14324 20047 14325 20087
rect 14464 20056 14465 20096
rect 14505 20056 14506 20096
rect 14464 20047 14506 20056
rect 14667 20096 14709 20105
rect 15339 20096 15381 20105
rect 15874 20096 15932 20097
rect 14667 20056 14668 20096
rect 14708 20056 14709 20096
rect 14667 20047 14709 20056
rect 14763 20087 14805 20096
rect 14763 20047 14764 20087
rect 14804 20047 14805 20087
rect 15339 20056 15340 20096
rect 15380 20056 15381 20096
rect 15339 20047 15381 20056
rect 15435 20087 15477 20096
rect 15435 20047 15436 20087
rect 15476 20047 15477 20087
rect 15874 20056 15883 20096
rect 15923 20056 15932 20096
rect 15874 20055 15932 20056
rect 16105 20096 16147 20105
rect 16105 20056 16106 20096
rect 16146 20056 16147 20096
rect 16105 20047 16147 20056
rect 16378 20096 16436 20097
rect 16378 20056 16387 20096
rect 16427 20056 16436 20096
rect 16378 20055 16436 20056
rect 16694 20096 16736 20105
rect 16694 20056 16695 20096
rect 16735 20056 16736 20096
rect 16868 20101 16926 20102
rect 16868 20061 16877 20101
rect 16917 20061 16926 20101
rect 16868 20060 16926 20061
rect 17177 20096 17219 20105
rect 16694 20047 16736 20056
rect 17177 20056 17178 20096
rect 17218 20056 17219 20096
rect 17177 20047 17219 20056
rect 17451 20096 17493 20105
rect 17451 20056 17452 20096
rect 17492 20056 17493 20096
rect 17451 20047 17493 20056
rect 17818 20096 17876 20097
rect 17818 20056 17827 20096
rect 17867 20056 17876 20096
rect 17818 20055 17876 20056
rect 18106 20096 18164 20097
rect 18106 20056 18115 20096
rect 18155 20056 18164 20096
rect 18106 20055 18164 20056
rect 18358 20096 18400 20105
rect 18358 20056 18359 20096
rect 18399 20056 18400 20096
rect 18358 20047 18400 20056
rect 18603 20096 18645 20105
rect 18603 20056 18604 20096
rect 18644 20056 18645 20096
rect 18603 20047 18645 20056
rect 19083 20096 19125 20105
rect 19083 20056 19084 20096
rect 19124 20056 19125 20096
rect 19083 20047 19125 20056
rect 19258 20096 19316 20097
rect 19258 20056 19267 20096
rect 19307 20056 19316 20096
rect 19258 20055 19316 20056
rect 19371 20096 19413 20105
rect 19371 20056 19372 20096
rect 19412 20056 19413 20096
rect 19371 20047 19413 20056
rect 19755 20096 19797 20105
rect 19755 20056 19756 20096
rect 19796 20056 19797 20096
rect 19755 20047 19797 20056
rect 19899 20096 19941 20105
rect 19899 20056 19900 20096
rect 19940 20056 19941 20096
rect 19899 20047 19941 20056
rect 20427 20096 20469 20105
rect 20427 20056 20428 20096
rect 20468 20056 20469 20096
rect 20427 20047 20469 20056
rect 20811 20096 20853 20105
rect 20811 20056 20812 20096
rect 20852 20056 20853 20096
rect 20811 20047 20853 20056
rect 21562 20096 21620 20097
rect 21562 20056 21571 20096
rect 21611 20056 21620 20096
rect 21562 20055 21620 20056
rect 21675 20096 21717 20105
rect 21675 20056 21676 20096
rect 21716 20056 21717 20096
rect 21675 20047 21717 20056
rect 22426 20096 22484 20097
rect 22426 20056 22435 20096
rect 22475 20056 22484 20096
rect 22426 20055 22484 20056
rect 23115 20096 23157 20105
rect 23115 20056 23116 20096
rect 23156 20056 23157 20096
rect 23115 20047 23157 20056
rect 23691 20096 23733 20105
rect 23691 20056 23692 20096
rect 23732 20056 23733 20096
rect 23691 20047 23733 20056
rect 23931 20096 23989 20097
rect 23931 20056 23940 20096
rect 23980 20056 23989 20096
rect 23931 20055 23989 20056
rect 24118 20096 24160 20105
rect 24118 20056 24119 20096
rect 24159 20056 24160 20096
rect 23806 20054 23864 20055
rect 14283 20038 14325 20047
rect 14763 20038 14805 20047
rect 15435 20038 15477 20047
rect 9915 20005 9957 20014
rect 10042 20012 10100 20013
rect 8619 19963 8661 19972
rect 10042 19972 10051 20012
rect 10091 19972 10100 20012
rect 10042 19971 10100 19972
rect 10251 20012 10293 20021
rect 10251 19972 10252 20012
rect 10292 19972 10293 20012
rect 10251 19963 10293 19972
rect 15994 20012 16052 20013
rect 15994 19972 16003 20012
rect 16043 19972 16052 20012
rect 15994 19971 16052 19972
rect 16203 20012 16245 20021
rect 16203 19972 16204 20012
rect 16244 19972 16245 20012
rect 16203 19963 16245 19972
rect 17643 20012 17685 20021
rect 17643 19972 17644 20012
rect 17684 19972 17685 20012
rect 17643 19963 17685 19972
rect 18219 20012 18261 20021
rect 18219 19972 18220 20012
rect 18260 19972 18261 20012
rect 18219 19963 18261 19972
rect 18490 20012 18548 20013
rect 18490 19972 18499 20012
rect 18539 19972 18548 20012
rect 18490 19971 18548 19972
rect 22042 20012 22100 20013
rect 22042 19972 22051 20012
rect 22091 19972 22100 20012
rect 22042 19971 22100 19972
rect 22618 20012 22676 20013
rect 22618 19972 22627 20012
rect 22667 19972 22676 20012
rect 22618 19971 22676 19972
rect 23025 20012 23067 20021
rect 23806 20014 23815 20054
rect 23855 20014 23864 20054
rect 24118 20047 24160 20056
rect 24363 20096 24405 20105
rect 24363 20056 24364 20096
rect 24404 20056 24405 20096
rect 24363 20047 24405 20056
rect 24747 20096 24789 20105
rect 24747 20056 24748 20096
rect 24788 20056 24789 20096
rect 24747 20047 24789 20056
rect 25018 20096 25076 20097
rect 25018 20056 25027 20096
rect 25067 20056 25076 20096
rect 25018 20055 25076 20056
rect 27610 20096 27668 20097
rect 27610 20056 27619 20096
rect 27659 20056 27668 20096
rect 27610 20055 27668 20056
rect 28203 20096 28245 20105
rect 30411 20096 30453 20105
rect 28203 20056 28204 20096
rect 28244 20056 28245 20096
rect 28203 20047 28245 20056
rect 29058 20087 29104 20096
rect 29058 20047 29059 20087
rect 29099 20047 29104 20087
rect 30411 20056 30412 20096
rect 30452 20056 30453 20096
rect 30411 20047 30453 20056
rect 29058 20038 29104 20047
rect 23806 20013 23864 20014
rect 23025 19972 23026 20012
rect 23066 19972 23067 20012
rect 23025 19963 23067 19972
rect 24250 20012 24308 20013
rect 24250 19972 24259 20012
rect 24299 19972 24308 20012
rect 24250 19971 24308 19972
rect 24459 20012 24501 20021
rect 24459 19972 24460 20012
rect 24500 19972 24501 20012
rect 24459 19963 24501 19972
rect 27994 20012 28052 20013
rect 27994 19972 28003 20012
rect 28043 19972 28052 20012
rect 27994 19971 28052 19972
rect 3186 19954 3232 19963
rect 6027 19928 6069 19937
rect 6027 19888 6028 19928
rect 6068 19888 6069 19928
rect 6027 19879 6069 19888
rect 17307 19928 17349 19937
rect 17307 19888 17308 19928
rect 17348 19888 17349 19928
rect 17307 19879 17349 19888
rect 19275 19928 19317 19937
rect 19275 19888 19276 19928
rect 19316 19888 19317 19928
rect 19275 19879 19317 19888
rect 21003 19928 21045 19937
rect 21003 19888 21004 19928
rect 21044 19888 21045 19928
rect 21003 19879 21045 19888
rect 21867 19928 21909 19937
rect 21867 19888 21868 19928
rect 21908 19888 21909 19928
rect 21867 19879 21909 19888
rect 25419 19928 25461 19937
rect 25419 19888 25420 19928
rect 25460 19888 25461 19928
rect 25419 19879 25461 19888
rect 29547 19928 29589 19937
rect 29547 19888 29548 19928
rect 29588 19888 29589 19928
rect 29547 19879 29589 19888
rect 29931 19928 29973 19937
rect 29931 19888 29932 19928
rect 29972 19888 29973 19928
rect 29931 19879 29973 19888
rect 2571 19844 2613 19853
rect 2571 19804 2572 19844
rect 2612 19804 2613 19844
rect 2571 19795 2613 19804
rect 3418 19844 3476 19845
rect 3418 19804 3427 19844
rect 3467 19804 3476 19844
rect 3418 19803 3476 19804
rect 4378 19844 4436 19845
rect 4378 19804 4387 19844
rect 4427 19804 4436 19844
rect 4378 19803 4436 19804
rect 8811 19844 8853 19853
rect 8811 19804 8812 19844
rect 8852 19804 8853 19844
rect 8811 19795 8853 19804
rect 9771 19844 9813 19853
rect 9771 19804 9772 19844
rect 9812 19804 9813 19844
rect 9771 19795 9813 19804
rect 11578 19844 11636 19845
rect 11578 19804 11587 19844
rect 11627 19804 11636 19844
rect 11578 19803 11636 19804
rect 12651 19844 12693 19853
rect 12651 19804 12652 19844
rect 12692 19804 12693 19844
rect 12651 19795 12693 19804
rect 15130 19844 15188 19845
rect 15130 19804 15139 19844
rect 15179 19804 15188 19844
rect 15130 19803 15188 19804
rect 16683 19844 16725 19853
rect 16683 19804 16684 19844
rect 16724 19804 16725 19844
rect 16683 19795 16725 19804
rect 17163 19844 17205 19853
rect 17163 19804 17164 19844
rect 17204 19804 17205 19844
rect 17163 19795 17205 19804
rect 20187 19844 20229 19853
rect 20187 19804 20188 19844
rect 20228 19804 20229 19844
rect 20187 19795 20229 19804
rect 22923 19844 22965 19853
rect 22923 19804 22924 19844
rect 22964 19804 22965 19844
rect 22923 19795 22965 19804
rect 25707 19844 25749 19853
rect 25707 19804 25708 19844
rect 25748 19804 25749 19844
rect 25707 19795 25749 19804
rect 576 19676 31392 19700
rect 576 19636 3112 19676
rect 3480 19636 10886 19676
rect 11254 19636 18660 19676
rect 19028 19636 26434 19676
rect 26802 19636 31392 19676
rect 576 19612 31392 19636
rect 3130 19508 3188 19509
rect 3130 19468 3139 19508
rect 3179 19468 3188 19508
rect 3130 19467 3188 19468
rect 3610 19508 3668 19509
rect 3610 19468 3619 19508
rect 3659 19468 3668 19508
rect 3610 19467 3668 19468
rect 7738 19508 7796 19509
rect 7738 19468 7747 19508
rect 7787 19468 7796 19508
rect 7738 19467 7796 19468
rect 9946 19508 10004 19509
rect 9946 19468 9955 19508
rect 9995 19468 10004 19508
rect 9946 19467 10004 19468
rect 11194 19508 11252 19509
rect 11194 19468 11203 19508
rect 11243 19468 11252 19508
rect 11194 19467 11252 19468
rect 13035 19508 13077 19517
rect 13035 19468 13036 19508
rect 13076 19468 13077 19508
rect 13035 19459 13077 19468
rect 14266 19508 14324 19509
rect 14266 19468 14275 19508
rect 14315 19468 14324 19508
rect 14266 19467 14324 19468
rect 15226 19508 15284 19509
rect 15226 19468 15235 19508
rect 15275 19468 15284 19508
rect 15226 19467 15284 19468
rect 16186 19508 16244 19509
rect 16186 19468 16195 19508
rect 16235 19468 16244 19508
rect 16186 19467 16244 19468
rect 16666 19508 16724 19509
rect 16666 19468 16675 19508
rect 16715 19468 16724 19508
rect 16666 19467 16724 19468
rect 17451 19508 17493 19517
rect 17451 19468 17452 19508
rect 17492 19468 17493 19508
rect 17451 19459 17493 19468
rect 20715 19508 20757 19517
rect 20715 19468 20716 19508
rect 20756 19468 20757 19508
rect 20715 19459 20757 19468
rect 22683 19508 22725 19517
rect 22683 19468 22684 19508
rect 22724 19468 22725 19508
rect 22683 19459 22725 19468
rect 28107 19508 28149 19517
rect 28107 19468 28108 19508
rect 28148 19468 28149 19508
rect 28107 19459 28149 19468
rect 12459 19424 12501 19433
rect 9723 19415 9765 19424
rect 9723 19375 9724 19415
rect 9764 19375 9765 19415
rect 12459 19384 12460 19424
rect 12500 19384 12501 19424
rect 12459 19375 12501 19384
rect 18603 19424 18645 19433
rect 18603 19384 18604 19424
rect 18644 19384 18645 19424
rect 18603 19375 18645 19384
rect 22347 19424 22389 19433
rect 22347 19384 22348 19424
rect 22388 19384 22389 19424
rect 22347 19375 22389 19384
rect 28779 19424 28821 19433
rect 28779 19384 28780 19424
rect 28820 19384 28821 19424
rect 28779 19375 28821 19384
rect 9723 19366 9765 19375
rect 1018 19340 1076 19341
rect 1018 19300 1027 19340
rect 1067 19300 1076 19340
rect 1018 19299 1076 19300
rect 1227 19340 1269 19349
rect 1227 19300 1228 19340
rect 1268 19300 1269 19340
rect 1227 19291 1269 19300
rect 1419 19340 1461 19349
rect 1419 19300 1420 19340
rect 1460 19300 1461 19340
rect 1419 19291 1461 19300
rect 1995 19340 2037 19349
rect 1995 19300 1996 19340
rect 2036 19300 2037 19340
rect 1995 19291 2037 19300
rect 2187 19340 2229 19349
rect 2187 19300 2188 19340
rect 2228 19300 2229 19340
rect 2187 19291 2229 19300
rect 4203 19340 4245 19349
rect 4203 19300 4204 19340
rect 4244 19300 4245 19340
rect 4203 19291 4245 19300
rect 5931 19340 5973 19349
rect 6722 19340 6764 19349
rect 5931 19300 5932 19340
rect 5972 19300 5973 19340
rect 5931 19291 5973 19300
rect 6162 19331 6208 19340
rect 6162 19291 6163 19331
rect 6203 19291 6208 19331
rect 6722 19300 6723 19340
rect 6763 19300 6764 19340
rect 6722 19291 6764 19300
rect 8698 19340 8756 19341
rect 8698 19300 8707 19340
rect 8747 19300 8756 19340
rect 8698 19299 8756 19300
rect 8907 19340 8949 19349
rect 8907 19300 8908 19340
rect 8948 19300 8949 19340
rect 8907 19291 8949 19300
rect 17722 19340 17780 19341
rect 17722 19300 17731 19340
rect 17771 19300 17780 19340
rect 17722 19299 17780 19300
rect 17931 19340 17973 19349
rect 25131 19340 25173 19349
rect 17931 19300 17932 19340
rect 17972 19300 17973 19340
rect 17931 19291 17973 19300
rect 23250 19331 23296 19340
rect 23250 19291 23251 19331
rect 23291 19291 23296 19331
rect 25131 19300 25132 19340
rect 25172 19300 25173 19340
rect 25131 19291 25173 19300
rect 26283 19340 26325 19349
rect 26283 19300 26284 19340
rect 26324 19300 26325 19340
rect 26283 19291 26325 19300
rect 27675 19340 27717 19349
rect 27675 19300 27676 19340
rect 27716 19300 27717 19340
rect 27675 19291 27717 19300
rect 6162 19282 6208 19291
rect 23250 19282 23296 19291
rect 7750 19267 7808 19268
rect 886 19256 928 19265
rect 886 19216 887 19256
rect 927 19216 928 19256
rect 886 19207 928 19216
rect 1131 19256 1173 19265
rect 1131 19216 1132 19256
rect 1172 19216 1173 19256
rect 1131 19207 1173 19216
rect 1594 19256 1652 19257
rect 1594 19216 1603 19256
rect 1643 19216 1652 19256
rect 1594 19215 1652 19216
rect 2283 19256 2325 19265
rect 2283 19216 2284 19256
rect 2324 19216 2325 19256
rect 2283 19207 2325 19216
rect 2402 19256 2444 19265
rect 2402 19216 2403 19256
rect 2443 19216 2444 19256
rect 2402 19207 2444 19216
rect 2512 19256 2570 19257
rect 2512 19216 2521 19256
rect 2561 19216 2570 19256
rect 2512 19215 2570 19216
rect 2763 19256 2805 19265
rect 2763 19216 2764 19256
rect 2804 19216 2805 19256
rect 2763 19207 2805 19216
rect 2882 19256 2924 19265
rect 2882 19216 2883 19256
rect 2923 19216 2924 19256
rect 2882 19207 2924 19216
rect 2994 19256 3036 19265
rect 2994 19216 2995 19256
rect 3035 19216 3036 19256
rect 2994 19207 3036 19216
rect 3427 19256 3485 19257
rect 3427 19216 3436 19256
rect 3476 19216 3485 19256
rect 3427 19215 3485 19216
rect 3907 19256 3965 19257
rect 3907 19216 3916 19256
rect 3956 19216 3965 19256
rect 3907 19215 3965 19216
rect 4299 19256 4341 19265
rect 4299 19216 4300 19256
rect 4340 19216 4341 19256
rect 4299 19207 4341 19216
rect 4418 19256 4460 19265
rect 4418 19216 4419 19256
rect 4459 19216 4460 19256
rect 4418 19207 4460 19216
rect 4528 19256 4586 19257
rect 4528 19216 4537 19256
rect 4577 19216 4586 19256
rect 4528 19215 4586 19216
rect 4779 19256 4821 19265
rect 4779 19216 4780 19256
rect 4820 19216 4821 19256
rect 4779 19207 4821 19216
rect 4898 19256 4940 19265
rect 4898 19216 4899 19256
rect 4939 19216 4940 19256
rect 4898 19207 4940 19216
rect 5008 19256 5066 19257
rect 5008 19216 5017 19256
rect 5057 19216 5066 19256
rect 5008 19215 5066 19216
rect 5259 19256 5301 19265
rect 5259 19216 5260 19256
rect 5300 19216 5301 19256
rect 5259 19207 5301 19216
rect 5578 19256 5636 19257
rect 5578 19216 5587 19256
rect 5627 19216 5636 19256
rect 5578 19215 5636 19216
rect 6027 19256 6069 19265
rect 6027 19216 6028 19256
rect 6068 19216 6069 19256
rect 6027 19207 6069 19216
rect 6256 19256 6314 19257
rect 6256 19216 6265 19256
rect 6305 19216 6314 19256
rect 6256 19215 6314 19216
rect 6603 19256 6645 19265
rect 6603 19216 6604 19256
rect 6644 19216 6645 19256
rect 6603 19207 6645 19216
rect 6832 19256 6890 19257
rect 6832 19216 6841 19256
rect 6881 19216 6890 19256
rect 6832 19215 6890 19216
rect 6981 19256 7039 19257
rect 6981 19216 6990 19256
rect 7030 19216 7039 19256
rect 6981 19215 7039 19216
rect 7088 19256 7146 19257
rect 7088 19216 7097 19256
rect 7137 19216 7146 19256
rect 7088 19215 7146 19216
rect 7220 19256 7278 19257
rect 7220 19216 7229 19256
rect 7269 19216 7278 19256
rect 7220 19215 7278 19216
rect 7354 19256 7412 19257
rect 7354 19216 7363 19256
rect 7403 19216 7412 19256
rect 7354 19215 7412 19216
rect 7530 19256 7588 19257
rect 7530 19216 7539 19256
rect 7579 19216 7588 19256
rect 7750 19227 7759 19267
rect 7799 19227 7808 19267
rect 7750 19226 7808 19227
rect 7882 19256 7940 19257
rect 7530 19215 7588 19216
rect 7882 19216 7891 19256
rect 7931 19216 7940 19256
rect 7882 19215 7940 19216
rect 7988 19256 8046 19257
rect 7988 19216 7997 19256
rect 8037 19216 8046 19256
rect 7988 19215 8046 19216
rect 8122 19256 8180 19257
rect 8122 19216 8131 19256
rect 8171 19216 8180 19256
rect 8122 19215 8180 19216
rect 8299 19256 8357 19257
rect 8299 19216 8308 19256
rect 8348 19216 8357 19256
rect 8299 19215 8357 19216
rect 8578 19256 8636 19257
rect 8578 19216 8587 19256
rect 8627 19216 8636 19256
rect 8578 19215 8636 19216
rect 8811 19256 8853 19265
rect 8811 19216 8812 19256
rect 8852 19216 8853 19256
rect 8811 19207 8853 19216
rect 9195 19256 9237 19265
rect 9195 19216 9196 19256
rect 9236 19216 9237 19256
rect 9195 19207 9237 19216
rect 9387 19256 9429 19265
rect 9387 19216 9388 19256
rect 9428 19216 9429 19256
rect 9387 19207 9429 19216
rect 9754 19256 9812 19257
rect 9754 19216 9763 19256
rect 9803 19216 9812 19256
rect 9754 19215 9812 19216
rect 10240 19256 10282 19265
rect 10240 19216 10241 19256
rect 10281 19216 10282 19256
rect 10240 19207 10282 19216
rect 10531 19256 10589 19257
rect 10531 19216 10540 19256
rect 10580 19216 10589 19256
rect 10531 19215 10589 19216
rect 10827 19256 10869 19265
rect 10827 19216 10828 19256
rect 10868 19216 10869 19256
rect 10827 19207 10869 19216
rect 11200 19256 11242 19265
rect 11200 19216 11201 19256
rect 11241 19216 11242 19256
rect 11200 19207 11242 19216
rect 11491 19256 11549 19257
rect 11491 19216 11500 19256
rect 11540 19216 11549 19256
rect 11491 19215 11549 19216
rect 11626 19256 11684 19257
rect 11626 19216 11635 19256
rect 11675 19216 11684 19256
rect 11626 19215 11684 19216
rect 11835 19256 11877 19265
rect 11835 19216 11836 19256
rect 11876 19216 11877 19256
rect 11835 19207 11877 19216
rect 12651 19256 12693 19265
rect 12651 19216 12652 19256
rect 12692 19216 12693 19256
rect 12651 19207 12693 19216
rect 13035 19256 13077 19265
rect 13035 19216 13036 19256
rect 13076 19216 13077 19256
rect 13035 19207 13077 19216
rect 13227 19256 13269 19265
rect 13227 19216 13228 19256
rect 13268 19216 13269 19256
rect 13227 19207 13269 19216
rect 13515 19256 13557 19265
rect 13515 19216 13516 19256
rect 13556 19216 13557 19256
rect 13515 19207 13557 19216
rect 13995 19256 14037 19265
rect 13995 19216 13996 19256
rect 14036 19216 14037 19256
rect 13995 19207 14037 19216
rect 14269 19256 14311 19265
rect 14269 19216 14270 19256
rect 14310 19216 14311 19256
rect 14269 19207 14311 19216
rect 14565 19256 14623 19257
rect 14565 19216 14574 19256
rect 14614 19216 14623 19256
rect 14565 19215 14623 19216
rect 14724 19256 14766 19265
rect 14724 19216 14725 19256
rect 14765 19216 14766 19256
rect 14724 19207 14766 19216
rect 14842 19256 14900 19257
rect 14842 19216 14851 19256
rect 14891 19216 14900 19256
rect 14842 19215 14900 19216
rect 14955 19256 14997 19265
rect 14955 19216 14956 19256
rect 14996 19216 14997 19256
rect 14955 19207 14997 19216
rect 15523 19256 15581 19257
rect 15523 19216 15532 19256
rect 15572 19216 15581 19256
rect 15523 19215 15581 19216
rect 16045 19256 16103 19257
rect 16045 19216 16054 19256
rect 16094 19216 16103 19256
rect 16045 19215 16103 19216
rect 16483 19256 16541 19257
rect 16483 19216 16492 19256
rect 16532 19216 16541 19256
rect 16483 19215 16541 19216
rect 16963 19256 17021 19257
rect 16963 19216 16972 19256
rect 17012 19216 17021 19256
rect 16963 19215 17021 19216
rect 17146 19256 17204 19257
rect 17146 19216 17155 19256
rect 17195 19216 17204 19256
rect 17146 19215 17204 19216
rect 17462 19256 17504 19265
rect 17462 19216 17463 19256
rect 17503 19216 17504 19256
rect 17462 19207 17504 19216
rect 17602 19256 17660 19257
rect 17602 19216 17611 19256
rect 17651 19216 17660 19256
rect 17602 19215 17660 19216
rect 17835 19256 17877 19265
rect 17835 19216 17836 19256
rect 17876 19216 17877 19256
rect 17835 19207 17877 19216
rect 18123 19256 18165 19265
rect 18123 19216 18124 19256
rect 18164 19216 18165 19256
rect 18123 19207 18165 19216
rect 18315 19256 18357 19265
rect 19275 19256 19317 19265
rect 18315 19216 18316 19256
rect 18356 19216 18357 19256
rect 18315 19207 18357 19216
rect 18987 19247 19029 19256
rect 18987 19207 18988 19247
rect 19028 19207 19029 19247
rect 19275 19216 19276 19256
rect 19316 19216 19317 19256
rect 19275 19207 19317 19216
rect 20235 19256 20277 19265
rect 20235 19216 20236 19256
rect 20276 19216 20277 19256
rect 20235 19207 20277 19216
rect 20523 19256 20565 19265
rect 20523 19216 20524 19256
rect 20564 19216 20565 19256
rect 20523 19207 20565 19216
rect 20842 19256 20900 19257
rect 20842 19216 20851 19256
rect 20891 19216 20900 19256
rect 20842 19215 20900 19216
rect 21003 19256 21045 19265
rect 21003 19216 21004 19256
rect 21044 19216 21045 19256
rect 21003 19207 21045 19216
rect 21754 19256 21812 19257
rect 21754 19216 21763 19256
rect 21803 19216 21812 19256
rect 21754 19215 21812 19216
rect 21867 19256 21909 19265
rect 21867 19216 21868 19256
rect 21908 19216 21909 19256
rect 21867 19207 21909 19216
rect 22347 19256 22389 19265
rect 22347 19216 22348 19256
rect 22388 19216 22389 19256
rect 22347 19207 22389 19216
rect 22539 19256 22581 19265
rect 22539 19216 22540 19256
rect 22580 19216 22581 19256
rect 22539 19207 22581 19216
rect 22779 19256 22821 19265
rect 22779 19216 22780 19256
rect 22820 19216 22821 19256
rect 22779 19207 22821 19216
rect 23115 19256 23157 19265
rect 23115 19216 23116 19256
rect 23156 19216 23157 19256
rect 23115 19207 23157 19216
rect 23344 19256 23402 19257
rect 23344 19216 23353 19256
rect 23393 19216 23402 19256
rect 23344 19215 23402 19216
rect 23499 19256 23541 19265
rect 23499 19216 23500 19256
rect 23540 19216 23541 19256
rect 23499 19207 23541 19216
rect 23691 19256 23733 19265
rect 23691 19216 23692 19256
rect 23732 19216 23733 19256
rect 23691 19207 23733 19216
rect 24075 19256 24117 19265
rect 24075 19216 24076 19256
rect 24116 19216 24117 19256
rect 24075 19207 24117 19216
rect 24194 19256 24236 19265
rect 24194 19216 24195 19256
rect 24235 19216 24236 19256
rect 24194 19207 24236 19216
rect 24304 19256 24362 19257
rect 24304 19216 24313 19256
rect 24353 19216 24362 19256
rect 24304 19215 24362 19216
rect 24459 19256 24501 19265
rect 24459 19216 24460 19256
rect 24500 19216 24501 19256
rect 24459 19207 24501 19216
rect 25323 19256 25365 19265
rect 25323 19216 25324 19256
rect 25364 19216 25365 19256
rect 25323 19207 25365 19216
rect 26176 19256 26218 19265
rect 26176 19216 26177 19256
rect 26217 19216 26218 19256
rect 26176 19207 26218 19216
rect 26379 19256 26421 19265
rect 26379 19216 26380 19256
rect 26420 19216 26421 19256
rect 26379 19207 26421 19216
rect 26667 19256 26709 19265
rect 28001 19261 28059 19262
rect 26667 19216 26668 19256
rect 26708 19216 26709 19256
rect 26667 19207 26709 19216
rect 27466 19256 27524 19257
rect 27466 19216 27475 19256
rect 27515 19216 27524 19256
rect 28001 19221 28010 19261
rect 28050 19221 28059 19261
rect 28001 19220 28059 19221
rect 28203 19256 28245 19265
rect 27466 19215 27524 19216
rect 28203 19216 28204 19256
rect 28244 19216 28245 19256
rect 28203 19207 28245 19216
rect 28395 19256 28437 19265
rect 28395 19216 28396 19256
rect 28436 19216 28437 19256
rect 28395 19207 28437 19216
rect 28587 19256 28629 19265
rect 28587 19216 28588 19256
rect 28628 19216 28629 19256
rect 28587 19207 28629 19216
rect 18987 19198 19029 19207
rect 1899 19172 1941 19181
rect 1899 19132 1900 19172
rect 1940 19132 1941 19172
rect 1899 19123 1941 19132
rect 3136 19172 3178 19181
rect 3136 19132 3137 19172
rect 3177 19132 3178 19172
rect 3136 19123 3178 19132
rect 3613 19172 3655 19181
rect 3613 19132 3614 19172
rect 3654 19132 3655 19172
rect 3613 19123 3655 19132
rect 5451 19172 5493 19181
rect 5451 19132 5452 19172
rect 5492 19132 5493 19172
rect 5451 19123 5493 19132
rect 6507 19172 6549 19181
rect 6507 19132 6508 19172
rect 6548 19132 6549 19172
rect 6507 19123 6549 19132
rect 9483 19172 9525 19181
rect 9483 19132 9484 19172
rect 9524 19132 9525 19172
rect 9483 19123 9525 19132
rect 10330 19172 10388 19173
rect 10330 19132 10339 19172
rect 10379 19132 10388 19172
rect 10330 19131 10388 19132
rect 13707 19172 13749 19181
rect 13707 19132 13708 19172
rect 13748 19132 13749 19172
rect 13707 19123 13749 19132
rect 15232 19172 15274 19181
rect 15232 19132 15233 19172
rect 15273 19132 15274 19172
rect 15232 19123 15274 19132
rect 16189 19172 16231 19181
rect 16189 19132 16190 19172
rect 16230 19132 16231 19172
rect 16189 19123 16231 19132
rect 16672 19172 16714 19181
rect 16672 19132 16673 19172
rect 16713 19132 16714 19172
rect 16672 19123 16714 19132
rect 17259 19172 17301 19181
rect 17259 19132 17260 19172
rect 17300 19132 17301 19172
rect 17259 19123 17301 19132
rect 18891 19172 18933 19181
rect 18891 19132 18892 19172
rect 18932 19132 18933 19172
rect 18891 19123 18933 19132
rect 27339 19172 27381 19181
rect 27339 19132 27340 19172
rect 27380 19132 27381 19172
rect 27339 19123 27381 19132
rect 2667 19088 2709 19097
rect 2667 19048 2668 19088
rect 2708 19048 2709 19088
rect 2667 19039 2709 19048
rect 3339 19088 3381 19097
rect 3339 19048 3340 19088
rect 3380 19048 3381 19088
rect 3339 19039 3381 19048
rect 3819 19088 3861 19097
rect 3819 19048 3820 19088
rect 3860 19048 3861 19088
rect 3819 19039 3861 19048
rect 4683 19088 4725 19097
rect 4683 19048 4684 19088
rect 4724 19048 4725 19088
rect 4683 19039 4725 19048
rect 6970 19088 7028 19089
rect 6970 19048 6979 19088
rect 7019 19048 7028 19088
rect 6970 19047 7028 19048
rect 9946 19088 10004 19089
rect 9946 19048 9955 19088
rect 9995 19048 10004 19088
rect 9946 19047 10004 19048
rect 10443 19088 10485 19097
rect 10443 19048 10444 19088
rect 10484 19048 10485 19088
rect 10443 19039 10485 19048
rect 10714 19088 10772 19089
rect 10714 19048 10723 19088
rect 10763 19048 10772 19088
rect 10714 19047 10772 19048
rect 11019 19088 11061 19097
rect 11019 19048 11020 19088
rect 11060 19048 11061 19088
rect 11019 19039 11061 19048
rect 11403 19088 11445 19097
rect 11403 19048 11404 19088
rect 11444 19048 11445 19088
rect 11403 19039 11445 19048
rect 12730 19088 12788 19089
rect 12730 19048 12739 19088
rect 12779 19048 12788 19088
rect 12730 19047 12788 19048
rect 13402 19088 13460 19089
rect 13402 19048 13411 19088
rect 13451 19048 13460 19088
rect 13402 19047 13460 19048
rect 14475 19088 14517 19097
rect 14475 19048 14476 19088
rect 14516 19048 14517 19088
rect 14475 19039 14517 19048
rect 15034 19088 15092 19089
rect 15034 19048 15043 19088
rect 15083 19048 15092 19088
rect 15034 19047 15092 19048
rect 15435 19088 15477 19097
rect 15435 19048 15436 19088
rect 15476 19048 15477 19088
rect 15435 19039 15477 19048
rect 15850 19088 15908 19089
rect 15850 19048 15859 19088
rect 15899 19048 15908 19088
rect 15850 19047 15908 19048
rect 16395 19088 16437 19097
rect 16395 19048 16396 19088
rect 16436 19048 16437 19088
rect 16395 19039 16437 19048
rect 16875 19088 16917 19097
rect 16875 19048 16876 19088
rect 16916 19048 16917 19088
rect 16875 19039 16917 19048
rect 18219 19088 18261 19097
rect 18219 19048 18220 19088
rect 18260 19048 18261 19088
rect 18219 19039 18261 19048
rect 19563 19088 19605 19097
rect 19563 19048 19564 19088
rect 19604 19048 19605 19088
rect 19563 19039 19605 19048
rect 21099 19088 21141 19097
rect 21099 19048 21100 19088
rect 21140 19048 21141 19088
rect 21099 19039 21141 19048
rect 22155 19088 22197 19097
rect 22155 19048 22156 19088
rect 22196 19048 22197 19088
rect 22155 19039 22197 19048
rect 23019 19088 23061 19097
rect 23019 19048 23020 19088
rect 23060 19048 23061 19088
rect 23019 19039 23061 19048
rect 23499 19088 23541 19097
rect 23499 19048 23500 19088
rect 23540 19048 23541 19088
rect 23499 19039 23541 19048
rect 23979 19088 24021 19097
rect 23979 19048 23980 19088
rect 24020 19048 24021 19088
rect 23979 19039 24021 19048
rect 25995 19088 26037 19097
rect 25995 19048 25996 19088
rect 26036 19048 26037 19088
rect 25995 19039 26037 19048
rect 28395 19088 28437 19097
rect 28395 19048 28396 19088
rect 28436 19048 28437 19088
rect 28395 19039 28437 19048
rect 29163 19088 29205 19097
rect 29163 19048 29164 19088
rect 29204 19048 29205 19088
rect 29163 19039 29205 19048
rect 29547 19088 29589 19097
rect 29547 19048 29548 19088
rect 29588 19048 29589 19088
rect 29547 19039 29589 19048
rect 576 18920 31392 18944
rect 576 18880 4352 18920
rect 4720 18880 12126 18920
rect 12494 18880 19900 18920
rect 20268 18880 27674 18920
rect 28042 18880 31392 18920
rect 576 18856 31392 18880
rect 6490 18794 6548 18795
rect 3226 18752 3284 18753
rect 3226 18712 3235 18752
rect 3275 18712 3284 18752
rect 3226 18711 3284 18712
rect 3339 18752 3381 18761
rect 3339 18712 3340 18752
rect 3380 18712 3381 18752
rect 3339 18703 3381 18712
rect 3723 18752 3765 18761
rect 3723 18712 3724 18752
rect 3764 18712 3765 18752
rect 3723 18703 3765 18712
rect 4779 18752 4821 18761
rect 6490 18754 6499 18794
rect 6539 18754 6548 18794
rect 6490 18753 6548 18754
rect 4779 18712 4780 18752
rect 4820 18712 4821 18752
rect 4779 18703 4821 18712
rect 5050 18752 5108 18753
rect 5050 18712 5059 18752
rect 5099 18712 5108 18752
rect 10723 18752 10781 18753
rect 5050 18711 5108 18712
rect 6615 18710 6657 18719
rect 10723 18712 10732 18752
rect 10772 18712 10781 18752
rect 10723 18711 10781 18712
rect 12682 18752 12740 18753
rect 12682 18712 12691 18752
rect 12731 18712 12740 18752
rect 12682 18711 12740 18712
rect 16090 18752 16148 18753
rect 16090 18712 16099 18752
rect 16139 18712 16148 18752
rect 16090 18711 16148 18712
rect 17242 18752 17300 18753
rect 17242 18712 17251 18752
rect 17291 18712 17300 18752
rect 17242 18711 17300 18712
rect 18298 18752 18356 18753
rect 18298 18712 18307 18752
rect 18347 18712 18356 18752
rect 18298 18711 18356 18712
rect 22539 18752 22581 18761
rect 22539 18712 22540 18752
rect 22580 18712 22581 18752
rect 778 18668 836 18669
rect 778 18628 787 18668
rect 827 18628 836 18668
rect 778 18627 836 18628
rect 1611 18668 1653 18677
rect 1611 18628 1612 18668
rect 1652 18628 1653 18668
rect 1611 18619 1653 18628
rect 3133 18668 3175 18677
rect 3133 18628 3134 18668
rect 3174 18628 3175 18668
rect 3133 18619 3175 18628
rect 4203 18668 4245 18677
rect 4203 18628 4204 18668
rect 4244 18628 4245 18668
rect 6615 18670 6616 18710
rect 6656 18670 6657 18710
rect 22539 18703 22581 18712
rect 25131 18752 25173 18761
rect 25131 18712 25132 18752
rect 25172 18712 25173 18752
rect 25131 18703 25173 18712
rect 27915 18752 27957 18761
rect 27915 18712 27916 18752
rect 27956 18712 27957 18752
rect 27915 18703 27957 18712
rect 6615 18661 6657 18670
rect 14557 18668 14599 18677
rect 4203 18619 4245 18628
rect 14557 18628 14558 18668
rect 14598 18628 14599 18668
rect 6826 18626 6884 18627
rect 973 18584 1031 18585
rect 973 18544 982 18584
rect 1022 18544 1031 18584
rect 973 18543 1031 18544
rect 1090 18584 1148 18585
rect 1090 18544 1099 18584
rect 1139 18544 1148 18584
rect 1090 18543 1148 18544
rect 1323 18584 1365 18593
rect 1323 18544 1324 18584
rect 1364 18544 1365 18584
rect 1323 18535 1365 18544
rect 1707 18584 1749 18593
rect 1707 18544 1708 18584
rect 1748 18544 1749 18584
rect 1707 18535 1749 18544
rect 1924 18584 1966 18593
rect 1924 18544 1925 18584
rect 1965 18544 1966 18584
rect 1924 18535 1966 18544
rect 2283 18584 2325 18593
rect 2283 18544 2284 18584
rect 2324 18544 2325 18584
rect 2283 18535 2325 18544
rect 2402 18584 2444 18593
rect 2402 18544 2403 18584
rect 2443 18544 2444 18584
rect 2402 18535 2444 18544
rect 2523 18584 2565 18593
rect 2523 18544 2524 18584
rect 2564 18544 2565 18584
rect 2523 18535 2565 18544
rect 2772 18584 2814 18593
rect 2772 18544 2773 18584
rect 2813 18544 2814 18584
rect 2772 18535 2814 18544
rect 2980 18584 3022 18593
rect 3627 18584 3669 18593
rect 2980 18544 2981 18584
rect 3021 18544 3022 18584
rect 2980 18535 3022 18544
rect 3435 18575 3477 18584
rect 3435 18535 3436 18575
rect 3476 18535 3477 18575
rect 3627 18544 3628 18584
rect 3668 18544 3669 18584
rect 3627 18535 3669 18544
rect 3802 18584 3860 18585
rect 3802 18544 3811 18584
rect 3851 18544 3860 18584
rect 3802 18543 3860 18544
rect 4107 18584 4149 18593
rect 4107 18544 4108 18584
rect 4148 18544 4149 18584
rect 4107 18535 4149 18544
rect 4282 18584 4340 18585
rect 4282 18544 4291 18584
rect 4331 18544 4340 18584
rect 4282 18543 4340 18544
rect 4971 18584 5013 18593
rect 4971 18544 4972 18584
rect 5012 18544 5013 18584
rect 4971 18535 5013 18544
rect 5355 18584 5397 18593
rect 5355 18544 5356 18584
rect 5396 18544 5397 18584
rect 5355 18535 5397 18544
rect 5643 18584 5685 18593
rect 5643 18544 5644 18584
rect 5684 18544 5685 18584
rect 5643 18535 5685 18544
rect 5860 18584 5902 18593
rect 5860 18544 5861 18584
rect 5901 18544 5902 18584
rect 5860 18535 5902 18544
rect 6027 18584 6069 18593
rect 6027 18544 6028 18584
rect 6068 18544 6069 18584
rect 6027 18535 6069 18544
rect 6218 18584 6260 18593
rect 6218 18544 6219 18584
rect 6259 18544 6260 18584
rect 6218 18535 6260 18544
rect 6542 18584 6584 18593
rect 6826 18586 6835 18626
rect 6875 18586 6884 18626
rect 14557 18619 14599 18628
rect 18010 18668 18068 18669
rect 18010 18628 18019 18668
rect 18059 18628 18068 18668
rect 18010 18627 18068 18628
rect 18490 18668 18548 18669
rect 18490 18628 18499 18668
rect 18539 18628 18548 18668
rect 18490 18627 18548 18628
rect 25306 18668 25364 18669
rect 25306 18628 25315 18668
rect 25355 18628 25364 18668
rect 25306 18627 25364 18628
rect 6826 18585 6884 18586
rect 7362 18584 7420 18585
rect 6542 18544 6543 18584
rect 6583 18544 6584 18584
rect 6542 18535 6584 18544
rect 6979 18573 7021 18582
rect 3435 18526 3477 18535
rect 6979 18533 6980 18573
rect 7020 18533 7021 18573
rect 6979 18524 7021 18533
rect 7083 18575 7125 18584
rect 7083 18535 7084 18575
rect 7124 18535 7125 18575
rect 7083 18526 7125 18535
rect 7266 18575 7312 18584
rect 7266 18535 7267 18575
rect 7307 18535 7312 18575
rect 7362 18544 7371 18584
rect 7411 18544 7420 18584
rect 7707 18584 7749 18593
rect 7362 18543 7420 18544
rect 7488 18573 7530 18582
rect 7266 18526 7312 18535
rect 7488 18533 7489 18573
rect 7529 18533 7530 18573
rect 7707 18544 7708 18584
rect 7748 18544 7749 18584
rect 7707 18535 7749 18544
rect 8022 18584 8064 18593
rect 8022 18544 8023 18584
rect 8063 18544 8064 18584
rect 8022 18535 8064 18544
rect 8162 18584 8204 18593
rect 8162 18544 8163 18584
rect 8203 18544 8204 18584
rect 8162 18535 8204 18544
rect 8427 18584 8469 18593
rect 8427 18544 8428 18584
rect 8468 18544 8469 18584
rect 8427 18535 8469 18544
rect 8656 18584 8714 18585
rect 8656 18544 8665 18584
rect 8705 18544 8714 18584
rect 8656 18543 8714 18544
rect 8907 18584 8949 18593
rect 8907 18544 8908 18584
rect 8948 18544 8949 18584
rect 8907 18535 8949 18544
rect 9099 18584 9141 18593
rect 9099 18544 9100 18584
rect 9140 18544 9141 18584
rect 9099 18535 9141 18544
rect 9679 18584 9737 18585
rect 9679 18544 9688 18584
rect 9728 18544 9737 18584
rect 9679 18543 9737 18544
rect 9867 18584 9909 18593
rect 9867 18544 9868 18584
rect 9908 18544 9909 18584
rect 9867 18535 9909 18544
rect 10059 18584 10101 18593
rect 10059 18544 10060 18584
rect 10100 18544 10101 18584
rect 10059 18535 10101 18544
rect 10330 18584 10388 18585
rect 10330 18544 10339 18584
rect 10379 18544 10388 18584
rect 10330 18543 10388 18544
rect 11098 18584 11156 18585
rect 11098 18544 11107 18584
rect 11147 18544 11156 18584
rect 11098 18543 11156 18544
rect 11499 18584 11541 18593
rect 11499 18544 11500 18584
rect 11540 18544 11541 18584
rect 11499 18535 11541 18544
rect 11792 18584 11834 18593
rect 11792 18544 11793 18584
rect 11833 18544 11834 18584
rect 11792 18535 11834 18544
rect 12106 18584 12164 18585
rect 12106 18544 12115 18584
rect 12155 18544 12164 18584
rect 12106 18543 12164 18544
rect 13131 18584 13173 18593
rect 13131 18544 13132 18584
rect 13172 18544 13173 18584
rect 12874 18542 12932 18543
rect 7488 18524 7530 18533
rect 1210 18500 1268 18501
rect 1210 18460 1219 18500
rect 1259 18460 1268 18500
rect 1210 18459 1268 18460
rect 1419 18500 1461 18509
rect 1419 18460 1420 18500
rect 1460 18460 1461 18500
rect 1419 18451 1461 18460
rect 1826 18500 1868 18509
rect 1826 18460 1827 18500
rect 1867 18460 1868 18500
rect 1826 18451 1868 18460
rect 2187 18500 2229 18509
rect 2187 18460 2188 18500
rect 2228 18460 2229 18500
rect 2187 18451 2229 18460
rect 2667 18500 2709 18509
rect 2667 18460 2668 18500
rect 2708 18460 2709 18500
rect 2667 18451 2709 18460
rect 2882 18500 2924 18509
rect 2882 18460 2883 18500
rect 2923 18460 2924 18500
rect 2882 18451 2924 18460
rect 5547 18500 5589 18509
rect 6699 18500 6741 18509
rect 5547 18460 5548 18500
rect 5588 18460 5589 18500
rect 5547 18451 5589 18460
rect 5778 18491 5824 18500
rect 5778 18451 5779 18491
rect 5819 18451 5824 18491
rect 6699 18460 6700 18500
rect 6740 18460 6741 18500
rect 6699 18451 6741 18460
rect 7851 18500 7893 18509
rect 7851 18460 7852 18500
rect 7892 18460 7893 18500
rect 7851 18451 7893 18460
rect 8331 18500 8373 18509
rect 12874 18502 12883 18542
rect 12923 18502 12932 18542
rect 13131 18535 13173 18544
rect 13498 18584 13556 18585
rect 13498 18544 13507 18584
rect 13547 18544 13556 18584
rect 13498 18543 13556 18544
rect 13899 18584 13941 18593
rect 13899 18544 13900 18584
rect 13940 18544 13941 18584
rect 13899 18535 13941 18544
rect 14038 18584 14080 18593
rect 14038 18544 14039 18584
rect 14079 18544 14080 18584
rect 14038 18535 14080 18544
rect 14283 18584 14325 18593
rect 14283 18544 14284 18584
rect 14324 18544 14325 18584
rect 14283 18535 14325 18544
rect 14763 18584 14805 18593
rect 15435 18584 15477 18593
rect 14763 18544 14764 18584
rect 14804 18544 14805 18584
rect 14763 18535 14805 18544
rect 14859 18575 14901 18584
rect 14859 18535 14860 18575
rect 14900 18535 14901 18575
rect 14859 18526 14901 18535
rect 15138 18575 15184 18584
rect 15138 18535 15139 18575
rect 15179 18535 15184 18575
rect 15435 18544 15436 18584
rect 15476 18544 15477 18584
rect 15435 18535 15477 18544
rect 15766 18584 15808 18593
rect 15766 18544 15767 18584
rect 15807 18544 15808 18584
rect 15766 18535 15808 18544
rect 16011 18584 16053 18593
rect 16011 18544 16012 18584
rect 16052 18544 16053 18584
rect 16011 18535 16053 18544
rect 16315 18584 16373 18585
rect 16315 18544 16324 18584
rect 16364 18544 16373 18584
rect 16315 18543 16373 18544
rect 16474 18584 16532 18585
rect 16474 18544 16483 18584
rect 16523 18544 16532 18584
rect 16474 18543 16532 18544
rect 16599 18584 16641 18593
rect 16599 18544 16600 18584
rect 16640 18544 16641 18584
rect 16599 18535 16641 18544
rect 16757 18584 16815 18585
rect 16757 18544 16766 18584
rect 16806 18544 16815 18584
rect 16757 18543 16815 18544
rect 16858 18584 16916 18585
rect 16858 18544 16867 18584
rect 16907 18544 16916 18584
rect 16858 18543 16916 18544
rect 17083 18584 17141 18585
rect 17083 18544 17092 18584
rect 17132 18544 17141 18584
rect 17083 18543 17141 18544
rect 17242 18584 17300 18585
rect 17242 18544 17251 18584
rect 17291 18544 17300 18584
rect 17242 18543 17300 18544
rect 17367 18584 17409 18593
rect 17367 18544 17368 18584
rect 17408 18544 17409 18584
rect 17632 18584 17690 18585
rect 17367 18535 17409 18544
rect 17526 18573 17584 18574
rect 15138 18526 15184 18535
rect 17526 18533 17535 18573
rect 17575 18533 17584 18573
rect 17632 18544 17641 18584
rect 17681 18544 17690 18584
rect 17632 18543 17690 18544
rect 18219 18584 18261 18593
rect 18219 18544 18220 18584
rect 18260 18544 18261 18584
rect 18219 18535 18261 18544
rect 18874 18584 18932 18585
rect 18874 18544 18883 18584
rect 18923 18544 18932 18584
rect 18874 18543 18932 18544
rect 21082 18584 21140 18585
rect 21082 18544 21091 18584
rect 21131 18544 21140 18584
rect 21082 18543 21140 18544
rect 22093 18584 22151 18585
rect 22093 18544 22102 18584
rect 22142 18544 22151 18584
rect 22539 18584 22581 18593
rect 22093 18543 22151 18544
rect 22327 18576 22385 18577
rect 22327 18536 22336 18576
rect 22376 18536 22385 18576
rect 22327 18535 22385 18536
rect 22539 18544 22540 18584
rect 22580 18544 22581 18584
rect 22539 18535 22581 18544
rect 22827 18584 22869 18593
rect 22827 18544 22828 18584
rect 22868 18544 22869 18584
rect 22827 18535 22869 18544
rect 23194 18584 23252 18585
rect 23194 18544 23203 18584
rect 23243 18544 23252 18584
rect 23194 18543 23252 18544
rect 25690 18584 25748 18585
rect 25690 18544 25699 18584
rect 25739 18544 25748 18584
rect 25690 18543 25748 18544
rect 27819 18584 27861 18593
rect 27819 18544 27820 18584
rect 27860 18544 27861 18584
rect 27819 18535 27861 18544
rect 27994 18584 28052 18585
rect 27994 18544 28003 18584
rect 28043 18544 28052 18584
rect 27994 18543 28052 18544
rect 28587 18584 28629 18593
rect 28587 18544 28588 18584
rect 28628 18544 28629 18584
rect 28587 18535 28629 18544
rect 28779 18584 28821 18593
rect 28779 18544 28780 18584
rect 28820 18544 28821 18584
rect 28779 18535 28821 18544
rect 29067 18584 29109 18593
rect 29067 18544 29068 18584
rect 29108 18544 29109 18584
rect 29067 18535 29109 18544
rect 17526 18532 17584 18533
rect 12874 18501 12932 18502
rect 9514 18500 9572 18501
rect 8331 18460 8332 18500
rect 8372 18460 8373 18500
rect 8331 18451 8373 18460
rect 8562 18491 8608 18500
rect 8562 18451 8563 18491
rect 8603 18451 8608 18491
rect 9514 18460 9523 18500
rect 9563 18460 9572 18500
rect 9514 18459 9572 18460
rect 13419 18500 13461 18509
rect 13419 18460 13420 18500
rect 13460 18460 13461 18500
rect 13419 18451 13461 18460
rect 14170 18500 14228 18501
rect 14170 18460 14179 18500
rect 14219 18460 14228 18500
rect 14170 18459 14228 18460
rect 14379 18500 14421 18509
rect 14379 18460 14380 18500
rect 14420 18460 14421 18500
rect 14379 18451 14421 18460
rect 15322 18500 15380 18501
rect 15322 18460 15331 18500
rect 15371 18460 15380 18500
rect 15322 18459 15380 18460
rect 15898 18500 15956 18501
rect 15898 18460 15907 18500
rect 15947 18460 15956 18500
rect 15898 18459 15956 18460
rect 21898 18500 21956 18501
rect 21898 18460 21907 18500
rect 21947 18460 21956 18500
rect 21898 18459 21956 18460
rect 24747 18500 24789 18509
rect 24747 18460 24748 18500
rect 24788 18460 24789 18500
rect 24747 18451 24789 18460
rect 27243 18500 27285 18509
rect 27243 18460 27244 18500
rect 27284 18460 27285 18500
rect 27243 18451 27285 18460
rect 5778 18442 5824 18451
rect 8562 18442 8608 18451
rect 6202 18416 6260 18417
rect 6202 18376 6211 18416
rect 6251 18376 6260 18416
rect 6202 18375 6260 18376
rect 7947 18416 7989 18425
rect 7947 18376 7948 18416
rect 7988 18376 7989 18416
rect 7947 18367 7989 18376
rect 9099 18416 9141 18425
rect 9099 18376 9100 18416
rect 9140 18376 9141 18416
rect 9099 18367 9141 18376
rect 10426 18416 10484 18417
rect 10426 18376 10435 18416
rect 10475 18376 10484 18416
rect 10426 18375 10484 18376
rect 20427 18416 20469 18425
rect 20427 18376 20428 18416
rect 20468 18376 20469 18416
rect 20427 18367 20469 18376
rect 20811 18416 20853 18425
rect 20811 18376 20812 18416
rect 20852 18376 20853 18416
rect 20811 18367 20853 18376
rect 28203 18416 28245 18425
rect 28203 18376 28204 18416
rect 28244 18376 28245 18416
rect 28203 18367 28245 18376
rect 28683 18416 28725 18425
rect 28683 18376 28684 18416
rect 28724 18376 28725 18416
rect 28683 18367 28725 18376
rect 5211 18332 5253 18341
rect 5211 18292 5212 18332
rect 5252 18292 5253 18332
rect 5211 18283 5253 18292
rect 6970 18332 7028 18333
rect 6970 18292 6979 18332
rect 7019 18292 7028 18332
rect 6970 18291 7028 18292
rect 9963 18332 10005 18341
rect 9963 18292 9964 18332
rect 10004 18292 10005 18332
rect 9963 18283 10005 18292
rect 11019 18332 11061 18341
rect 11019 18292 11020 18332
rect 11060 18292 11061 18332
rect 11019 18283 11061 18292
rect 11979 18332 12021 18341
rect 11979 18292 11980 18332
rect 12020 18292 12021 18332
rect 11979 18283 12021 18292
rect 12987 18332 13029 18341
rect 12987 18292 12988 18332
rect 13028 18292 13029 18332
rect 12987 18283 13029 18292
rect 14554 18332 14612 18333
rect 14554 18292 14563 18332
rect 14603 18292 14612 18332
rect 14554 18291 14612 18292
rect 16875 18332 16917 18341
rect 16875 18292 16876 18332
rect 16916 18292 16917 18332
rect 16875 18283 16917 18292
rect 21291 18332 21333 18341
rect 21291 18292 21292 18332
rect 21332 18292 21333 18332
rect 21291 18283 21333 18292
rect 27627 18332 27669 18341
rect 27627 18292 27628 18332
rect 27668 18292 27669 18332
rect 27627 18283 27669 18292
rect 28923 18332 28965 18341
rect 28923 18292 28924 18332
rect 28964 18292 28965 18332
rect 28923 18283 28965 18292
rect 576 18164 31392 18188
rect 576 18124 3112 18164
rect 3480 18124 10886 18164
rect 11254 18124 18660 18164
rect 19028 18124 26434 18164
rect 26802 18124 31392 18164
rect 576 18100 31392 18124
rect 730 17996 788 17997
rect 730 17956 739 17996
rect 779 17956 788 17996
rect 730 17955 788 17956
rect 1995 17996 2037 18005
rect 1995 17956 1996 17996
rect 2036 17956 2037 17996
rect 1995 17947 2037 17956
rect 3322 17996 3380 17997
rect 3322 17956 3331 17996
rect 3371 17956 3380 17996
rect 3322 17955 3380 17956
rect 3802 17996 3860 17997
rect 3802 17956 3811 17996
rect 3851 17956 3860 17996
rect 3802 17955 3860 17956
rect 5434 17996 5492 17997
rect 5434 17956 5443 17996
rect 5483 17956 5492 17996
rect 5434 17955 5492 17956
rect 11578 17996 11636 17997
rect 11578 17956 11587 17996
rect 11627 17956 11636 17996
rect 11578 17955 11636 17956
rect 15915 17996 15957 18005
rect 15915 17956 15916 17996
rect 15956 17956 15957 17996
rect 15915 17947 15957 17956
rect 23578 17996 23636 17997
rect 23578 17956 23587 17996
rect 23627 17956 23636 17996
rect 23578 17955 23636 17956
rect 1707 17912 1749 17921
rect 1707 17872 1708 17912
rect 1748 17872 1749 17912
rect 1707 17863 1749 17872
rect 5067 17912 5109 17921
rect 5067 17872 5068 17912
rect 5108 17872 5109 17912
rect 5067 17863 5109 17872
rect 6411 17912 6453 17921
rect 9675 17912 9717 17921
rect 6411 17872 6412 17912
rect 6452 17872 6453 17912
rect 6411 17863 6453 17872
rect 7019 17903 7061 17912
rect 7019 17863 7020 17903
rect 7060 17863 7061 17903
rect 9675 17872 9676 17912
rect 9716 17872 9717 17912
rect 9675 17863 9717 17872
rect 17931 17912 17973 17921
rect 17931 17872 17932 17912
rect 17972 17872 17973 17912
rect 17931 17863 17973 17872
rect 21195 17912 21237 17921
rect 21195 17872 21196 17912
rect 21236 17872 21237 17912
rect 21195 17863 21237 17872
rect 24267 17912 24309 17921
rect 24267 17872 24268 17912
rect 24308 17872 24309 17912
rect 24267 17863 24309 17872
rect 25131 17912 25173 17921
rect 25131 17872 25132 17912
rect 25172 17872 25173 17912
rect 25131 17863 25173 17872
rect 26859 17912 26901 17921
rect 26859 17872 26860 17912
rect 26900 17872 26901 17912
rect 26859 17863 26901 17872
rect 27627 17912 27669 17921
rect 27627 17872 27628 17912
rect 27668 17872 27669 17912
rect 27627 17863 27669 17872
rect 28011 17912 28053 17921
rect 28011 17872 28012 17912
rect 28052 17872 28053 17912
rect 28011 17863 28053 17872
rect 7019 17854 7061 17863
rect 1227 17828 1269 17837
rect 1227 17788 1228 17828
rect 1268 17788 1269 17828
rect 1227 17779 1269 17788
rect 1803 17828 1845 17837
rect 1803 17788 1804 17828
rect 1844 17788 1845 17828
rect 1803 17779 1845 17788
rect 2594 17828 2636 17837
rect 2594 17788 2595 17828
rect 2635 17788 2636 17828
rect 2594 17779 2636 17788
rect 3074 17828 3116 17837
rect 3074 17788 3075 17828
rect 3115 17788 3116 17828
rect 5163 17828 5205 17837
rect 3074 17779 3116 17788
rect 4971 17786 5013 17795
rect 939 17744 981 17753
rect 939 17704 940 17744
rect 980 17704 981 17744
rect 939 17695 981 17704
rect 1027 17744 1085 17745
rect 1027 17704 1036 17744
rect 1076 17704 1085 17744
rect 1027 17703 1085 17704
rect 1402 17744 1460 17745
rect 1402 17704 1411 17744
rect 1451 17704 1460 17744
rect 1402 17703 1460 17704
rect 1995 17744 2037 17753
rect 1995 17704 1996 17744
rect 2036 17704 2037 17744
rect 1995 17695 2037 17704
rect 2187 17744 2229 17753
rect 2187 17704 2188 17744
rect 2228 17704 2229 17744
rect 2187 17695 2229 17704
rect 2475 17744 2517 17753
rect 2475 17704 2476 17744
rect 2516 17704 2517 17744
rect 2475 17695 2517 17704
rect 2704 17744 2762 17745
rect 2704 17704 2713 17744
rect 2753 17704 2762 17744
rect 2704 17703 2762 17704
rect 2955 17744 2997 17753
rect 4971 17746 4972 17786
rect 5012 17746 5013 17786
rect 5163 17788 5164 17828
rect 5204 17788 5205 17828
rect 5163 17779 5205 17788
rect 6507 17828 6549 17837
rect 6507 17788 6508 17828
rect 6548 17788 6549 17828
rect 6507 17779 6549 17788
rect 12290 17828 12332 17837
rect 12290 17788 12291 17828
rect 12331 17788 12332 17828
rect 12290 17779 12332 17788
rect 13154 17828 13196 17837
rect 13154 17788 13155 17828
rect 13195 17788 13196 17828
rect 13154 17779 13196 17788
rect 13498 17828 13556 17829
rect 13498 17788 13507 17828
rect 13547 17788 13556 17828
rect 13498 17787 13556 17788
rect 14667 17828 14709 17837
rect 14667 17788 14668 17828
rect 14708 17788 14709 17828
rect 14667 17779 14709 17788
rect 18891 17828 18933 17837
rect 18891 17788 18892 17828
rect 18932 17788 18933 17828
rect 18891 17779 18933 17788
rect 20811 17828 20853 17837
rect 20811 17788 20812 17828
rect 20852 17788 20853 17828
rect 20811 17779 20853 17788
rect 22234 17828 22292 17829
rect 22234 17788 22243 17828
rect 22283 17788 22292 17828
rect 22234 17787 22292 17788
rect 23787 17828 23829 17837
rect 23787 17788 23788 17828
rect 23828 17788 23829 17828
rect 23787 17779 23829 17788
rect 24363 17828 24405 17837
rect 24363 17788 24364 17828
rect 24404 17788 24405 17828
rect 24363 17779 24405 17788
rect 2955 17704 2956 17744
rect 2996 17704 2997 17744
rect 2955 17695 2997 17704
rect 3184 17744 3242 17745
rect 3184 17704 3193 17744
rect 3233 17704 3242 17744
rect 3184 17703 3242 17704
rect 3619 17744 3677 17745
rect 3619 17704 3628 17744
rect 3668 17704 3677 17744
rect 3619 17703 3677 17704
rect 4099 17744 4157 17745
rect 4099 17704 4108 17744
rect 4148 17704 4157 17744
rect 4099 17703 4157 17704
rect 4714 17744 4772 17745
rect 4714 17704 4723 17744
rect 4763 17704 4772 17744
rect 4714 17703 4772 17704
rect 4836 17744 4894 17745
rect 4836 17704 4845 17744
rect 4885 17704 4894 17744
rect 4971 17737 5013 17746
rect 5547 17755 5589 17764
rect 5290 17744 5348 17745
rect 4836 17703 4894 17704
rect 5290 17704 5299 17744
rect 5339 17704 5348 17744
rect 5290 17703 5348 17704
rect 5434 17744 5492 17745
rect 5434 17704 5443 17744
rect 5483 17704 5492 17744
rect 5547 17715 5548 17755
rect 5588 17715 5589 17755
rect 13995 17755 14037 17764
rect 5547 17706 5589 17715
rect 5826 17744 5884 17745
rect 5434 17703 5492 17704
rect 5826 17704 5835 17744
rect 5875 17704 5884 17744
rect 5826 17703 5884 17704
rect 5962 17744 6020 17745
rect 5962 17704 5971 17744
rect 6011 17704 6020 17744
rect 5962 17703 6020 17704
rect 6180 17744 6238 17745
rect 6180 17704 6189 17744
rect 6229 17704 6238 17744
rect 6180 17703 6238 17704
rect 6350 17744 6392 17753
rect 6350 17704 6351 17744
rect 6391 17704 6392 17744
rect 5730 17693 5776 17702
rect 6350 17695 6392 17704
rect 6634 17744 6692 17745
rect 6634 17704 6643 17744
rect 6683 17704 6692 17744
rect 6634 17703 6692 17704
rect 6970 17744 7028 17745
rect 6970 17704 6979 17744
rect 7019 17704 7028 17744
rect 6970 17703 7028 17704
rect 7291 17744 7349 17745
rect 7291 17704 7300 17744
rect 7340 17704 7349 17744
rect 7291 17703 7349 17704
rect 7450 17744 7508 17745
rect 7450 17704 7459 17744
rect 7499 17704 7508 17744
rect 7450 17703 7508 17704
rect 7575 17744 7617 17753
rect 7575 17704 7576 17744
rect 7616 17704 7617 17744
rect 7575 17695 7617 17704
rect 7706 17744 7764 17745
rect 7706 17704 7715 17744
rect 7755 17704 7764 17744
rect 7706 17703 7764 17704
rect 7834 17744 7892 17745
rect 7834 17704 7843 17744
rect 7883 17704 7892 17744
rect 7834 17703 7892 17704
rect 8215 17744 8273 17745
rect 8215 17704 8224 17744
rect 8264 17704 8273 17744
rect 8215 17703 8273 17704
rect 9007 17744 9065 17745
rect 9007 17704 9016 17744
rect 9056 17704 9065 17744
rect 9007 17703 9065 17704
rect 9195 17744 9237 17753
rect 9195 17704 9196 17744
rect 9236 17704 9237 17744
rect 9195 17695 9237 17704
rect 9562 17744 9620 17745
rect 9562 17704 9571 17744
rect 9611 17704 9620 17744
rect 9562 17703 9620 17704
rect 9946 17744 10004 17745
rect 9946 17704 9955 17744
rect 9995 17704 10004 17744
rect 9946 17703 10004 17704
rect 10251 17744 10293 17753
rect 10251 17704 10252 17744
rect 10292 17704 10293 17744
rect 10251 17695 10293 17704
rect 10539 17744 10581 17753
rect 10539 17704 10540 17744
rect 10580 17704 10581 17744
rect 10539 17695 10581 17704
rect 10731 17744 10773 17753
rect 10731 17704 10732 17744
rect 10772 17704 10773 17744
rect 10731 17695 10773 17704
rect 11095 17744 11153 17745
rect 11095 17704 11104 17744
rect 11144 17704 11153 17744
rect 11095 17703 11153 17704
rect 11787 17744 11829 17753
rect 11787 17704 11788 17744
rect 11828 17704 11829 17744
rect 11787 17695 11829 17704
rect 11875 17744 11933 17745
rect 11875 17704 11884 17744
rect 11924 17704 11933 17744
rect 11875 17703 11933 17704
rect 12171 17744 12213 17753
rect 12171 17704 12172 17744
rect 12212 17704 12213 17744
rect 12171 17695 12213 17704
rect 12411 17744 12453 17753
rect 12411 17704 12412 17744
rect 12452 17704 12453 17744
rect 12411 17695 12453 17704
rect 12555 17744 12597 17753
rect 12555 17704 12556 17744
rect 12596 17704 12597 17744
rect 12555 17695 12597 17704
rect 12747 17744 12789 17753
rect 12747 17704 12748 17744
rect 12788 17704 12789 17744
rect 12747 17695 12789 17704
rect 13035 17744 13077 17753
rect 13035 17704 13036 17744
rect 13076 17704 13077 17744
rect 13035 17695 13077 17704
rect 13264 17744 13322 17745
rect 13264 17704 13273 17744
rect 13313 17704 13322 17744
rect 13264 17703 13322 17704
rect 13380 17744 13422 17753
rect 13380 17704 13381 17744
rect 13421 17704 13422 17744
rect 13380 17695 13422 17704
rect 13611 17744 13653 17753
rect 13611 17704 13612 17744
rect 13652 17704 13653 17744
rect 13611 17695 13653 17704
rect 13882 17744 13940 17745
rect 13882 17704 13891 17744
rect 13931 17704 13940 17744
rect 13995 17715 13996 17755
rect 14036 17715 14037 17755
rect 13995 17706 14037 17715
rect 14140 17744 14198 17745
rect 13882 17703 13940 17704
rect 14140 17704 14149 17744
rect 14189 17704 14198 17744
rect 14140 17703 14198 17704
rect 14269 17744 14311 17753
rect 14269 17704 14270 17744
rect 14310 17704 14311 17744
rect 14269 17695 14311 17704
rect 14443 17744 14501 17745
rect 14443 17704 14452 17744
rect 14492 17704 14501 17744
rect 14443 17703 14501 17704
rect 14772 17744 14814 17753
rect 15003 17744 15045 17753
rect 14772 17704 14773 17744
rect 14813 17704 14814 17744
rect 14772 17695 14814 17704
rect 14898 17735 14944 17744
rect 14898 17695 14899 17735
rect 14939 17695 14944 17735
rect 15003 17704 15004 17744
rect 15044 17704 15045 17744
rect 15003 17695 15045 17704
rect 15355 17744 15413 17745
rect 15355 17704 15364 17744
rect 15404 17704 15413 17744
rect 15355 17703 15413 17704
rect 15514 17744 15572 17745
rect 15514 17704 15523 17744
rect 15563 17704 15572 17744
rect 15514 17703 15572 17704
rect 15639 17744 15681 17753
rect 15639 17704 15640 17744
rect 15680 17704 15681 17744
rect 15639 17695 15681 17704
rect 15802 17744 15860 17745
rect 15802 17704 15811 17744
rect 15851 17704 15860 17744
rect 15802 17703 15860 17704
rect 15924 17744 15982 17745
rect 15924 17704 15933 17744
rect 15973 17704 15982 17744
rect 15924 17703 15982 17704
rect 16102 17744 16144 17753
rect 16102 17704 16103 17744
rect 16143 17704 16144 17744
rect 16102 17695 16144 17704
rect 16282 17744 16340 17745
rect 16282 17704 16291 17744
rect 16331 17704 16340 17744
rect 16282 17703 16340 17704
rect 16587 17744 16629 17753
rect 16587 17704 16588 17744
rect 16628 17704 16629 17744
rect 16587 17695 16629 17704
rect 16762 17744 16820 17745
rect 16762 17704 16771 17744
rect 16811 17704 16820 17744
rect 16762 17703 16820 17704
rect 17263 17744 17321 17745
rect 17263 17704 17272 17744
rect 17312 17704 17321 17744
rect 17263 17703 17321 17704
rect 17401 17744 17459 17745
rect 17401 17704 17410 17744
rect 17450 17704 17459 17744
rect 17401 17703 17459 17704
rect 17932 17744 17974 17753
rect 17932 17704 17933 17744
rect 17973 17704 17974 17744
rect 17932 17695 17974 17704
rect 18123 17744 18165 17753
rect 18123 17704 18124 17744
rect 18164 17704 18165 17744
rect 18123 17695 18165 17704
rect 18394 17744 18452 17745
rect 18394 17704 18403 17744
rect 18443 17704 18452 17744
rect 18394 17703 18452 17704
rect 18507 17744 18549 17753
rect 18507 17704 18508 17744
rect 18548 17704 18549 17744
rect 18507 17695 18549 17704
rect 18987 17744 19029 17753
rect 18987 17704 18988 17744
rect 19028 17704 19029 17744
rect 18987 17695 19029 17704
rect 19459 17744 19517 17745
rect 19459 17704 19468 17744
rect 19508 17704 19517 17744
rect 19459 17703 19517 17704
rect 19978 17744 20036 17745
rect 19978 17704 19987 17744
rect 20027 17704 20036 17744
rect 19978 17703 20036 17704
rect 20331 17744 20373 17753
rect 21867 17744 21909 17753
rect 20331 17704 20332 17744
rect 20372 17704 20373 17744
rect 20331 17695 20373 17704
rect 21579 17735 21621 17744
rect 21579 17695 21580 17735
rect 21620 17695 21621 17735
rect 21867 17704 21868 17744
rect 21908 17704 21909 17744
rect 21867 17695 21909 17704
rect 22102 17744 22144 17753
rect 22102 17704 22103 17744
rect 22143 17704 22144 17744
rect 22102 17695 22144 17704
rect 22347 17744 22389 17753
rect 22347 17704 22348 17744
rect 22388 17704 22389 17744
rect 22347 17695 22389 17704
rect 23215 17744 23273 17745
rect 23215 17704 23224 17744
rect 23264 17704 23273 17744
rect 23215 17703 23273 17704
rect 23398 17744 23440 17753
rect 23398 17704 23399 17744
rect 23439 17704 23440 17744
rect 23398 17695 23440 17704
rect 23578 17744 23636 17745
rect 23578 17704 23587 17744
rect 23627 17704 23636 17744
rect 23578 17703 23636 17704
rect 23962 17744 24020 17745
rect 23962 17704 23971 17744
rect 24011 17704 24020 17744
rect 23962 17703 24020 17704
rect 24730 17744 24788 17745
rect 24730 17704 24739 17744
rect 24779 17704 24788 17744
rect 24730 17703 24788 17704
rect 25711 17744 25769 17745
rect 25711 17704 25720 17744
rect 25760 17704 25769 17744
rect 25711 17703 25769 17704
rect 25995 17744 26037 17753
rect 25995 17704 25996 17744
rect 26036 17704 26037 17744
rect 25995 17695 26037 17704
rect 26667 17744 26709 17753
rect 26667 17704 26668 17744
rect 26708 17704 26709 17744
rect 26667 17695 26709 17704
rect 27243 17744 27285 17753
rect 27243 17704 27244 17744
rect 27284 17704 27285 17744
rect 27243 17695 27285 17704
rect 27435 17744 27477 17753
rect 27435 17704 27436 17744
rect 27476 17704 27477 17744
rect 27435 17695 27477 17704
rect 736 17660 778 17669
rect 736 17620 737 17660
rect 777 17620 778 17660
rect 736 17611 778 17620
rect 3328 17660 3370 17669
rect 3328 17620 3329 17660
rect 3369 17620 3370 17660
rect 3328 17611 3370 17620
rect 3808 17660 3850 17669
rect 3808 17620 3809 17660
rect 3849 17620 3850 17660
rect 5730 17653 5731 17693
rect 5771 17653 5776 17693
rect 14898 17686 14944 17695
rect 21579 17686 21621 17695
rect 5730 17644 5776 17653
rect 6795 17660 6837 17669
rect 3808 17611 3850 17620
rect 6795 17620 6796 17660
rect 6836 17620 6837 17660
rect 6795 17611 6837 17620
rect 11581 17660 11623 17669
rect 11581 17620 11582 17660
rect 11622 17620 11623 17660
rect 11581 17611 11623 17620
rect 13690 17660 13748 17661
rect 13690 17620 13699 17660
rect 13739 17620 13748 17660
rect 13690 17619 13748 17620
rect 16683 17660 16725 17669
rect 16683 17620 16684 17660
rect 16724 17620 16725 17660
rect 16683 17611 16725 17620
rect 17595 17660 17637 17669
rect 17595 17620 17596 17660
rect 17636 17620 17637 17660
rect 17595 17611 17637 17620
rect 20475 17660 20517 17669
rect 20475 17620 20476 17660
rect 20516 17620 20517 17660
rect 20475 17611 20517 17620
rect 21483 17660 21525 17669
rect 21483 17620 21484 17660
rect 21524 17620 21525 17660
rect 21483 17611 21525 17620
rect 2379 17576 2421 17585
rect 2379 17536 2380 17576
rect 2420 17536 2421 17576
rect 2379 17527 2421 17536
rect 2859 17576 2901 17585
rect 2859 17536 2860 17576
rect 2900 17536 2901 17576
rect 2859 17527 2901 17536
rect 3531 17576 3573 17585
rect 3531 17536 3532 17576
rect 3572 17536 3573 17576
rect 3531 17527 3573 17536
rect 4011 17576 4053 17585
rect 4011 17536 4012 17576
rect 4052 17536 4053 17576
rect 4011 17527 4053 17536
rect 4522 17576 4580 17577
rect 4522 17536 4531 17576
rect 4571 17536 4580 17576
rect 4522 17535 4580 17536
rect 7354 17576 7412 17577
rect 7354 17536 7363 17576
rect 7403 17536 7412 17576
rect 7354 17535 7412 17536
rect 8379 17576 8421 17585
rect 8379 17536 8380 17576
rect 8420 17536 8421 17576
rect 8379 17527 8421 17536
rect 8842 17576 8900 17577
rect 8842 17536 8851 17576
rect 8891 17536 8900 17576
rect 8842 17535 8900 17536
rect 10155 17576 10197 17585
rect 10155 17536 10156 17576
rect 10196 17536 10197 17576
rect 10155 17527 10197 17536
rect 10635 17576 10677 17585
rect 10635 17536 10636 17576
rect 10676 17536 10677 17576
rect 10635 17527 10677 17536
rect 11259 17576 11301 17585
rect 11259 17536 11260 17576
rect 11300 17536 11301 17576
rect 11259 17527 11301 17536
rect 12075 17576 12117 17585
rect 12075 17536 12076 17576
rect 12116 17536 12117 17576
rect 12075 17527 12117 17536
rect 12555 17576 12597 17585
rect 12555 17536 12556 17576
rect 12596 17536 12597 17576
rect 12555 17527 12597 17536
rect 12939 17576 12981 17585
rect 12939 17536 12940 17576
rect 12980 17536 12981 17576
rect 12939 17527 12981 17536
rect 14266 17576 14324 17577
rect 14266 17536 14275 17576
rect 14315 17536 14324 17576
rect 14266 17535 14324 17536
rect 16203 17576 16245 17585
rect 16203 17536 16204 17576
rect 16244 17536 16245 17576
rect 16203 17527 16245 17536
rect 17098 17576 17156 17577
rect 17098 17536 17107 17576
rect 17147 17536 17156 17576
rect 17098 17535 17156 17536
rect 20139 17576 20181 17585
rect 20139 17536 20140 17576
rect 20180 17536 20181 17576
rect 20139 17527 20181 17536
rect 20571 17576 20613 17585
rect 20571 17536 20572 17576
rect 20612 17536 20613 17576
rect 20571 17527 20613 17536
rect 22426 17576 22484 17577
rect 22426 17536 22435 17576
rect 22475 17536 22484 17576
rect 22426 17535 22484 17536
rect 23050 17576 23108 17577
rect 23050 17536 23059 17576
rect 23099 17536 23108 17576
rect 23050 17535 23108 17536
rect 24939 17576 24981 17585
rect 24939 17536 24940 17576
rect 24980 17536 24981 17576
rect 24939 17527 24981 17536
rect 25546 17576 25604 17577
rect 25546 17536 25555 17576
rect 25595 17536 25604 17576
rect 25546 17535 25604 17536
rect 27339 17576 27381 17585
rect 27339 17536 27340 17576
rect 27380 17536 27381 17576
rect 27339 17527 27381 17536
rect 576 17408 31392 17432
rect 576 17368 4352 17408
rect 4720 17368 12126 17408
rect 12494 17368 19900 17408
rect 20268 17368 27674 17408
rect 28042 17368 31392 17408
rect 576 17344 31392 17368
rect 1611 17240 1653 17249
rect 1611 17200 1612 17240
rect 1652 17200 1653 17240
rect 1611 17191 1653 17200
rect 3147 17240 3189 17249
rect 3147 17200 3148 17240
rect 3188 17200 3189 17240
rect 3147 17191 3189 17200
rect 3531 17240 3573 17249
rect 3531 17200 3532 17240
rect 3572 17200 3573 17240
rect 3531 17191 3573 17200
rect 4875 17240 4917 17249
rect 4875 17200 4876 17240
rect 4916 17200 4917 17240
rect 6298 17240 6356 17241
rect 4875 17191 4917 17200
rect 5367 17198 5409 17207
rect 6298 17200 6307 17240
rect 6347 17200 6356 17240
rect 6298 17199 6356 17200
rect 10923 17240 10965 17249
rect 10923 17200 10924 17240
rect 10964 17200 10965 17240
rect 928 17156 970 17165
rect 928 17116 929 17156
rect 969 17116 970 17156
rect 928 17107 970 17116
rect 1721 17156 1763 17165
rect 1721 17116 1722 17156
rect 1762 17116 1763 17156
rect 1721 17107 1763 17116
rect 1899 17156 1941 17165
rect 1899 17116 1900 17156
rect 1940 17116 1941 17156
rect 1899 17107 1941 17116
rect 4203 17156 4245 17165
rect 4203 17116 4204 17156
rect 4244 17116 4245 17156
rect 5367 17158 5368 17198
rect 5408 17158 5409 17198
rect 10923 17191 10965 17200
rect 11674 17240 11732 17241
rect 11674 17200 11683 17240
rect 11723 17200 11732 17240
rect 11674 17199 11732 17200
rect 11962 17240 12020 17241
rect 11962 17200 11971 17240
rect 12011 17200 12020 17240
rect 11962 17199 12020 17200
rect 12826 17240 12884 17241
rect 12826 17200 12835 17240
rect 12875 17200 12884 17240
rect 12826 17199 12884 17200
rect 14074 17240 14132 17241
rect 14074 17200 14083 17240
rect 14123 17200 14132 17240
rect 14074 17199 14132 17200
rect 15418 17240 15476 17241
rect 15418 17200 15427 17240
rect 15467 17200 15476 17240
rect 15418 17199 15476 17200
rect 17067 17240 17109 17249
rect 17067 17200 17068 17240
rect 17108 17200 17109 17240
rect 17067 17191 17109 17200
rect 18315 17240 18357 17249
rect 18315 17200 18316 17240
rect 18356 17200 18357 17240
rect 18315 17191 18357 17200
rect 5367 17149 5409 17158
rect 8043 17156 8085 17165
rect 13046 17156 13088 17165
rect 4203 17107 4245 17116
rect 8043 17116 8044 17156
rect 8084 17116 8085 17156
rect 8043 17107 8085 17116
rect 12258 17147 12304 17156
rect 12258 17107 12259 17147
rect 12299 17107 12304 17147
rect 13046 17116 13047 17156
rect 13087 17116 13088 17156
rect 13046 17107 13088 17116
rect 17482 17156 17540 17157
rect 17482 17116 17491 17156
rect 17531 17116 17540 17156
rect 17482 17115 17540 17116
rect 21003 17156 21045 17165
rect 21003 17116 21004 17156
rect 21044 17116 21045 17156
rect 14746 17114 14804 17115
rect 12258 17098 12304 17107
rect 13642 17105 13700 17110
rect 1131 17072 1173 17081
rect 1402 17072 1460 17073
rect 1131 17032 1132 17072
rect 1172 17032 1173 17072
rect 1131 17023 1173 17032
rect 1227 17063 1269 17072
rect 1227 17023 1228 17063
rect 1268 17023 1269 17063
rect 1402 17032 1411 17072
rect 1451 17032 1460 17072
rect 1402 17031 1460 17032
rect 1515 17072 1557 17081
rect 1515 17032 1516 17072
rect 1556 17032 1557 17072
rect 1515 17023 1557 17032
rect 1995 17072 2037 17081
rect 2235 17072 2277 17081
rect 1995 17032 1996 17072
rect 2036 17032 2037 17072
rect 1995 17023 2037 17032
rect 2130 17063 2176 17072
rect 2130 17023 2131 17063
rect 2171 17023 2176 17063
rect 2235 17032 2236 17072
rect 2276 17032 2277 17072
rect 2235 17023 2277 17032
rect 2338 17072 2396 17073
rect 2338 17032 2347 17072
rect 2387 17032 2396 17072
rect 2338 17031 2396 17032
rect 2571 17072 2613 17081
rect 2571 17032 2572 17072
rect 2612 17032 2613 17072
rect 2571 17023 2613 17032
rect 3051 17072 3093 17081
rect 3051 17032 3052 17072
rect 3092 17032 3093 17072
rect 3051 17023 3093 17032
rect 3226 17072 3284 17073
rect 3226 17032 3235 17072
rect 3275 17032 3284 17072
rect 3226 17031 3284 17032
rect 3435 17072 3477 17081
rect 3435 17032 3436 17072
rect 3476 17032 3477 17072
rect 3435 17023 3477 17032
rect 3627 17072 3669 17081
rect 3627 17032 3628 17072
rect 3668 17032 3669 17072
rect 3627 17023 3669 17032
rect 3915 17072 3957 17081
rect 3915 17032 3916 17072
rect 3956 17032 3957 17072
rect 3915 17023 3957 17032
rect 4102 17072 4144 17081
rect 4102 17032 4103 17072
rect 4143 17032 4144 17072
rect 4102 17023 4144 17032
rect 4282 17072 4340 17073
rect 4282 17032 4291 17072
rect 4331 17032 4340 17072
rect 4282 17031 4340 17032
rect 4774 17072 4816 17081
rect 4774 17032 4775 17072
rect 4815 17032 4816 17072
rect 4774 17023 4816 17032
rect 4954 17072 5012 17073
rect 4954 17032 4963 17072
rect 5003 17032 5012 17072
rect 4954 17031 5012 17032
rect 5115 17072 5157 17081
rect 5115 17032 5116 17072
rect 5156 17032 5157 17072
rect 5698 17072 5756 17073
rect 5115 17023 5157 17032
rect 5287 17030 5329 17039
rect 5698 17032 5707 17072
rect 5747 17032 5756 17072
rect 5698 17031 5756 17032
rect 6146 17072 6188 17081
rect 6146 17032 6147 17072
rect 6187 17032 6188 17072
rect 1227 17014 1269 17023
rect 2130 17014 2176 17023
rect 2452 16988 2494 16997
rect 2452 16948 2453 16988
rect 2493 16948 2494 16988
rect 2452 16939 2494 16948
rect 2667 16988 2709 16997
rect 2667 16948 2668 16988
rect 2708 16948 2709 16988
rect 5287 16990 5288 17030
rect 5328 16990 5329 17030
rect 5578 17030 5636 17031
rect 5287 16981 5329 16990
rect 5461 16988 5503 16997
rect 5578 16990 5587 17030
rect 5627 16990 5636 17030
rect 6010 17030 6068 17031
rect 5578 16989 5636 16990
rect 2667 16939 2709 16948
rect 5461 16948 5462 16988
rect 5502 16948 5503 16988
rect 5461 16939 5503 16948
rect 5835 16988 5877 16997
rect 6010 16990 6019 17030
rect 6059 16990 6068 17030
rect 6146 17023 6188 17032
rect 6459 17072 6501 17081
rect 6459 17032 6460 17072
rect 6500 17032 6501 17072
rect 6459 17023 6501 17032
rect 6603 17072 6645 17081
rect 6603 17032 6604 17072
rect 6644 17032 6645 17072
rect 6603 17023 6645 17032
rect 7179 17072 7221 17081
rect 7851 17072 7893 17081
rect 7179 17032 7180 17072
rect 7220 17032 7221 17072
rect 7179 17023 7221 17032
rect 7314 17063 7360 17072
rect 7314 17023 7315 17063
rect 7355 17023 7360 17063
rect 7314 17014 7360 17023
rect 7419 17030 7461 17039
rect 6010 16989 6068 16990
rect 5835 16948 5836 16988
rect 5876 16948 5877 16988
rect 5835 16939 5877 16948
rect 7083 16988 7125 16997
rect 7083 16948 7084 16988
rect 7124 16948 7125 16988
rect 7419 16990 7420 17030
rect 7460 16990 7461 17030
rect 7851 17032 7852 17072
rect 7892 17032 7893 17072
rect 7851 17023 7893 17032
rect 8170 17072 8228 17073
rect 8170 17032 8179 17072
rect 8219 17032 8228 17072
rect 8170 17031 8228 17032
rect 8379 17072 8421 17081
rect 8379 17032 8380 17072
rect 8420 17032 8421 17072
rect 8379 17023 8421 17032
rect 8694 17072 8736 17081
rect 8694 17032 8695 17072
rect 8735 17032 8736 17072
rect 8694 17023 8736 17032
rect 8836 17072 8894 17073
rect 8836 17032 8845 17072
rect 8885 17032 8894 17072
rect 8836 17031 8894 17032
rect 8962 17072 9020 17073
rect 8962 17032 8971 17072
rect 9011 17032 9020 17072
rect 8962 17031 9020 17032
rect 9256 17072 9298 17081
rect 9256 17032 9257 17072
rect 9297 17032 9298 17072
rect 9256 17023 9298 17032
rect 9418 17072 9476 17073
rect 9418 17032 9427 17072
rect 9467 17032 9476 17072
rect 9418 17031 9476 17032
rect 9671 17072 9713 17081
rect 9671 17032 9672 17072
rect 9712 17032 9713 17072
rect 9671 17023 9713 17032
rect 9867 17072 9909 17081
rect 9867 17032 9868 17072
rect 9908 17032 9909 17072
rect 9867 17023 9909 17032
rect 10639 17072 10697 17073
rect 10639 17032 10648 17072
rect 10688 17032 10697 17072
rect 10639 17031 10697 17032
rect 11019 17072 11061 17081
rect 11019 17032 11020 17072
rect 11060 17032 11061 17072
rect 11019 17023 11061 17032
rect 11248 17072 11306 17073
rect 11248 17032 11257 17072
rect 11297 17032 11306 17072
rect 11248 17031 11306 17032
rect 11362 17072 11420 17073
rect 11362 17032 11371 17072
rect 11411 17032 11420 17072
rect 11362 17031 11420 17032
rect 11595 17072 11637 17081
rect 11595 17032 11596 17072
rect 11636 17032 11637 17072
rect 11595 17023 11637 17032
rect 11962 17072 12020 17073
rect 12346 17072 12404 17073
rect 11962 17032 11971 17072
rect 12011 17032 12020 17072
rect 11962 17031 12020 17032
rect 12075 17063 12117 17072
rect 12075 17023 12076 17063
rect 12116 17023 12117 17063
rect 12346 17032 12355 17072
rect 12395 17032 12404 17072
rect 12730 17072 12788 17073
rect 12346 17031 12404 17032
rect 12523 17061 12581 17062
rect 12075 17014 12117 17023
rect 12523 17021 12532 17061
rect 12572 17021 12581 17061
rect 12730 17032 12739 17072
rect 12779 17032 12788 17072
rect 12730 17031 12788 17032
rect 13323 17072 13365 17081
rect 13323 17032 13324 17072
rect 13364 17032 13365 17072
rect 13642 17065 13651 17105
rect 13691 17065 13700 17105
rect 13642 17064 13700 17065
rect 13995 17072 14037 17081
rect 13323 17023 13365 17032
rect 13995 17032 13996 17072
rect 14036 17032 14037 17072
rect 13995 17023 14037 17032
rect 14283 17072 14325 17081
rect 14746 17074 14755 17114
rect 14795 17074 14804 17114
rect 21003 17107 21045 17116
rect 21963 17156 22005 17165
rect 21963 17116 21964 17156
rect 22004 17116 22005 17156
rect 21963 17107 22005 17116
rect 28090 17156 28148 17157
rect 28090 17116 28099 17156
rect 28139 17116 28148 17156
rect 28090 17115 28148 17116
rect 23121 17105 23179 17110
rect 14746 17073 14804 17074
rect 14283 17032 14284 17072
rect 14324 17032 14325 17072
rect 14283 17023 14325 17032
rect 14458 17072 14516 17073
rect 14458 17032 14467 17072
rect 14507 17032 14516 17072
rect 14458 17031 14516 17032
rect 14880 17072 14922 17081
rect 14880 17032 14881 17072
rect 14921 17032 14922 17072
rect 14880 17023 14922 17032
rect 15178 17072 15236 17073
rect 15178 17032 15187 17072
rect 15227 17032 15236 17072
rect 15536 17072 15578 17081
rect 15178 17031 15236 17032
rect 15355 17061 15397 17070
rect 12523 17020 12581 17021
rect 15355 17021 15356 17061
rect 15396 17021 15397 17061
rect 15536 17032 15537 17072
rect 15577 17032 15578 17072
rect 15536 17023 15578 17032
rect 15658 17072 15716 17073
rect 15658 17032 15667 17072
rect 15707 17032 15716 17072
rect 15658 17031 15716 17032
rect 15802 17072 15860 17073
rect 15802 17032 15811 17072
rect 15851 17032 15860 17072
rect 16429 17072 16487 17073
rect 15802 17031 15860 17032
rect 15915 17061 15957 17070
rect 15355 17012 15397 17021
rect 15915 17021 15916 17061
rect 15956 17021 15957 17061
rect 16429 17032 16438 17072
rect 16478 17032 16487 17072
rect 16429 17031 16487 17032
rect 16587 17072 16629 17081
rect 16587 17032 16588 17072
rect 16628 17032 16629 17072
rect 16587 17023 16629 17032
rect 16779 17072 16821 17081
rect 16779 17032 16780 17072
rect 16820 17032 16821 17072
rect 16779 17023 16821 17032
rect 16972 17072 17014 17081
rect 16972 17032 16973 17072
rect 17013 17032 17014 17072
rect 16972 17023 17014 17032
rect 17156 17072 17198 17081
rect 17156 17032 17157 17072
rect 17197 17032 17198 17072
rect 17156 17023 17198 17032
rect 17677 17072 17735 17073
rect 17677 17032 17686 17072
rect 17726 17032 17735 17072
rect 17677 17031 17735 17032
rect 17931 17072 17973 17081
rect 17931 17032 17932 17072
rect 17972 17032 17973 17072
rect 17931 17023 17973 17032
rect 18123 17072 18165 17081
rect 18123 17032 18124 17072
rect 18164 17032 18165 17072
rect 18123 17023 18165 17032
rect 18490 17072 18548 17073
rect 19467 17072 19509 17081
rect 18490 17032 18499 17072
rect 18539 17032 18548 17072
rect 18490 17031 18548 17032
rect 18987 17063 19029 17072
rect 18987 17023 18988 17063
rect 19028 17023 19029 17063
rect 19467 17032 19468 17072
rect 19508 17032 19509 17072
rect 19467 17023 19509 17032
rect 19947 17072 19989 17081
rect 19947 17032 19948 17072
rect 19988 17032 19989 17072
rect 19947 17023 19989 17032
rect 20057 17072 20115 17073
rect 20057 17032 20066 17072
rect 20106 17032 20115 17072
rect 20057 17031 20115 17032
rect 20619 17072 20661 17081
rect 20619 17032 20620 17072
rect 20660 17032 20661 17072
rect 20619 17023 20661 17032
rect 20890 17072 20948 17073
rect 20890 17032 20899 17072
rect 20939 17032 20948 17072
rect 20890 17031 20948 17032
rect 22084 17072 22142 17073
rect 22084 17032 22093 17072
rect 22133 17032 22142 17072
rect 22084 17031 22142 17032
rect 22347 17072 22389 17081
rect 22347 17032 22348 17072
rect 22388 17032 22389 17072
rect 22347 17023 22389 17032
rect 23019 17072 23061 17081
rect 23019 17032 23020 17072
rect 23060 17032 23061 17072
rect 23121 17065 23130 17105
rect 23170 17065 23179 17105
rect 23121 17064 23179 17065
rect 23403 17072 23445 17081
rect 23019 17023 23061 17032
rect 23403 17032 23404 17072
rect 23444 17032 23445 17072
rect 23403 17023 23445 17032
rect 23962 17072 24020 17073
rect 24939 17072 24981 17081
rect 23962 17032 23971 17072
rect 24011 17032 24020 17072
rect 23962 17031 24020 17032
rect 24459 17063 24501 17072
rect 24459 17023 24460 17063
rect 24500 17023 24501 17063
rect 24939 17032 24940 17072
rect 24980 17032 24981 17072
rect 24939 17023 24981 17032
rect 25419 17072 25461 17081
rect 25419 17032 25420 17072
rect 25460 17032 25461 17072
rect 25419 17023 25461 17032
rect 25520 17072 25562 17081
rect 25520 17032 25521 17072
rect 25561 17032 25562 17072
rect 25520 17023 25562 17032
rect 27706 17072 27764 17073
rect 27706 17032 27715 17072
rect 27755 17032 27764 17072
rect 27706 17031 27764 17032
rect 15915 17012 15957 17021
rect 18987 17014 19029 17023
rect 24459 17014 24501 17023
rect 7419 16981 7461 16990
rect 8523 16988 8565 16997
rect 7083 16939 7125 16948
rect 8523 16948 8524 16988
rect 8564 16948 8565 16988
rect 8523 16939 8565 16948
rect 9099 16988 9141 16997
rect 9099 16948 9100 16988
rect 9140 16948 9141 16988
rect 9099 16939 9141 16948
rect 10474 16988 10532 16989
rect 11482 16988 11540 16989
rect 10474 16948 10483 16988
rect 10523 16948 10532 16988
rect 10474 16947 10532 16948
rect 11154 16979 11200 16988
rect 11154 16939 11155 16979
rect 11195 16939 11200 16979
rect 11482 16948 11491 16988
rect 11531 16948 11540 16988
rect 11482 16947 11540 16948
rect 13419 16988 13461 16997
rect 13419 16948 13420 16988
rect 13460 16948 13461 16988
rect 13419 16939 13461 16948
rect 15051 16988 15093 16997
rect 15051 16948 15052 16988
rect 15092 16948 15093 16988
rect 15051 16939 15093 16948
rect 16234 16988 16292 16989
rect 16234 16948 16243 16988
rect 16283 16948 16292 16988
rect 16234 16947 16292 16948
rect 19563 16988 19605 16997
rect 19563 16948 19564 16988
rect 19604 16948 19605 16988
rect 19563 16939 19605 16948
rect 25035 16988 25077 16997
rect 25035 16948 25036 16988
rect 25076 16948 25077 16988
rect 25035 16939 25077 16948
rect 11154 16930 11200 16939
rect 8619 16904 8661 16913
rect 5931 16862 5973 16871
rect 922 16820 980 16821
rect 922 16780 931 16820
rect 971 16780 980 16820
rect 922 16779 980 16780
rect 3771 16820 3813 16829
rect 3771 16780 3772 16820
rect 3812 16780 3813 16820
rect 5931 16822 5932 16862
rect 5972 16822 5973 16862
rect 8619 16864 8620 16904
rect 8660 16864 8661 16904
rect 8619 16855 8661 16864
rect 9195 16904 9237 16913
rect 9195 16864 9196 16904
rect 9236 16864 9237 16904
rect 9195 16855 9237 16864
rect 9867 16904 9909 16913
rect 9867 16864 9868 16904
rect 9908 16864 9909 16904
rect 9867 16855 9909 16864
rect 14955 16904 14997 16913
rect 14955 16864 14956 16904
rect 14996 16864 14997 16904
rect 14955 16855 14997 16864
rect 16587 16904 16629 16913
rect 16587 16864 16588 16904
rect 16628 16864 16629 16904
rect 16587 16855 16629 16864
rect 21291 16904 21333 16913
rect 21291 16864 21292 16904
rect 21332 16864 21333 16904
rect 21291 16855 21333 16864
rect 22731 16904 22773 16913
rect 22731 16864 22732 16904
rect 22772 16864 22773 16904
rect 22731 16855 22773 16864
rect 5931 16813 5973 16822
rect 13035 16820 13077 16829
rect 3771 16771 3813 16780
rect 13035 16780 13036 16820
rect 13076 16780 13077 16820
rect 13035 16771 13077 16780
rect 13803 16820 13845 16829
rect 13803 16780 13804 16820
rect 13844 16780 13845 16820
rect 13803 16771 13845 16780
rect 14458 16820 14516 16821
rect 14458 16780 14467 16820
rect 14507 16780 14516 16820
rect 14458 16779 14516 16780
rect 17931 16820 17973 16829
rect 17931 16780 17932 16820
rect 17972 16780 17973 16820
rect 17931 16771 17973 16780
rect 21675 16820 21717 16829
rect 21675 16780 21676 16820
rect 21716 16780 21717 16820
rect 21675 16771 21717 16780
rect 23739 16820 23781 16829
rect 23739 16780 23740 16820
rect 23780 16780 23781 16820
rect 23739 16771 23781 16780
rect 25803 16820 25845 16829
rect 25803 16780 25804 16820
rect 25844 16780 25845 16820
rect 25803 16771 25845 16780
rect 26187 16820 26229 16829
rect 26187 16780 26188 16820
rect 26228 16780 26229 16820
rect 26187 16771 26229 16780
rect 576 16652 31392 16676
rect 576 16612 3112 16652
rect 3480 16612 10886 16652
rect 11254 16612 18660 16652
rect 19028 16612 26434 16652
rect 26802 16612 31392 16652
rect 576 16588 31392 16612
rect 2554 16484 2612 16485
rect 2554 16444 2563 16484
rect 2603 16444 2612 16484
rect 2554 16443 2612 16444
rect 10810 16484 10868 16485
rect 10810 16444 10819 16484
rect 10859 16444 10868 16484
rect 10810 16443 10868 16444
rect 15435 16484 15477 16493
rect 15435 16444 15436 16484
rect 15476 16444 15477 16484
rect 15435 16435 15477 16444
rect 15610 16484 15668 16485
rect 15610 16444 15619 16484
rect 15659 16444 15668 16484
rect 15610 16443 15668 16444
rect 21579 16484 21621 16493
rect 21579 16444 21580 16484
rect 21620 16444 21621 16484
rect 21579 16435 21621 16444
rect 22443 16484 22485 16493
rect 22443 16444 22444 16484
rect 22484 16444 22485 16484
rect 22443 16435 22485 16444
rect 23883 16484 23925 16493
rect 23883 16444 23884 16484
rect 23924 16444 23925 16484
rect 23883 16435 23925 16444
rect 5643 16400 5685 16409
rect 5643 16360 5644 16400
rect 5684 16360 5685 16400
rect 5643 16351 5685 16360
rect 6795 16400 6837 16409
rect 6795 16360 6796 16400
rect 6836 16360 6837 16400
rect 6795 16351 6837 16360
rect 8134 16400 8176 16409
rect 8134 16360 8135 16400
rect 8175 16360 8176 16400
rect 8134 16351 8176 16360
rect 8794 16400 8852 16401
rect 11211 16400 11253 16409
rect 8794 16360 8803 16400
rect 8843 16360 8852 16400
rect 8794 16359 8852 16360
rect 10603 16391 10645 16400
rect 10603 16351 10604 16391
rect 10644 16351 10645 16391
rect 11211 16360 11212 16400
rect 11252 16360 11253 16400
rect 11211 16351 11253 16360
rect 13035 16400 13077 16409
rect 13035 16360 13036 16400
rect 13076 16360 13077 16400
rect 13035 16351 13077 16360
rect 17355 16400 17397 16409
rect 17355 16360 17356 16400
rect 17396 16360 17397 16400
rect 17355 16351 17397 16360
rect 20427 16400 20469 16409
rect 20427 16360 20428 16400
rect 20468 16360 20469 16400
rect 20427 16351 20469 16360
rect 21754 16400 21812 16401
rect 21754 16360 21763 16400
rect 21803 16360 21812 16400
rect 21754 16359 21812 16360
rect 24267 16400 24309 16409
rect 24267 16360 24268 16400
rect 24308 16360 24309 16400
rect 24267 16351 24309 16360
rect 29067 16400 29109 16409
rect 29067 16360 29068 16400
rect 29108 16360 29109 16400
rect 29067 16351 29109 16360
rect 10603 16342 10645 16351
rect 1131 16316 1173 16325
rect 795 16274 837 16283
rect 795 16234 796 16274
rect 836 16234 837 16274
rect 1131 16276 1132 16316
rect 1172 16276 1173 16316
rect 1131 16267 1173 16276
rect 1306 16316 1364 16317
rect 1306 16276 1315 16316
rect 1355 16276 1364 16316
rect 1306 16275 1364 16276
rect 1882 16316 1940 16317
rect 1882 16276 1891 16316
rect 1931 16276 1940 16316
rect 1882 16275 1940 16276
rect 3610 16316 3668 16317
rect 3610 16276 3619 16316
rect 3659 16276 3668 16316
rect 3610 16275 3668 16276
rect 3819 16316 3861 16325
rect 3819 16276 3820 16316
rect 3860 16276 3861 16316
rect 3819 16267 3861 16276
rect 4706 16316 4748 16325
rect 4706 16276 4707 16316
rect 4747 16276 4748 16316
rect 4706 16267 4748 16276
rect 4971 16316 5013 16325
rect 4971 16276 4972 16316
rect 5012 16276 5013 16316
rect 4971 16267 5013 16276
rect 5186 16316 5228 16325
rect 5186 16276 5187 16316
rect 5227 16276 5228 16316
rect 5186 16267 5228 16276
rect 5739 16316 5781 16325
rect 5739 16276 5740 16316
rect 5780 16276 5781 16316
rect 5739 16267 5781 16276
rect 6338 16316 6380 16325
rect 6338 16276 6339 16316
rect 6379 16276 6380 16316
rect 6338 16267 6380 16276
rect 6891 16316 6933 16325
rect 6891 16276 6892 16316
rect 6932 16276 6933 16316
rect 6891 16267 6933 16276
rect 8235 16316 8277 16325
rect 8235 16276 8236 16316
rect 8276 16276 8277 16316
rect 7018 16274 7076 16275
rect 795 16225 837 16234
rect 922 16232 980 16233
rect 922 16192 931 16232
rect 971 16192 980 16232
rect 922 16191 980 16192
rect 1035 16232 1077 16241
rect 1035 16192 1036 16232
rect 1076 16192 1077 16232
rect 1035 16183 1077 16192
rect 1690 16232 1748 16233
rect 1690 16192 1699 16232
rect 1739 16192 1748 16232
rect 1690 16191 1748 16192
rect 2080 16232 2122 16241
rect 2080 16192 2081 16232
rect 2121 16192 2122 16232
rect 2080 16183 2122 16192
rect 2369 16232 2427 16233
rect 2369 16192 2378 16232
rect 2418 16192 2427 16232
rect 2369 16191 2427 16192
rect 2851 16232 2909 16233
rect 2851 16192 2860 16232
rect 2900 16192 2909 16232
rect 2851 16191 2909 16192
rect 3343 16232 3401 16233
rect 3343 16192 3352 16232
rect 3392 16192 3401 16232
rect 3343 16191 3401 16192
rect 3483 16232 3525 16241
rect 3483 16192 3484 16232
rect 3524 16192 3525 16232
rect 3483 16183 3525 16192
rect 3723 16232 3765 16241
rect 3723 16192 3724 16232
rect 3764 16192 3765 16232
rect 3723 16183 3765 16192
rect 4107 16232 4149 16241
rect 4107 16192 4108 16232
rect 4148 16192 4149 16232
rect 4107 16183 4149 16192
rect 4226 16232 4268 16241
rect 4226 16192 4227 16232
rect 4267 16192 4268 16232
rect 4226 16183 4268 16192
rect 4336 16232 4394 16233
rect 4336 16192 4345 16232
rect 4385 16192 4394 16232
rect 4336 16191 4394 16192
rect 4587 16232 4629 16241
rect 4587 16192 4588 16232
rect 4628 16192 4629 16232
rect 4587 16183 4629 16192
rect 4816 16232 4874 16233
rect 4816 16192 4825 16232
rect 4865 16192 4874 16232
rect 4816 16191 4874 16192
rect 5076 16232 5118 16241
rect 5076 16192 5077 16232
rect 5117 16192 5118 16232
rect 5076 16183 5118 16192
rect 5298 16232 5340 16241
rect 5298 16192 5299 16232
rect 5339 16192 5340 16232
rect 5298 16183 5340 16192
rect 5582 16232 5624 16241
rect 5582 16192 5583 16232
rect 5623 16192 5624 16232
rect 5582 16183 5624 16192
rect 5866 16232 5924 16233
rect 5866 16192 5875 16232
rect 5915 16192 5924 16232
rect 5866 16191 5924 16192
rect 6219 16232 6261 16241
rect 6219 16192 6220 16232
rect 6260 16192 6261 16232
rect 6219 16183 6261 16192
rect 6448 16232 6506 16233
rect 6448 16192 6457 16232
rect 6497 16192 6506 16232
rect 6448 16191 6506 16192
rect 6734 16232 6776 16241
rect 7018 16234 7027 16274
rect 7067 16234 7076 16274
rect 8235 16267 8277 16276
rect 9003 16316 9045 16325
rect 11307 16316 11349 16325
rect 9003 16276 9004 16316
rect 9044 16276 9045 16316
rect 9003 16267 9045 16276
rect 10290 16307 10336 16316
rect 10290 16267 10291 16307
rect 10331 16267 10336 16307
rect 11307 16276 11308 16316
rect 11348 16276 11349 16316
rect 11307 16267 11349 16276
rect 11883 16316 11925 16325
rect 12939 16316 12981 16325
rect 11883 16276 11884 16316
rect 11924 16276 11925 16316
rect 11434 16274 11492 16275
rect 10290 16258 10336 16267
rect 7018 16233 7076 16234
rect 6734 16192 6735 16232
rect 6775 16192 6776 16232
rect 6734 16183 6776 16192
rect 7195 16232 7253 16233
rect 7195 16192 7204 16232
rect 7244 16192 7253 16232
rect 7195 16191 7253 16192
rect 7354 16232 7412 16233
rect 7354 16192 7363 16232
rect 7403 16192 7412 16232
rect 7354 16191 7412 16192
rect 7479 16232 7521 16241
rect 7479 16192 7480 16232
rect 7520 16192 7521 16232
rect 7479 16183 7521 16192
rect 7603 16232 7661 16233
rect 7603 16192 7612 16232
rect 7652 16192 7661 16232
rect 7603 16191 7661 16192
rect 7745 16232 7803 16233
rect 7745 16192 7754 16232
rect 7794 16192 7803 16232
rect 7745 16191 7803 16192
rect 7908 16232 7966 16233
rect 7908 16192 7917 16232
rect 7957 16192 7966 16232
rect 7908 16191 7966 16192
rect 8078 16232 8120 16241
rect 8078 16192 8079 16232
rect 8119 16192 8120 16232
rect 8078 16183 8120 16192
rect 8362 16232 8420 16233
rect 8362 16192 8371 16232
rect 8411 16192 8420 16232
rect 8362 16191 8420 16192
rect 8619 16232 8661 16241
rect 8619 16192 8620 16232
rect 8660 16192 8661 16232
rect 8619 16183 8661 16192
rect 8794 16232 8852 16233
rect 8794 16192 8803 16232
rect 8843 16192 8852 16232
rect 8794 16191 8852 16192
rect 9322 16232 9380 16233
rect 9322 16192 9331 16232
rect 9371 16192 9380 16232
rect 9322 16191 9380 16192
rect 10155 16232 10197 16241
rect 10155 16192 10156 16232
rect 10196 16192 10197 16232
rect 10155 16183 10197 16192
rect 10384 16232 10442 16233
rect 10384 16192 10393 16232
rect 10433 16192 10442 16232
rect 10384 16191 10442 16192
rect 10618 16232 10676 16233
rect 10618 16192 10627 16232
rect 10667 16192 10676 16232
rect 10618 16191 10676 16192
rect 10971 16232 11013 16241
rect 10971 16192 10972 16232
rect 11012 16192 11013 16232
rect 10971 16183 11013 16192
rect 11150 16232 11192 16241
rect 11434 16234 11443 16274
rect 11483 16234 11492 16274
rect 11883 16267 11925 16276
rect 12594 16307 12640 16316
rect 12594 16267 12595 16307
rect 12635 16267 12640 16307
rect 12939 16276 12940 16316
rect 12980 16276 12981 16316
rect 12939 16267 12981 16276
rect 17259 16316 17301 16325
rect 17259 16276 17260 16316
rect 17300 16276 17301 16316
rect 13114 16274 13172 16275
rect 12594 16258 12640 16267
rect 11434 16233 11492 16234
rect 11150 16192 11151 16232
rect 11191 16192 11192 16232
rect 11150 16183 11192 16192
rect 11547 16232 11589 16241
rect 11547 16192 11548 16232
rect 11588 16192 11589 16232
rect 11547 16183 11589 16192
rect 11726 16232 11768 16241
rect 11726 16192 11727 16232
rect 11767 16192 11768 16232
rect 11726 16183 11768 16192
rect 12004 16232 12046 16241
rect 12004 16192 12005 16232
rect 12045 16192 12046 16232
rect 12004 16183 12046 16192
rect 12459 16232 12501 16241
rect 12459 16192 12460 16232
rect 12500 16192 12501 16232
rect 12459 16183 12501 16192
rect 12699 16232 12741 16241
rect 13114 16234 13123 16274
rect 13163 16234 13172 16274
rect 17259 16267 17301 16276
rect 17818 16316 17876 16317
rect 17818 16276 17827 16316
rect 17867 16276 17876 16316
rect 17818 16275 17876 16276
rect 18027 16316 18069 16325
rect 18027 16276 18028 16316
rect 18068 16276 18069 16316
rect 18027 16267 18069 16276
rect 19371 16316 19413 16325
rect 19371 16276 19372 16316
rect 19412 16276 19413 16316
rect 19018 16274 19076 16275
rect 13899 16243 13941 16252
rect 13114 16233 13172 16234
rect 12699 16192 12700 16232
rect 12740 16192 12741 16232
rect 12699 16183 12741 16192
rect 12802 16232 12860 16233
rect 12802 16192 12811 16232
rect 12851 16192 12860 16232
rect 12802 16191 12860 16192
rect 13268 16232 13310 16241
rect 13268 16192 13269 16232
rect 13309 16192 13310 16232
rect 13606 16232 13664 16233
rect 13268 16183 13310 16192
rect 13402 16205 13460 16206
rect 13402 16165 13411 16205
rect 13451 16165 13460 16205
rect 13606 16192 13615 16232
rect 13655 16192 13664 16232
rect 13606 16191 13664 16192
rect 13786 16232 13844 16233
rect 13786 16192 13795 16232
rect 13835 16192 13844 16232
rect 13899 16203 13900 16243
rect 13940 16203 13941 16243
rect 15291 16243 15333 16252
rect 13899 16194 13941 16203
rect 14036 16232 14094 16233
rect 13786 16191 13844 16192
rect 14036 16192 14045 16232
rect 14085 16192 14094 16232
rect 14036 16191 14094 16192
rect 14170 16232 14228 16233
rect 14170 16192 14179 16232
rect 14219 16192 14228 16232
rect 14170 16191 14228 16192
rect 14347 16232 14405 16233
rect 14347 16192 14356 16232
rect 14396 16192 14405 16232
rect 14347 16191 14405 16192
rect 14875 16232 14933 16233
rect 14875 16192 14884 16232
rect 14924 16192 14933 16232
rect 14875 16191 14933 16192
rect 15034 16232 15092 16233
rect 15034 16192 15043 16232
rect 15083 16192 15092 16232
rect 15034 16191 15092 16192
rect 15159 16232 15201 16241
rect 15159 16192 15160 16232
rect 15200 16192 15201 16232
rect 15291 16203 15292 16243
rect 15332 16203 15333 16243
rect 15291 16194 15333 16203
rect 15418 16232 15476 16233
rect 15159 16183 15201 16192
rect 15418 16192 15427 16232
rect 15467 16192 15476 16232
rect 15418 16191 15476 16192
rect 15622 16232 15680 16233
rect 15622 16192 15631 16232
rect 15671 16192 15680 16232
rect 15622 16191 15680 16192
rect 15728 16232 15786 16233
rect 15728 16192 15737 16232
rect 15777 16192 15786 16232
rect 15728 16191 15786 16192
rect 15894 16232 15952 16233
rect 15894 16192 15903 16232
rect 15943 16192 15952 16232
rect 15894 16191 15952 16192
rect 16002 16232 16060 16233
rect 16002 16192 16011 16232
rect 16051 16192 16060 16232
rect 16002 16191 16060 16192
rect 16128 16232 16186 16233
rect 16128 16192 16137 16232
rect 16177 16192 16186 16232
rect 16128 16191 16186 16192
rect 16378 16232 16436 16233
rect 16378 16192 16387 16232
rect 16427 16192 16436 16232
rect 16378 16191 16436 16192
rect 16496 16232 16554 16233
rect 16496 16192 16505 16232
rect 16545 16192 16554 16232
rect 16496 16191 16554 16192
rect 16664 16232 16706 16241
rect 16664 16192 16665 16232
rect 16705 16192 16706 16232
rect 16664 16183 16706 16192
rect 16762 16232 16820 16233
rect 16762 16192 16771 16232
rect 16811 16192 16820 16232
rect 16762 16191 16820 16192
rect 16896 16232 16954 16233
rect 16896 16192 16905 16232
rect 16945 16192 16954 16232
rect 16896 16191 16954 16192
rect 17115 16232 17157 16241
rect 17115 16192 17116 16232
rect 17156 16192 17157 16232
rect 17115 16183 17157 16192
rect 17430 16232 17472 16241
rect 17430 16192 17431 16232
rect 17471 16192 17472 16232
rect 17430 16183 17472 16192
rect 17578 16232 17636 16233
rect 17578 16192 17587 16232
rect 17627 16192 17636 16232
rect 17578 16191 17636 16192
rect 17691 16232 17733 16241
rect 17691 16192 17692 16232
rect 17732 16192 17733 16232
rect 17691 16183 17733 16192
rect 17931 16232 17973 16241
rect 19018 16234 19027 16274
rect 19067 16234 19076 16274
rect 19371 16267 19413 16276
rect 26859 16316 26901 16325
rect 26859 16276 26860 16316
rect 26900 16276 26901 16316
rect 26859 16267 26901 16276
rect 28683 16274 28725 16283
rect 19018 16233 19076 16234
rect 17931 16192 17932 16232
rect 17972 16192 17973 16232
rect 17931 16183 17973 16192
rect 18511 16232 18569 16233
rect 18511 16192 18520 16232
rect 18560 16192 18569 16232
rect 18511 16191 18569 16192
rect 19563 16232 19605 16241
rect 20139 16232 20181 16241
rect 19563 16192 19564 16232
rect 19604 16192 19605 16232
rect 19563 16183 19605 16192
rect 19842 16223 19888 16232
rect 19842 16183 19843 16223
rect 19883 16183 19888 16223
rect 20139 16192 20140 16232
rect 20180 16192 20181 16232
rect 20139 16183 20181 16192
rect 20907 16232 20949 16241
rect 20907 16192 20908 16232
rect 20948 16192 20949 16232
rect 20907 16183 20949 16192
rect 21178 16232 21236 16233
rect 21178 16192 21187 16232
rect 21227 16192 21236 16232
rect 21178 16191 21236 16192
rect 21963 16232 22005 16241
rect 21963 16192 21964 16232
rect 22004 16192 22005 16232
rect 21963 16183 22005 16192
rect 22084 16232 22126 16241
rect 22084 16192 22085 16232
rect 22125 16192 22126 16232
rect 22084 16183 22126 16192
rect 22486 16232 22528 16241
rect 22731 16232 22773 16241
rect 22486 16192 22487 16232
rect 22527 16192 22528 16232
rect 22486 16183 22528 16192
rect 22626 16223 22672 16232
rect 22626 16183 22627 16223
rect 22667 16183 22672 16223
rect 22731 16192 22732 16232
rect 22772 16192 22773 16232
rect 22731 16183 22773 16192
rect 23211 16232 23253 16241
rect 23211 16192 23212 16232
rect 23252 16192 23253 16232
rect 23211 16183 23253 16192
rect 23482 16232 23540 16233
rect 23482 16192 23491 16232
rect 23531 16192 23540 16232
rect 23482 16191 23540 16192
rect 24118 16232 24160 16241
rect 24363 16232 24405 16241
rect 24118 16192 24119 16232
rect 24159 16192 24160 16232
rect 24118 16183 24160 16192
rect 24258 16223 24304 16232
rect 24258 16183 24259 16223
rect 24299 16183 24304 16223
rect 24363 16192 24364 16232
rect 24404 16192 24405 16232
rect 24363 16183 24405 16192
rect 24555 16232 24597 16241
rect 24555 16192 24556 16232
rect 24596 16192 24597 16232
rect 24555 16183 24597 16192
rect 26091 16232 26133 16241
rect 26091 16192 26092 16232
rect 26132 16192 26133 16232
rect 26091 16183 26133 16192
rect 26362 16232 26420 16233
rect 26362 16192 26371 16232
rect 26411 16192 26420 16232
rect 26362 16191 26420 16192
rect 26475 16232 26517 16241
rect 26475 16192 26476 16232
rect 26516 16192 26517 16232
rect 26475 16183 26517 16192
rect 26955 16232 26997 16241
rect 26955 16192 26956 16232
rect 26996 16192 26997 16232
rect 26955 16183 26997 16192
rect 27427 16232 27485 16233
rect 27427 16192 27436 16232
rect 27476 16192 27485 16232
rect 27427 16191 27485 16192
rect 27946 16232 28004 16233
rect 27946 16192 27955 16232
rect 27995 16192 28004 16232
rect 27946 16191 28004 16192
rect 28299 16232 28341 16241
rect 28299 16192 28300 16232
rect 28340 16192 28341 16232
rect 28299 16183 28341 16192
rect 28491 16232 28533 16241
rect 28491 16192 28492 16232
rect 28532 16192 28533 16232
rect 28683 16234 28684 16274
rect 28724 16234 28725 16274
rect 28683 16225 28725 16234
rect 28875 16232 28917 16241
rect 28491 16183 28533 16192
rect 28875 16192 28876 16232
rect 28916 16192 28917 16232
rect 28875 16183 28917 16192
rect 19842 16174 19888 16183
rect 22626 16174 22672 16183
rect 24258 16174 24304 16183
rect 13402 16164 13460 16165
rect 2560 16148 2602 16157
rect 2560 16108 2561 16148
rect 2601 16108 2602 16148
rect 2560 16099 2602 16108
rect 4491 16148 4533 16157
rect 4491 16108 4492 16148
rect 4532 16108 4533 16148
rect 4491 16099 4533 16108
rect 6123 16148 6165 16157
rect 6123 16108 6124 16148
rect 6164 16108 6165 16148
rect 6123 16099 6165 16108
rect 9531 16148 9573 16157
rect 9531 16108 9532 16148
rect 9572 16108 9573 16148
rect 19131 16148 19173 16157
rect 9531 16099 9573 16108
rect 11799 16106 11841 16115
rect 1402 16064 1460 16065
rect 1402 16024 1411 16064
rect 1451 16024 1460 16064
rect 1402 16023 1460 16024
rect 2170 16064 2228 16065
rect 2170 16024 2179 16064
rect 2219 16024 2228 16064
rect 2170 16023 2228 16024
rect 2283 16064 2325 16073
rect 2283 16024 2284 16064
rect 2324 16024 2325 16064
rect 2283 16015 2325 16024
rect 2763 16064 2805 16073
rect 2763 16024 2764 16064
rect 2804 16024 2805 16064
rect 2763 16015 2805 16024
rect 3178 16064 3236 16065
rect 3178 16024 3187 16064
rect 3227 16024 3236 16064
rect 3178 16023 3236 16024
rect 4011 16064 4053 16073
rect 4011 16024 4012 16064
rect 4052 16024 4053 16064
rect 4011 16015 4053 16024
rect 7258 16064 7316 16065
rect 7258 16024 7267 16064
rect 7307 16024 7316 16064
rect 7258 16023 7316 16024
rect 9243 16064 9285 16073
rect 9243 16024 9244 16064
rect 9284 16024 9285 16064
rect 5530 16022 5588 16023
rect 5530 15982 5539 16022
rect 5579 15982 5588 16022
rect 5530 15981 5588 15982
rect 6682 16022 6740 16023
rect 6682 15982 6691 16022
rect 6731 15982 6740 16022
rect 9243 16015 9285 16024
rect 10059 16064 10101 16073
rect 10059 16024 10060 16064
rect 10100 16024 10101 16064
rect 11799 16066 11800 16106
rect 11840 16066 11841 16106
rect 19131 16108 19132 16148
rect 19172 16108 19173 16148
rect 19131 16099 19173 16108
rect 19947 16148 19989 16157
rect 19947 16108 19948 16148
rect 19988 16108 19989 16148
rect 19947 16099 19989 16108
rect 21291 16148 21333 16157
rect 21291 16108 21292 16148
rect 21332 16108 21333 16148
rect 21291 16099 21333 16108
rect 23595 16148 23637 16157
rect 23595 16108 23596 16148
rect 23636 16108 23637 16148
rect 23595 16099 23637 16108
rect 25227 16148 25269 16157
rect 25227 16108 25228 16148
rect 25268 16108 25269 16148
rect 25227 16099 25269 16108
rect 11799 16057 11841 16066
rect 12363 16064 12405 16073
rect 10059 16015 10101 16024
rect 12363 16024 12364 16064
rect 12404 16024 12405 16064
rect 12363 16015 12405 16024
rect 13594 16064 13652 16065
rect 13594 16024 13603 16064
rect 13643 16024 13652 16064
rect 13594 16023 13652 16024
rect 14266 16064 14324 16065
rect 14266 16024 14275 16064
rect 14315 16024 14324 16064
rect 14266 16023 14324 16024
rect 16858 16064 16916 16065
rect 16858 16024 16867 16064
rect 16907 16024 16916 16064
rect 16858 16023 16916 16024
rect 18346 16064 18404 16065
rect 18346 16024 18355 16064
rect 18395 16024 18404 16064
rect 18346 16023 18404 16024
rect 18826 16064 18884 16065
rect 18826 16024 18835 16064
rect 18875 16024 18884 16064
rect 18826 16023 18884 16024
rect 19707 16064 19749 16073
rect 19707 16024 19708 16064
rect 19748 16024 19749 16064
rect 19707 16015 19749 16024
rect 22059 16064 22101 16073
rect 22059 16024 22060 16064
rect 22100 16024 22101 16064
rect 22059 16015 22101 16024
rect 25419 16064 25461 16073
rect 25419 16024 25420 16064
rect 25460 16024 25461 16064
rect 25419 16015 25461 16024
rect 28107 16064 28149 16073
rect 28107 16024 28108 16064
rect 28148 16024 28149 16064
rect 28107 16015 28149 16024
rect 28395 16064 28437 16073
rect 28395 16024 28396 16064
rect 28436 16024 28437 16064
rect 28395 16015 28437 16024
rect 28779 16064 28821 16073
rect 28779 16024 28780 16064
rect 28820 16024 28821 16064
rect 28779 16015 28821 16024
rect 6682 15981 6740 15982
rect 576 15896 31392 15920
rect 576 15856 4352 15896
rect 4720 15856 12126 15896
rect 12494 15856 19900 15896
rect 20268 15856 27674 15896
rect 28042 15856 31392 15896
rect 576 15832 31392 15856
rect 1498 15728 1556 15729
rect 1498 15688 1507 15728
rect 1547 15688 1556 15728
rect 1498 15687 1556 15688
rect 1611 15728 1653 15737
rect 1611 15688 1612 15728
rect 1652 15688 1653 15728
rect 1611 15679 1653 15688
rect 1978 15728 2036 15729
rect 1978 15688 1987 15728
rect 2027 15688 2036 15728
rect 1978 15687 2036 15688
rect 2955 15728 2997 15737
rect 2955 15688 2956 15728
rect 2996 15688 2997 15728
rect 2955 15679 2997 15688
rect 3435 15728 3477 15737
rect 3435 15688 3436 15728
rect 3476 15688 3477 15728
rect 3435 15679 3477 15688
rect 3994 15728 4052 15729
rect 3994 15688 4003 15728
rect 4043 15688 4052 15728
rect 3994 15687 4052 15688
rect 4474 15728 4532 15729
rect 4474 15688 4483 15728
rect 4523 15688 4532 15728
rect 4474 15687 4532 15688
rect 4875 15728 4917 15737
rect 4875 15688 4876 15728
rect 4916 15688 4917 15728
rect 4875 15679 4917 15688
rect 5739 15728 5781 15737
rect 5739 15688 5740 15728
rect 5780 15688 5781 15728
rect 5739 15679 5781 15688
rect 6298 15728 6356 15729
rect 6298 15688 6307 15728
rect 6347 15688 6356 15728
rect 6298 15687 6356 15688
rect 7755 15728 7797 15737
rect 7755 15688 7756 15728
rect 7796 15688 7797 15728
rect 7755 15679 7797 15688
rect 8139 15728 8181 15737
rect 8139 15688 8140 15728
rect 8180 15688 8181 15728
rect 8139 15679 8181 15688
rect 10731 15728 10773 15737
rect 10731 15688 10732 15728
rect 10772 15688 10773 15728
rect 10731 15679 10773 15688
rect 12027 15728 12069 15737
rect 12027 15688 12028 15728
rect 12068 15688 12069 15728
rect 12027 15679 12069 15688
rect 13803 15728 13845 15737
rect 13803 15688 13804 15728
rect 13844 15688 13845 15728
rect 13803 15679 13845 15688
rect 14859 15728 14901 15737
rect 14859 15688 14860 15728
rect 14900 15688 14901 15728
rect 14859 15679 14901 15688
rect 16011 15728 16053 15737
rect 16011 15688 16012 15728
rect 16052 15688 16053 15728
rect 16011 15679 16053 15688
rect 16858 15728 16916 15729
rect 16858 15688 16867 15728
rect 16907 15688 16916 15728
rect 16858 15687 16916 15688
rect 17818 15728 17876 15729
rect 17818 15688 17827 15728
rect 17867 15688 17876 15728
rect 17818 15687 17876 15688
rect 17931 15728 17973 15737
rect 17931 15688 17932 15728
rect 17972 15688 17973 15728
rect 17931 15679 17973 15688
rect 21771 15728 21813 15737
rect 21771 15688 21772 15728
rect 21812 15688 21813 15728
rect 21771 15679 21813 15688
rect 22330 15728 22388 15729
rect 22330 15688 22339 15728
rect 22379 15688 22388 15728
rect 22330 15687 22388 15688
rect 23787 15728 23829 15737
rect 23787 15688 23788 15728
rect 23828 15688 23829 15728
rect 23787 15679 23829 15688
rect 24939 15728 24981 15737
rect 24939 15688 24940 15728
rect 24980 15688 24981 15728
rect 24939 15679 24981 15688
rect 25210 15728 25268 15729
rect 25210 15688 25219 15728
rect 25259 15688 25268 15728
rect 25210 15687 25268 15688
rect 25899 15728 25941 15737
rect 25899 15688 25900 15728
rect 25940 15688 25941 15728
rect 25899 15679 25941 15688
rect 28971 15728 29013 15737
rect 28971 15688 28972 15728
rect 29012 15688 29013 15728
rect 28971 15679 29013 15688
rect 3232 15644 3274 15653
rect 3232 15604 3233 15644
rect 3273 15604 3274 15644
rect 3232 15595 3274 15604
rect 3706 15644 3764 15645
rect 3706 15604 3715 15644
rect 3755 15604 3764 15644
rect 3706 15603 3764 15604
rect 7179 15644 7221 15653
rect 7179 15604 7180 15644
rect 7220 15604 7221 15644
rect 7179 15595 7221 15604
rect 8986 15644 9044 15645
rect 12352 15644 12394 15653
rect 8986 15604 8995 15644
rect 9035 15604 9044 15644
rect 8986 15603 9044 15604
rect 10818 15635 10864 15644
rect 10818 15595 10819 15635
rect 10859 15595 10864 15635
rect 12352 15604 12353 15644
rect 12393 15604 12394 15644
rect 12352 15595 12394 15604
rect 15627 15644 15669 15653
rect 15627 15604 15628 15644
rect 15668 15604 15669 15644
rect 13210 15602 13268 15603
rect 10818 15586 10864 15595
rect 922 15560 980 15561
rect 922 15520 931 15560
rect 971 15520 980 15560
rect 922 15519 980 15520
rect 1227 15560 1269 15569
rect 1227 15520 1228 15560
rect 1268 15520 1269 15560
rect 1227 15511 1269 15520
rect 1408 15560 1450 15569
rect 1899 15560 1941 15569
rect 1408 15520 1409 15560
rect 1449 15520 1450 15560
rect 1408 15511 1450 15520
rect 1707 15551 1749 15560
rect 1707 15511 1708 15551
rect 1748 15511 1749 15551
rect 1899 15520 1900 15560
rect 1940 15520 1941 15560
rect 1899 15511 1941 15520
rect 2187 15560 2229 15569
rect 2187 15520 2188 15560
rect 2228 15520 2229 15560
rect 2187 15511 2229 15520
rect 2326 15560 2368 15569
rect 2326 15520 2327 15560
rect 2367 15520 2368 15560
rect 2326 15511 2368 15520
rect 2458 15560 2516 15561
rect 2458 15520 2467 15560
rect 2507 15520 2516 15560
rect 2458 15519 2516 15520
rect 2571 15560 2613 15569
rect 2571 15520 2572 15560
rect 2612 15520 2613 15560
rect 2571 15511 2613 15520
rect 2859 15560 2901 15569
rect 2859 15520 2860 15560
rect 2900 15520 2901 15560
rect 2859 15511 2901 15520
rect 3051 15560 3093 15569
rect 3915 15560 3957 15569
rect 3051 15520 3052 15560
rect 3092 15520 3093 15560
rect 3051 15511 3093 15520
rect 3531 15551 3573 15560
rect 3531 15511 3532 15551
rect 3572 15511 3573 15551
rect 3915 15520 3916 15560
rect 3956 15520 3957 15560
rect 3915 15511 3957 15520
rect 4150 15560 4192 15569
rect 4150 15520 4151 15560
rect 4191 15520 4192 15560
rect 4150 15511 4192 15520
rect 4395 15560 4437 15569
rect 4395 15520 4396 15560
rect 4436 15520 4437 15560
rect 4395 15511 4437 15520
rect 4971 15560 5013 15569
rect 4971 15520 4972 15560
rect 5012 15520 5013 15560
rect 4971 15511 5013 15520
rect 5202 15560 5244 15569
rect 5202 15520 5203 15560
rect 5243 15520 5244 15560
rect 5202 15511 5244 15520
rect 5355 15560 5397 15569
rect 5355 15520 5356 15560
rect 5396 15520 5397 15560
rect 5355 15511 5397 15520
rect 5547 15560 5589 15569
rect 5547 15520 5548 15560
rect 5588 15520 5589 15560
rect 5547 15511 5589 15520
rect 5835 15560 5877 15569
rect 5835 15520 5836 15560
rect 5876 15520 5877 15560
rect 5835 15511 5877 15520
rect 6066 15560 6108 15569
rect 6066 15520 6067 15560
rect 6107 15520 6108 15560
rect 6066 15511 6108 15520
rect 6202 15560 6260 15561
rect 6202 15520 6211 15560
rect 6251 15520 6260 15560
rect 6202 15519 6260 15520
rect 6518 15560 6560 15569
rect 6518 15520 6519 15560
rect 6559 15520 6560 15560
rect 6518 15511 6560 15520
rect 6795 15560 6837 15569
rect 6795 15520 6796 15560
rect 6836 15520 6837 15560
rect 6795 15511 6837 15520
rect 6970 15560 7028 15561
rect 6970 15520 6979 15560
rect 7019 15520 7028 15560
rect 6970 15519 7028 15520
rect 7275 15560 7317 15569
rect 7275 15520 7276 15560
rect 7316 15520 7317 15560
rect 7275 15511 7317 15520
rect 7492 15560 7534 15569
rect 7492 15520 7493 15560
rect 7533 15520 7534 15560
rect 7492 15511 7534 15520
rect 7659 15560 7701 15569
rect 7659 15520 7660 15560
rect 7700 15520 7701 15560
rect 7659 15511 7701 15520
rect 7834 15560 7892 15561
rect 7834 15520 7843 15560
rect 7883 15520 7892 15560
rect 7834 15519 7892 15520
rect 8043 15560 8085 15569
rect 8043 15520 8044 15560
rect 8084 15520 8085 15560
rect 8427 15560 8469 15569
rect 8043 15511 8085 15520
rect 8235 15518 8277 15527
rect 1707 15502 1749 15511
rect 3531 15502 3573 15511
rect 2667 15476 2709 15485
rect 2667 15436 2668 15476
rect 2708 15436 2709 15476
rect 2667 15427 2709 15436
rect 4282 15476 4340 15477
rect 4282 15436 4291 15476
rect 4331 15436 4340 15476
rect 4282 15435 4340 15436
rect 5090 15476 5132 15485
rect 5090 15436 5091 15476
rect 5131 15436 5132 15476
rect 5090 15427 5132 15436
rect 5954 15476 5996 15485
rect 5954 15436 5955 15476
rect 5995 15436 5996 15476
rect 5954 15427 5996 15436
rect 7394 15476 7436 15485
rect 7394 15436 7395 15476
rect 7435 15436 7436 15476
rect 8235 15478 8236 15518
rect 8276 15478 8277 15518
rect 8427 15520 8428 15560
rect 8468 15520 8469 15560
rect 8427 15511 8469 15520
rect 8674 15560 8732 15561
rect 8674 15520 8683 15560
rect 8723 15520 8732 15560
rect 8674 15519 8732 15520
rect 8907 15560 8949 15569
rect 8907 15520 8908 15560
rect 8948 15520 8949 15560
rect 8907 15511 8949 15520
rect 9274 15560 9332 15561
rect 9274 15520 9283 15560
rect 9323 15520 9332 15560
rect 9274 15519 9332 15520
rect 9562 15560 9620 15561
rect 9562 15520 9571 15560
rect 9611 15520 9620 15560
rect 9562 15519 9620 15520
rect 10059 15560 10101 15569
rect 10059 15520 10060 15560
rect 10100 15520 10101 15560
rect 10059 15511 10101 15520
rect 10276 15560 10318 15569
rect 10276 15520 10277 15560
rect 10317 15520 10318 15560
rect 10276 15511 10318 15520
rect 10514 15560 10572 15561
rect 10514 15520 10523 15560
rect 10563 15520 10572 15560
rect 10514 15519 10572 15520
rect 10678 15560 10736 15561
rect 10678 15520 10687 15560
rect 10727 15520 10736 15560
rect 10678 15519 10736 15520
rect 10902 15560 10960 15561
rect 10902 15520 10911 15560
rect 10951 15520 10960 15560
rect 10902 15519 10960 15520
rect 11083 15560 11141 15561
rect 11083 15520 11092 15560
rect 11132 15520 11141 15560
rect 11083 15519 11141 15520
rect 11451 15560 11493 15569
rect 11451 15520 11452 15560
rect 11492 15520 11493 15560
rect 11451 15511 11493 15520
rect 11906 15560 11948 15569
rect 11906 15520 11907 15560
rect 11947 15520 11948 15560
rect 11770 15518 11828 15519
rect 8235 15469 8277 15478
rect 8794 15476 8852 15477
rect 7394 15427 7436 15436
rect 8794 15436 8803 15476
rect 8843 15436 8852 15476
rect 8794 15435 8852 15436
rect 9178 15476 9236 15477
rect 9178 15436 9187 15476
rect 9227 15436 9236 15476
rect 9178 15435 9236 15436
rect 9723 15476 9765 15485
rect 9723 15436 9724 15476
rect 9764 15436 9765 15476
rect 9723 15427 9765 15436
rect 9963 15476 10005 15485
rect 9963 15436 9964 15476
rect 10004 15436 10005 15476
rect 9963 15427 10005 15436
rect 10178 15476 10220 15485
rect 10178 15436 10179 15476
rect 10219 15436 10220 15476
rect 10178 15427 10220 15436
rect 11595 15476 11637 15485
rect 11770 15478 11779 15518
rect 11819 15478 11828 15518
rect 11906 15511 11948 15520
rect 12171 15560 12213 15569
rect 12171 15520 12172 15560
rect 12212 15520 12213 15560
rect 12171 15511 12213 15520
rect 12555 15560 12597 15569
rect 13210 15562 13219 15602
rect 13259 15562 13268 15602
rect 15627 15595 15669 15604
rect 17248 15644 17290 15653
rect 17248 15604 17249 15644
rect 17289 15604 17290 15644
rect 17248 15595 17290 15604
rect 17725 15644 17767 15653
rect 17725 15604 17726 15644
rect 17766 15604 17767 15644
rect 17725 15595 17767 15604
rect 21003 15644 21045 15653
rect 21003 15604 21004 15644
rect 21044 15604 21045 15644
rect 21003 15595 21045 15604
rect 21113 15644 21155 15653
rect 21113 15604 21114 15644
rect 21154 15604 21155 15644
rect 21113 15595 21155 15604
rect 22841 15644 22883 15653
rect 22841 15604 22842 15644
rect 22882 15604 22883 15644
rect 22841 15595 22883 15604
rect 23194 15644 23252 15645
rect 23194 15604 23203 15644
rect 23243 15604 23252 15644
rect 23194 15603 23252 15604
rect 23292 15571 23350 15572
rect 13210 15561 13268 15562
rect 13419 15560 13461 15569
rect 12555 15520 12556 15560
rect 12596 15520 12597 15560
rect 12555 15511 12597 15520
rect 12651 15551 12693 15560
rect 12651 15511 12652 15551
rect 12692 15511 12693 15551
rect 12651 15502 12693 15511
rect 12795 15518 12837 15527
rect 13419 15520 13420 15560
rect 13460 15520 13461 15560
rect 11770 15477 11828 15478
rect 12795 15478 12796 15518
rect 12836 15478 12837 15518
rect 13114 15518 13172 15519
rect 11595 15436 11596 15476
rect 11636 15436 11637 15476
rect 12795 15469 12837 15478
rect 12937 15476 12979 15485
rect 13114 15478 13123 15518
rect 13163 15478 13172 15518
rect 13419 15511 13461 15520
rect 13611 15560 13653 15569
rect 13611 15520 13612 15560
rect 13652 15520 13653 15560
rect 13611 15511 13653 15520
rect 13899 15560 13941 15569
rect 13899 15520 13900 15560
rect 13940 15520 13941 15560
rect 13899 15511 13941 15520
rect 14128 15560 14186 15561
rect 14128 15520 14137 15560
rect 14177 15520 14186 15560
rect 14128 15519 14186 15520
rect 14244 15560 14302 15561
rect 14244 15520 14253 15560
rect 14293 15520 14302 15560
rect 14244 15519 14302 15520
rect 14400 15560 14442 15569
rect 14400 15520 14401 15560
rect 14441 15520 14442 15560
rect 14400 15511 14442 15520
rect 14692 15560 14734 15569
rect 14692 15520 14693 15560
rect 14733 15520 14734 15560
rect 14692 15511 14734 15520
rect 15034 15560 15092 15561
rect 15034 15520 15043 15560
rect 15083 15520 15092 15560
rect 15034 15519 15092 15520
rect 15531 15560 15573 15569
rect 15531 15520 15532 15560
rect 15572 15520 15573 15560
rect 15531 15511 15573 15520
rect 15723 15560 15765 15569
rect 15723 15520 15724 15560
rect 15764 15520 15765 15560
rect 15723 15511 15765 15520
rect 15915 15560 15957 15569
rect 15915 15520 15916 15560
rect 15956 15520 15957 15560
rect 15915 15511 15957 15520
rect 16107 15560 16149 15569
rect 16107 15520 16108 15560
rect 16148 15520 16149 15560
rect 16107 15511 16149 15520
rect 16666 15560 16724 15561
rect 16666 15520 16675 15560
rect 16715 15520 16724 15560
rect 16666 15519 16724 15520
rect 17451 15560 17493 15569
rect 18222 15560 18264 15569
rect 17451 15520 17452 15560
rect 17492 15520 17493 15560
rect 17451 15511 17493 15520
rect 17547 15551 17589 15560
rect 17547 15511 17548 15551
rect 17588 15511 17589 15551
rect 17547 15502 17589 15511
rect 18027 15551 18069 15560
rect 18027 15511 18028 15551
rect 18068 15511 18069 15551
rect 18222 15520 18223 15560
rect 18263 15520 18264 15560
rect 18222 15511 18264 15520
rect 18336 15560 18394 15561
rect 18336 15520 18345 15560
rect 18385 15520 18394 15560
rect 18336 15519 18394 15520
rect 18507 15560 18549 15569
rect 18507 15520 18508 15560
rect 18548 15520 18549 15560
rect 18507 15511 18549 15520
rect 18742 15560 18784 15569
rect 18742 15520 18743 15560
rect 18783 15520 18784 15560
rect 18742 15511 18784 15520
rect 18987 15560 19029 15569
rect 18987 15520 18988 15560
rect 19028 15520 19029 15560
rect 18987 15511 19029 15520
rect 19234 15560 19292 15561
rect 19234 15520 19243 15560
rect 19283 15520 19292 15560
rect 19234 15519 19292 15520
rect 19467 15560 19509 15569
rect 19467 15520 19468 15560
rect 19508 15520 19509 15560
rect 19467 15511 19509 15520
rect 19707 15560 19749 15569
rect 19707 15520 19708 15560
rect 19748 15520 19749 15560
rect 19707 15511 19749 15520
rect 19886 15560 19928 15569
rect 19886 15520 19887 15560
rect 19927 15520 19928 15560
rect 19886 15511 19928 15520
rect 20427 15560 20469 15569
rect 20427 15520 20428 15560
rect 20468 15520 20469 15560
rect 20170 15518 20228 15519
rect 18027 15502 18069 15511
rect 13114 15477 13172 15478
rect 11595 15427 11637 15436
rect 12937 15436 12938 15476
rect 12978 15436 12979 15476
rect 12937 15427 12979 15436
rect 14018 15476 14060 15485
rect 14018 15436 14019 15476
rect 14059 15436 14060 15476
rect 14018 15427 14060 15436
rect 14571 15476 14613 15485
rect 14571 15436 14572 15476
rect 14612 15436 14613 15476
rect 18874 15476 18932 15477
rect 14571 15427 14613 15436
rect 15082 15448 15140 15449
rect 15082 15408 15091 15448
rect 15131 15408 15140 15448
rect 18874 15436 18883 15476
rect 18923 15436 18932 15476
rect 18874 15435 18932 15436
rect 19083 15476 19125 15485
rect 19083 15436 19084 15476
rect 19124 15436 19125 15476
rect 19083 15427 19125 15436
rect 19354 15476 19412 15477
rect 19354 15436 19363 15476
rect 19403 15436 19412 15476
rect 19354 15435 19412 15436
rect 19563 15476 19605 15485
rect 19563 15436 19564 15476
rect 19604 15436 19605 15476
rect 19563 15427 19605 15436
rect 20043 15476 20085 15485
rect 20170 15478 20179 15518
rect 20219 15478 20228 15518
rect 20427 15511 20469 15520
rect 20667 15560 20709 15569
rect 20667 15520 20668 15560
rect 20708 15520 20709 15560
rect 20667 15511 20709 15520
rect 20794 15560 20852 15561
rect 20794 15520 20803 15560
rect 20843 15520 20852 15560
rect 20794 15519 20852 15520
rect 20907 15560 20949 15569
rect 20907 15520 20908 15560
rect 20948 15520 20949 15560
rect 20907 15511 20949 15520
rect 21483 15560 21525 15569
rect 21483 15520 21484 15560
rect 21524 15520 21525 15560
rect 21483 15511 21525 15520
rect 21814 15560 21872 15561
rect 21814 15520 21823 15560
rect 21863 15520 21872 15560
rect 21814 15519 21872 15520
rect 22018 15560 22076 15561
rect 22018 15520 22027 15560
rect 22067 15520 22076 15560
rect 22018 15519 22076 15520
rect 22251 15560 22293 15569
rect 22251 15520 22252 15560
rect 22292 15520 22293 15560
rect 22251 15511 22293 15520
rect 22522 15560 22580 15561
rect 22522 15520 22531 15560
rect 22571 15520 22580 15560
rect 22522 15519 22580 15520
rect 22635 15560 22677 15569
rect 22635 15520 22636 15560
rect 22676 15520 22677 15560
rect 23292 15531 23301 15571
rect 23341 15531 23350 15571
rect 23292 15530 23350 15531
rect 23499 15560 23541 15569
rect 22635 15511 22677 15520
rect 23499 15520 23500 15560
rect 23540 15520 23541 15560
rect 23499 15511 23541 15520
rect 23830 15560 23872 15569
rect 24075 15560 24117 15569
rect 23830 15520 23831 15560
rect 23871 15520 23872 15560
rect 23830 15511 23872 15520
rect 23970 15551 24016 15560
rect 23970 15511 23971 15551
rect 24011 15511 24016 15551
rect 24075 15520 24076 15560
rect 24116 15520 24117 15560
rect 24075 15511 24117 15520
rect 24538 15560 24596 15561
rect 24538 15520 24547 15560
rect 24587 15520 24596 15560
rect 24538 15519 24596 15520
rect 24651 15560 24693 15569
rect 24651 15520 24652 15560
rect 24692 15520 24693 15560
rect 24651 15511 24693 15520
rect 25419 15560 25461 15569
rect 25419 15520 25420 15560
rect 25460 15520 25461 15560
rect 25419 15511 25461 15520
rect 25707 15560 25749 15569
rect 25707 15520 25708 15560
rect 25748 15520 25749 15560
rect 25707 15511 25749 15520
rect 27802 15560 27860 15561
rect 27802 15520 27811 15560
rect 27851 15520 27860 15560
rect 27802 15519 27860 15520
rect 28186 15560 28244 15561
rect 28875 15560 28917 15569
rect 28186 15520 28195 15560
rect 28235 15520 28244 15560
rect 28186 15519 28244 15520
rect 28386 15551 28432 15560
rect 28386 15511 28387 15551
rect 28427 15511 28432 15551
rect 28875 15520 28876 15560
rect 28916 15520 28917 15560
rect 28875 15511 28917 15520
rect 29067 15560 29109 15569
rect 29067 15520 29068 15560
rect 29108 15520 29109 15560
rect 29067 15511 29109 15520
rect 29259 15560 29301 15569
rect 29259 15520 29260 15560
rect 29300 15520 29301 15560
rect 29259 15511 29301 15520
rect 23970 15502 24016 15511
rect 28386 15502 28432 15511
rect 20170 15477 20228 15478
rect 20043 15436 20044 15476
rect 20084 15436 20085 15476
rect 20043 15427 20085 15436
rect 20331 15476 20373 15485
rect 20331 15436 20332 15476
rect 20372 15436 20373 15476
rect 20331 15427 20373 15436
rect 20546 15476 20588 15485
rect 20546 15436 20547 15476
rect 20587 15436 20588 15476
rect 20546 15427 20588 15436
rect 21705 15476 21747 15485
rect 21705 15436 21706 15476
rect 21746 15436 21747 15476
rect 21705 15427 21747 15436
rect 22138 15476 22196 15477
rect 22138 15436 22147 15476
rect 22187 15436 22196 15476
rect 22138 15435 22196 15436
rect 26266 15476 26324 15477
rect 26266 15436 26275 15476
rect 26315 15436 26324 15476
rect 26266 15435 26324 15436
rect 28539 15476 28581 15485
rect 28539 15436 28540 15476
rect 28580 15436 28581 15476
rect 28539 15427 28581 15436
rect 15082 15407 15140 15408
rect 1227 15392 1269 15401
rect 1227 15352 1228 15392
rect 1268 15352 1269 15392
rect 1227 15343 1269 15352
rect 11691 15392 11733 15401
rect 11691 15352 11692 15392
rect 11732 15352 11733 15392
rect 11691 15343 11733 15352
rect 13035 15392 13077 15401
rect 13035 15352 13036 15392
rect 13076 15352 13077 15392
rect 13035 15343 13077 15352
rect 13515 15392 13557 15401
rect 13515 15352 13516 15392
rect 13556 15352 13557 15392
rect 13515 15343 13557 15352
rect 14475 15392 14517 15401
rect 14475 15352 14476 15392
rect 14516 15352 14517 15392
rect 14475 15343 14517 15352
rect 16646 15392 16688 15401
rect 16646 15352 16647 15392
rect 16687 15352 16688 15392
rect 16646 15343 16688 15352
rect 19947 15392 19989 15401
rect 19947 15352 19948 15392
rect 19988 15352 19989 15392
rect 19947 15343 19989 15352
rect 21579 15392 21621 15401
rect 21579 15352 21580 15392
rect 21620 15352 21621 15392
rect 21579 15343 21621 15352
rect 3226 15308 3284 15309
rect 3226 15268 3235 15308
rect 3275 15268 3284 15308
rect 3226 15267 3284 15268
rect 5451 15308 5493 15317
rect 5451 15268 5452 15308
rect 5492 15268 5493 15308
rect 5451 15259 5493 15268
rect 6507 15308 6549 15317
rect 6507 15268 6508 15308
rect 6548 15268 6549 15308
rect 6507 15259 6549 15268
rect 6970 15308 7028 15309
rect 6970 15268 6979 15308
rect 7019 15268 7028 15308
rect 6970 15267 7028 15268
rect 8571 15308 8613 15317
rect 8571 15268 8572 15308
rect 8612 15268 8613 15308
rect 8571 15259 8613 15268
rect 10522 15308 10580 15309
rect 10522 15268 10531 15308
rect 10571 15268 10580 15308
rect 10522 15267 10580 15268
rect 12346 15308 12404 15309
rect 12346 15268 12355 15308
rect 12395 15268 12404 15308
rect 12346 15267 12404 15268
rect 17242 15308 17300 15309
rect 17242 15268 17251 15308
rect 17291 15268 17300 15308
rect 17242 15267 17300 15268
rect 18219 15308 18261 15317
rect 18219 15268 18220 15308
rect 18260 15268 18261 15308
rect 18219 15259 18261 15268
rect 22827 15308 22869 15317
rect 22827 15268 22828 15308
rect 22868 15268 22869 15308
rect 22827 15259 22869 15268
rect 23979 15308 24021 15317
rect 23979 15268 23980 15308
rect 24020 15268 24021 15308
rect 23979 15259 24021 15268
rect 576 15140 31392 15164
rect 576 15100 3112 15140
rect 3480 15100 10886 15140
rect 11254 15100 18660 15140
rect 19028 15100 26434 15140
rect 26802 15100 31392 15140
rect 576 15076 31392 15100
rect 4666 14972 4724 14973
rect 4666 14932 4675 14972
rect 4715 14932 4724 14972
rect 4666 14931 4724 14932
rect 5067 14972 5109 14981
rect 5067 14932 5068 14972
rect 5108 14932 5109 14972
rect 5067 14923 5109 14932
rect 9963 14972 10005 14981
rect 9963 14932 9964 14972
rect 10004 14932 10005 14972
rect 9963 14923 10005 14932
rect 12843 14972 12885 14981
rect 12843 14932 12844 14972
rect 12884 14932 12885 14972
rect 12843 14923 12885 14932
rect 13611 14972 13653 14981
rect 13611 14932 13612 14972
rect 13652 14932 13653 14972
rect 13611 14923 13653 14932
rect 14955 14972 14997 14981
rect 14955 14932 14956 14972
rect 14996 14932 14997 14972
rect 14955 14923 14997 14932
rect 17434 14972 17492 14973
rect 17434 14932 17443 14972
rect 17483 14932 17492 14972
rect 17434 14931 17492 14932
rect 17931 14972 17973 14981
rect 17931 14932 17932 14972
rect 17972 14932 17973 14972
rect 17931 14923 17973 14932
rect 18603 14972 18645 14981
rect 18603 14932 18604 14972
rect 18644 14932 18645 14972
rect 18603 14923 18645 14932
rect 19083 14972 19125 14981
rect 19083 14932 19084 14972
rect 19124 14932 19125 14972
rect 19083 14923 19125 14932
rect 20523 14972 20565 14981
rect 20523 14932 20524 14972
rect 20564 14932 20565 14972
rect 20523 14923 20565 14932
rect 21963 14972 22005 14981
rect 21963 14932 21964 14972
rect 22004 14932 22005 14972
rect 21963 14923 22005 14932
rect 23499 14972 23541 14981
rect 23499 14932 23500 14972
rect 23540 14932 23541 14972
rect 23499 14923 23541 14932
rect 28011 14972 28053 14981
rect 28011 14932 28012 14972
rect 28052 14932 28053 14972
rect 28011 14923 28053 14932
rect 28971 14972 29013 14981
rect 28971 14932 28972 14972
rect 29012 14932 29013 14972
rect 28971 14923 29013 14932
rect 3147 14888 3189 14897
rect 3147 14848 3148 14888
rect 3188 14848 3189 14888
rect 3147 14839 3189 14848
rect 3994 14888 4052 14889
rect 3994 14848 4003 14888
rect 4043 14848 4052 14888
rect 3994 14847 4052 14848
rect 8938 14888 8996 14889
rect 8938 14848 8947 14888
rect 8987 14848 8996 14888
rect 8938 14847 8996 14848
rect 11019 14888 11061 14897
rect 11019 14848 11020 14888
rect 11060 14848 11061 14888
rect 11019 14839 11061 14848
rect 15418 14888 15476 14889
rect 15418 14848 15427 14888
rect 15467 14848 15476 14888
rect 15418 14847 15476 14848
rect 19467 14888 19509 14897
rect 19467 14848 19468 14888
rect 19508 14848 19509 14888
rect 19467 14839 19509 14848
rect 20811 14888 20853 14897
rect 20811 14848 20812 14888
rect 20852 14848 20853 14888
rect 20811 14839 20853 14848
rect 23979 14888 24021 14897
rect 23979 14848 23980 14888
rect 24020 14848 24021 14888
rect 23979 14839 24021 14848
rect 26955 14888 26997 14897
rect 26955 14848 26956 14888
rect 26996 14848 26997 14888
rect 26955 14839 26997 14848
rect 29835 14888 29877 14897
rect 29835 14848 29836 14888
rect 29876 14848 29877 14888
rect 29835 14839 29877 14848
rect 1018 14804 1076 14805
rect 1018 14764 1027 14804
rect 1067 14764 1076 14804
rect 1018 14763 1076 14764
rect 2938 14804 2996 14805
rect 2938 14764 2947 14804
rect 2987 14764 2996 14804
rect 2938 14763 2996 14764
rect 5979 14804 6021 14813
rect 5979 14764 5980 14804
rect 6020 14764 6021 14804
rect 5979 14755 6021 14764
rect 6394 14804 6452 14805
rect 6394 14764 6403 14804
rect 6443 14764 6452 14804
rect 6394 14763 6452 14764
rect 6603 14804 6645 14813
rect 6603 14764 6604 14804
rect 6644 14764 6645 14804
rect 6603 14755 6645 14764
rect 7642 14804 7700 14805
rect 7642 14764 7651 14804
rect 7691 14764 7700 14804
rect 7642 14763 7700 14764
rect 7851 14804 7893 14813
rect 7851 14764 7852 14804
rect 7892 14764 7893 14804
rect 7851 14755 7893 14764
rect 9562 14804 9620 14805
rect 9562 14764 9571 14804
rect 9611 14764 9620 14804
rect 9562 14763 9620 14764
rect 9771 14804 9813 14813
rect 9771 14764 9772 14804
rect 9812 14764 9813 14804
rect 9147 14753 9189 14762
rect 9771 14755 9813 14764
rect 10562 14804 10604 14813
rect 10562 14764 10563 14804
rect 10603 14764 10604 14804
rect 11115 14804 11157 14813
rect 10562 14755 10604 14764
rect 10951 14762 10993 14771
rect 2554 14720 2612 14721
rect 2554 14680 2563 14720
rect 2603 14680 2612 14720
rect 2554 14679 2612 14680
rect 3147 14720 3189 14729
rect 3147 14680 3148 14720
rect 3188 14680 3189 14720
rect 3147 14671 3189 14680
rect 3264 14720 3322 14721
rect 3264 14680 3273 14720
rect 3313 14680 3322 14720
rect 3264 14679 3322 14680
rect 3435 14720 3477 14729
rect 3435 14680 3436 14720
rect 3476 14680 3477 14720
rect 3435 14671 3477 14680
rect 3819 14720 3861 14729
rect 3819 14680 3820 14720
rect 3860 14680 3861 14720
rect 3819 14671 3861 14680
rect 3994 14720 4052 14721
rect 3994 14680 4003 14720
rect 4043 14680 4052 14720
rect 3994 14679 4052 14680
rect 4480 14720 4522 14729
rect 4480 14680 4481 14720
rect 4521 14680 4522 14720
rect 4480 14671 4522 14680
rect 4587 14720 4629 14729
rect 4587 14680 4588 14720
rect 4628 14680 4629 14720
rect 4587 14671 4629 14680
rect 4971 14720 5013 14729
rect 4971 14680 4972 14720
rect 5012 14680 5013 14720
rect 4971 14671 5013 14680
rect 5163 14720 5205 14729
rect 5163 14680 5164 14720
rect 5204 14680 5205 14720
rect 5163 14671 5205 14680
rect 5302 14720 5344 14729
rect 5302 14680 5303 14720
rect 5343 14680 5344 14720
rect 5302 14671 5344 14680
rect 5434 14720 5492 14721
rect 5434 14680 5443 14720
rect 5483 14680 5492 14720
rect 5434 14679 5492 14680
rect 5547 14720 5589 14729
rect 5547 14680 5548 14720
rect 5588 14680 5589 14720
rect 5547 14671 5589 14680
rect 5815 14720 5873 14721
rect 5815 14680 5824 14720
rect 5864 14680 5873 14720
rect 5815 14679 5873 14680
rect 6262 14720 6304 14729
rect 6262 14680 6263 14720
rect 6303 14680 6304 14720
rect 6262 14671 6304 14680
rect 6507 14720 6549 14729
rect 6507 14680 6508 14720
rect 6548 14680 6549 14720
rect 6507 14671 6549 14680
rect 6972 14720 7014 14729
rect 6972 14680 6973 14720
rect 7013 14680 7014 14720
rect 6972 14671 7014 14680
rect 7083 14720 7125 14729
rect 7083 14680 7084 14720
rect 7124 14680 7125 14720
rect 7083 14671 7125 14680
rect 7510 14720 7552 14729
rect 7510 14680 7511 14720
rect 7551 14680 7552 14720
rect 7510 14671 7552 14680
rect 7755 14720 7797 14729
rect 7755 14680 7756 14720
rect 7796 14680 7797 14720
rect 7755 14671 7797 14680
rect 8023 14720 8081 14721
rect 8023 14680 8032 14720
rect 8072 14680 8081 14720
rect 8023 14679 8081 14680
rect 8845 14720 8903 14721
rect 8845 14680 8854 14720
rect 8894 14680 8903 14720
rect 9147 14713 9148 14753
rect 9188 14713 9189 14753
rect 9147 14704 9189 14713
rect 9243 14720 9285 14729
rect 8845 14679 8903 14680
rect 9243 14680 9244 14720
rect 9284 14680 9285 14720
rect 9243 14671 9285 14680
rect 9447 14720 9489 14729
rect 9447 14680 9448 14720
rect 9488 14680 9489 14720
rect 9447 14671 9489 14680
rect 9675 14720 9717 14729
rect 9675 14680 9676 14720
rect 9716 14680 9717 14720
rect 9675 14671 9717 14680
rect 9963 14720 10005 14729
rect 9963 14680 9964 14720
rect 10004 14680 10005 14720
rect 9963 14671 10005 14680
rect 10155 14720 10197 14729
rect 10155 14680 10156 14720
rect 10196 14680 10197 14720
rect 10155 14671 10197 14680
rect 10443 14720 10485 14729
rect 10443 14680 10444 14720
rect 10484 14680 10485 14720
rect 10443 14671 10485 14680
rect 10660 14720 10702 14729
rect 10951 14722 10952 14762
rect 10992 14722 10993 14762
rect 11115 14764 11116 14804
rect 11156 14764 11157 14804
rect 11115 14755 11157 14764
rect 11787 14804 11829 14813
rect 11787 14764 11788 14804
rect 11828 14764 11829 14804
rect 11787 14755 11829 14764
rect 12651 14804 12693 14813
rect 12651 14764 12652 14804
rect 12692 14764 12693 14804
rect 12651 14755 12693 14764
rect 14554 14804 14612 14805
rect 14554 14764 14563 14804
rect 14603 14764 14612 14804
rect 14554 14763 14612 14764
rect 22370 14804 22412 14813
rect 22370 14764 22371 14804
rect 22411 14764 22412 14804
rect 15711 14753 15753 14762
rect 10660 14680 10661 14720
rect 10701 14680 10702 14720
rect 10660 14671 10702 14680
rect 10788 14720 10846 14721
rect 10788 14680 10797 14720
rect 10837 14680 10846 14720
rect 10951 14713 10993 14722
rect 11451 14720 11493 14729
rect 10788 14679 10846 14680
rect 11451 14680 11452 14720
rect 11492 14680 11493 14720
rect 11242 14678 11300 14679
rect 11242 14638 11251 14678
rect 11291 14638 11300 14678
rect 11451 14671 11493 14680
rect 11578 14720 11636 14721
rect 11578 14680 11587 14720
rect 11627 14680 11636 14720
rect 11578 14679 11636 14680
rect 11691 14720 11733 14729
rect 11691 14680 11692 14720
rect 11732 14680 11733 14720
rect 11691 14671 11733 14680
rect 11979 14720 12021 14729
rect 11979 14680 11980 14720
rect 12020 14680 12021 14720
rect 11979 14671 12021 14680
rect 12171 14720 12213 14729
rect 12171 14680 12172 14720
rect 12212 14680 12213 14720
rect 12171 14671 12213 14680
rect 12886 14720 12928 14729
rect 13131 14720 13173 14729
rect 12886 14680 12887 14720
rect 12927 14680 12928 14720
rect 12886 14671 12928 14680
rect 13026 14711 13072 14720
rect 13026 14671 13027 14711
rect 13067 14671 13072 14711
rect 13131 14680 13132 14720
rect 13172 14680 13173 14720
rect 13131 14671 13173 14680
rect 13306 14720 13364 14721
rect 13306 14680 13315 14720
rect 13355 14680 13364 14720
rect 13306 14679 13364 14680
rect 13419 14720 13461 14729
rect 13419 14680 13420 14720
rect 13460 14680 13461 14720
rect 13419 14671 13461 14680
rect 13899 14720 13941 14729
rect 13899 14680 13900 14720
rect 13940 14680 13941 14720
rect 13899 14671 13941 14680
rect 14018 14720 14060 14729
rect 14018 14680 14019 14720
rect 14059 14680 14060 14720
rect 14018 14671 14060 14680
rect 14128 14720 14186 14721
rect 14667 14720 14709 14729
rect 14128 14680 14137 14720
rect 14177 14680 14186 14720
rect 14128 14679 14186 14680
rect 14370 14711 14416 14720
rect 14370 14671 14371 14711
rect 14411 14671 14416 14711
rect 14667 14680 14668 14720
rect 14708 14680 14709 14720
rect 14667 14671 14709 14680
rect 14955 14720 14997 14729
rect 14955 14680 14956 14720
rect 14996 14680 14997 14720
rect 14955 14671 14997 14680
rect 15147 14720 15189 14729
rect 15147 14680 15148 14720
rect 15188 14680 15189 14720
rect 15711 14713 15712 14753
rect 15752 14713 15753 14753
rect 18786 14753 18832 14762
rect 15711 14704 15753 14713
rect 15802 14720 15860 14721
rect 15147 14671 15189 14680
rect 15802 14680 15811 14720
rect 15851 14680 15860 14720
rect 15802 14679 15860 14680
rect 16096 14720 16138 14729
rect 16096 14680 16097 14720
rect 16137 14680 16138 14720
rect 16096 14671 16138 14680
rect 16387 14720 16445 14721
rect 16387 14680 16396 14720
rect 16436 14680 16445 14720
rect 16387 14679 16445 14680
rect 16587 14720 16629 14729
rect 16587 14680 16588 14720
rect 16628 14680 16629 14720
rect 16587 14671 16629 14680
rect 16779 14720 16821 14729
rect 16779 14680 16780 14720
rect 16820 14680 16821 14720
rect 16779 14671 16821 14680
rect 17259 14720 17301 14729
rect 17259 14680 17260 14720
rect 17300 14680 17301 14720
rect 17259 14671 17301 14680
rect 17434 14720 17492 14721
rect 17434 14680 17443 14720
rect 17483 14680 17492 14720
rect 17434 14679 17492 14680
rect 17931 14720 17973 14729
rect 17931 14680 17932 14720
rect 17972 14680 17973 14720
rect 17931 14671 17973 14680
rect 18123 14720 18165 14729
rect 18123 14680 18124 14720
rect 18164 14680 18165 14720
rect 18123 14671 18165 14680
rect 18411 14720 18453 14729
rect 18411 14680 18412 14720
rect 18452 14680 18453 14720
rect 18411 14671 18453 14680
rect 18646 14720 18688 14729
rect 18646 14680 18647 14720
rect 18687 14680 18688 14720
rect 18786 14713 18787 14753
rect 18827 14713 18832 14753
rect 21339 14753 21381 14762
rect 22370 14755 22412 14764
rect 23019 14804 23061 14813
rect 23019 14764 23020 14804
rect 23060 14764 23061 14804
rect 23019 14755 23061 14764
rect 23153 14804 23195 14813
rect 23153 14764 23154 14804
rect 23194 14764 23195 14804
rect 23153 14755 23195 14764
rect 26571 14804 26613 14813
rect 26571 14764 26572 14804
rect 26612 14764 26613 14804
rect 18786 14704 18832 14713
rect 18878 14720 18936 14721
rect 18646 14671 18688 14680
rect 18878 14680 18887 14720
rect 18927 14680 18936 14720
rect 18878 14679 18936 14680
rect 19083 14720 19125 14729
rect 19083 14680 19084 14720
rect 19124 14680 19125 14720
rect 19083 14671 19125 14680
rect 19275 14720 19317 14729
rect 19275 14680 19276 14720
rect 19316 14680 19317 14720
rect 19275 14671 19317 14680
rect 20218 14720 20276 14721
rect 20218 14680 20227 14720
rect 20267 14680 20276 14720
rect 20218 14679 20276 14680
rect 20534 14720 20576 14729
rect 20534 14680 20535 14720
rect 20575 14680 20576 14720
rect 20534 14671 20576 14680
rect 20715 14720 20757 14729
rect 20715 14680 20716 14720
rect 20756 14680 20757 14720
rect 20715 14671 20757 14680
rect 20842 14720 20900 14721
rect 20842 14680 20851 14720
rect 20891 14680 20900 14720
rect 20842 14679 20900 14680
rect 20956 14720 21014 14721
rect 20956 14680 20965 14720
rect 21005 14680 21014 14720
rect 21339 14713 21340 14753
rect 21380 14713 21381 14753
rect 23542 14753 23584 14762
rect 26571 14755 26613 14764
rect 21339 14704 21381 14713
rect 21435 14720 21477 14729
rect 20956 14679 21014 14680
rect 21435 14680 21436 14720
rect 21476 14680 21477 14720
rect 21435 14671 21477 14680
rect 21675 14720 21717 14729
rect 21675 14680 21676 14720
rect 21716 14680 21717 14720
rect 21675 14671 21717 14680
rect 21807 14720 21865 14721
rect 21807 14680 21816 14720
rect 21856 14680 21865 14720
rect 21807 14679 21865 14680
rect 21916 14720 21974 14721
rect 21916 14680 21925 14720
rect 21965 14680 21974 14720
rect 21916 14679 21974 14680
rect 22251 14720 22293 14729
rect 22251 14680 22252 14720
rect 22292 14680 22293 14720
rect 22251 14671 22293 14680
rect 22468 14720 22510 14729
rect 22468 14680 22469 14720
rect 22509 14680 22510 14720
rect 22468 14671 22510 14680
rect 22666 14720 22724 14721
rect 22666 14680 22675 14720
rect 22715 14680 22724 14720
rect 22666 14679 22724 14680
rect 22923 14720 22965 14729
rect 22923 14680 22924 14720
rect 22964 14680 22965 14720
rect 22923 14671 22965 14680
rect 23254 14720 23312 14721
rect 23254 14680 23263 14720
rect 23303 14680 23312 14720
rect 23542 14713 23543 14753
rect 23583 14713 23584 14753
rect 23787 14720 23829 14729
rect 23542 14704 23584 14713
rect 23682 14711 23728 14720
rect 23254 14679 23312 14680
rect 23682 14671 23683 14711
rect 23723 14671 23728 14711
rect 23787 14680 23788 14720
rect 23828 14680 23829 14720
rect 23787 14671 23829 14680
rect 24132 14720 24190 14721
rect 24132 14680 24141 14720
rect 24181 14680 24190 14720
rect 24132 14679 24190 14680
rect 24248 14720 24306 14721
rect 24248 14680 24257 14720
rect 24297 14680 24306 14720
rect 24248 14679 24306 14680
rect 24360 14720 24418 14721
rect 24360 14680 24369 14720
rect 24409 14680 24418 14720
rect 24360 14679 24418 14680
rect 25018 14720 25076 14721
rect 25018 14680 25027 14720
rect 25067 14680 25076 14720
rect 25018 14679 25076 14680
rect 27339 14720 27381 14729
rect 27339 14680 27340 14720
rect 27380 14680 27381 14720
rect 27339 14671 27381 14680
rect 28138 14720 28196 14721
rect 28138 14680 28147 14720
rect 28187 14680 28196 14720
rect 28138 14679 28196 14680
rect 29643 14720 29685 14729
rect 29643 14680 29644 14720
rect 29684 14680 29685 14720
rect 29643 14671 29685 14680
rect 13026 14662 13072 14671
rect 14370 14662 14416 14671
rect 23682 14662 23728 14671
rect 11242 14637 11300 14638
rect 5626 14636 5684 14637
rect 5626 14596 5635 14636
rect 5675 14596 5684 14636
rect 5626 14595 5684 14596
rect 12075 14636 12117 14645
rect 12075 14596 12076 14636
rect 12116 14596 12117 14636
rect 12075 14587 12117 14596
rect 13622 14636 13664 14645
rect 13622 14596 13623 14636
rect 13663 14596 13664 14636
rect 13622 14587 13664 14596
rect 20331 14636 20373 14645
rect 20331 14596 20332 14636
rect 20372 14596 20373 14636
rect 20331 14587 20373 14596
rect 24634 14636 24692 14637
rect 24634 14596 24643 14636
rect 24683 14596 24692 14636
rect 24634 14595 24692 14596
rect 28347 14636 28389 14645
rect 28347 14596 28348 14636
rect 28388 14596 28389 14636
rect 28347 14587 28389 14596
rect 651 14552 693 14561
rect 651 14512 652 14552
rect 692 14512 693 14552
rect 651 14503 693 14512
rect 6778 14552 6836 14553
rect 6778 14512 6787 14552
rect 6827 14512 6836 14552
rect 6778 14511 6836 14512
rect 8187 14552 8229 14561
rect 8187 14512 8188 14552
rect 8228 14512 8229 14552
rect 8187 14503 8229 14512
rect 8650 14552 8708 14553
rect 8650 14512 8659 14552
rect 8699 14512 8708 14552
rect 8650 14511 8708 14512
rect 10347 14552 10389 14561
rect 10347 14512 10348 14552
rect 10388 14512 10389 14552
rect 10347 14503 10389 14512
rect 12411 14552 12453 14561
rect 12411 14512 12412 14552
rect 12452 14512 12453 14552
rect 12411 14503 12453 14512
rect 13803 14552 13845 14561
rect 13803 14512 13804 14552
rect 13844 14512 13845 14552
rect 13803 14503 13845 14512
rect 15946 14552 16004 14553
rect 15946 14512 15955 14552
rect 15995 14512 16004 14552
rect 15946 14511 16004 14512
rect 16186 14552 16244 14553
rect 16186 14512 16195 14552
rect 16235 14512 16244 14552
rect 16186 14511 16244 14512
rect 16299 14552 16341 14561
rect 16299 14512 16300 14552
rect 16340 14512 16341 14552
rect 16299 14503 16341 14512
rect 16683 14552 16725 14561
rect 16683 14512 16684 14552
rect 16724 14512 16725 14552
rect 16683 14503 16725 14512
rect 18267 14552 18309 14561
rect 18267 14512 18268 14552
rect 18308 14512 18309 14552
rect 18267 14503 18309 14512
rect 19851 14552 19893 14561
rect 19851 14512 19852 14552
rect 19892 14512 19893 14552
rect 19851 14503 19893 14512
rect 21178 14552 21236 14553
rect 21178 14512 21187 14552
rect 21227 14512 21236 14552
rect 21178 14511 21236 14512
rect 22155 14552 22197 14561
rect 22155 14512 22156 14552
rect 22196 14512 22197 14552
rect 22155 14503 22197 14512
rect 22779 14552 22821 14561
rect 22779 14512 22780 14552
rect 22820 14512 22821 14552
rect 22779 14503 22821 14512
rect 23019 14552 23061 14561
rect 23019 14512 23020 14552
rect 23060 14512 23061 14552
rect 23019 14503 23061 14512
rect 576 14384 31392 14408
rect 576 14344 4352 14384
rect 4720 14344 12126 14384
rect 12494 14344 19900 14384
rect 20268 14344 27674 14384
rect 28042 14344 31392 14384
rect 576 14320 31392 14344
rect 730 14216 788 14217
rect 730 14176 739 14216
rect 779 14176 788 14216
rect 730 14175 788 14176
rect 1227 14216 1269 14225
rect 1227 14176 1228 14216
rect 1268 14176 1269 14216
rect 1227 14167 1269 14176
rect 3051 14216 3093 14225
rect 3051 14176 3052 14216
rect 3092 14176 3093 14216
rect 3051 14167 3093 14176
rect 3723 14216 3765 14225
rect 3723 14176 3724 14216
rect 3764 14176 3765 14216
rect 3723 14167 3765 14176
rect 4186 14216 4244 14217
rect 4186 14176 4195 14216
rect 4235 14176 4244 14216
rect 4186 14175 4244 14176
rect 4971 14216 5013 14225
rect 4971 14176 4972 14216
rect 5012 14176 5013 14216
rect 4971 14167 5013 14176
rect 5818 14216 5876 14217
rect 5818 14176 5827 14216
rect 5867 14176 5876 14216
rect 5818 14175 5876 14176
rect 6123 14216 6165 14225
rect 6123 14176 6124 14216
rect 6164 14176 6165 14216
rect 6123 14167 6165 14176
rect 7179 14216 7221 14225
rect 7179 14176 7180 14216
rect 7220 14176 7221 14216
rect 7179 14167 7221 14176
rect 7371 14216 7413 14225
rect 7371 14176 7372 14216
rect 7412 14176 7413 14216
rect 7371 14167 7413 14176
rect 8026 14216 8084 14217
rect 8026 14176 8035 14216
rect 8075 14176 8084 14216
rect 8026 14175 8084 14176
rect 9322 14216 9380 14217
rect 9322 14176 9331 14216
rect 9371 14176 9380 14216
rect 9322 14175 9380 14176
rect 9754 14216 9812 14217
rect 9754 14176 9763 14216
rect 9803 14176 9812 14216
rect 9754 14175 9812 14176
rect 10539 14216 10581 14225
rect 10539 14176 10540 14216
rect 10580 14176 10581 14216
rect 10539 14167 10581 14176
rect 12586 14216 12644 14217
rect 12586 14176 12595 14216
rect 12635 14176 12644 14216
rect 12586 14175 12644 14176
rect 13978 14216 14036 14217
rect 13978 14176 13987 14216
rect 14027 14176 14036 14216
rect 13978 14175 14036 14176
rect 15226 14216 15284 14217
rect 15226 14176 15235 14216
rect 15275 14176 15284 14216
rect 15226 14175 15284 14176
rect 15994 14216 16052 14217
rect 15994 14176 16003 14216
rect 16043 14176 16052 14216
rect 15994 14175 16052 14176
rect 16570 14216 16628 14217
rect 16570 14176 16579 14216
rect 16619 14176 16628 14216
rect 16570 14175 16628 14176
rect 18891 14216 18933 14225
rect 18891 14176 18892 14216
rect 18932 14176 18933 14216
rect 18891 14167 18933 14176
rect 19371 14216 19413 14225
rect 19371 14176 19372 14216
rect 19412 14176 19413 14216
rect 19371 14167 19413 14176
rect 21946 14216 22004 14217
rect 21946 14176 21955 14216
rect 21995 14176 22004 14216
rect 21946 14175 22004 14176
rect 22251 14216 22293 14225
rect 22251 14176 22252 14216
rect 22292 14176 22293 14216
rect 22251 14167 22293 14176
rect 24154 14216 24212 14217
rect 24154 14176 24163 14216
rect 24203 14176 24212 14216
rect 24154 14175 24212 14176
rect 24747 14216 24789 14225
rect 24747 14176 24748 14216
rect 24788 14176 24789 14216
rect 24747 14167 24789 14176
rect 29451 14216 29493 14225
rect 29451 14176 29452 14216
rect 29492 14176 29493 14216
rect 29451 14167 29493 14176
rect 10262 14132 10304 14141
rect 5058 14123 5104 14132
rect 5058 14083 5059 14123
rect 5099 14083 5104 14123
rect 10262 14092 10263 14132
rect 10303 14092 10304 14132
rect 10262 14083 10304 14092
rect 12507 14132 12549 14141
rect 12507 14092 12508 14132
rect 12548 14092 12549 14132
rect 12507 14083 12549 14092
rect 15901 14132 15943 14141
rect 15901 14092 15902 14132
rect 15942 14092 15943 14132
rect 15901 14083 15943 14092
rect 19947 14132 19989 14141
rect 19947 14092 19948 14132
rect 19988 14092 19989 14132
rect 19947 14083 19989 14092
rect 21370 14132 21428 14133
rect 21370 14092 21379 14132
rect 21419 14092 21428 14132
rect 21370 14091 21428 14092
rect 22539 14132 22581 14141
rect 22539 14092 22540 14132
rect 22580 14092 22581 14132
rect 22539 14083 22581 14092
rect 24634 14132 24692 14133
rect 24634 14092 24643 14132
rect 24683 14092 24692 14132
rect 24634 14091 24692 14092
rect 5058 14074 5104 14083
rect 843 14048 885 14057
rect 843 14008 844 14048
rect 884 14008 885 14048
rect 843 13999 885 14008
rect 1899 14048 1941 14057
rect 1899 14008 1900 14048
rect 1940 14008 1941 14048
rect 1899 13999 1941 14008
rect 2752 14048 2794 14057
rect 2752 14008 2753 14048
rect 2793 14008 2794 14048
rect 2752 13999 2794 14008
rect 2859 14048 2901 14057
rect 2859 14008 2860 14048
rect 2900 14008 2901 14048
rect 2859 13999 2901 14008
rect 3243 14048 3285 14057
rect 3243 14008 3244 14048
rect 3284 14008 3285 14048
rect 3243 13999 3285 14008
rect 3531 14048 3573 14057
rect 3531 14008 3532 14048
rect 3572 14008 3573 14048
rect 4226 14048 4268 14057
rect 3531 13999 3573 14008
rect 4027 14037 4069 14046
rect 4027 13997 4028 14037
rect 4068 13997 4069 14037
rect 4226 14008 4227 14048
rect 4267 14008 4268 14048
rect 4226 13999 4268 14008
rect 4330 14048 4388 14049
rect 4330 14008 4339 14048
rect 4379 14008 4388 14048
rect 4330 14007 4388 14008
rect 4474 14048 4532 14049
rect 4474 14008 4483 14048
rect 4523 14008 4532 14048
rect 4474 14007 4532 14008
rect 4596 14048 4654 14049
rect 4596 14008 4605 14048
rect 4645 14008 4654 14048
rect 4596 14007 4654 14008
rect 4762 14048 4820 14049
rect 5146 14048 5204 14049
rect 4762 14008 4771 14048
rect 4811 14008 4820 14048
rect 4762 14007 4820 14008
rect 4875 14039 4917 14048
rect 4875 13999 4876 14039
rect 4916 13999 4917 14039
rect 5146 14008 5155 14048
rect 5195 14008 5204 14048
rect 5146 14007 5204 14008
rect 5323 14048 5381 14049
rect 5323 14008 5332 14048
rect 5372 14008 5381 14048
rect 5323 14007 5381 14008
rect 5494 14048 5536 14057
rect 5494 14008 5495 14048
rect 5535 14008 5536 14048
rect 5494 13999 5536 14008
rect 5739 14048 5781 14057
rect 5739 14008 5740 14048
rect 5780 14008 5781 14048
rect 5739 13999 5781 14008
rect 6027 14048 6069 14057
rect 6027 14008 6028 14048
rect 6068 14008 6069 14048
rect 6027 13999 6069 14008
rect 6219 14048 6261 14057
rect 6219 14008 6220 14048
rect 6260 14008 6261 14048
rect 6219 13999 6261 14008
rect 6370 14048 6428 14049
rect 6370 14008 6379 14048
rect 6419 14008 6428 14048
rect 6370 14007 6428 14008
rect 6490 14048 6548 14049
rect 6490 14008 6499 14048
rect 6539 14008 6548 14048
rect 6490 14007 6548 14008
rect 6603 14048 6645 14057
rect 6603 14008 6604 14048
rect 6644 14008 6645 14048
rect 6603 13999 6645 14008
rect 6891 14048 6933 14057
rect 6891 14008 6892 14048
rect 6932 14008 6933 14048
rect 6891 13999 6933 14008
rect 7132 14048 7190 14049
rect 7751 14048 7809 14049
rect 7132 14008 7141 14048
rect 7181 14008 7190 14048
rect 7132 14007 7190 14008
rect 7532 14039 7574 14048
rect 7005 14006 7063 14007
rect 4027 13988 4069 13997
rect 4875 13990 4917 13999
rect 5626 13964 5684 13965
rect 5626 13924 5635 13964
rect 5675 13924 5684 13964
rect 5626 13923 5684 13924
rect 6699 13964 6741 13973
rect 7005 13966 7014 14006
rect 7054 13966 7063 14006
rect 7532 13999 7533 14039
rect 7573 13999 7574 14039
rect 7532 13990 7574 13999
rect 7650 14039 7696 14048
rect 7650 13999 7651 14039
rect 7691 13999 7696 14039
rect 7751 14008 7760 14048
rect 7800 14008 7809 14048
rect 7751 14007 7809 14008
rect 8187 14048 8229 14057
rect 8187 14008 8188 14048
rect 8228 14008 8229 14048
rect 8187 13999 8229 14008
rect 8331 14048 8373 14057
rect 9178 14048 9236 14049
rect 8331 14008 8332 14048
rect 8372 14008 8373 14048
rect 8331 13999 8373 14008
rect 9087 14039 9129 14048
rect 9087 13999 9088 14039
rect 9128 13999 9129 14039
rect 9178 14008 9187 14048
rect 9227 14008 9236 14048
rect 9178 14007 9236 14008
rect 9430 14048 9472 14057
rect 9430 14008 9431 14048
rect 9471 14008 9472 14048
rect 9430 13999 9472 14008
rect 9675 14048 9717 14057
rect 9675 14008 9676 14048
rect 9716 14008 9717 14048
rect 9675 13999 9717 14008
rect 9946 14048 10004 14049
rect 9946 14008 9955 14048
rect 9995 14008 10004 14048
rect 9946 14007 10004 14008
rect 10059 14048 10101 14057
rect 10059 14008 10060 14048
rect 10100 14008 10101 14048
rect 10059 13999 10101 14008
rect 10443 14048 10485 14057
rect 10443 14008 10444 14048
rect 10484 14008 10485 14048
rect 10443 13999 10485 14008
rect 10633 14048 10675 14057
rect 10971 14048 11013 14057
rect 10633 14008 10634 14048
rect 10674 14008 10675 14048
rect 10633 13999 10675 14008
rect 10818 14039 10864 14048
rect 10818 13999 10819 14039
rect 10859 13999 10864 14039
rect 10971 14008 10972 14048
rect 11012 14008 11013 14048
rect 10971 13999 11013 14008
rect 11403 14048 11445 14057
rect 11403 14008 11404 14048
rect 11444 14008 11445 14048
rect 11403 13999 11445 14008
rect 11518 14048 11560 14057
rect 11518 14008 11519 14048
rect 11559 14008 11560 14048
rect 11518 13999 11560 14008
rect 11691 14048 11733 14057
rect 11691 14008 11692 14048
rect 11732 14008 11733 14048
rect 11691 13999 11733 14008
rect 11883 14048 11925 14057
rect 11883 14008 11884 14048
rect 11924 14008 11925 14048
rect 11883 13999 11925 14008
rect 12267 14048 12309 14057
rect 12267 14008 12268 14048
rect 12308 14008 12309 14048
rect 12267 13999 12309 14008
rect 12730 14048 12788 14049
rect 13323 14048 13365 14057
rect 12730 14008 12739 14048
rect 12779 14008 12788 14048
rect 12730 14007 12788 14008
rect 12843 14039 12885 14048
rect 12843 13999 12844 14039
rect 12884 13999 12885 14039
rect 13323 14008 13324 14048
rect 13364 14008 13365 14048
rect 13323 13999 13365 14008
rect 13498 14048 13556 14049
rect 13498 14008 13507 14048
rect 13547 14008 13556 14048
rect 13884 14048 13942 14049
rect 14475 14048 14517 14057
rect 13498 14007 13556 14008
rect 13659 14006 13701 14015
rect 13884 14008 13893 14048
rect 13933 14008 13942 14048
rect 13884 14007 13942 14008
rect 14178 14039 14224 14048
rect 7650 13990 7696 13999
rect 9087 13990 9129 13999
rect 10818 13990 10864 13999
rect 12843 13990 12885 13999
rect 7005 13965 7063 13966
rect 13659 13966 13660 14006
rect 13700 13966 13701 14006
rect 14178 13999 14179 14039
rect 14219 13999 14224 14039
rect 14475 14008 14476 14048
rect 14516 14008 14517 14048
rect 14475 13999 14517 14008
rect 14902 14048 14944 14057
rect 14902 14008 14903 14048
rect 14943 14008 14944 14048
rect 14902 13999 14944 14008
rect 15147 14048 15189 14057
rect 15147 14008 15148 14048
rect 15188 14008 15189 14048
rect 15147 13999 15189 14008
rect 15531 14048 15573 14057
rect 15531 14008 15532 14048
rect 15572 14008 15573 14048
rect 15531 13999 15573 14008
rect 15760 14048 15818 14049
rect 15760 14008 15769 14048
rect 15809 14008 15818 14048
rect 15760 14007 15818 14008
rect 16107 14048 16149 14057
rect 16875 14048 16917 14057
rect 16107 14008 16108 14048
rect 16148 14008 16149 14048
rect 16107 13999 16149 14008
rect 16203 14039 16245 14048
rect 16203 13999 16204 14039
rect 16244 13999 16245 14039
rect 16875 14008 16876 14048
rect 16916 14008 16917 14048
rect 16875 13999 16917 14008
rect 17643 14048 17685 14057
rect 17643 14008 17644 14048
rect 17684 14008 17685 14048
rect 17643 13999 17685 14008
rect 18267 14048 18309 14057
rect 18267 14008 18268 14048
rect 18308 14008 18309 14048
rect 18267 13999 18309 14008
rect 18568 14048 18610 14057
rect 18568 14008 18569 14048
rect 18609 14008 18610 14048
rect 18568 13999 18610 14008
rect 18730 14048 18788 14049
rect 18730 14008 18739 14048
rect 18779 14008 18788 14048
rect 18730 14007 18788 14008
rect 18987 14048 19029 14057
rect 18987 14008 18988 14048
rect 19028 14008 19029 14048
rect 18987 13999 19029 14008
rect 19216 14048 19274 14049
rect 19216 14008 19225 14048
rect 19265 14008 19274 14048
rect 19696 14048 19754 14049
rect 19216 14007 19274 14008
rect 19467 14006 19509 14015
rect 19696 14008 19705 14048
rect 19745 14008 19754 14048
rect 19696 14007 19754 14008
rect 19851 14048 19893 14057
rect 19851 14008 19852 14048
rect 19892 14008 19893 14048
rect 14178 13990 14224 13999
rect 16203 13990 16245 13999
rect 6699 13924 6700 13964
rect 6740 13924 6741 13964
rect 6699 13915 6741 13924
rect 9562 13964 9620 13965
rect 9562 13924 9571 13964
rect 9611 13924 9620 13964
rect 13659 13957 13701 13966
rect 13786 13964 13844 13965
rect 9562 13923 9620 13924
rect 13786 13924 13795 13964
rect 13835 13924 13844 13964
rect 13786 13923 13844 13924
rect 15034 13964 15092 13965
rect 15034 13924 15043 13964
rect 15083 13924 15092 13964
rect 15034 13923 15092 13924
rect 15435 13964 15477 13973
rect 15435 13924 15436 13964
rect 15476 13924 15477 13964
rect 15435 13915 15477 13924
rect 15650 13964 15692 13973
rect 15650 13924 15651 13964
rect 15691 13924 15692 13964
rect 15650 13915 15692 13924
rect 16785 13964 16827 13973
rect 16785 13924 16786 13964
rect 16826 13924 16827 13964
rect 16785 13915 16827 13924
rect 17553 13964 17595 13973
rect 17553 13924 17554 13964
rect 17594 13924 17595 13964
rect 17553 13915 17595 13924
rect 18411 13964 18453 13973
rect 18411 13924 18412 13964
rect 18452 13924 18453 13964
rect 18411 13915 18453 13924
rect 19106 13964 19148 13973
rect 19106 13924 19107 13964
rect 19147 13924 19148 13964
rect 19467 13966 19468 14006
rect 19508 13966 19509 14006
rect 19851 13999 19893 14008
rect 20139 14048 20181 14057
rect 20139 14008 20140 14048
rect 20180 14008 20181 14048
rect 20139 13999 20181 14008
rect 20331 14048 20373 14057
rect 20331 14008 20332 14048
rect 20372 14008 20373 14048
rect 20331 13999 20373 14008
rect 20506 14048 20564 14049
rect 20506 14008 20515 14048
rect 20555 14008 20564 14048
rect 20506 14007 20564 14008
rect 20619 14048 20661 14057
rect 20619 14008 20620 14048
rect 20660 14008 20661 14048
rect 20619 13999 20661 14008
rect 20811 14048 20853 14057
rect 20811 14008 20812 14048
rect 20852 14008 20853 14048
rect 20811 13999 20853 14008
rect 21142 14048 21200 14049
rect 21522 14048 21580 14049
rect 21771 14048 21813 14057
rect 21142 14008 21151 14048
rect 21191 14008 21200 14048
rect 21142 14007 21200 14008
rect 21432 14039 21474 14048
rect 21432 13999 21433 14039
rect 21473 13999 21474 14039
rect 21522 14008 21531 14048
rect 21571 14008 21580 14048
rect 21522 14007 21580 14008
rect 21666 14039 21712 14048
rect 21432 13990 21474 13999
rect 21666 13999 21667 14039
rect 21707 13999 21712 14039
rect 21771 14008 21772 14048
rect 21812 14008 21813 14048
rect 21771 13999 21813 14008
rect 22059 14048 22101 14057
rect 22059 14008 22060 14048
rect 22100 14008 22101 14048
rect 22059 13999 22101 14008
rect 22443 14048 22485 14057
rect 22443 14008 22444 14048
rect 22484 14008 22485 14048
rect 22443 13999 22485 14008
rect 22635 14048 22677 14057
rect 22635 14008 22636 14048
rect 22676 14008 22677 14048
rect 22635 13999 22677 14008
rect 22788 14048 22846 14049
rect 22788 14008 22797 14048
rect 22837 14008 22846 14048
rect 23403 14048 23445 14057
rect 22788 14007 22846 14008
rect 22923 14006 22965 14015
rect 23403 14008 23404 14048
rect 23444 14008 23445 14048
rect 21666 13990 21712 13999
rect 19467 13957 19509 13966
rect 19586 13964 19628 13973
rect 22923 13966 22924 14006
rect 22964 13966 22965 14006
rect 19106 13915 19148 13924
rect 19586 13924 19587 13964
rect 19627 13924 19628 13964
rect 19586 13915 19628 13924
rect 21042 13955 21088 13964
rect 22923 13957 22965 13966
rect 23242 14006 23300 14007
rect 23242 13966 23251 14006
rect 23291 13966 23300 14006
rect 23403 13999 23445 14008
rect 23734 14048 23792 14049
rect 23734 14008 23743 14048
rect 23783 14008 23792 14048
rect 23734 14007 23792 14008
rect 24075 14048 24117 14057
rect 24075 14008 24076 14048
rect 24116 14008 24117 14048
rect 24075 13999 24117 14008
rect 24363 14048 24405 14057
rect 24363 14008 24364 14048
rect 24404 14008 24405 14048
rect 24363 13999 24405 14008
rect 24544 14048 24586 14057
rect 25707 14048 25749 14057
rect 24544 14008 24545 14048
rect 24585 14008 24586 14048
rect 24544 13999 24586 14008
rect 24843 14039 24885 14048
rect 24843 13999 24844 14039
rect 24884 13999 24885 14039
rect 25707 14008 25708 14048
rect 25748 14008 25749 14048
rect 25707 13999 25749 14008
rect 26571 14048 26613 14057
rect 26571 14008 26572 14048
rect 26612 14008 26613 14048
rect 26571 13999 26613 14008
rect 26763 14048 26805 14057
rect 26763 14008 26764 14048
rect 26804 14008 26805 14048
rect 26763 13999 26805 14008
rect 26955 14048 26997 14057
rect 26955 14008 26956 14048
rect 26996 14008 26997 14048
rect 26955 13999 26997 14008
rect 27514 14048 27572 14049
rect 27514 14008 27523 14048
rect 27563 14008 27572 14048
rect 27514 14007 27572 14008
rect 24843 13990 24885 13999
rect 23242 13965 23300 13966
rect 23110 13964 23168 13965
rect 27147 13964 27189 13973
rect 21042 13915 21043 13955
rect 21083 13915 21088 13955
rect 23110 13924 23119 13964
rect 23159 13924 23168 13964
rect 23110 13923 23168 13924
rect 23634 13955 23680 13964
rect 21042 13906 21088 13915
rect 23634 13915 23635 13955
rect 23675 13915 23680 13955
rect 27147 13924 27148 13964
rect 27188 13924 27189 13964
rect 27147 13915 27189 13924
rect 23634 13906 23680 13915
rect 1035 13880 1077 13889
rect 1035 13840 1036 13880
rect 1076 13840 1077 13880
rect 1035 13831 1077 13840
rect 2091 13880 2133 13889
rect 2091 13840 2092 13880
rect 2132 13840 2133 13880
rect 2091 13831 2133 13840
rect 11403 13880 11445 13889
rect 11403 13840 11404 13880
rect 11444 13840 11445 13880
rect 11403 13831 11445 13840
rect 13131 13880 13173 13889
rect 13131 13840 13132 13880
rect 13172 13840 13173 13880
rect 13131 13831 13173 13840
rect 13498 13880 13556 13881
rect 13498 13840 13507 13880
rect 13547 13840 13556 13880
rect 13498 13839 13556 13840
rect 14475 13880 14517 13889
rect 14475 13840 14476 13880
rect 14516 13840 14517 13880
rect 14475 13831 14517 13840
rect 18507 13880 18549 13889
rect 18507 13840 18508 13880
rect 18548 13840 18549 13880
rect 18507 13831 18549 13840
rect 21195 13880 21237 13889
rect 21195 13840 21196 13880
rect 21236 13840 21237 13880
rect 21195 13831 21237 13840
rect 23019 13880 23061 13889
rect 23019 13840 23020 13880
rect 23060 13840 23061 13880
rect 23019 13831 23061 13840
rect 23787 13880 23829 13889
rect 23787 13840 23788 13880
rect 23828 13840 23829 13880
rect 23787 13831 23829 13840
rect 26763 13880 26805 13889
rect 26763 13840 26764 13880
rect 26804 13840 26805 13880
rect 26763 13831 26805 13840
rect 29643 13880 29685 13889
rect 29643 13840 29644 13880
rect 29684 13840 29685 13880
rect 29643 13831 29685 13840
rect 8139 13796 8181 13805
rect 8139 13756 8140 13796
rect 8180 13756 8181 13796
rect 8139 13747 8181 13756
rect 8794 13796 8852 13797
rect 8794 13756 8803 13796
rect 8843 13756 8852 13796
rect 8794 13755 8852 13756
rect 10251 13796 10293 13805
rect 10251 13756 10252 13796
rect 10292 13756 10293 13796
rect 10251 13747 10293 13756
rect 12507 13796 12549 13805
rect 12507 13756 12508 13796
rect 12548 13756 12549 13796
rect 12507 13747 12549 13756
rect 14266 13796 14324 13797
rect 14266 13756 14275 13796
rect 14315 13756 14324 13796
rect 14266 13755 14324 13756
rect 17451 13796 17493 13805
rect 17451 13756 17452 13796
rect 17492 13756 17493 13796
rect 17451 13747 17493 13756
rect 20619 13796 20661 13805
rect 20619 13756 20620 13796
rect 20660 13756 20661 13796
rect 20619 13747 20661 13756
rect 20907 13796 20949 13805
rect 20907 13756 20908 13796
rect 20948 13756 20949 13796
rect 20907 13747 20949 13756
rect 23499 13796 23541 13805
rect 23499 13756 23500 13796
rect 23540 13756 23541 13796
rect 23499 13747 23541 13756
rect 25035 13796 25077 13805
rect 25035 13756 25036 13796
rect 25076 13756 25077 13796
rect 25035 13747 25077 13756
rect 25899 13796 25941 13805
rect 25899 13756 25900 13796
rect 25940 13756 25941 13796
rect 25899 13747 25941 13756
rect 29067 13796 29109 13805
rect 29067 13756 29068 13796
rect 29108 13756 29109 13796
rect 29067 13747 29109 13756
rect 576 13628 31392 13652
rect 576 13588 3112 13628
rect 3480 13588 10886 13628
rect 11254 13588 18660 13628
rect 19028 13588 26434 13628
rect 26802 13588 31392 13628
rect 576 13564 31392 13588
rect 2554 13460 2612 13461
rect 2554 13420 2563 13460
rect 2603 13420 2612 13460
rect 2554 13419 2612 13420
rect 3819 13460 3861 13469
rect 3819 13420 3820 13460
rect 3860 13420 3861 13460
rect 3819 13411 3861 13420
rect 9130 13460 9188 13461
rect 9130 13420 9139 13460
rect 9179 13420 9188 13460
rect 9130 13419 9188 13420
rect 12346 13460 12404 13461
rect 12346 13420 12355 13460
rect 12395 13420 12404 13460
rect 12346 13419 12404 13420
rect 15723 13460 15765 13469
rect 15723 13420 15724 13460
rect 15764 13420 15765 13460
rect 15723 13411 15765 13420
rect 18394 13460 18452 13461
rect 18394 13420 18403 13460
rect 18443 13420 18452 13460
rect 18394 13419 18452 13420
rect 19083 13460 19125 13469
rect 19083 13420 19084 13460
rect 19124 13420 19125 13460
rect 19083 13411 19125 13420
rect 19467 13460 19509 13469
rect 19467 13420 19468 13460
rect 19508 13420 19509 13460
rect 19467 13411 19509 13420
rect 20235 13460 20277 13469
rect 20235 13420 20236 13460
rect 20276 13420 20277 13460
rect 20235 13411 20277 13420
rect 20890 13460 20948 13461
rect 20890 13420 20899 13460
rect 20939 13420 20948 13460
rect 20890 13419 20948 13420
rect 21754 13460 21812 13461
rect 21754 13420 21763 13460
rect 21803 13420 21812 13460
rect 21754 13419 21812 13420
rect 22827 13460 22869 13469
rect 22827 13420 22828 13460
rect 22868 13420 22869 13460
rect 22827 13411 22869 13420
rect 23403 13460 23445 13469
rect 23403 13420 23404 13460
rect 23444 13420 23445 13460
rect 23403 13411 23445 13420
rect 24027 13460 24069 13469
rect 24027 13420 24028 13460
rect 24068 13420 24069 13460
rect 24027 13411 24069 13420
rect 24651 13460 24693 13469
rect 24651 13420 24652 13460
rect 24692 13420 24693 13460
rect 24651 13411 24693 13420
rect 28779 13460 28821 13469
rect 28779 13420 28780 13460
rect 28820 13420 28821 13460
rect 28779 13411 28821 13420
rect 4762 13376 4820 13377
rect 4762 13336 4771 13376
rect 4811 13336 4820 13376
rect 4762 13335 4820 13336
rect 9370 13376 9428 13377
rect 9370 13336 9379 13376
rect 9419 13336 9428 13376
rect 9370 13335 9428 13336
rect 18123 13376 18165 13385
rect 18123 13336 18124 13376
rect 18164 13336 18165 13376
rect 18123 13327 18165 13336
rect 19851 13376 19893 13385
rect 19851 13336 19852 13376
rect 19892 13336 19893 13376
rect 19851 13327 19893 13336
rect 21195 13376 21237 13385
rect 21195 13336 21196 13376
rect 21236 13336 21237 13376
rect 21195 13327 21237 13336
rect 22347 13376 22389 13385
rect 22347 13336 22348 13376
rect 22388 13336 22389 13376
rect 22347 13327 22389 13336
rect 5338 13292 5396 13293
rect 5338 13252 5347 13292
rect 5387 13252 5396 13292
rect 5338 13251 5396 13252
rect 5547 13292 5589 13301
rect 5547 13252 5548 13292
rect 5588 13252 5589 13292
rect 5818 13292 5876 13293
rect 5547 13243 5589 13252
rect 5691 13250 5733 13259
rect 5818 13252 5827 13292
rect 5867 13252 5876 13292
rect 5818 13251 5876 13252
rect 6298 13292 6356 13293
rect 6298 13252 6307 13292
rect 6347 13252 6356 13292
rect 6298 13251 6356 13252
rect 6507 13292 6549 13301
rect 6507 13252 6508 13292
rect 6548 13252 6549 13292
rect 939 13208 981 13217
rect 939 13168 940 13208
rect 980 13168 981 13208
rect 939 13159 981 13168
rect 2266 13208 2324 13209
rect 2266 13168 2275 13208
rect 2315 13168 2324 13208
rect 2266 13167 2324 13168
rect 2379 13208 2421 13217
rect 2379 13168 2380 13208
rect 2420 13168 2421 13208
rect 2379 13159 2421 13168
rect 2938 13208 2996 13209
rect 2938 13168 2947 13208
rect 2987 13168 2996 13208
rect 2938 13167 2996 13168
rect 3243 13208 3285 13217
rect 3243 13168 3244 13208
rect 3284 13168 3285 13208
rect 3243 13159 3285 13168
rect 3514 13208 3572 13209
rect 3514 13168 3523 13208
rect 3563 13168 3572 13208
rect 3514 13167 3572 13168
rect 3627 13208 3669 13217
rect 3627 13168 3628 13208
rect 3668 13168 3669 13208
rect 3627 13159 3669 13168
rect 4474 13208 4532 13209
rect 4474 13168 4483 13208
rect 4523 13168 4532 13208
rect 4474 13167 4532 13168
rect 4587 13208 4629 13217
rect 4587 13168 4588 13208
rect 4628 13168 4629 13208
rect 4587 13159 4629 13168
rect 5218 13208 5276 13209
rect 5218 13168 5227 13208
rect 5267 13168 5276 13208
rect 5218 13167 5276 13168
rect 5451 13208 5493 13217
rect 5451 13168 5452 13208
rect 5492 13168 5493 13208
rect 5691 13210 5692 13250
rect 5732 13210 5733 13250
rect 6507 13243 6549 13252
rect 7851 13292 7893 13301
rect 7851 13252 7852 13292
rect 7892 13252 7893 13292
rect 7851 13243 7893 13252
rect 10257 13292 10299 13301
rect 10257 13252 10258 13292
rect 10298 13252 10299 13292
rect 9663 13241 9705 13250
rect 10257 13243 10299 13252
rect 10906 13292 10964 13293
rect 10906 13252 10915 13292
rect 10955 13252 10964 13292
rect 10906 13251 10964 13252
rect 13083 13292 13125 13301
rect 13083 13252 13084 13292
rect 13124 13252 13125 13292
rect 13083 13243 13125 13252
rect 13634 13292 13676 13301
rect 13634 13252 13635 13292
rect 13675 13252 13676 13292
rect 13634 13243 13676 13252
rect 17186 13292 17228 13301
rect 17186 13252 17187 13292
rect 17227 13252 17228 13292
rect 17186 13243 17228 13252
rect 25978 13292 26036 13293
rect 25978 13252 25987 13292
rect 26027 13252 26036 13292
rect 25978 13251 26036 13252
rect 17945 13250 18003 13251
rect 28618 13250 28676 13251
rect 5691 13201 5733 13210
rect 5929 13208 5971 13217
rect 5451 13159 5493 13168
rect 5929 13168 5930 13208
rect 5970 13168 5971 13208
rect 5929 13159 5971 13168
rect 6166 13208 6208 13217
rect 6166 13168 6167 13208
rect 6207 13168 6208 13208
rect 6166 13159 6208 13168
rect 6411 13208 6453 13217
rect 6411 13168 6412 13208
rect 6452 13168 6453 13208
rect 6411 13159 6453 13168
rect 6682 13208 6740 13209
rect 6682 13168 6691 13208
rect 6731 13168 6740 13208
rect 6682 13167 6740 13168
rect 6795 13208 6837 13217
rect 6795 13168 6796 13208
rect 6836 13168 6837 13208
rect 6795 13159 6837 13168
rect 7341 13208 7383 13217
rect 7341 13168 7342 13208
rect 7382 13168 7383 13208
rect 7947 13208 7989 13217
rect 7341 13159 7383 13168
rect 7450 13180 7508 13181
rect 7450 13140 7459 13180
rect 7499 13140 7508 13180
rect 7947 13168 7948 13208
rect 7988 13168 7989 13208
rect 7947 13159 7989 13168
rect 8419 13208 8477 13209
rect 8419 13168 8428 13208
rect 8468 13168 8477 13208
rect 8419 13167 8477 13168
rect 8907 13208 8965 13209
rect 8907 13168 8916 13208
rect 8956 13168 8965 13208
rect 9663 13201 9664 13241
rect 9704 13201 9705 13241
rect 17850 13241 17892 13250
rect 9663 13192 9705 13201
rect 9754 13208 9812 13209
rect 8907 13167 8965 13168
rect 9754 13168 9763 13208
rect 9803 13168 9812 13208
rect 9754 13167 9812 13168
rect 10342 13208 10400 13209
rect 10342 13168 10351 13208
rect 10391 13168 10400 13208
rect 10342 13167 10400 13168
rect 10774 13208 10816 13217
rect 10774 13168 10775 13208
rect 10815 13168 10816 13208
rect 10774 13159 10816 13168
rect 11019 13208 11061 13217
rect 11019 13168 11020 13208
rect 11060 13168 11061 13208
rect 11019 13159 11061 13168
rect 11695 13208 11753 13209
rect 11695 13168 11704 13208
rect 11744 13168 11753 13208
rect 11695 13167 11753 13168
rect 12205 13208 12263 13209
rect 12205 13168 12214 13208
rect 12254 13168 12263 13208
rect 12205 13167 12263 13168
rect 12643 13208 12701 13209
rect 12643 13168 12652 13208
rect 12692 13168 12701 13208
rect 12643 13167 12701 13168
rect 12919 13208 12977 13209
rect 12919 13168 12928 13208
rect 12968 13168 12977 13208
rect 12919 13167 12977 13168
rect 13515 13208 13557 13217
rect 13515 13168 13516 13208
rect 13556 13168 13557 13208
rect 13515 13159 13557 13168
rect 13744 13208 13802 13209
rect 13744 13168 13753 13208
rect 13793 13168 13802 13208
rect 13744 13167 13802 13168
rect 14187 13208 14229 13217
rect 14187 13168 14188 13208
rect 14228 13168 14229 13208
rect 14187 13159 14229 13168
rect 14306 13208 14348 13217
rect 14306 13168 14307 13208
rect 14347 13168 14348 13208
rect 14306 13159 14348 13168
rect 14416 13208 14474 13209
rect 14416 13168 14425 13208
rect 14465 13168 14474 13208
rect 14416 13167 14474 13168
rect 14710 13208 14752 13217
rect 14710 13168 14711 13208
rect 14751 13168 14752 13208
rect 14710 13159 14752 13168
rect 14842 13208 14900 13209
rect 14842 13168 14851 13208
rect 14891 13168 14900 13208
rect 14842 13167 14900 13168
rect 14955 13208 14997 13217
rect 14955 13168 14956 13208
rect 14996 13168 14997 13208
rect 14955 13159 14997 13168
rect 15226 13208 15284 13209
rect 15226 13168 15235 13208
rect 15275 13168 15284 13208
rect 15226 13167 15284 13168
rect 15545 13208 15587 13217
rect 16395 13208 16437 13217
rect 15545 13168 15546 13208
rect 15586 13168 15587 13208
rect 15545 13159 15587 13168
rect 16107 13199 16149 13208
rect 16107 13159 16108 13199
rect 16148 13159 16149 13199
rect 16395 13168 16396 13208
rect 16436 13168 16437 13208
rect 16395 13159 16437 13168
rect 17067 13208 17109 13217
rect 17067 13168 17068 13208
rect 17108 13168 17109 13208
rect 17067 13159 17109 13168
rect 17296 13208 17354 13209
rect 17296 13168 17305 13208
rect 17345 13168 17354 13208
rect 17296 13167 17354 13168
rect 17731 13208 17789 13209
rect 17731 13168 17740 13208
rect 17780 13168 17789 13208
rect 17850 13201 17851 13241
rect 17891 13201 17892 13241
rect 17945 13210 17954 13250
rect 17994 13210 18003 13250
rect 21089 13241 21131 13250
rect 17945 13209 18003 13210
rect 17850 13192 17892 13201
rect 18795 13208 18837 13217
rect 17731 13167 17789 13168
rect 18795 13168 18796 13208
rect 18836 13168 18837 13208
rect 18795 13159 18837 13168
rect 19083 13208 19125 13217
rect 19083 13168 19084 13208
rect 19124 13168 19125 13208
rect 19083 13159 19125 13168
rect 19275 13208 19317 13217
rect 19275 13168 19276 13208
rect 19316 13168 19317 13208
rect 19275 13159 19317 13168
rect 19467 13208 19509 13217
rect 19467 13168 19468 13208
rect 19508 13168 19509 13208
rect 19467 13159 19509 13168
rect 19659 13208 19701 13217
rect 19659 13168 19660 13208
rect 19700 13168 19701 13208
rect 19659 13159 19701 13168
rect 19851 13208 19893 13217
rect 19851 13168 19852 13208
rect 19892 13168 19893 13208
rect 19851 13159 19893 13168
rect 20043 13208 20085 13217
rect 20043 13168 20044 13208
rect 20084 13168 20085 13208
rect 20043 13159 20085 13168
rect 20235 13208 20277 13217
rect 20235 13168 20236 13208
rect 20276 13168 20277 13208
rect 20235 13159 20277 13168
rect 20523 13208 20565 13217
rect 20523 13168 20524 13208
rect 20564 13168 20565 13208
rect 20523 13159 20565 13168
rect 20715 13208 20757 13217
rect 20715 13168 20716 13208
rect 20756 13168 20757 13208
rect 20715 13159 20757 13168
rect 20906 13208 20948 13217
rect 20906 13168 20907 13208
rect 20947 13168 20948 13208
rect 21089 13201 21090 13241
rect 21130 13201 21131 13241
rect 23739 13241 23781 13250
rect 21089 13192 21131 13201
rect 21271 13208 21313 13217
rect 20906 13159 20948 13168
rect 21271 13168 21272 13208
rect 21312 13168 21313 13208
rect 21271 13159 21313 13168
rect 21387 13208 21429 13217
rect 21387 13168 21388 13208
rect 21428 13168 21429 13208
rect 21387 13159 21429 13168
rect 21574 13208 21616 13217
rect 21574 13168 21575 13208
rect 21615 13168 21616 13208
rect 21574 13159 21616 13168
rect 21770 13208 21812 13217
rect 21770 13168 21771 13208
rect 21811 13168 21812 13208
rect 21770 13159 21812 13168
rect 21994 13208 22052 13209
rect 21994 13168 22003 13208
rect 22043 13168 22052 13208
rect 21994 13167 22052 13168
rect 22251 13208 22293 13217
rect 22251 13168 22252 13208
rect 22292 13168 22293 13208
rect 22251 13159 22293 13168
rect 22378 13208 22436 13209
rect 22378 13168 22387 13208
rect 22427 13168 22436 13208
rect 22378 13167 22436 13168
rect 22492 13208 22550 13209
rect 22492 13168 22501 13208
rect 22541 13168 22550 13208
rect 22492 13167 22550 13168
rect 22731 13208 22773 13217
rect 22731 13168 22732 13208
rect 22772 13168 22773 13208
rect 22731 13159 22773 13168
rect 22916 13205 22958 13214
rect 22916 13165 22917 13205
rect 22957 13165 22958 13205
rect 23098 13208 23156 13209
rect 23098 13168 23107 13208
rect 23147 13168 23156 13208
rect 23098 13167 23156 13168
rect 23595 13208 23637 13217
rect 23595 13168 23596 13208
rect 23636 13168 23637 13208
rect 23739 13201 23740 13241
rect 23780 13201 23781 13241
rect 23739 13192 23781 13201
rect 24171 13208 24213 13217
rect 16107 13150 16149 13159
rect 22916 13156 22958 13165
rect 23595 13159 23637 13168
rect 24171 13168 24172 13208
rect 24212 13168 24213 13208
rect 24171 13159 24213 13168
rect 24363 13208 24405 13217
rect 24363 13168 24364 13208
rect 24404 13168 24405 13208
rect 24363 13159 24405 13168
rect 24538 13208 24596 13209
rect 24538 13168 24547 13208
rect 24587 13168 24596 13208
rect 24538 13167 24596 13168
rect 24651 13208 24693 13217
rect 24651 13168 24652 13208
rect 24692 13168 24693 13208
rect 24651 13159 24693 13168
rect 25018 13208 25076 13209
rect 25018 13168 25027 13208
rect 25067 13168 25076 13208
rect 25018 13167 25076 13168
rect 25131 13208 25173 13217
rect 28618 13210 28627 13250
rect 28667 13210 28676 13250
rect 28618 13209 28676 13210
rect 25131 13168 25132 13208
rect 25172 13168 25173 13208
rect 25131 13159 25173 13168
rect 27514 13208 27572 13209
rect 27514 13168 27523 13208
rect 27563 13168 27572 13208
rect 27514 13167 27572 13168
rect 28779 13208 28821 13217
rect 28779 13168 28780 13208
rect 28820 13168 28821 13208
rect 28779 13159 28821 13168
rect 28971 13208 29013 13217
rect 28971 13168 28972 13208
rect 29012 13168 29013 13208
rect 28971 13159 29013 13168
rect 7450 13139 7508 13140
rect 3147 13124 3189 13133
rect 3147 13084 3148 13124
rect 3188 13084 3189 13124
rect 3147 13075 3189 13084
rect 3830 13124 3872 13133
rect 3830 13084 3831 13124
rect 3871 13084 3872 13124
rect 3830 13075 3872 13084
rect 7001 13124 7043 13133
rect 7001 13084 7002 13124
rect 7042 13084 7043 13124
rect 7001 13075 7043 13084
rect 11098 13124 11156 13125
rect 11098 13084 11107 13124
rect 11147 13084 11156 13124
rect 11098 13083 11156 13084
rect 11530 13124 11588 13125
rect 11530 13084 11539 13124
rect 11579 13084 11588 13124
rect 11530 13083 11588 13084
rect 12352 13124 12394 13133
rect 12352 13084 12353 13124
rect 12393 13084 12394 13124
rect 12352 13075 12394 13084
rect 13419 13124 13461 13133
rect 13419 13084 13420 13124
rect 13460 13084 13461 13124
rect 13419 13075 13461 13084
rect 15034 13124 15092 13125
rect 15034 13084 15043 13124
rect 15083 13084 15092 13124
rect 15034 13083 15092 13084
rect 16011 13124 16053 13133
rect 16011 13084 16012 13124
rect 16052 13084 16053 13124
rect 16011 13075 16053 13084
rect 16971 13124 17013 13133
rect 16971 13084 16972 13124
rect 17012 13084 17013 13124
rect 16971 13075 17013 13084
rect 23211 13124 23253 13133
rect 23211 13084 23212 13124
rect 23252 13084 23253 13124
rect 23211 13075 23253 13084
rect 23417 13124 23459 13133
rect 23417 13084 23418 13124
rect 23458 13084 23459 13124
rect 23417 13075 23459 13084
rect 23931 13124 23973 13133
rect 23931 13084 23932 13124
rect 23972 13084 23973 13124
rect 23931 13075 23973 13084
rect 25594 13124 25652 13125
rect 25594 13084 25603 13124
rect 25643 13084 25652 13124
rect 25594 13083 25652 13084
rect 27898 13124 27956 13125
rect 27898 13084 27907 13124
rect 27947 13084 27956 13124
rect 27898 13083 27956 13084
rect 1611 13040 1653 13049
rect 1611 13000 1612 13040
rect 1652 13000 1653 13040
rect 1611 12991 1653 13000
rect 6010 13040 6068 13041
rect 6010 13000 6019 13040
rect 6059 13000 6068 13040
rect 6010 12999 6068 13000
rect 6891 13040 6933 13049
rect 6891 13000 6892 13040
rect 6932 13000 6933 13040
rect 6891 12991 6933 13000
rect 10042 13040 10100 13041
rect 10042 13000 10051 13040
rect 10091 13000 10100 13040
rect 10042 12999 10100 13000
rect 12010 13040 12068 13041
rect 12010 13000 12019 13040
rect 12059 13000 12068 13040
rect 12010 12999 12068 13000
rect 12555 13040 12597 13049
rect 12555 13000 12556 13040
rect 12596 13000 12597 13040
rect 9898 12998 9956 12999
rect 9898 12958 9907 12998
rect 9947 12958 9956 12998
rect 12555 12991 12597 13000
rect 14091 13040 14133 13049
rect 14091 13000 14092 13040
rect 14132 13000 14133 13040
rect 14091 12991 14133 13000
rect 15322 13040 15380 13041
rect 15322 13000 15331 13040
rect 15371 13000 15380 13040
rect 15322 12999 15380 13000
rect 15435 13040 15477 13049
rect 15435 13000 15436 13040
rect 15476 13000 15477 13040
rect 15435 12991 15477 13000
rect 22107 13040 22149 13049
rect 22107 13000 22108 13040
rect 22148 13000 22149 13040
rect 22107 12991 22149 13000
rect 25419 13040 25461 13049
rect 25419 13000 25420 13040
rect 25460 13000 25461 13040
rect 25419 12991 25461 13000
rect 28426 13040 28484 13041
rect 28426 13000 28435 13040
rect 28475 13000 28484 13040
rect 28426 12999 28484 13000
rect 9898 12957 9956 12958
rect 576 12872 31392 12896
rect 576 12832 4352 12872
rect 4720 12832 12126 12872
rect 12494 12832 19900 12872
rect 20268 12832 27674 12872
rect 28042 12832 31392 12872
rect 576 12808 31392 12832
rect 826 12704 884 12705
rect 826 12664 835 12704
rect 875 12664 884 12704
rect 826 12663 884 12664
rect 1803 12704 1845 12713
rect 1803 12664 1804 12704
rect 1844 12664 1845 12704
rect 1803 12655 1845 12664
rect 2026 12704 2084 12705
rect 2026 12664 2035 12704
rect 2075 12664 2084 12704
rect 2026 12663 2084 12664
rect 3034 12704 3092 12705
rect 3034 12664 3043 12704
rect 3083 12664 3092 12704
rect 3034 12663 3092 12664
rect 3562 12704 3620 12705
rect 3562 12664 3571 12704
rect 3611 12664 3620 12704
rect 3562 12663 3620 12664
rect 4587 12704 4629 12713
rect 4587 12664 4588 12704
rect 4628 12664 4629 12704
rect 4587 12655 4629 12664
rect 6027 12704 6069 12713
rect 6027 12664 6028 12704
rect 6068 12664 6069 12704
rect 6027 12655 6069 12664
rect 6298 12704 6356 12705
rect 6298 12664 6307 12704
rect 6347 12664 6356 12704
rect 6298 12663 6356 12664
rect 6411 12704 6453 12713
rect 6411 12664 6412 12704
rect 6452 12664 6453 12704
rect 6411 12655 6453 12664
rect 9274 12704 9332 12705
rect 9274 12664 9283 12704
rect 9323 12664 9332 12704
rect 9274 12663 9332 12664
rect 9754 12704 9812 12705
rect 9754 12664 9763 12704
rect 9803 12664 9812 12704
rect 9754 12663 9812 12664
rect 10858 12704 10916 12705
rect 10858 12664 10867 12704
rect 10907 12664 10916 12704
rect 10858 12663 10916 12664
rect 11403 12704 11445 12713
rect 11403 12664 11404 12704
rect 11444 12664 11445 12704
rect 11403 12655 11445 12664
rect 13419 12704 13461 12713
rect 13419 12664 13420 12704
rect 13460 12664 13461 12704
rect 13419 12655 13461 12664
rect 15082 12704 15140 12705
rect 15082 12664 15091 12704
rect 15131 12664 15140 12704
rect 15082 12663 15140 12664
rect 16011 12704 16053 12713
rect 16011 12664 16012 12704
rect 16052 12664 16053 12704
rect 16011 12655 16053 12664
rect 16282 12704 16340 12705
rect 16282 12664 16291 12704
rect 16331 12664 16340 12704
rect 16282 12663 16340 12664
rect 16875 12704 16917 12713
rect 16875 12664 16876 12704
rect 16916 12664 16917 12704
rect 16875 12655 16917 12664
rect 17643 12704 17685 12713
rect 17643 12664 17644 12704
rect 17684 12664 17685 12704
rect 17643 12655 17685 12664
rect 18202 12704 18260 12705
rect 18202 12664 18211 12704
rect 18251 12664 18260 12704
rect 18202 12663 18260 12664
rect 19066 12704 19124 12705
rect 19066 12664 19075 12704
rect 19115 12664 19124 12704
rect 19066 12663 19124 12664
rect 20602 12704 20660 12705
rect 20602 12664 20611 12704
rect 20651 12664 20660 12704
rect 20602 12663 20660 12664
rect 21099 12704 21141 12713
rect 21099 12664 21100 12704
rect 21140 12664 21141 12704
rect 21099 12655 21141 12664
rect 23787 12704 23829 12713
rect 23787 12664 23788 12704
rect 23828 12664 23829 12704
rect 23787 12655 23829 12664
rect 24939 12704 24981 12713
rect 24939 12664 24940 12704
rect 24980 12664 24981 12704
rect 24939 12655 24981 12664
rect 25498 12704 25556 12705
rect 25498 12664 25507 12704
rect 25547 12664 25556 12704
rect 25498 12663 25556 12664
rect 26859 12704 26901 12713
rect 26859 12664 26860 12704
rect 26900 12664 26901 12704
rect 26859 12655 26901 12664
rect 28203 12704 28245 12713
rect 28203 12664 28204 12704
rect 28244 12664 28245 12704
rect 28203 12655 28245 12664
rect 6688 12620 6730 12629
rect 6688 12580 6689 12620
rect 6729 12580 6730 12620
rect 6688 12571 6730 12580
rect 8331 12620 8373 12629
rect 8331 12580 8332 12620
rect 8372 12580 8373 12620
rect 8331 12571 8373 12580
rect 8715 12620 8757 12629
rect 8715 12580 8716 12620
rect 8756 12580 8757 12620
rect 8715 12571 8757 12580
rect 11200 12620 11242 12629
rect 11200 12580 11201 12620
rect 11241 12580 11242 12620
rect 11200 12571 11242 12580
rect 11962 12620 12020 12621
rect 16189 12620 16231 12629
rect 11962 12580 11971 12620
rect 12011 12580 12020 12620
rect 11962 12579 12020 12580
rect 14178 12611 14224 12620
rect 14178 12571 14179 12611
rect 14219 12571 14224 12611
rect 16189 12580 16190 12620
rect 16230 12580 16231 12620
rect 16189 12571 16231 12580
rect 16395 12620 16437 12629
rect 16395 12580 16396 12620
rect 16436 12580 16437 12620
rect 16395 12571 16437 12580
rect 17437 12620 17479 12629
rect 17437 12580 17438 12620
rect 17478 12580 17479 12620
rect 17437 12571 17479 12580
rect 21466 12620 21524 12621
rect 21466 12580 21475 12620
rect 21515 12580 21524 12620
rect 21466 12579 21524 12580
rect 26966 12620 27008 12629
rect 26966 12580 26967 12620
rect 27007 12580 27008 12620
rect 26966 12571 27008 12580
rect 27613 12620 27655 12629
rect 27613 12580 27614 12620
rect 27654 12580 27655 12620
rect 27613 12571 27655 12580
rect 14178 12562 14224 12571
rect 939 12536 981 12545
rect 939 12496 940 12536
rect 980 12496 981 12536
rect 939 12487 981 12496
rect 1323 12536 1365 12545
rect 1323 12496 1324 12536
rect 1364 12496 1365 12536
rect 1323 12487 1365 12496
rect 1707 12536 1749 12545
rect 1707 12496 1708 12536
rect 1748 12496 1749 12536
rect 1707 12487 1749 12496
rect 2170 12536 2228 12537
rect 2722 12536 2780 12537
rect 2170 12496 2179 12536
rect 2219 12496 2228 12536
rect 2170 12495 2228 12496
rect 2283 12527 2325 12536
rect 2283 12487 2284 12527
rect 2324 12487 2325 12527
rect 2722 12496 2731 12536
rect 2771 12496 2780 12536
rect 2722 12495 2780 12496
rect 2955 12536 2997 12545
rect 2955 12496 2956 12536
rect 2996 12496 2997 12536
rect 2955 12487 2997 12496
rect 3757 12536 3815 12537
rect 3757 12496 3766 12536
rect 3806 12496 3815 12536
rect 3757 12495 3815 12496
rect 4186 12536 4244 12537
rect 4186 12496 4195 12536
rect 4235 12496 4244 12536
rect 4186 12495 4244 12496
rect 4299 12536 4341 12545
rect 4299 12496 4300 12536
rect 4340 12496 4341 12536
rect 4299 12487 4341 12496
rect 4738 12536 4796 12537
rect 4738 12496 4747 12536
rect 4787 12496 4796 12536
rect 4738 12495 4796 12496
rect 4971 12536 5013 12545
rect 4971 12496 4972 12536
rect 5012 12496 5013 12536
rect 4971 12487 5013 12496
rect 5626 12536 5684 12537
rect 5626 12496 5635 12536
rect 5675 12496 5684 12536
rect 5626 12495 5684 12496
rect 5739 12536 5781 12545
rect 5739 12496 5740 12536
rect 5780 12496 5781 12536
rect 5739 12487 5781 12496
rect 6208 12536 6250 12545
rect 6891 12536 6933 12545
rect 7179 12536 7221 12545
rect 6208 12496 6209 12536
rect 6249 12496 6250 12536
rect 6208 12487 6250 12496
rect 6507 12527 6549 12536
rect 6507 12487 6508 12527
rect 6548 12487 6549 12527
rect 6891 12496 6892 12536
rect 6932 12496 6933 12536
rect 6891 12487 6933 12496
rect 6987 12527 7029 12536
rect 6987 12487 6988 12527
rect 7028 12487 7029 12527
rect 7179 12496 7180 12536
rect 7220 12496 7221 12536
rect 7179 12487 7221 12496
rect 7366 12536 7424 12537
rect 7366 12496 7375 12536
rect 7415 12496 7424 12536
rect 7366 12495 7424 12496
rect 7851 12536 7893 12545
rect 7851 12496 7852 12536
rect 7892 12496 7893 12536
rect 7851 12487 7893 12496
rect 8041 12536 8083 12545
rect 8041 12496 8042 12536
rect 8082 12496 8083 12536
rect 8041 12487 8083 12496
rect 8235 12536 8277 12545
rect 8235 12496 8236 12536
rect 8276 12496 8277 12536
rect 8235 12487 8277 12496
rect 8427 12536 8469 12545
rect 8427 12496 8428 12536
rect 8468 12496 8469 12536
rect 8427 12487 8469 12496
rect 8608 12536 8650 12545
rect 8608 12496 8609 12536
rect 8649 12496 8650 12536
rect 8608 12487 8650 12496
rect 8811 12536 8853 12545
rect 8811 12496 8812 12536
rect 8852 12496 8853 12536
rect 8811 12487 8853 12496
rect 9003 12536 9045 12545
rect 9003 12496 9004 12536
rect 9044 12496 9045 12536
rect 9003 12487 9045 12496
rect 9435 12536 9493 12537
rect 9435 12496 9444 12536
rect 9484 12496 9493 12536
rect 9435 12495 9493 12496
rect 9579 12536 9621 12545
rect 9579 12496 9580 12536
rect 9620 12496 9621 12536
rect 9579 12487 9621 12496
rect 9915 12536 9957 12545
rect 9915 12496 9916 12536
rect 9956 12496 9957 12536
rect 9915 12487 9957 12496
rect 10059 12536 10101 12545
rect 10059 12496 10060 12536
rect 10100 12496 10101 12536
rect 10059 12487 10101 12496
rect 11053 12536 11111 12537
rect 12171 12536 12213 12545
rect 11053 12496 11062 12536
rect 11102 12496 11111 12536
rect 11053 12495 11111 12496
rect 11499 12527 11541 12536
rect 11499 12487 11500 12527
rect 11540 12487 11541 12527
rect 12171 12496 12172 12536
rect 12212 12496 12213 12536
rect 12171 12487 12213 12496
rect 12730 12536 12788 12537
rect 12730 12496 12739 12536
rect 12779 12496 12788 12536
rect 12730 12495 12788 12496
rect 12837 12536 12895 12537
rect 12837 12496 12846 12536
rect 12886 12496 12895 12536
rect 12837 12495 12895 12496
rect 13515 12536 13557 12545
rect 13515 12496 13516 12536
rect 13556 12496 13557 12536
rect 13515 12487 13557 12496
rect 13744 12536 13802 12537
rect 13744 12496 13753 12536
rect 13793 12496 13802 12536
rect 13744 12495 13802 12496
rect 13882 12536 13940 12537
rect 14266 12536 14324 12537
rect 13882 12496 13891 12536
rect 13931 12496 13940 12536
rect 13882 12495 13940 12496
rect 13995 12527 14037 12536
rect 13995 12487 13996 12527
rect 14036 12487 14037 12527
rect 14266 12496 14275 12536
rect 14315 12496 14324 12536
rect 15277 12536 15335 12537
rect 14266 12495 14324 12496
rect 14443 12525 14501 12526
rect 2283 12478 2325 12487
rect 6507 12478 6549 12487
rect 6987 12478 7029 12487
rect 11499 12478 11541 12487
rect 13995 12478 14037 12487
rect 14443 12485 14452 12525
rect 14492 12485 14501 12525
rect 15277 12496 15286 12536
rect 15326 12496 15335 12536
rect 15277 12495 15335 12496
rect 15610 12536 15668 12537
rect 15610 12496 15619 12536
rect 15659 12496 15668 12536
rect 15610 12495 15668 12496
rect 15723 12536 15765 12545
rect 16971 12536 17013 12545
rect 15723 12496 15724 12536
rect 15764 12496 15765 12536
rect 15723 12487 15765 12496
rect 16491 12527 16533 12536
rect 16491 12487 16492 12527
rect 16532 12487 16533 12527
rect 16971 12496 16972 12536
rect 17012 12496 17013 12536
rect 16971 12487 17013 12496
rect 17200 12536 17258 12537
rect 18507 12536 18549 12545
rect 17200 12496 17209 12536
rect 17249 12496 17258 12536
rect 17200 12495 17258 12496
rect 17739 12527 17781 12536
rect 17739 12487 17740 12527
rect 17780 12487 17781 12527
rect 18507 12496 18508 12536
rect 18548 12496 18549 12536
rect 18507 12487 18549 12496
rect 19275 12536 19317 12545
rect 19275 12496 19276 12536
rect 19316 12496 19317 12536
rect 19275 12487 19317 12496
rect 19563 12536 19605 12545
rect 19563 12496 19564 12536
rect 19604 12496 19605 12536
rect 19563 12487 19605 12496
rect 19755 12536 19797 12545
rect 19755 12496 19756 12536
rect 19796 12496 19797 12536
rect 19755 12487 19797 12496
rect 20139 12536 20181 12545
rect 20139 12496 20140 12536
rect 20180 12496 20181 12536
rect 20139 12487 20181 12496
rect 20331 12536 20373 12545
rect 20331 12496 20332 12536
rect 20372 12496 20373 12536
rect 20331 12487 20373 12496
rect 20715 12536 20757 12545
rect 20715 12496 20716 12536
rect 20756 12496 20757 12536
rect 20715 12487 20757 12496
rect 21099 12536 21141 12545
rect 21099 12496 21100 12536
rect 21140 12496 21141 12536
rect 21099 12487 21141 12496
rect 21291 12536 21333 12545
rect 21291 12496 21292 12536
rect 21332 12496 21333 12536
rect 21291 12487 21333 12496
rect 21850 12536 21908 12537
rect 21850 12496 21859 12536
rect 21899 12496 21908 12536
rect 21850 12495 21908 12496
rect 24651 12536 24693 12545
rect 24651 12496 24652 12536
rect 24692 12496 24693 12536
rect 24651 12487 24693 12496
rect 24939 12536 24981 12545
rect 24939 12496 24940 12536
rect 24980 12496 24981 12536
rect 24939 12487 24981 12496
rect 25129 12536 25171 12545
rect 25129 12496 25130 12536
rect 25170 12496 25171 12536
rect 25129 12487 25171 12496
rect 25402 12536 25460 12537
rect 25402 12496 25411 12536
rect 25451 12496 25460 12536
rect 25402 12495 25460 12496
rect 25718 12536 25760 12545
rect 26043 12536 26085 12545
rect 25718 12496 25719 12536
rect 25759 12496 25760 12536
rect 25718 12487 25760 12496
rect 25890 12527 25936 12536
rect 25890 12487 25891 12527
rect 25931 12487 25936 12527
rect 26043 12496 26044 12536
rect 26084 12496 26085 12536
rect 26043 12487 26085 12496
rect 26650 12536 26708 12537
rect 26650 12496 26659 12536
rect 26699 12496 26708 12536
rect 26650 12495 26708 12496
rect 26763 12536 26805 12545
rect 26763 12496 26764 12536
rect 26804 12496 26805 12536
rect 26763 12487 26805 12496
rect 27094 12536 27136 12545
rect 27094 12496 27095 12536
rect 27135 12496 27136 12536
rect 27094 12487 27136 12496
rect 27339 12536 27381 12545
rect 27339 12496 27340 12536
rect 27380 12496 27381 12536
rect 27339 12487 27381 12496
rect 27819 12536 27861 12545
rect 28107 12536 28149 12545
rect 27819 12496 27820 12536
rect 27860 12496 27861 12536
rect 27819 12487 27861 12496
rect 27915 12527 27957 12536
rect 27915 12487 27916 12527
rect 27956 12487 27957 12527
rect 28107 12496 28108 12536
rect 28148 12496 28149 12536
rect 28107 12487 28149 12496
rect 28280 12536 28322 12545
rect 28280 12496 28281 12536
rect 28321 12496 28322 12536
rect 28280 12487 28322 12496
rect 14443 12484 14501 12485
rect 16491 12478 16533 12487
rect 17739 12478 17781 12487
rect 25890 12478 25936 12487
rect 27915 12478 27957 12487
rect 2842 12452 2900 12453
rect 2842 12412 2851 12452
rect 2891 12412 2900 12452
rect 2842 12411 2900 12412
rect 4858 12452 4916 12453
rect 4858 12412 4867 12452
rect 4907 12412 4916 12452
rect 4858 12411 4916 12412
rect 5067 12452 5109 12461
rect 17090 12452 17132 12461
rect 5067 12412 5068 12452
rect 5108 12412 5109 12452
rect 5067 12403 5109 12412
rect 13650 12443 13696 12452
rect 13650 12403 13651 12443
rect 13691 12403 13696 12443
rect 17090 12412 17091 12452
rect 17131 12412 17132 12452
rect 17090 12403 17132 12412
rect 18417 12452 18459 12461
rect 18417 12412 18418 12452
rect 18458 12412 18459 12452
rect 18417 12403 18459 12412
rect 23403 12452 23445 12461
rect 23403 12412 23404 12452
rect 23444 12412 23445 12452
rect 23403 12403 23445 12412
rect 27220 12452 27262 12461
rect 27220 12412 27221 12452
rect 27261 12412 27262 12452
rect 27220 12403 27262 12412
rect 27435 12452 27477 12461
rect 27435 12412 27436 12452
rect 27476 12412 27477 12452
rect 27435 12403 27477 12412
rect 13650 12394 13696 12403
rect 1131 12368 1173 12377
rect 1131 12328 1132 12368
rect 1172 12328 1173 12368
rect 1131 12319 1173 12328
rect 2571 12368 2613 12377
rect 2571 12328 2572 12368
rect 2612 12328 2613 12368
rect 2571 12319 2613 12328
rect 7275 12368 7317 12377
rect 7275 12328 7276 12368
rect 7316 12328 7317 12368
rect 7275 12319 7317 12328
rect 21195 12368 21237 12377
rect 21195 12328 21196 12368
rect 21236 12328 21237 12368
rect 21195 12319 21237 12328
rect 28491 12368 28533 12377
rect 28491 12328 28492 12368
rect 28532 12328 28533 12368
rect 28491 12319 28533 12328
rect 28875 12368 28917 12377
rect 28875 12328 28876 12368
rect 28916 12328 28917 12368
rect 28875 12319 28917 12328
rect 6682 12284 6740 12285
rect 6682 12244 6691 12284
rect 6731 12244 6740 12284
rect 6682 12243 6740 12244
rect 7851 12284 7893 12293
rect 7851 12244 7852 12284
rect 7892 12244 7893 12284
rect 7851 12235 7893 12244
rect 9147 12284 9189 12293
rect 9147 12244 9148 12284
rect 9188 12244 9189 12284
rect 9147 12235 9189 12244
rect 11194 12284 11252 12285
rect 11194 12244 11203 12284
rect 11243 12244 11252 12284
rect 11194 12243 11252 12244
rect 13018 12284 13076 12285
rect 13018 12244 13027 12284
rect 13067 12244 13076 12284
rect 13018 12243 13076 12244
rect 13882 12284 13940 12285
rect 13882 12244 13891 12284
rect 13931 12244 13940 12284
rect 13882 12243 13940 12244
rect 17434 12284 17492 12285
rect 17434 12244 17443 12284
rect 17483 12244 17492 12284
rect 17434 12243 17492 12244
rect 19851 12284 19893 12293
rect 19851 12244 19852 12284
rect 19892 12244 19893 12284
rect 19851 12235 19893 12244
rect 20139 12284 20181 12293
rect 20139 12244 20140 12284
rect 20180 12244 20181 12284
rect 20139 12235 20181 12244
rect 20907 12284 20949 12293
rect 20907 12244 20908 12284
rect 20948 12244 20949 12284
rect 20907 12235 20949 12244
rect 23979 12284 24021 12293
rect 23979 12244 23980 12284
rect 24020 12244 24021 12284
rect 23979 12235 24021 12244
rect 25707 12284 25749 12293
rect 25707 12244 25708 12284
rect 25748 12244 25749 12284
rect 25707 12235 25749 12244
rect 27610 12284 27668 12285
rect 27610 12244 27619 12284
rect 27659 12244 27668 12284
rect 27610 12243 27668 12244
rect 576 12116 31392 12140
rect 576 12076 3112 12116
rect 3480 12076 10886 12116
rect 11254 12076 18660 12116
rect 19028 12076 26434 12116
rect 26802 12076 31392 12116
rect 576 12052 31392 12076
rect 3339 11948 3381 11957
rect 3339 11908 3340 11948
rect 3380 11908 3381 11948
rect 3339 11899 3381 11908
rect 6874 11948 6932 11949
rect 6874 11908 6883 11948
rect 6923 11908 6932 11948
rect 6874 11907 6932 11908
rect 8331 11948 8373 11957
rect 8331 11908 8332 11948
rect 8372 11908 8373 11948
rect 8331 11899 8373 11908
rect 10443 11948 10485 11957
rect 10443 11908 10444 11948
rect 10484 11908 10485 11948
rect 10443 11899 10485 11908
rect 12747 11948 12789 11957
rect 12747 11908 12748 11948
rect 12788 11908 12789 11948
rect 12747 11899 12789 11908
rect 13995 11948 14037 11957
rect 13995 11908 13996 11948
rect 14036 11908 14037 11948
rect 13995 11899 14037 11908
rect 14763 11948 14805 11957
rect 14763 11908 14764 11948
rect 14804 11908 14805 11948
rect 14763 11899 14805 11908
rect 15723 11948 15765 11957
rect 15723 11908 15724 11948
rect 15764 11908 15765 11948
rect 15723 11899 15765 11908
rect 17434 11948 17492 11949
rect 17434 11908 17443 11948
rect 17483 11908 17492 11948
rect 17434 11907 17492 11908
rect 19371 11948 19413 11957
rect 19371 11908 19372 11948
rect 19412 11908 19413 11948
rect 19371 11899 19413 11908
rect 22731 11948 22773 11957
rect 22731 11908 22732 11948
rect 22772 11908 22773 11948
rect 22731 11899 22773 11908
rect 24075 11948 24117 11957
rect 24075 11908 24076 11948
rect 24116 11908 24117 11948
rect 24075 11899 24117 11908
rect 25515 11948 25557 11957
rect 25515 11908 25516 11948
rect 25556 11908 25557 11948
rect 25515 11899 25557 11908
rect 27627 11864 27669 11873
rect 16459 11855 16501 11864
rect 16459 11815 16460 11855
rect 16500 11815 16501 11855
rect 27627 11824 27628 11864
rect 27668 11824 27669 11864
rect 27627 11815 27669 11824
rect 28107 11864 28149 11873
rect 28107 11824 28108 11864
rect 28148 11824 28149 11864
rect 28107 11815 28149 11824
rect 16459 11806 16501 11815
rect 970 11780 1028 11781
rect 970 11740 979 11780
rect 1019 11740 1028 11780
rect 970 11739 1028 11740
rect 2379 11780 2421 11789
rect 2379 11740 2380 11780
rect 2420 11740 2421 11780
rect 2379 11731 2421 11740
rect 3610 11780 3668 11781
rect 3610 11740 3619 11780
rect 3659 11740 3668 11780
rect 3610 11739 3668 11740
rect 3819 11780 3861 11789
rect 3819 11740 3820 11780
rect 3860 11740 3861 11780
rect 2890 11738 2948 11739
rect 1165 11696 1223 11697
rect 1165 11656 1174 11696
rect 1214 11656 1223 11696
rect 1165 11655 1223 11656
rect 1498 11696 1556 11697
rect 1498 11656 1507 11696
rect 1547 11656 1556 11696
rect 1498 11655 1556 11656
rect 1611 11696 1653 11705
rect 1611 11656 1612 11696
rect 1652 11656 1653 11696
rect 1611 11647 1653 11656
rect 2038 11696 2080 11705
rect 2038 11656 2039 11696
rect 2079 11656 2080 11696
rect 2038 11647 2080 11656
rect 2170 11696 2228 11697
rect 2170 11656 2179 11696
rect 2219 11656 2228 11696
rect 2170 11655 2228 11656
rect 2283 11696 2325 11705
rect 2890 11698 2899 11738
rect 2939 11698 2948 11738
rect 3819 11731 3861 11740
rect 6219 11780 6261 11789
rect 6897 11780 6939 11789
rect 6219 11740 6220 11780
rect 6260 11740 6261 11780
rect 6219 11731 6261 11740
rect 6450 11771 6496 11780
rect 6450 11731 6451 11771
rect 6491 11731 6496 11771
rect 6897 11740 6898 11780
rect 6938 11740 6939 11780
rect 6897 11731 6939 11740
rect 11217 11780 11259 11789
rect 11217 11740 11218 11780
rect 11258 11740 11259 11780
rect 11217 11731 11259 11740
rect 11722 11780 11780 11781
rect 11722 11740 11731 11780
rect 11771 11740 11780 11780
rect 11722 11739 11780 11740
rect 13634 11780 13676 11789
rect 13634 11740 13635 11780
rect 13675 11740 13676 11780
rect 13634 11731 13676 11740
rect 15435 11780 15477 11789
rect 15435 11740 15436 11780
rect 15476 11740 15477 11780
rect 15435 11731 15477 11740
rect 15825 11780 15867 11789
rect 15825 11740 15826 11780
rect 15866 11740 15867 11780
rect 15825 11731 15867 11740
rect 16971 11780 17013 11789
rect 16971 11740 16972 11780
rect 17012 11740 17013 11780
rect 16971 11731 17013 11740
rect 18874 11780 18932 11781
rect 18874 11740 18883 11780
rect 18923 11740 18932 11780
rect 18874 11739 18932 11740
rect 23434 11780 23492 11781
rect 23434 11740 23443 11780
rect 23483 11740 23492 11780
rect 23434 11739 23492 11740
rect 27418 11780 27476 11781
rect 27418 11740 27427 11780
rect 27467 11740 27476 11780
rect 27418 11739 27476 11740
rect 6450 11722 6496 11731
rect 24036 11729 24082 11738
rect 2890 11697 2948 11698
rect 2283 11656 2284 11696
rect 2324 11656 2325 11696
rect 2283 11647 2325 11656
rect 3032 11696 3090 11697
rect 3032 11656 3041 11696
rect 3081 11656 3090 11696
rect 3032 11655 3090 11656
rect 3350 11696 3392 11705
rect 3350 11656 3351 11696
rect 3391 11656 3392 11696
rect 3350 11647 3392 11656
rect 3483 11696 3525 11705
rect 3483 11656 3484 11696
rect 3524 11656 3525 11696
rect 3483 11647 3525 11656
rect 3723 11696 3765 11705
rect 3723 11656 3724 11696
rect 3764 11656 3765 11696
rect 3723 11647 3765 11656
rect 4299 11696 4341 11705
rect 4299 11656 4300 11696
rect 4340 11656 4341 11696
rect 4299 11647 4341 11656
rect 4971 11696 5013 11705
rect 4971 11656 4972 11696
rect 5012 11656 5013 11696
rect 4971 11647 5013 11656
rect 5098 11696 5156 11697
rect 5098 11656 5107 11696
rect 5147 11656 5156 11696
rect 5098 11655 5156 11656
rect 5494 11696 5536 11705
rect 5494 11656 5495 11696
rect 5535 11656 5536 11696
rect 5494 11647 5536 11656
rect 5626 11696 5684 11697
rect 5626 11656 5635 11696
rect 5675 11656 5684 11696
rect 5626 11655 5684 11656
rect 5739 11696 5781 11705
rect 5739 11656 5740 11696
rect 5780 11656 5781 11696
rect 5739 11647 5781 11656
rect 6315 11696 6357 11705
rect 6315 11656 6316 11696
rect 6356 11656 6357 11696
rect 6315 11647 6357 11656
rect 6544 11696 6602 11697
rect 6544 11656 6553 11696
rect 6593 11656 6602 11696
rect 6544 11655 6602 11656
rect 6987 11696 7029 11705
rect 6987 11656 6988 11696
rect 7028 11656 7029 11696
rect 6987 11647 7029 11656
rect 7755 11696 7797 11705
rect 7755 11656 7756 11696
rect 7796 11656 7797 11696
rect 7755 11647 7797 11656
rect 8043 11696 8085 11705
rect 8043 11656 8044 11696
rect 8084 11656 8085 11696
rect 8043 11647 8085 11656
rect 8412 11696 8454 11705
rect 8412 11656 8413 11696
rect 8453 11656 8454 11696
rect 8412 11647 8454 11656
rect 8523 11696 8565 11705
rect 8523 11656 8524 11696
rect 8564 11656 8565 11696
rect 8523 11647 8565 11656
rect 9003 11696 9045 11705
rect 9003 11656 9004 11696
rect 9044 11656 9045 11696
rect 9003 11647 9045 11656
rect 9387 11696 9429 11705
rect 9387 11656 9388 11696
rect 9428 11656 9429 11696
rect 9387 11647 9429 11656
rect 9771 11696 9813 11705
rect 9771 11656 9772 11696
rect 9812 11656 9813 11696
rect 9771 11647 9813 11656
rect 9946 11696 10004 11697
rect 9946 11656 9955 11696
rect 9995 11656 10004 11696
rect 9946 11655 10004 11656
rect 10141 11696 10199 11697
rect 10141 11656 10150 11696
rect 10190 11656 10199 11696
rect 10141 11655 10199 11656
rect 10454 11696 10496 11705
rect 10454 11656 10455 11696
rect 10495 11656 10496 11696
rect 10454 11647 10496 11656
rect 10635 11696 10677 11705
rect 10635 11656 10636 11696
rect 10676 11656 10677 11696
rect 10635 11647 10677 11656
rect 10827 11696 10869 11705
rect 10827 11656 10828 11696
rect 10868 11656 10869 11696
rect 10827 11647 10869 11656
rect 11307 11696 11349 11705
rect 11307 11656 11308 11696
rect 11348 11656 11349 11696
rect 11307 11647 11349 11656
rect 11979 11696 12021 11705
rect 11979 11656 11980 11696
rect 12020 11656 12021 11696
rect 11979 11647 12021 11656
rect 12363 11696 12405 11705
rect 12363 11656 12364 11696
rect 12404 11656 12405 11696
rect 12363 11647 12405 11656
rect 12795 11696 12837 11705
rect 12795 11656 12796 11696
rect 12836 11656 12837 11696
rect 12795 11647 12837 11656
rect 12939 11696 12981 11705
rect 12939 11656 12940 11696
rect 12980 11656 12981 11696
rect 12939 11647 12981 11656
rect 13515 11696 13557 11705
rect 13515 11656 13516 11696
rect 13556 11656 13557 11696
rect 13515 11647 13557 11656
rect 13732 11696 13774 11705
rect 13732 11656 13733 11696
rect 13773 11656 13774 11696
rect 13732 11647 13774 11656
rect 13899 11696 13941 11705
rect 13899 11656 13900 11696
rect 13940 11656 13941 11696
rect 13899 11647 13941 11656
rect 14091 11696 14133 11705
rect 14091 11656 14092 11696
rect 14132 11656 14133 11696
rect 14091 11647 14133 11656
rect 14266 11696 14324 11697
rect 14266 11656 14275 11696
rect 14315 11656 14324 11696
rect 14266 11655 14324 11656
rect 14379 11696 14421 11705
rect 14379 11656 14380 11696
rect 14420 11656 14421 11696
rect 14379 11647 14421 11656
rect 14763 11696 14805 11705
rect 14763 11656 14764 11696
rect 14804 11656 14805 11696
rect 14763 11647 14805 11656
rect 14955 11696 14997 11705
rect 14955 11656 14956 11696
rect 14996 11656 14997 11696
rect 14955 11647 14997 11656
rect 15094 11696 15136 11705
rect 15094 11656 15095 11696
rect 15135 11656 15136 11696
rect 15094 11647 15136 11656
rect 15226 11696 15284 11697
rect 15226 11656 15235 11696
rect 15275 11656 15284 11696
rect 15226 11655 15284 11656
rect 15340 11696 15382 11705
rect 15340 11656 15341 11696
rect 15381 11656 15382 11696
rect 15340 11647 15382 11656
rect 15915 11696 15957 11705
rect 15915 11656 15916 11696
rect 15956 11656 15957 11696
rect 15915 11647 15957 11656
rect 16474 11696 16532 11697
rect 16474 11656 16483 11696
rect 16523 11656 16532 11696
rect 16474 11655 16532 11656
rect 16683 11696 16725 11705
rect 16683 11656 16684 11696
rect 16724 11656 16725 11696
rect 16683 11647 16725 11656
rect 17067 11696 17109 11705
rect 17067 11656 17068 11696
rect 17108 11656 17109 11696
rect 17067 11647 17109 11656
rect 17186 11696 17228 11705
rect 17186 11656 17187 11696
rect 17227 11656 17228 11696
rect 17186 11647 17228 11656
rect 17296 11696 17354 11697
rect 17296 11656 17305 11696
rect 17345 11656 17354 11696
rect 17296 11655 17354 11656
rect 17440 11696 17482 11705
rect 17440 11656 17441 11696
rect 17481 11656 17482 11696
rect 17440 11647 17482 11656
rect 17731 11696 17789 11697
rect 17731 11656 17740 11696
rect 17780 11656 17789 11696
rect 17731 11655 17789 11656
rect 18507 11696 18549 11705
rect 18507 11656 18508 11696
rect 18548 11656 18549 11696
rect 18507 11647 18549 11656
rect 18742 11696 18784 11705
rect 18742 11656 18743 11696
rect 18783 11656 18784 11696
rect 18742 11647 18784 11656
rect 18987 11696 19029 11705
rect 18987 11656 18988 11696
rect 19028 11656 19029 11696
rect 18987 11647 19029 11656
rect 19467 11696 19509 11705
rect 19467 11656 19468 11696
rect 19508 11656 19509 11696
rect 19467 11647 19509 11656
rect 20026 11696 20084 11697
rect 20026 11656 20035 11696
rect 20075 11656 20084 11696
rect 20026 11655 20084 11656
rect 20139 11696 20181 11705
rect 20139 11656 20140 11696
rect 20180 11656 20181 11696
rect 20139 11647 20181 11656
rect 21178 11696 21236 11697
rect 21178 11656 21187 11696
rect 21227 11656 21236 11696
rect 21178 11655 21236 11656
rect 23599 11696 23657 11697
rect 23599 11656 23608 11696
rect 23648 11656 23657 11696
rect 23599 11655 23657 11656
rect 23787 11696 23829 11705
rect 23787 11656 23788 11696
rect 23828 11656 23829 11696
rect 23787 11647 23829 11656
rect 23901 11696 23959 11697
rect 23901 11656 23910 11696
rect 23950 11656 23959 11696
rect 24036 11689 24037 11729
rect 24077 11689 24082 11729
rect 27627 11729 27669 11738
rect 24036 11680 24082 11689
rect 24267 11696 24309 11705
rect 23901 11655 23959 11656
rect 24267 11656 24268 11696
rect 24308 11656 24309 11696
rect 24267 11647 24309 11656
rect 27034 11696 27092 11697
rect 27034 11656 27043 11696
rect 27083 11656 27092 11696
rect 27627 11689 27628 11729
rect 27668 11689 27669 11729
rect 27915 11729 27957 11738
rect 27627 11680 27669 11689
rect 27725 11696 27767 11705
rect 27034 11655 27092 11656
rect 27725 11656 27726 11696
rect 27766 11656 27767 11696
rect 27915 11689 27916 11729
rect 27956 11689 27957 11729
rect 27915 11680 27957 11689
rect 27725 11647 27767 11656
rect 5818 11612 5876 11613
rect 5818 11572 5827 11612
rect 5867 11572 5876 11612
rect 5818 11571 5876 11572
rect 9867 11612 9909 11621
rect 9867 11572 9868 11612
rect 9908 11572 9909 11612
rect 9867 11563 9909 11572
rect 10251 11612 10293 11621
rect 10251 11572 10252 11612
rect 10292 11572 10293 11612
rect 10251 11563 10293 11572
rect 10731 11612 10773 11621
rect 10731 11572 10732 11612
rect 10772 11572 10773 11612
rect 10731 11563 10773 11572
rect 14475 11612 14517 11621
rect 14475 11572 14476 11612
rect 14516 11572 14517 11612
rect 14475 11563 14517 11572
rect 14582 11612 14624 11621
rect 14582 11572 14583 11612
rect 14623 11572 14624 11612
rect 14582 11563 14624 11572
rect 17643 11612 17685 11621
rect 17643 11572 17644 11612
rect 17684 11572 17685 11612
rect 17643 11563 17685 11572
rect 18106 11612 18164 11613
rect 18106 11572 18115 11612
rect 18155 11572 18164 11612
rect 18106 11571 18164 11572
rect 20794 11612 20852 11613
rect 20794 11572 20803 11612
rect 20843 11572 20852 11612
rect 20794 11571 20852 11572
rect 25114 11612 25172 11613
rect 25114 11572 25123 11612
rect 25163 11572 25172 11612
rect 25114 11571 25172 11572
rect 1899 11528 1941 11537
rect 1899 11488 1900 11528
rect 1940 11488 1941 11528
rect 1899 11479 1941 11488
rect 2698 11528 2756 11529
rect 2698 11488 2707 11528
rect 2747 11488 2756 11528
rect 2698 11487 2756 11488
rect 3130 11528 3188 11529
rect 3130 11488 3139 11528
rect 3179 11488 3188 11528
rect 3130 11487 3188 11488
rect 4186 11528 4244 11529
rect 4186 11488 4195 11528
rect 4235 11488 4244 11528
rect 4186 11487 4244 11488
rect 4491 11528 4533 11537
rect 4491 11488 4492 11528
rect 4532 11488 4533 11528
rect 4491 11479 4533 11488
rect 5259 11528 5301 11537
rect 5259 11488 5260 11528
rect 5300 11488 5301 11528
rect 5259 11479 5301 11488
rect 7546 11528 7604 11529
rect 7546 11488 7555 11528
rect 7595 11488 7604 11528
rect 7546 11487 7604 11488
rect 9483 11528 9525 11537
rect 9483 11488 9484 11528
rect 9524 11488 9525 11528
rect 9483 11479 9525 11488
rect 11002 11528 11060 11529
rect 11002 11488 11011 11528
rect 11051 11488 11060 11528
rect 11002 11487 11060 11488
rect 13419 11528 13461 11537
rect 13419 11488 13420 11528
rect 13460 11488 13461 11528
rect 13419 11479 13461 11488
rect 14362 11528 14420 11529
rect 14362 11488 14371 11528
rect 14411 11488 14420 11528
rect 14362 11487 14420 11488
rect 19066 11528 19124 11529
rect 19066 11488 19075 11528
rect 19115 11488 19124 11528
rect 19066 11487 19124 11488
rect 20427 11528 20469 11537
rect 20427 11488 20428 11528
rect 20468 11488 20469 11528
rect 20427 11479 20469 11488
rect 23115 11528 23157 11537
rect 23115 11488 23116 11528
rect 23156 11488 23157 11528
rect 23115 11479 23157 11488
rect 24939 11528 24981 11537
rect 24939 11488 24940 11528
rect 24980 11488 24981 11528
rect 24939 11479 24981 11488
rect 576 11360 31392 11384
rect 576 11320 4352 11360
rect 4720 11320 12126 11360
rect 12494 11320 19900 11360
rect 20268 11320 27674 11360
rect 28042 11320 31392 11360
rect 576 11296 31392 11320
rect 747 11192 789 11201
rect 747 11152 748 11192
rect 788 11152 789 11192
rect 747 11143 789 11152
rect 1611 11192 1653 11201
rect 1611 11152 1612 11192
rect 1652 11152 1653 11192
rect 1611 11143 1653 11152
rect 2379 11192 2421 11201
rect 2379 11152 2380 11192
rect 2420 11152 2421 11192
rect 2379 11143 2421 11152
rect 2763 11192 2805 11201
rect 2763 11152 2764 11192
rect 2804 11152 2805 11192
rect 2763 11143 2805 11152
rect 3226 11192 3284 11193
rect 3226 11152 3235 11192
rect 3275 11152 3284 11192
rect 3226 11151 3284 11152
rect 4186 11192 4244 11193
rect 4186 11152 4195 11192
rect 4235 11152 4244 11192
rect 4186 11151 4244 11152
rect 4474 11192 4532 11193
rect 4474 11152 4483 11192
rect 4523 11152 4532 11192
rect 4474 11151 4532 11152
rect 5451 11192 5493 11201
rect 5451 11152 5452 11192
rect 5492 11152 5493 11192
rect 5451 11143 5493 11152
rect 6490 11192 6548 11193
rect 6490 11152 6499 11192
rect 6539 11152 6548 11192
rect 6490 11151 6548 11152
rect 7323 11192 7365 11201
rect 7323 11152 7324 11192
rect 7364 11152 7365 11192
rect 7323 11143 7365 11152
rect 7546 11192 7604 11193
rect 7546 11152 7555 11192
rect 7595 11152 7604 11192
rect 7546 11151 7604 11152
rect 8523 11192 8565 11201
rect 8523 11152 8524 11192
rect 8564 11152 8565 11192
rect 8523 11143 8565 11152
rect 9099 11192 9141 11201
rect 9099 11152 9100 11192
rect 9140 11152 9141 11192
rect 9099 11143 9141 11152
rect 9867 11192 9909 11201
rect 9867 11152 9868 11192
rect 9908 11152 9909 11192
rect 9867 11143 9909 11152
rect 10138 11192 10196 11193
rect 10138 11152 10147 11192
rect 10187 11152 10196 11192
rect 10138 11151 10196 11152
rect 12346 11192 12404 11193
rect 12346 11152 12355 11192
rect 12395 11152 12404 11192
rect 12346 11151 12404 11152
rect 12922 11192 12980 11193
rect 12922 11152 12931 11192
rect 12971 11152 12980 11192
rect 12922 11151 12980 11152
rect 13210 11192 13268 11193
rect 13210 11152 13219 11192
rect 13259 11152 13268 11192
rect 13210 11151 13268 11152
rect 13978 11192 14036 11193
rect 13978 11152 13987 11192
rect 14027 11152 14036 11192
rect 13978 11151 14036 11152
rect 14746 11192 14804 11193
rect 14746 11152 14755 11192
rect 14795 11152 14804 11192
rect 14746 11151 14804 11152
rect 16474 11192 16532 11193
rect 16474 11152 16483 11192
rect 16523 11152 16532 11192
rect 16474 11151 16532 11152
rect 17739 11192 17781 11201
rect 17739 11152 17740 11192
rect 17780 11152 17781 11192
rect 17739 11143 17781 11152
rect 18010 11192 18068 11193
rect 18010 11152 18019 11192
rect 18059 11152 18068 11192
rect 18010 11151 18068 11152
rect 18490 11192 18548 11193
rect 18490 11152 18499 11192
rect 18539 11152 18548 11192
rect 18490 11151 18548 11152
rect 20026 11192 20084 11193
rect 20026 11152 20035 11192
rect 20075 11152 20084 11192
rect 20026 11151 20084 11152
rect 21771 11192 21813 11201
rect 21771 11152 21772 11192
rect 21812 11152 21813 11192
rect 21771 11143 21813 11152
rect 23355 11192 23397 11201
rect 23355 11152 23356 11192
rect 23396 11152 23397 11192
rect 23355 11143 23397 11152
rect 23979 11192 24021 11201
rect 23979 11152 23980 11192
rect 24020 11152 24021 11192
rect 23979 11143 24021 11152
rect 24603 11192 24645 11201
rect 24603 11152 24604 11192
rect 24644 11152 24645 11192
rect 24603 11143 24645 11152
rect 27706 11192 27764 11193
rect 27706 11152 27715 11192
rect 27755 11152 27764 11192
rect 27706 11151 27764 11152
rect 4587 11108 4629 11117
rect 4587 11068 4588 11108
rect 4628 11068 4629 11108
rect 4587 11059 4629 11068
rect 7769 11108 7811 11117
rect 7769 11068 7770 11108
rect 7810 11068 7811 11108
rect 7769 11059 7811 11068
rect 8427 11108 8469 11117
rect 8427 11068 8428 11108
rect 8468 11068 8469 11108
rect 8427 11059 8469 11068
rect 9562 11108 9620 11109
rect 9562 11068 9571 11108
rect 9611 11068 9620 11108
rect 9562 11067 9620 11068
rect 10347 11108 10389 11117
rect 10347 11068 10348 11108
rect 10388 11068 10389 11108
rect 10347 11059 10389 11068
rect 19707 11108 19749 11117
rect 19707 11068 19708 11108
rect 19748 11068 19749 11108
rect 19707 11059 19749 11068
rect 651 11024 693 11033
rect 651 10984 652 11024
rect 692 10984 693 11024
rect 651 10975 693 10984
rect 826 11024 884 11025
rect 826 10984 835 11024
rect 875 10984 884 11024
rect 826 10983 884 10984
rect 1323 11024 1365 11033
rect 1323 10984 1324 11024
rect 1364 10984 1365 11024
rect 1323 10975 1365 10984
rect 1450 11024 1508 11025
rect 1450 10984 1459 11024
rect 1499 10984 1508 11024
rect 1450 10983 1508 10984
rect 1978 11024 2036 11025
rect 1978 10984 1987 11024
rect 2027 10984 2036 11024
rect 1978 10983 2036 10984
rect 2091 11024 2133 11033
rect 2091 10984 2092 11024
rect 2132 10984 2133 11024
rect 2091 10975 2133 10984
rect 2763 11024 2805 11033
rect 2763 10984 2764 11024
rect 2804 10984 2805 11024
rect 2763 10975 2805 10984
rect 2955 11024 2997 11033
rect 2955 10984 2956 11024
rect 2996 10984 2997 11024
rect 2955 10975 2997 10984
rect 3339 11024 3381 11033
rect 3339 10984 3340 11024
rect 3380 10984 3381 11024
rect 3339 10975 3381 10984
rect 3723 11024 3765 11033
rect 3723 10984 3724 11024
rect 3764 10984 3765 11024
rect 3723 10975 3765 10984
rect 3862 11024 3904 11033
rect 3862 10984 3863 11024
rect 3903 10984 3904 11024
rect 3862 10975 3904 10984
rect 4107 11024 4149 11033
rect 4107 10984 4108 11024
rect 4148 10984 4149 11024
rect 4107 10975 4149 10984
rect 4378 11024 4436 11025
rect 4378 10984 4387 11024
rect 4427 10984 4436 11024
rect 4378 10983 4436 10984
rect 4694 11024 4736 11033
rect 4694 10984 4695 11024
rect 4735 10984 4736 11024
rect 4694 10975 4736 10984
rect 5050 11024 5108 11025
rect 5050 10984 5059 11024
rect 5099 10984 5108 11024
rect 5050 10983 5108 10984
rect 5163 11024 5205 11033
rect 5163 10984 5164 11024
rect 5204 10984 5205 11024
rect 5163 10975 5205 10984
rect 5595 11024 5637 11033
rect 5595 10984 5596 11024
rect 5636 10984 5637 11024
rect 5595 10975 5637 10984
rect 5896 11024 5938 11033
rect 5896 10984 5897 11024
rect 5937 10984 5938 11024
rect 5896 10975 5938 10984
rect 6050 11024 6092 11033
rect 6050 10984 6051 11024
rect 6091 10984 6092 11024
rect 6050 10975 6092 10984
rect 6603 11024 6645 11033
rect 6603 10984 6604 11024
rect 6644 10984 6645 11024
rect 6603 10975 6645 10984
rect 6987 11024 7029 11033
rect 6987 10984 6988 11024
rect 7028 10984 7029 11024
rect 6987 10975 7029 10984
rect 7179 11024 7221 11033
rect 7179 10984 7180 11024
rect 7220 10984 7221 11024
rect 7179 10975 7221 10984
rect 7450 11024 7508 11025
rect 7450 10984 7459 11024
rect 7499 10984 7508 11024
rect 7450 10983 7508 10984
rect 7947 11024 7989 11033
rect 7947 10984 7948 11024
rect 7988 10984 7989 11024
rect 7947 10975 7989 10984
rect 8139 11024 8181 11033
rect 8139 10984 8140 11024
rect 8180 10984 8181 11024
rect 8139 10975 8181 10984
rect 8314 11024 8372 11025
rect 8314 10984 8323 11024
rect 8363 10984 8372 11024
rect 8314 10983 8372 10984
rect 8630 11024 8672 11033
rect 8630 10984 8631 11024
rect 8671 10984 8672 11024
rect 8630 10975 8672 10984
rect 8811 11024 8853 11033
rect 8811 10984 8812 11024
rect 8852 10984 8853 11024
rect 8811 10975 8853 10984
rect 8945 11024 9003 11025
rect 8945 10984 8954 11024
rect 8994 10984 9003 11024
rect 8945 10983 9003 10984
rect 9238 11024 9280 11033
rect 9238 10984 9239 11024
rect 9279 10984 9280 11024
rect 9238 10975 9280 10984
rect 9483 11024 9525 11033
rect 9483 10984 9484 11024
rect 9524 10984 9525 11024
rect 9483 10975 9525 10984
rect 10059 11024 10101 11033
rect 10059 10984 10060 11024
rect 10100 10984 10101 11024
rect 10059 10975 10101 10984
rect 10522 11024 10580 11025
rect 10522 10984 10531 11024
rect 10571 10984 10580 11024
rect 10522 10983 10580 10984
rect 11119 11024 11177 11025
rect 11119 10984 11128 11024
rect 11168 10984 11177 11024
rect 11119 10983 11177 10984
rect 11691 11024 11733 11033
rect 11691 10984 11692 11024
rect 11732 10984 11733 11024
rect 11691 10975 11733 10984
rect 11866 11024 11924 11025
rect 11866 10984 11875 11024
rect 11915 10984 11924 11024
rect 12268 11024 12310 11033
rect 11866 10983 11924 10984
rect 12027 10982 12069 10991
rect 3994 10940 4052 10941
rect 3994 10900 4003 10940
rect 4043 10900 4052 10940
rect 3994 10899 4052 10900
rect 5739 10940 5781 10949
rect 5739 10900 5740 10940
rect 5780 10900 5781 10940
rect 5739 10891 5781 10900
rect 9370 10940 9428 10941
rect 9370 10900 9379 10940
rect 9419 10900 9428 10940
rect 10954 10940 11012 10941
rect 9370 10899 9428 10900
rect 10571 10898 10613 10907
rect 10954 10900 10963 10940
rect 11003 10900 11012 10940
rect 10954 10899 11012 10900
rect 11307 10940 11349 10949
rect 11307 10900 11308 10940
rect 11348 10900 11349 10940
rect 12027 10942 12028 10982
rect 12068 10942 12069 10982
rect 12268 10984 12269 11024
rect 12309 10984 12310 11024
rect 12268 10975 12310 10984
rect 12603 11024 12645 11033
rect 12603 10984 12604 11024
rect 12644 10984 12645 11024
rect 12603 10975 12645 10984
rect 12843 11024 12885 11033
rect 12843 10984 12844 11024
rect 12884 10984 12885 11024
rect 12843 10975 12885 10984
rect 13419 11024 13461 11033
rect 13419 10984 13420 11024
rect 13460 10984 13461 11024
rect 13419 10975 13461 10984
rect 13707 11024 13749 11033
rect 13707 10984 13708 11024
rect 13748 10984 13749 11024
rect 13707 10975 13749 10984
rect 14091 11024 14133 11033
rect 14091 10984 14092 11024
rect 14132 10984 14133 11024
rect 14091 10975 14133 10984
rect 14475 11024 14517 11033
rect 14475 10984 14476 11024
rect 14516 10984 14517 11024
rect 14475 10975 14517 10984
rect 14955 11024 14997 11033
rect 14955 10984 14956 11024
rect 14996 10984 14997 11024
rect 14955 10975 14997 10984
rect 15243 11024 15285 11033
rect 15243 10984 15244 11024
rect 15284 10984 15285 11024
rect 15243 10975 15285 10984
rect 16011 11024 16053 11033
rect 16011 10984 16012 11024
rect 16052 10984 16053 11024
rect 16011 10975 16053 10984
rect 16138 11024 16196 11025
rect 16138 10984 16147 11024
rect 16187 10984 16196 11024
rect 16138 10983 16196 10984
rect 16779 11024 16821 11033
rect 16779 10984 16780 11024
rect 16820 10984 16821 11024
rect 16779 10975 16821 10984
rect 17242 11024 17300 11025
rect 17242 10984 17251 11024
rect 17291 10984 17300 11024
rect 17242 10983 17300 10984
rect 17547 11024 17589 11033
rect 17547 10984 17548 11024
rect 17588 10984 17589 11024
rect 17547 10975 17589 10984
rect 17931 11024 17973 11033
rect 17931 10984 17932 11024
rect 17972 10984 17973 11024
rect 17931 10975 17973 10984
rect 18166 11024 18208 11033
rect 18166 10984 18167 11024
rect 18207 10984 18208 11024
rect 18166 10975 18208 10984
rect 18411 11024 18453 11033
rect 18411 10984 18412 11024
rect 18452 10984 18453 11024
rect 18411 10975 18453 10984
rect 19021 11024 19079 11025
rect 20331 11024 20373 11033
rect 19021 10984 19030 11024
rect 19070 10984 19079 11024
rect 19021 10983 19079 10984
rect 19554 11015 19600 11024
rect 19554 10975 19555 11015
rect 19595 10975 19600 11015
rect 20331 10984 20332 11024
rect 20372 10984 20373 11024
rect 20331 10975 20373 10984
rect 20907 11024 20949 11033
rect 20907 10984 20908 11024
rect 20948 10984 20949 11024
rect 20907 10975 20949 10984
rect 22443 11024 22485 11033
rect 22443 10984 22444 11024
rect 22484 10984 22485 11024
rect 22443 10975 22485 10984
rect 22731 11024 22773 11033
rect 22731 10984 22732 11024
rect 22772 10984 22773 11024
rect 22731 10975 22773 10984
rect 22923 11024 22965 11033
rect 24171 11024 24213 11033
rect 26938 11024 26996 11025
rect 22923 10984 22924 11024
rect 22964 10984 22965 11024
rect 22923 10975 22965 10984
rect 23202 11015 23248 11024
rect 23202 10975 23203 11015
rect 23243 10975 23248 11015
rect 24171 10984 24172 11024
rect 24212 10984 24213 11024
rect 24171 10975 24213 10984
rect 24450 11015 24496 11024
rect 24450 10975 24451 11015
rect 24491 10975 24496 11015
rect 26938 10984 26947 11024
rect 26987 10984 26996 11024
rect 26938 10983 26996 10984
rect 27531 11024 27573 11033
rect 27531 10984 27532 11024
rect 27572 10984 27573 11024
rect 27531 10975 27573 10984
rect 27723 11024 27765 11033
rect 27723 10984 27724 11024
rect 27764 10984 27765 11024
rect 27723 10975 27765 10984
rect 19554 10966 19600 10975
rect 23202 10966 23248 10975
rect 24450 10966 24496 10975
rect 12027 10933 12069 10942
rect 12154 10940 12212 10941
rect 5835 10856 5877 10865
rect 5835 10816 5836 10856
rect 5876 10816 5877 10856
rect 10571 10858 10572 10898
rect 10612 10858 10613 10898
rect 11307 10891 11349 10900
rect 12154 10900 12163 10940
rect 12203 10900 12212 10940
rect 12154 10899 12212 10900
rect 12730 10940 12788 10941
rect 12730 10900 12739 10940
rect 12779 10900 12788 10940
rect 12730 10899 12788 10900
rect 16689 10940 16731 10949
rect 16689 10900 16690 10940
rect 16730 10900 16731 10940
rect 16689 10891 16731 10900
rect 18298 10940 18356 10941
rect 18298 10900 18307 10940
rect 18347 10900 18356 10940
rect 18298 10899 18356 10900
rect 18826 10940 18884 10941
rect 18826 10900 18835 10940
rect 18875 10900 18884 10940
rect 18826 10899 18884 10900
rect 20241 10940 20283 10949
rect 20241 10900 20242 10940
rect 20282 10900 20283 10940
rect 20241 10891 20283 10900
rect 25402 10940 25460 10941
rect 25402 10900 25411 10940
rect 25451 10900 25460 10940
rect 25402 10899 25460 10900
rect 27322 10940 27380 10941
rect 27322 10900 27331 10940
rect 27371 10900 27380 10940
rect 27322 10899 27380 10900
rect 10571 10849 10613 10858
rect 11866 10856 11924 10857
rect 5835 10807 5877 10816
rect 11866 10816 11875 10856
rect 11915 10816 11924 10856
rect 11866 10815 11924 10816
rect 16186 10856 16244 10857
rect 16186 10816 16195 10856
rect 16235 10816 16244 10856
rect 16186 10815 16244 10816
rect 17547 10856 17589 10865
rect 17547 10816 17548 10856
rect 17588 10816 17589 10856
rect 17547 10807 17589 10816
rect 19371 10856 19413 10865
rect 19371 10816 19372 10856
rect 19412 10816 19413 10856
rect 19371 10807 19413 10816
rect 22714 10856 22772 10857
rect 22714 10816 22723 10856
rect 22763 10816 22772 10856
rect 22714 10815 22772 10816
rect 7755 10772 7797 10781
rect 7755 10732 7756 10772
rect 7796 10732 7797 10772
rect 7755 10723 7797 10732
rect 8043 10772 8085 10781
rect 8043 10732 8044 10772
rect 8084 10732 8085 10772
rect 8043 10723 8085 10732
rect 11547 10772 11589 10781
rect 11547 10732 11548 10772
rect 11588 10732 11589 10772
rect 11547 10723 11589 10732
rect 21579 10772 21621 10781
rect 21579 10732 21580 10772
rect 21620 10732 21621 10772
rect 21579 10723 21621 10732
rect 25035 10772 25077 10781
rect 25035 10732 25036 10772
rect 25076 10732 25077 10772
rect 25035 10723 25077 10732
rect 576 10604 31392 10628
rect 576 10564 3112 10604
rect 3480 10564 10886 10604
rect 11254 10564 18660 10604
rect 19028 10564 26434 10604
rect 26802 10564 31392 10604
rect 576 10540 31392 10564
rect 1755 10436 1797 10445
rect 1755 10396 1756 10436
rect 1796 10396 1797 10436
rect 1755 10387 1797 10396
rect 3130 10436 3188 10437
rect 3130 10396 3139 10436
rect 3179 10396 3188 10436
rect 3130 10395 3188 10396
rect 3531 10436 3573 10445
rect 3531 10396 3532 10436
rect 3572 10396 3573 10436
rect 3531 10387 3573 10396
rect 4474 10436 4532 10437
rect 4474 10396 4483 10436
rect 4523 10396 4532 10436
rect 4474 10395 4532 10396
rect 6586 10436 6644 10437
rect 6586 10396 6595 10436
rect 6635 10396 6644 10436
rect 6586 10395 6644 10396
rect 8715 10436 8757 10445
rect 8715 10396 8716 10436
rect 8756 10396 8757 10436
rect 8715 10387 8757 10396
rect 9195 10436 9237 10445
rect 9195 10396 9196 10436
rect 9236 10396 9237 10436
rect 9195 10387 9237 10396
rect 12058 10436 12116 10437
rect 12058 10396 12067 10436
rect 12107 10396 12116 10436
rect 12058 10395 12116 10396
rect 13690 10436 13748 10437
rect 13690 10396 13699 10436
rect 13739 10396 13748 10436
rect 13690 10395 13748 10396
rect 14187 10436 14229 10445
rect 14187 10396 14188 10436
rect 14228 10396 14229 10436
rect 14187 10387 14229 10396
rect 16186 10436 16244 10437
rect 16186 10396 16195 10436
rect 16235 10396 16244 10436
rect 16186 10395 16244 10396
rect 16587 10436 16629 10445
rect 16587 10396 16588 10436
rect 16628 10396 16629 10436
rect 16587 10387 16629 10396
rect 21483 10436 21525 10445
rect 21483 10396 21484 10436
rect 21524 10396 21525 10436
rect 21483 10387 21525 10396
rect 24075 10436 24117 10445
rect 24075 10396 24076 10436
rect 24116 10396 24117 10436
rect 24075 10387 24117 10396
rect 922 10352 980 10353
rect 922 10312 931 10352
rect 971 10312 980 10352
rect 922 10311 980 10312
rect 2523 10352 2565 10361
rect 2523 10312 2524 10352
rect 2564 10312 2565 10352
rect 2523 10303 2565 10312
rect 4011 10352 4053 10361
rect 4011 10312 4012 10352
rect 4052 10312 4053 10352
rect 4011 10303 4053 10312
rect 5355 10352 5397 10361
rect 5355 10312 5356 10352
rect 5396 10312 5397 10352
rect 5355 10303 5397 10312
rect 8026 10352 8084 10353
rect 8026 10312 8035 10352
rect 8075 10312 8084 10352
rect 8026 10311 8084 10312
rect 15531 10352 15573 10361
rect 15531 10312 15532 10352
rect 15572 10312 15573 10352
rect 15531 10303 15573 10312
rect 17739 10352 17781 10361
rect 17739 10312 17740 10352
rect 17780 10312 17781 10352
rect 17739 10303 17781 10312
rect 21867 10352 21909 10361
rect 21867 10312 21868 10352
rect 21908 10312 21909 10352
rect 21867 10303 21909 10312
rect 23674 10352 23732 10353
rect 23674 10312 23683 10352
rect 23723 10312 23732 10352
rect 23674 10311 23732 10312
rect 27147 10352 27189 10361
rect 27147 10312 27148 10352
rect 27188 10312 27189 10352
rect 27147 10303 27189 10312
rect 1978 10268 2036 10269
rect 1978 10228 1987 10268
rect 2027 10228 2036 10268
rect 1978 10227 2036 10228
rect 2187 10268 2229 10277
rect 2187 10228 2188 10268
rect 2228 10228 2229 10268
rect 2187 10219 2229 10228
rect 4762 10268 4820 10269
rect 4762 10228 4771 10268
rect 4811 10228 4820 10268
rect 4762 10227 4820 10228
rect 4971 10268 5013 10277
rect 4971 10228 4972 10268
rect 5012 10228 5013 10268
rect 4971 10219 5013 10228
rect 5259 10268 5301 10277
rect 5259 10228 5260 10268
rect 5300 10228 5301 10268
rect 5259 10219 5301 10228
rect 7275 10268 7317 10277
rect 7275 10228 7276 10268
rect 7316 10228 7317 10268
rect 7275 10219 7317 10228
rect 11674 10268 11732 10269
rect 11674 10228 11683 10268
rect 11723 10228 11732 10268
rect 11674 10227 11732 10228
rect 12634 10268 12692 10269
rect 12634 10228 12643 10268
rect 12683 10228 12692 10268
rect 12634 10227 12692 10228
rect 12843 10268 12885 10277
rect 12843 10228 12844 10268
rect 12884 10228 12885 10268
rect 11106 10217 11152 10226
rect 12843 10219 12885 10228
rect 13227 10268 13269 10277
rect 16689 10268 16731 10277
rect 13227 10228 13228 10268
rect 13268 10228 13269 10268
rect 13227 10219 13269 10228
rect 13458 10259 13504 10268
rect 13458 10219 13459 10259
rect 13499 10219 13504 10259
rect 747 10184 789 10193
rect 747 10144 748 10184
rect 788 10144 789 10184
rect 747 10135 789 10144
rect 922 10184 980 10185
rect 922 10144 931 10184
rect 971 10144 980 10184
rect 922 10143 980 10144
rect 1131 10184 1173 10193
rect 1131 10144 1132 10184
rect 1172 10144 1173 10184
rect 1131 10135 1173 10144
rect 1515 10184 1557 10193
rect 1515 10144 1516 10184
rect 1556 10144 1557 10184
rect 1515 10135 1557 10144
rect 1846 10184 1888 10193
rect 1846 10144 1847 10184
rect 1887 10144 1888 10184
rect 1846 10135 1888 10144
rect 2091 10184 2133 10193
rect 2091 10144 2092 10184
rect 2132 10144 2133 10184
rect 2091 10135 2133 10144
rect 2379 10184 2421 10193
rect 2379 10144 2380 10184
rect 2420 10144 2421 10184
rect 2379 10135 2421 10144
rect 2842 10184 2900 10185
rect 2842 10144 2851 10184
rect 2891 10144 2900 10184
rect 2842 10143 2900 10144
rect 2955 10184 2997 10193
rect 2955 10144 2956 10184
rect 2996 10144 2997 10184
rect 2955 10135 2997 10144
rect 3435 10184 3477 10193
rect 3435 10144 3436 10184
rect 3476 10144 3477 10184
rect 3435 10135 3477 10144
rect 3627 10184 3669 10193
rect 3627 10144 3628 10184
rect 3668 10144 3669 10184
rect 3627 10135 3669 10144
rect 3915 10184 3957 10193
rect 3915 10144 3916 10184
rect 3956 10144 3957 10184
rect 3915 10135 3957 10144
rect 4107 10184 4149 10193
rect 4107 10144 4108 10184
rect 4148 10144 4149 10184
rect 4107 10135 4149 10144
rect 4299 10184 4341 10193
rect 4299 10144 4300 10184
rect 4340 10144 4341 10184
rect 4299 10135 4341 10144
rect 4490 10184 4532 10193
rect 4490 10144 4491 10184
rect 4531 10144 4532 10184
rect 4490 10135 4532 10144
rect 4630 10184 4672 10193
rect 4630 10144 4631 10184
rect 4671 10144 4672 10184
rect 4630 10135 4672 10144
rect 4875 10184 4917 10193
rect 4875 10144 4876 10184
rect 4916 10144 4917 10184
rect 4875 10135 4917 10144
rect 5122 10184 5180 10185
rect 5122 10144 5131 10184
rect 5171 10144 5180 10184
rect 5122 10143 5180 10144
rect 5416 10184 5458 10193
rect 5416 10144 5417 10184
rect 5457 10144 5458 10184
rect 5416 10135 5458 10144
rect 5578 10184 5636 10185
rect 5578 10144 5587 10184
rect 5627 10144 5636 10184
rect 5578 10143 5636 10144
rect 5739 10184 5781 10193
rect 5739 10144 5740 10184
rect 5780 10144 5781 10184
rect 5739 10135 5781 10144
rect 5936 10184 5978 10193
rect 5936 10144 5937 10184
rect 5977 10144 5978 10184
rect 5936 10135 5978 10144
rect 6298 10184 6356 10185
rect 6298 10144 6307 10184
rect 6347 10144 6356 10184
rect 6298 10143 6356 10144
rect 6411 10184 6453 10193
rect 6411 10144 6412 10184
rect 6452 10144 6453 10184
rect 6411 10135 6453 10144
rect 6948 10184 7006 10185
rect 6948 10144 6957 10184
rect 6997 10144 7006 10184
rect 6948 10143 7006 10144
rect 7104 10184 7146 10193
rect 7104 10144 7105 10184
rect 7145 10144 7146 10184
rect 7104 10135 7146 10144
rect 7396 10184 7438 10193
rect 7396 10144 7397 10184
rect 7437 10144 7438 10184
rect 7396 10135 7438 10144
rect 7738 10184 7796 10185
rect 7738 10144 7747 10184
rect 7787 10144 7796 10184
rect 7738 10143 7796 10144
rect 7851 10184 7893 10193
rect 7851 10144 7852 10184
rect 7892 10144 7893 10184
rect 7851 10135 7893 10144
rect 8506 10184 8564 10185
rect 8506 10144 8515 10184
rect 8555 10144 8564 10184
rect 8506 10143 8564 10144
rect 8619 10184 8661 10193
rect 8619 10144 8620 10184
rect 8660 10144 8661 10184
rect 8619 10135 8661 10144
rect 9243 10184 9285 10193
rect 9243 10144 9244 10184
rect 9284 10144 9285 10184
rect 9243 10135 9285 10144
rect 9387 10184 9429 10193
rect 9387 10144 9388 10184
rect 9428 10144 9429 10184
rect 9387 10135 9429 10144
rect 10044 10184 10086 10193
rect 10044 10144 10045 10184
rect 10085 10144 10086 10184
rect 10044 10135 10086 10144
rect 10155 10184 10197 10193
rect 10155 10144 10156 10184
rect 10196 10144 10197 10184
rect 10155 10135 10197 10144
rect 10635 10184 10677 10193
rect 10635 10144 10636 10184
rect 10676 10144 10677 10184
rect 10635 10135 10677 10144
rect 10774 10184 10816 10193
rect 10774 10144 10775 10184
rect 10815 10144 10816 10184
rect 11106 10177 11107 10217
rect 11147 10177 11152 10217
rect 13458 10210 13504 10219
rect 14187 10226 14229 10235
rect 11106 10168 11152 10177
rect 11542 10184 11584 10193
rect 10774 10135 10816 10144
rect 11542 10144 11543 10184
rect 11583 10144 11584 10184
rect 11542 10135 11584 10144
rect 11787 10184 11829 10193
rect 11787 10144 11788 10184
rect 11828 10144 11829 10184
rect 11787 10135 11829 10144
rect 12061 10184 12103 10193
rect 12061 10144 12062 10184
rect 12102 10144 12103 10184
rect 12061 10135 12103 10144
rect 12355 10184 12413 10185
rect 12355 10144 12364 10184
rect 12404 10144 12413 10184
rect 12355 10143 12413 10144
rect 12514 10184 12572 10185
rect 12514 10144 12523 10184
rect 12563 10144 12572 10184
rect 12514 10143 12572 10144
rect 12747 10184 12789 10193
rect 12747 10144 12748 10184
rect 12788 10144 12789 10184
rect 12747 10135 12789 10144
rect 13323 10184 13365 10193
rect 14187 10186 14188 10226
rect 14228 10186 14229 10226
rect 13323 10144 13324 10184
rect 13364 10144 13365 10184
rect 13323 10135 13365 10144
rect 13552 10184 13610 10185
rect 13552 10144 13561 10184
rect 13601 10144 13610 10184
rect 13552 10143 13610 10144
rect 13987 10184 14045 10185
rect 13987 10144 13996 10184
rect 14036 10144 14045 10184
rect 14187 10177 14229 10186
rect 14379 10226 14421 10235
rect 16689 10228 16690 10268
rect 16730 10228 16731 10268
rect 14379 10186 14380 10226
rect 14420 10186 14421 10226
rect 14379 10177 14421 10186
rect 15255 10217 15297 10226
rect 16689 10219 16731 10228
rect 19563 10268 19605 10277
rect 19563 10228 19564 10268
rect 19604 10228 19605 10268
rect 19563 10219 19605 10228
rect 24177 10268 24219 10277
rect 24177 10228 24178 10268
rect 24218 10228 24219 10268
rect 24177 10219 24219 10228
rect 24874 10268 24932 10269
rect 24874 10228 24883 10268
rect 24923 10228 24932 10268
rect 24874 10227 24932 10228
rect 14602 10184 14660 10185
rect 13987 10143 14045 10144
rect 14602 10144 14611 10184
rect 14651 10144 14660 10184
rect 14602 10143 14660 10144
rect 14704 10184 14762 10185
rect 14704 10144 14713 10184
rect 14753 10144 14762 10184
rect 14704 10143 14762 10144
rect 15130 10184 15188 10185
rect 15130 10144 15139 10184
rect 15179 10144 15188 10184
rect 15255 10177 15256 10217
rect 15296 10177 15297 10217
rect 15255 10168 15297 10177
rect 16011 10184 16053 10193
rect 15130 10143 15188 10144
rect 16011 10144 16012 10184
rect 16052 10144 16053 10184
rect 16011 10135 16053 10144
rect 16138 10184 16196 10185
rect 16138 10144 16147 10184
rect 16187 10144 16196 10184
rect 16138 10143 16196 10144
rect 16779 10184 16821 10193
rect 16779 10144 16780 10184
rect 16820 10144 16821 10184
rect 16779 10135 16821 10144
rect 17259 10184 17301 10193
rect 17259 10144 17260 10184
rect 17300 10144 17301 10184
rect 17259 10135 17301 10144
rect 17393 10184 17451 10185
rect 17393 10144 17402 10184
rect 17442 10144 17451 10184
rect 17393 10143 17451 10144
rect 17931 10184 17973 10193
rect 17931 10144 17932 10184
rect 17972 10144 17973 10184
rect 17931 10135 17973 10144
rect 18219 10184 18261 10193
rect 18219 10144 18220 10184
rect 18260 10144 18261 10184
rect 18219 10135 18261 10144
rect 18394 10184 18452 10185
rect 18394 10144 18403 10184
rect 18443 10144 18452 10184
rect 18394 10143 18452 10144
rect 18890 10184 18932 10193
rect 18890 10144 18891 10184
rect 18931 10144 18932 10184
rect 18890 10135 18932 10144
rect 19018 10184 19076 10185
rect 19018 10144 19027 10184
rect 19067 10144 19076 10184
rect 19018 10143 19076 10144
rect 19930 10184 19988 10185
rect 19930 10144 19939 10184
rect 19979 10144 19988 10184
rect 19930 10143 19988 10144
rect 22059 10184 22101 10193
rect 22059 10144 22060 10184
rect 22100 10144 22101 10184
rect 22059 10135 22101 10144
rect 23019 10184 23061 10193
rect 23019 10144 23020 10184
rect 23060 10144 23061 10184
rect 23019 10135 23061 10144
rect 23386 10184 23444 10185
rect 23386 10144 23395 10184
rect 23435 10144 23444 10184
rect 23386 10143 23444 10144
rect 23499 10184 23541 10193
rect 23499 10144 23500 10184
rect 23540 10144 23541 10184
rect 23499 10135 23541 10144
rect 24267 10184 24309 10193
rect 24267 10144 24268 10184
rect 24308 10144 24309 10184
rect 24267 10135 24309 10144
rect 25039 10184 25097 10185
rect 25039 10144 25048 10184
rect 25088 10144 25097 10184
rect 25039 10143 25097 10144
rect 25419 10184 25461 10193
rect 25419 10144 25420 10184
rect 25460 10144 25461 10184
rect 25419 10135 25461 10144
rect 26955 10184 26997 10193
rect 26955 10144 26956 10184
rect 26996 10144 26997 10184
rect 26955 10135 26997 10144
rect 10971 10100 11013 10109
rect 7193 10058 7235 10067
rect 5739 10016 5781 10025
rect 5739 9976 5740 10016
rect 5780 9976 5781 10016
rect 7193 10018 7194 10058
rect 7234 10018 7235 10058
rect 10971 10060 10972 10100
rect 11012 10060 11013 10100
rect 10971 10051 11013 10060
rect 13693 10100 13735 10109
rect 13693 10060 13694 10100
rect 13734 10060 13735 10100
rect 13693 10051 13735 10060
rect 14907 10100 14949 10109
rect 14907 10060 14908 10100
rect 14948 10060 14949 10100
rect 14907 10051 14949 10060
rect 17595 10100 17637 10109
rect 17595 10060 17596 10100
rect 17636 10060 17637 10100
rect 17595 10051 17637 10060
rect 18315 10100 18357 10109
rect 18315 10060 18316 10100
rect 18356 10060 18357 10100
rect 18315 10051 18357 10060
rect 7193 10009 7235 10018
rect 9850 10016 9908 10017
rect 5739 9967 5781 9976
rect 9850 9976 9859 10016
rect 9899 9976 9908 10016
rect 9850 9975 9908 9976
rect 11259 10016 11301 10025
rect 11259 9976 11260 10016
rect 11300 9976 11301 10016
rect 11259 9967 11301 9976
rect 11866 10016 11924 10017
rect 11866 9976 11875 10016
rect 11915 9976 11924 10016
rect 11866 9975 11924 9976
rect 12267 10016 12309 10025
rect 12267 9976 12268 10016
rect 12308 9976 12309 10016
rect 12267 9967 12309 9976
rect 13899 10016 13941 10025
rect 18010 10016 18068 10017
rect 13899 9976 13900 10016
rect 13940 9976 13941 10016
rect 13899 9967 13941 9976
rect 15042 10007 15088 10016
rect 15042 9967 15043 10007
rect 15083 9967 15088 10007
rect 18010 9976 18019 10016
rect 18059 9976 18068 10016
rect 18010 9975 18068 9976
rect 19179 10016 19221 10025
rect 19179 9976 19180 10016
rect 19220 9976 19221 10016
rect 19179 9967 19221 9976
rect 22347 10016 22389 10025
rect 22347 9976 22348 10016
rect 22388 9976 22389 10016
rect 22347 9967 22389 9976
rect 26091 10016 26133 10025
rect 26091 9976 26092 10016
rect 26132 9976 26133 10016
rect 26091 9967 26133 9976
rect 26283 10016 26325 10025
rect 26283 9976 26284 10016
rect 26324 9976 26325 10016
rect 26283 9967 26325 9976
rect 15042 9958 15088 9967
rect 576 9848 31392 9872
rect 576 9808 4352 9848
rect 4720 9808 12126 9848
rect 12494 9808 19900 9848
rect 20268 9808 27674 9848
rect 28042 9808 31392 9848
rect 576 9784 31392 9808
rect 1114 9680 1172 9681
rect 1114 9640 1123 9680
rect 1163 9640 1172 9680
rect 1114 9639 1172 9640
rect 1498 9680 1556 9681
rect 1498 9640 1507 9680
rect 1547 9640 1556 9680
rect 1498 9639 1556 9640
rect 4779 9680 4821 9689
rect 4779 9640 4780 9680
rect 4820 9640 4821 9680
rect 4779 9631 4821 9640
rect 4954 9680 5012 9681
rect 4954 9640 4963 9680
rect 5003 9640 5012 9680
rect 4954 9639 5012 9640
rect 6315 9680 6357 9689
rect 6315 9640 6316 9680
rect 6356 9640 6357 9680
rect 6315 9631 6357 9640
rect 7179 9680 7221 9689
rect 7179 9640 7180 9680
rect 7220 9640 7221 9680
rect 7179 9631 7221 9640
rect 7563 9680 7605 9689
rect 7563 9640 7564 9680
rect 7604 9640 7605 9680
rect 7563 9631 7605 9640
rect 8314 9680 8372 9681
rect 8314 9640 8323 9680
rect 8363 9640 8372 9680
rect 8314 9639 8372 9640
rect 9466 9680 9524 9681
rect 9466 9640 9475 9680
rect 9515 9640 9524 9680
rect 9466 9639 9524 9640
rect 11499 9680 11541 9689
rect 11499 9640 11500 9680
rect 11540 9640 11541 9680
rect 11499 9631 11541 9640
rect 12363 9680 12405 9689
rect 12363 9640 12364 9680
rect 12404 9640 12405 9680
rect 12363 9631 12405 9640
rect 13114 9680 13172 9681
rect 13114 9640 13123 9680
rect 13163 9640 13172 9680
rect 13114 9639 13172 9640
rect 13786 9680 13844 9681
rect 13786 9640 13795 9680
rect 13835 9640 13844 9680
rect 13786 9639 13844 9640
rect 13899 9680 13941 9689
rect 13899 9640 13900 9680
rect 13940 9640 13941 9680
rect 13899 9631 13941 9640
rect 14266 9680 14324 9681
rect 14266 9640 14275 9680
rect 14315 9640 14324 9680
rect 14266 9639 14324 9640
rect 15034 9680 15092 9681
rect 15034 9640 15043 9680
rect 15083 9640 15092 9680
rect 15034 9639 15092 9640
rect 16282 9680 16340 9681
rect 16282 9640 16291 9680
rect 16331 9640 16340 9680
rect 16282 9639 16340 9640
rect 18411 9680 18453 9689
rect 18411 9640 18412 9680
rect 18452 9640 18453 9680
rect 18411 9631 18453 9640
rect 18778 9680 18836 9681
rect 18778 9640 18787 9680
rect 18827 9640 18836 9680
rect 18778 9639 18836 9640
rect 19546 9680 19604 9681
rect 19546 9640 19555 9680
rect 19595 9640 19604 9680
rect 19546 9639 19604 9640
rect 21082 9680 21140 9681
rect 21082 9640 21091 9680
rect 21131 9640 21140 9680
rect 21082 9639 21140 9640
rect 22810 9680 22868 9681
rect 22810 9640 22819 9680
rect 22859 9640 22868 9680
rect 22810 9639 22868 9640
rect 24171 9680 24213 9689
rect 24171 9640 24172 9680
rect 24212 9640 24213 9680
rect 24171 9631 24213 9640
rect 25035 9680 25077 9689
rect 25035 9640 25036 9680
rect 25076 9640 25077 9680
rect 25035 9631 25077 9640
rect 26187 9680 26229 9689
rect 26187 9640 26188 9680
rect 26228 9640 26229 9680
rect 26187 9631 26229 9640
rect 1721 9596 1763 9605
rect 1721 9556 1722 9596
rect 1762 9556 1763 9596
rect 1721 9547 1763 9556
rect 2170 9596 2228 9597
rect 2170 9556 2179 9596
rect 2219 9556 2228 9596
rect 2170 9555 2228 9556
rect 7467 9596 7509 9605
rect 7467 9556 7468 9596
rect 7508 9556 7509 9596
rect 7467 9547 7509 9556
rect 8811 9596 8853 9605
rect 8811 9556 8812 9596
rect 8852 9556 8853 9596
rect 8811 9547 8853 9556
rect 10635 9596 10677 9605
rect 10635 9556 10636 9596
rect 10676 9556 10677 9596
rect 10635 9547 10677 9556
rect 22138 9596 22196 9597
rect 22138 9556 22147 9596
rect 22187 9556 22196 9596
rect 22138 9555 22196 9556
rect 651 9512 693 9521
rect 651 9472 652 9512
rect 692 9472 693 9512
rect 651 9463 693 9472
rect 939 9512 981 9521
rect 939 9472 940 9512
rect 980 9472 981 9512
rect 939 9463 981 9472
rect 1131 9512 1173 9521
rect 1131 9472 1132 9512
rect 1172 9472 1173 9512
rect 1131 9463 1173 9472
rect 1402 9512 1460 9513
rect 1402 9472 1411 9512
rect 1451 9472 1460 9512
rect 1402 9471 1460 9472
rect 1515 9512 1557 9521
rect 1515 9472 1516 9512
rect 1556 9472 1557 9512
rect 1515 9463 1557 9472
rect 1846 9512 1888 9521
rect 1846 9472 1847 9512
rect 1887 9472 1888 9512
rect 1846 9463 1888 9472
rect 2091 9512 2133 9521
rect 2091 9472 2092 9512
rect 2132 9472 2133 9512
rect 2091 9463 2133 9472
rect 3051 9512 3093 9521
rect 3051 9472 3052 9512
rect 3092 9472 3093 9512
rect 3051 9463 3093 9472
rect 3435 9512 3477 9521
rect 3435 9472 3436 9512
rect 3476 9472 3477 9512
rect 3435 9463 3477 9472
rect 3723 9512 3765 9521
rect 3723 9472 3724 9512
rect 3764 9472 3765 9512
rect 3723 9463 3765 9472
rect 4378 9512 4436 9513
rect 4378 9472 4387 9512
rect 4427 9472 4436 9512
rect 4378 9471 4436 9472
rect 4491 9512 4533 9521
rect 4491 9472 4492 9512
rect 4532 9472 4533 9512
rect 4491 9463 4533 9472
rect 5259 9512 5301 9521
rect 5259 9472 5260 9512
rect 5300 9472 5301 9512
rect 5259 9463 5301 9472
rect 5835 9512 5877 9521
rect 5835 9472 5836 9512
rect 5876 9472 5877 9512
rect 5835 9463 5877 9472
rect 6219 9512 6261 9521
rect 6219 9472 6220 9512
rect 6260 9472 6261 9512
rect 6219 9463 6261 9472
rect 6778 9512 6836 9513
rect 6778 9472 6787 9512
rect 6827 9472 6836 9512
rect 6778 9471 6836 9472
rect 6891 9512 6933 9521
rect 6891 9472 6892 9512
rect 6932 9472 6933 9512
rect 6891 9463 6933 9472
rect 7354 9512 7412 9513
rect 7354 9472 7363 9512
rect 7403 9472 7412 9512
rect 7354 9471 7412 9472
rect 7670 9512 7712 9521
rect 7670 9472 7671 9512
rect 7711 9472 7712 9512
rect 7670 9463 7712 9472
rect 8235 9512 8277 9521
rect 8235 9472 8236 9512
rect 8276 9472 8277 9512
rect 8235 9463 8277 9472
rect 8698 9512 8756 9513
rect 8698 9472 8707 9512
rect 8747 9472 8756 9512
rect 8698 9471 8756 9472
rect 9014 9512 9056 9521
rect 9014 9472 9015 9512
rect 9055 9472 9056 9512
rect 9014 9463 9056 9472
rect 9142 9512 9184 9521
rect 9142 9472 9143 9512
rect 9183 9472 9184 9512
rect 9142 9463 9184 9472
rect 9387 9512 9429 9521
rect 9387 9472 9388 9512
rect 9428 9472 9429 9512
rect 9387 9463 9429 9472
rect 9730 9512 9788 9513
rect 9730 9472 9739 9512
rect 9779 9472 9788 9512
rect 9730 9471 9788 9472
rect 9963 9512 10005 9521
rect 9963 9472 9964 9512
rect 10004 9472 10005 9512
rect 9963 9463 10005 9472
rect 10426 9512 10484 9513
rect 10426 9472 10435 9512
rect 10475 9472 10484 9512
rect 10426 9471 10484 9472
rect 10731 9512 10773 9521
rect 10731 9472 10732 9512
rect 10772 9472 10773 9512
rect 10731 9463 10773 9472
rect 11019 9512 11061 9521
rect 11019 9472 11020 9512
rect 11060 9472 11061 9512
rect 11019 9463 11061 9472
rect 11403 9512 11445 9521
rect 11403 9472 11404 9512
rect 11444 9472 11445 9512
rect 11403 9463 11445 9472
rect 11962 9512 12020 9513
rect 11962 9472 11971 9512
rect 12011 9472 12020 9512
rect 11962 9471 12020 9472
rect 12075 9512 12117 9521
rect 12075 9472 12076 9512
rect 12116 9472 12117 9512
rect 12075 9463 12117 9472
rect 12507 9512 12549 9521
rect 12507 9472 12508 9512
rect 12548 9472 12549 9512
rect 12962 9512 13004 9521
rect 12507 9463 12549 9472
rect 12815 9470 12857 9479
rect 1978 9428 2036 9429
rect 1978 9388 1987 9428
rect 2027 9388 2036 9428
rect 1978 9387 2036 9388
rect 5169 9428 5211 9437
rect 5169 9388 5170 9428
rect 5210 9388 5211 9428
rect 5169 9379 5211 9388
rect 9274 9428 9332 9429
rect 9274 9388 9283 9428
rect 9323 9388 9332 9428
rect 9274 9387 9332 9388
rect 9850 9428 9908 9429
rect 9850 9388 9859 9428
rect 9899 9388 9908 9428
rect 9850 9387 9908 9388
rect 10059 9428 10101 9437
rect 10059 9388 10060 9428
rect 10100 9388 10101 9428
rect 10059 9379 10101 9388
rect 12651 9428 12693 9437
rect 12651 9388 12652 9428
rect 12692 9388 12693 9428
rect 12815 9430 12816 9470
rect 12856 9430 12857 9470
rect 12962 9472 12963 9512
rect 13003 9472 13004 9512
rect 12962 9463 13004 9472
rect 13275 9512 13317 9521
rect 13275 9472 13276 9512
rect 13316 9472 13317 9512
rect 13275 9463 13317 9472
rect 13419 9512 13461 9521
rect 13419 9472 13420 9512
rect 13460 9472 13461 9512
rect 13419 9463 13461 9472
rect 13693 9512 13735 9521
rect 14475 9512 14517 9521
rect 13693 9472 13694 9512
rect 13734 9472 13735 9512
rect 13693 9463 13735 9472
rect 13995 9503 14037 9512
rect 13995 9463 13996 9503
rect 14036 9463 14037 9503
rect 14475 9472 14476 9512
rect 14516 9472 14517 9512
rect 14475 9463 14517 9472
rect 14763 9512 14805 9521
rect 14763 9472 14764 9512
rect 14804 9472 14805 9512
rect 14763 9463 14805 9472
rect 15243 9512 15285 9521
rect 15243 9472 15244 9512
rect 15284 9472 15285 9512
rect 15243 9463 15285 9472
rect 15531 9512 15573 9521
rect 15531 9472 15532 9512
rect 15572 9472 15573 9512
rect 15531 9463 15573 9472
rect 15766 9512 15808 9521
rect 15766 9472 15767 9512
rect 15807 9472 15808 9512
rect 15766 9463 15808 9472
rect 16011 9512 16053 9521
rect 16011 9472 16012 9512
rect 16052 9472 16053 9512
rect 16011 9463 16053 9472
rect 16443 9512 16485 9521
rect 16443 9472 16444 9512
rect 16484 9472 16485 9512
rect 16443 9463 16485 9472
rect 16587 9512 16629 9521
rect 16587 9472 16588 9512
rect 16628 9472 16629 9512
rect 16587 9463 16629 9472
rect 17211 9512 17253 9521
rect 17211 9472 17212 9512
rect 17252 9472 17253 9512
rect 17211 9463 17253 9472
rect 17355 9512 17397 9521
rect 17355 9472 17356 9512
rect 17396 9472 17397 9512
rect 17355 9463 17397 9472
rect 17547 9512 17589 9521
rect 17547 9472 17548 9512
rect 17588 9472 17589 9512
rect 17547 9463 17589 9472
rect 17722 9512 17780 9513
rect 17722 9472 17731 9512
rect 17771 9472 17780 9512
rect 17722 9471 17780 9472
rect 17931 9512 17973 9521
rect 17931 9472 17932 9512
rect 17972 9472 17973 9512
rect 17931 9463 17973 9472
rect 18315 9512 18357 9521
rect 18315 9472 18316 9512
rect 18356 9472 18357 9512
rect 18315 9463 18357 9472
rect 18972 9512 19014 9521
rect 18972 9472 18973 9512
rect 19013 9472 19014 9512
rect 18972 9463 19014 9472
rect 19083 9512 19125 9521
rect 19083 9472 19084 9512
rect 19124 9472 19125 9512
rect 19083 9463 19125 9472
rect 19707 9512 19749 9521
rect 19707 9472 19708 9512
rect 19748 9472 19749 9512
rect 19707 9463 19749 9472
rect 19851 9512 19893 9521
rect 19851 9472 19852 9512
rect 19892 9472 19893 9512
rect 19851 9463 19893 9472
rect 20619 9512 20661 9521
rect 20619 9472 20620 9512
rect 20660 9472 20661 9512
rect 20619 9463 20661 9472
rect 21387 9512 21429 9521
rect 21387 9472 21388 9512
rect 21428 9472 21429 9512
rect 21387 9463 21429 9472
rect 22539 9512 22581 9521
rect 22539 9472 22540 9512
rect 22580 9472 22581 9512
rect 22539 9463 22581 9472
rect 23110 9512 23168 9513
rect 23110 9472 23119 9512
rect 23159 9472 23168 9512
rect 23110 9471 23168 9472
rect 23770 9512 23828 9513
rect 23770 9472 23779 9512
rect 23819 9472 23828 9512
rect 23770 9471 23828 9472
rect 23883 9512 23925 9521
rect 23883 9472 23884 9512
rect 23924 9472 23925 9512
rect 23883 9463 23925 9472
rect 24634 9512 24692 9513
rect 24634 9472 24643 9512
rect 24683 9472 24692 9512
rect 24634 9471 24692 9472
rect 24747 9512 24789 9521
rect 24747 9472 24748 9512
rect 24788 9472 24789 9512
rect 24747 9463 24789 9472
rect 25402 9512 25460 9513
rect 25402 9472 25411 9512
rect 25451 9472 25460 9512
rect 25402 9471 25460 9472
rect 26091 9512 26133 9521
rect 26091 9472 26092 9512
rect 26132 9472 26133 9512
rect 26091 9463 26133 9472
rect 26266 9512 26324 9513
rect 26266 9472 26275 9512
rect 26315 9472 26324 9512
rect 26266 9471 26324 9472
rect 13995 9454 14037 9463
rect 12815 9421 12857 9430
rect 15898 9428 15956 9429
rect 12651 9379 12693 9388
rect 15898 9388 15907 9428
rect 15947 9388 15956 9428
rect 15898 9387 15956 9388
rect 16107 9428 16149 9437
rect 16107 9388 16108 9428
rect 16148 9388 16149 9428
rect 16107 9379 16149 9388
rect 20529 9428 20571 9437
rect 20529 9388 20530 9428
rect 20570 9388 20571 9428
rect 20529 9379 20571 9388
rect 21297 9428 21339 9437
rect 21297 9388 21298 9428
rect 21338 9388 21339 9428
rect 21297 9379 21339 9388
rect 23025 9428 23067 9437
rect 23025 9388 23026 9428
rect 23066 9388 23067 9428
rect 23025 9379 23067 9388
rect 26475 9428 26517 9437
rect 26475 9388 26476 9428
rect 26516 9388 26517 9428
rect 26475 9379 26517 9388
rect 4666 9344 4724 9345
rect 4666 9304 4675 9344
rect 4715 9304 4724 9344
rect 4666 9303 4724 9304
rect 12747 9344 12789 9353
rect 12747 9304 12748 9344
rect 12788 9304 12789 9344
rect 12747 9295 12789 9304
rect 17002 9344 17060 9345
rect 17002 9304 17011 9344
rect 17051 9304 17060 9344
rect 17002 9303 17060 9304
rect 26715 9344 26757 9353
rect 26715 9304 26716 9344
rect 26756 9304 26757 9344
rect 26715 9295 26757 9304
rect 795 9260 837 9269
rect 795 9220 796 9260
rect 836 9220 837 9260
rect 795 9211 837 9220
rect 1707 9260 1749 9269
rect 1707 9220 1708 9260
rect 1748 9220 1749 9260
rect 1707 9211 1749 9220
rect 2379 9260 2421 9269
rect 2379 9220 2380 9260
rect 2420 9220 2421 9260
rect 2379 9211 2421 9220
rect 4059 9260 4101 9269
rect 4059 9220 4060 9260
rect 4100 9220 4101 9260
rect 4059 9211 4101 9220
rect 7066 9260 7124 9261
rect 7066 9220 7075 9260
rect 7115 9220 7124 9260
rect 7066 9219 7124 9220
rect 8043 9260 8085 9269
rect 8043 9220 8044 9260
rect 8084 9220 8085 9260
rect 8043 9211 8085 9220
rect 9003 9260 9045 9269
rect 9003 9220 9004 9260
rect 9044 9220 9045 9260
rect 9003 9211 9045 9220
rect 17722 9260 17780 9261
rect 17722 9220 17731 9260
rect 17771 9220 17780 9260
rect 17722 9219 17780 9220
rect 20427 9260 20469 9269
rect 20427 9220 20428 9260
rect 20468 9220 20469 9260
rect 20427 9211 20469 9220
rect 25611 9260 25653 9269
rect 25611 9220 25612 9260
rect 25652 9220 25653 9260
rect 25611 9211 25653 9220
rect 576 9092 31392 9116
rect 576 9052 3112 9092
rect 3480 9052 10886 9092
rect 11254 9052 18660 9092
rect 19028 9052 26434 9092
rect 26802 9052 31392 9092
rect 576 9028 31392 9052
rect 2859 8924 2901 8933
rect 2859 8884 2860 8924
rect 2900 8884 2901 8924
rect 2859 8875 2901 8884
rect 3610 8924 3668 8925
rect 3610 8884 3619 8924
rect 3659 8884 3668 8924
rect 3610 8883 3668 8884
rect 5547 8924 5589 8933
rect 5547 8884 5548 8924
rect 5588 8884 5589 8924
rect 5547 8875 5589 8884
rect 6027 8924 6069 8933
rect 6027 8884 6028 8924
rect 6068 8884 6069 8924
rect 6027 8875 6069 8884
rect 7947 8924 7989 8933
rect 7947 8884 7948 8924
rect 7988 8884 7989 8924
rect 7947 8875 7989 8884
rect 12651 8924 12693 8933
rect 12651 8884 12652 8924
rect 12692 8884 12693 8924
rect 12651 8875 12693 8884
rect 16282 8924 16340 8925
rect 16282 8884 16291 8924
rect 16331 8884 16340 8924
rect 16282 8883 16340 8884
rect 17530 8924 17588 8925
rect 17530 8884 17539 8924
rect 17579 8884 17588 8924
rect 17530 8883 17588 8884
rect 18586 8924 18644 8925
rect 18586 8884 18595 8924
rect 18635 8884 18644 8924
rect 18586 8883 18644 8884
rect 20122 8924 20180 8925
rect 20122 8884 20131 8924
rect 20171 8884 20180 8924
rect 20122 8883 20180 8884
rect 21243 8924 21285 8933
rect 21243 8884 21244 8924
rect 21284 8884 21285 8924
rect 21243 8875 21285 8884
rect 21867 8924 21909 8933
rect 21867 8884 21868 8924
rect 21908 8884 21909 8924
rect 21867 8875 21909 8884
rect 23403 8924 23445 8933
rect 23403 8884 23404 8924
rect 23444 8884 23445 8924
rect 23403 8875 23445 8884
rect 25707 8924 25749 8933
rect 25707 8884 25708 8924
rect 25748 8884 25749 8924
rect 25707 8875 25749 8884
rect 5115 8840 5157 8849
rect 6490 8840 6548 8841
rect 5115 8800 5116 8840
rect 5156 8800 5157 8840
rect 5115 8791 5157 8800
rect 6267 8831 6309 8840
rect 6267 8791 6268 8831
rect 6308 8791 6309 8831
rect 6490 8800 6499 8840
rect 6539 8800 6548 8840
rect 6490 8799 6548 8800
rect 9850 8840 9908 8841
rect 9850 8800 9859 8840
rect 9899 8800 9908 8840
rect 9850 8799 9908 8800
rect 13306 8840 13364 8841
rect 13306 8800 13315 8840
rect 13355 8800 13364 8840
rect 13306 8799 13364 8800
rect 14091 8840 14133 8849
rect 14091 8800 14092 8840
rect 14132 8800 14133 8840
rect 14091 8791 14133 8800
rect 24538 8840 24596 8841
rect 24538 8800 24547 8840
rect 24587 8800 24596 8840
rect 24538 8799 24596 8800
rect 26859 8840 26901 8849
rect 26859 8800 26860 8840
rect 26900 8800 26901 8840
rect 26859 8791 26901 8800
rect 6267 8782 6309 8791
rect 939 8756 981 8765
rect 939 8716 940 8756
rect 980 8716 981 8756
rect 939 8707 981 8716
rect 7258 8756 7316 8757
rect 7258 8716 7267 8756
rect 7307 8716 7316 8756
rect 7258 8715 7316 8716
rect 8337 8756 8379 8765
rect 10155 8756 10197 8765
rect 8337 8716 8338 8756
rect 8378 8716 8379 8756
rect 8337 8707 8379 8716
rect 9138 8747 9184 8756
rect 9138 8707 9139 8747
rect 9179 8707 9184 8747
rect 10155 8716 10156 8756
rect 10196 8716 10197 8756
rect 10155 8707 10197 8716
rect 10731 8756 10773 8765
rect 10731 8716 10732 8756
rect 10772 8716 10773 8756
rect 10731 8707 10773 8716
rect 13611 8756 13653 8765
rect 13611 8716 13612 8756
rect 13652 8716 13653 8756
rect 13611 8707 13653 8716
rect 14187 8756 14229 8765
rect 14187 8716 14188 8756
rect 14228 8716 14229 8756
rect 14187 8707 14229 8716
rect 15537 8756 15579 8765
rect 15537 8716 15538 8756
rect 15578 8716 15579 8756
rect 15537 8707 15579 8716
rect 16954 8756 17012 8757
rect 16954 8716 16963 8756
rect 17003 8716 17012 8756
rect 16954 8715 17012 8716
rect 18874 8756 18932 8757
rect 18874 8716 18883 8756
rect 18923 8716 18932 8756
rect 18874 8715 18932 8716
rect 19450 8756 19508 8757
rect 19450 8716 19459 8756
rect 19499 8716 19508 8756
rect 19450 8715 19508 8716
rect 23505 8756 23547 8765
rect 23505 8716 23506 8756
rect 23546 8716 23547 8756
rect 9138 8698 9184 8707
rect 18411 8705 18453 8714
rect 1306 8672 1364 8673
rect 1306 8632 1315 8672
rect 1355 8632 1364 8672
rect 1306 8631 1364 8632
rect 3579 8672 3621 8681
rect 3579 8632 3580 8672
rect 3620 8632 3621 8672
rect 3579 8623 3621 8632
rect 3723 8672 3765 8681
rect 3723 8632 3724 8672
rect 3764 8632 3765 8672
rect 3723 8623 3765 8632
rect 4491 8672 4533 8681
rect 4491 8632 4492 8672
rect 4532 8632 4533 8672
rect 4491 8623 4533 8632
rect 4779 8672 4821 8681
rect 4779 8632 4780 8672
rect 4820 8632 4821 8672
rect 4779 8623 4821 8632
rect 5242 8672 5300 8673
rect 5242 8632 5251 8672
rect 5291 8632 5300 8672
rect 5242 8631 5300 8632
rect 5355 8672 5397 8681
rect 5355 8632 5356 8672
rect 5396 8632 5397 8672
rect 5355 8623 5397 8632
rect 5722 8672 5780 8673
rect 5722 8632 5731 8672
rect 5771 8632 5780 8672
rect 5722 8631 5780 8632
rect 6298 8672 6356 8673
rect 6298 8632 6307 8672
rect 6347 8632 6356 8672
rect 6298 8631 6356 8632
rect 6646 8672 6688 8681
rect 6646 8632 6647 8672
rect 6687 8632 6688 8672
rect 6646 8623 6688 8632
rect 6778 8672 6836 8673
rect 6778 8632 6787 8672
rect 6827 8632 6836 8672
rect 6778 8631 6836 8632
rect 6891 8672 6933 8681
rect 6891 8632 6892 8672
rect 6932 8632 6933 8672
rect 6891 8623 6933 8632
rect 7126 8672 7168 8681
rect 7126 8632 7127 8672
rect 7167 8632 7168 8672
rect 7126 8623 7168 8632
rect 7371 8672 7413 8681
rect 7371 8632 7372 8672
rect 7412 8632 7413 8672
rect 7371 8623 7413 8632
rect 7642 8672 7700 8673
rect 7642 8632 7651 8672
rect 7691 8632 7700 8672
rect 7642 8631 7700 8632
rect 7961 8672 8003 8681
rect 7961 8632 7962 8672
rect 8002 8632 8003 8672
rect 7961 8623 8003 8632
rect 8427 8672 8469 8681
rect 8427 8632 8428 8672
rect 8468 8632 8469 8672
rect 8427 8623 8469 8632
rect 9003 8672 9045 8681
rect 9003 8632 9004 8672
rect 9044 8632 9045 8672
rect 9003 8623 9045 8632
rect 9232 8672 9290 8673
rect 9232 8632 9241 8672
rect 9281 8632 9290 8672
rect 9232 8631 9290 8632
rect 9562 8672 9620 8673
rect 9562 8632 9571 8672
rect 9611 8632 9620 8672
rect 9562 8631 9620 8632
rect 9675 8672 9717 8681
rect 9675 8632 9676 8672
rect 9716 8632 9717 8672
rect 9675 8623 9717 8632
rect 10330 8672 10388 8673
rect 10330 8632 10339 8672
rect 10379 8632 10388 8672
rect 10330 8631 10388 8632
rect 10923 8672 10965 8681
rect 10923 8632 10924 8672
rect 10964 8632 10965 8672
rect 10923 8623 10965 8632
rect 11115 8672 11157 8681
rect 11115 8632 11116 8672
rect 11156 8632 11157 8672
rect 11115 8623 11157 8632
rect 11307 8672 11349 8681
rect 11307 8632 11308 8672
rect 11348 8632 11349 8672
rect 11307 8623 11349 8632
rect 11595 8672 11637 8681
rect 11595 8632 11596 8672
rect 11636 8632 11637 8672
rect 11595 8623 11637 8632
rect 12459 8672 12501 8681
rect 12459 8632 12460 8672
rect 12500 8632 12501 8672
rect 12459 8623 12501 8632
rect 13137 8672 13179 8681
rect 13137 8632 13138 8672
rect 13178 8632 13179 8672
rect 13137 8623 13179 8632
rect 13258 8672 13316 8673
rect 13258 8632 13267 8672
rect 13307 8632 13316 8672
rect 13258 8631 13316 8632
rect 13786 8672 13844 8673
rect 13786 8632 13795 8672
rect 13835 8632 13844 8672
rect 13786 8631 13844 8632
rect 14523 8672 14565 8681
rect 14523 8632 14524 8672
rect 14564 8632 14565 8672
rect 14523 8623 14565 8632
rect 14667 8672 14709 8681
rect 14667 8632 14668 8672
rect 14708 8632 14709 8672
rect 14667 8623 14709 8632
rect 15627 8672 15669 8681
rect 15627 8632 15628 8672
rect 15668 8632 15669 8672
rect 15627 8623 15669 8632
rect 16251 8672 16293 8681
rect 16251 8632 16252 8672
rect 16292 8632 16293 8672
rect 16251 8623 16293 8632
rect 16395 8672 16437 8681
rect 16395 8632 16396 8672
rect 16436 8632 16437 8672
rect 16395 8623 16437 8632
rect 16822 8672 16864 8681
rect 16822 8632 16823 8672
rect 16863 8632 16864 8672
rect 16822 8623 16864 8632
rect 17052 8672 17110 8673
rect 17052 8632 17061 8672
rect 17101 8632 17110 8672
rect 17052 8631 17110 8632
rect 17355 8672 17397 8681
rect 17355 8632 17356 8672
rect 17396 8632 17397 8672
rect 17355 8623 17397 8632
rect 17530 8672 17588 8673
rect 17530 8632 17539 8672
rect 17579 8632 17588 8672
rect 17530 8631 17588 8632
rect 17931 8672 17973 8681
rect 17931 8632 17932 8672
rect 17972 8632 17973 8672
rect 18411 8665 18412 8705
rect 18452 8665 18453 8705
rect 22242 8705 22288 8714
rect 23505 8707 23547 8716
rect 25041 8756 25083 8765
rect 25041 8716 25042 8756
rect 25082 8716 25083 8756
rect 25041 8707 25083 8716
rect 26594 8756 26636 8765
rect 26594 8716 26595 8756
rect 26635 8716 26636 8756
rect 26594 8707 26636 8716
rect 26715 8714 26757 8723
rect 18411 8656 18453 8665
rect 18507 8672 18549 8681
rect 17931 8623 17973 8632
rect 18507 8632 18508 8672
rect 18548 8632 18549 8672
rect 18507 8623 18549 8632
rect 19258 8672 19316 8673
rect 19258 8632 19267 8672
rect 19307 8632 19316 8672
rect 19258 8631 19316 8632
rect 19947 8672 19989 8681
rect 19947 8632 19948 8672
rect 19988 8632 19989 8672
rect 19947 8623 19989 8632
rect 20074 8672 20132 8673
rect 20074 8632 20083 8672
rect 20123 8632 20132 8672
rect 20074 8631 20132 8632
rect 20619 8672 20661 8681
rect 20619 8632 20620 8672
rect 20660 8632 20661 8672
rect 20619 8623 20661 8632
rect 21003 8672 21045 8681
rect 21003 8632 21004 8672
rect 21044 8632 21045 8672
rect 21003 8623 21045 8632
rect 21669 8672 21727 8673
rect 21669 8632 21678 8672
rect 21718 8632 21727 8672
rect 21669 8631 21727 8632
rect 21867 8672 21909 8681
rect 21867 8632 21868 8672
rect 21908 8632 21909 8672
rect 21867 8623 21909 8632
rect 22040 8672 22082 8681
rect 22040 8632 22041 8672
rect 22081 8632 22082 8672
rect 22242 8665 22243 8705
rect 22283 8665 22288 8705
rect 22242 8656 22288 8665
rect 22683 8672 22725 8681
rect 22040 8623 22082 8632
rect 22683 8632 22684 8672
rect 22724 8632 22725 8672
rect 22683 8623 22725 8632
rect 22865 8672 22923 8673
rect 22865 8632 22874 8672
rect 22914 8632 22923 8672
rect 22865 8631 22923 8632
rect 23595 8672 23637 8681
rect 23595 8632 23596 8672
rect 23636 8632 23637 8672
rect 23595 8623 23637 8632
rect 24369 8672 24411 8681
rect 24369 8632 24370 8672
rect 24410 8632 24411 8672
rect 24369 8623 24411 8632
rect 24490 8672 24548 8673
rect 24490 8632 24499 8672
rect 24539 8632 24548 8672
rect 24490 8631 24548 8632
rect 25131 8672 25173 8681
rect 25131 8632 25132 8672
rect 25172 8632 25173 8672
rect 25131 8623 25173 8632
rect 25755 8672 25797 8681
rect 25755 8632 25756 8672
rect 25796 8632 25797 8672
rect 25755 8623 25797 8632
rect 25899 8672 25941 8681
rect 25899 8632 25900 8672
rect 25940 8632 25941 8672
rect 25899 8623 25941 8632
rect 26475 8672 26517 8681
rect 26475 8632 26476 8672
rect 26516 8632 26517 8672
rect 26715 8674 26716 8714
rect 26756 8674 26757 8714
rect 26715 8665 26757 8674
rect 26859 8672 26901 8681
rect 26475 8623 26517 8632
rect 26859 8632 26860 8672
rect 26900 8632 26901 8672
rect 26859 8623 26901 8632
rect 27051 8672 27093 8681
rect 27051 8632 27052 8672
rect 27092 8632 27093 8672
rect 27051 8623 27093 8632
rect 27243 8672 27285 8681
rect 27243 8632 27244 8672
rect 27284 8632 27285 8672
rect 27243 8623 27285 8632
rect 27435 8672 27477 8681
rect 27435 8632 27436 8672
rect 27476 8632 27477 8672
rect 27435 8623 27477 8632
rect 5561 8588 5603 8597
rect 5561 8548 5562 8588
rect 5602 8548 5603 8588
rect 5561 8539 5603 8548
rect 6038 8588 6080 8597
rect 6038 8548 6039 8588
rect 6079 8548 6080 8588
rect 6038 8539 6080 8548
rect 7450 8588 7508 8589
rect 7450 8548 7459 8588
rect 7499 8548 7508 8588
rect 7450 8547 7508 8548
rect 10635 8588 10677 8597
rect 10635 8548 10636 8588
rect 10676 8548 10677 8588
rect 10635 8539 10677 8548
rect 17146 8588 17204 8589
rect 17146 8548 17155 8588
rect 17195 8548 17204 8588
rect 17146 8547 17204 8548
rect 18970 8588 19028 8589
rect 18970 8548 18979 8588
rect 19019 8548 19028 8588
rect 18970 8547 19028 8548
rect 21373 8588 21415 8597
rect 21373 8548 21374 8588
rect 21414 8548 21415 8588
rect 21373 8539 21415 8548
rect 21466 8588 21524 8589
rect 21466 8548 21475 8588
rect 21515 8548 21524 8588
rect 21466 8547 21524 8548
rect 26379 8588 26421 8597
rect 26379 8548 26380 8588
rect 26420 8548 26421 8588
rect 26379 8539 26421 8548
rect 3243 8504 3285 8513
rect 3243 8464 3244 8504
rect 3284 8464 3285 8504
rect 3243 8455 3285 8464
rect 5818 8504 5876 8505
rect 5818 8464 5827 8504
rect 5867 8464 5876 8504
rect 5818 8463 5876 8464
rect 6970 8504 7028 8505
rect 6970 8464 6979 8504
rect 7019 8464 7028 8504
rect 6970 8463 7028 8464
rect 7738 8504 7796 8505
rect 7738 8464 7747 8504
rect 7787 8464 7796 8504
rect 7738 8463 7796 8464
rect 8122 8504 8180 8505
rect 8122 8464 8131 8504
rect 8171 8464 8180 8504
rect 8122 8463 8180 8464
rect 8907 8504 8949 8513
rect 8907 8464 8908 8504
rect 8948 8464 8949 8504
rect 8907 8455 8949 8464
rect 9963 8504 10005 8513
rect 9963 8464 9964 8504
rect 10004 8464 10005 8504
rect 9963 8455 10005 8464
rect 11098 8504 11156 8505
rect 11098 8464 11107 8504
rect 11147 8464 11156 8504
rect 11098 8463 11156 8464
rect 11787 8504 11829 8513
rect 11787 8464 11788 8504
rect 11828 8464 11829 8504
rect 11787 8455 11829 8464
rect 12346 8504 12404 8505
rect 12346 8464 12355 8504
rect 12395 8464 12404 8504
rect 12346 8463 12404 8464
rect 14362 8504 14420 8505
rect 14362 8464 14371 8504
rect 14411 8464 14420 8504
rect 14362 8463 14420 8464
rect 15322 8504 15380 8505
rect 15322 8464 15331 8504
rect 15371 8464 15380 8504
rect 15322 8463 15380 8464
rect 17787 8504 17829 8513
rect 17787 8464 17788 8504
rect 17828 8464 17829 8504
rect 17787 8455 17829 8464
rect 21579 8504 21621 8513
rect 21579 8464 21580 8504
rect 21620 8464 21621 8504
rect 21579 8455 21621 8464
rect 22395 8504 22437 8513
rect 22395 8464 22396 8504
rect 22436 8464 22437 8504
rect 22395 8455 22437 8464
rect 23019 8504 23061 8513
rect 23019 8464 23020 8504
rect 23060 8464 23061 8504
rect 23019 8455 23061 8464
rect 24826 8504 24884 8505
rect 24826 8464 24835 8504
rect 24875 8464 24884 8504
rect 24826 8463 24884 8464
rect 27243 8504 27285 8513
rect 27243 8464 27244 8504
rect 27284 8464 27285 8504
rect 27243 8455 27285 8464
rect 576 8336 31392 8360
rect 576 8296 4352 8336
rect 4720 8296 12126 8336
rect 12494 8296 19900 8336
rect 20268 8296 27674 8336
rect 28042 8296 31392 8336
rect 576 8272 31392 8296
rect 1210 8168 1268 8169
rect 1210 8128 1219 8168
rect 1259 8128 1268 8168
rect 1210 8127 1268 8128
rect 3531 8168 3573 8177
rect 3531 8128 3532 8168
rect 3572 8128 3573 8168
rect 3531 8119 3573 8128
rect 3867 8168 3909 8177
rect 3867 8128 3868 8168
rect 3908 8128 3909 8168
rect 3867 8119 3909 8128
rect 4395 8168 4437 8177
rect 4395 8128 4396 8168
rect 4436 8128 4437 8168
rect 4395 8119 4437 8128
rect 5259 8168 5301 8177
rect 5259 8128 5260 8168
rect 5300 8128 5301 8168
rect 5259 8119 5301 8128
rect 5626 8168 5684 8169
rect 5626 8128 5635 8168
rect 5675 8128 5684 8168
rect 5626 8127 5684 8128
rect 6795 8168 6837 8177
rect 6795 8128 6796 8168
rect 6836 8128 6837 8168
rect 6795 8119 6837 8128
rect 7755 8168 7797 8177
rect 7755 8128 7756 8168
rect 7796 8128 7797 8168
rect 7755 8119 7797 8128
rect 8715 8168 8757 8177
rect 8715 8128 8716 8168
rect 8756 8128 8757 8168
rect 8715 8119 8757 8128
rect 9483 8168 9525 8177
rect 9483 8128 9484 8168
rect 9524 8128 9525 8168
rect 9483 8119 9525 8128
rect 9754 8168 9812 8169
rect 9754 8128 9763 8168
rect 9803 8128 9812 8168
rect 9754 8127 9812 8128
rect 10635 8168 10677 8177
rect 10635 8128 10636 8168
rect 10676 8128 10677 8168
rect 10635 8119 10677 8128
rect 11386 8168 11444 8169
rect 11386 8128 11395 8168
rect 11435 8128 11444 8168
rect 11386 8127 11444 8128
rect 12106 8168 12164 8169
rect 12106 8128 12115 8168
rect 12155 8128 12164 8168
rect 12106 8127 12164 8128
rect 13611 8168 13653 8177
rect 13611 8128 13612 8168
rect 13652 8128 13653 8168
rect 13611 8119 13653 8128
rect 14187 8168 14229 8177
rect 14187 8128 14188 8168
rect 14228 8128 14229 8168
rect 14187 8119 14229 8128
rect 14859 8168 14901 8177
rect 14859 8128 14860 8168
rect 14900 8128 14901 8168
rect 14859 8119 14901 8128
rect 16395 8168 16437 8177
rect 16395 8128 16396 8168
rect 16436 8128 16437 8168
rect 16395 8119 16437 8128
rect 16666 8168 16724 8169
rect 16666 8128 16675 8168
rect 16715 8128 16724 8168
rect 16666 8127 16724 8128
rect 17626 8168 17684 8169
rect 17626 8128 17635 8168
rect 17675 8128 17684 8168
rect 17626 8127 17684 8128
rect 18891 8168 18933 8177
rect 18891 8128 18892 8168
rect 18932 8128 18933 8168
rect 18891 8119 18933 8128
rect 21195 8168 21237 8177
rect 21195 8128 21196 8168
rect 21236 8128 21237 8168
rect 21195 8119 21237 8128
rect 21562 8168 21620 8169
rect 21562 8128 21571 8168
rect 21611 8128 21620 8168
rect 21562 8127 21620 8128
rect 23290 8168 23348 8169
rect 23290 8128 23299 8168
rect 23339 8128 23348 8168
rect 23290 8127 23348 8128
rect 25786 8168 25844 8169
rect 25786 8128 25795 8168
rect 25835 8128 25844 8168
rect 25786 8127 25844 8128
rect 25899 8168 25941 8177
rect 25899 8128 25900 8168
rect 25940 8128 25941 8168
rect 25899 8119 25941 8128
rect 26266 8168 26324 8169
rect 26266 8128 26275 8168
rect 26315 8128 26324 8168
rect 26266 8127 26324 8128
rect 5056 8084 5098 8093
rect 5056 8044 5057 8084
rect 5097 8044 5098 8084
rect 5056 8035 5098 8044
rect 10432 8084 10474 8093
rect 10432 8044 10433 8084
rect 10473 8044 10474 8084
rect 10432 8035 10474 8044
rect 15147 8084 15189 8093
rect 15147 8044 15148 8084
rect 15188 8044 15189 8084
rect 15147 8035 15189 8044
rect 23200 8084 23242 8093
rect 23200 8044 23201 8084
rect 23241 8044 23242 8084
rect 23200 8035 23242 8044
rect 23691 8084 23733 8093
rect 23691 8044 23692 8084
rect 23732 8044 23733 8084
rect 23691 8035 23733 8044
rect 26379 8084 26421 8093
rect 26379 8044 26380 8084
rect 26420 8044 26421 8084
rect 26379 8035 26421 8044
rect 651 8000 693 8009
rect 651 7960 652 8000
rect 692 7960 693 8000
rect 651 7951 693 7960
rect 843 8000 885 8009
rect 843 7960 844 8000
rect 884 7960 885 8000
rect 843 7951 885 7960
rect 1035 8000 1077 8009
rect 1035 7960 1036 8000
rect 1076 7960 1077 8000
rect 1035 7951 1077 7960
rect 1226 8000 1268 8009
rect 1226 7960 1227 8000
rect 1267 7960 1268 8000
rect 1226 7951 1268 7960
rect 1402 8000 1444 8009
rect 1402 7960 1403 8000
rect 1443 7960 1444 8000
rect 1402 7951 1444 7960
rect 1611 8000 1653 8009
rect 1611 7960 1612 8000
rect 1652 7960 1653 8000
rect 1611 7951 1653 7960
rect 2091 8000 2133 8009
rect 2091 7960 2092 8000
rect 2132 7960 2133 8000
rect 2091 7951 2133 7960
rect 2283 8000 2325 8009
rect 2283 7960 2284 8000
rect 2324 7960 2325 8000
rect 2283 7951 2325 7960
rect 2602 8000 2660 8001
rect 2602 7960 2611 8000
rect 2651 7960 2660 8000
rect 2602 7959 2660 7960
rect 2797 8000 2855 8001
rect 2797 7960 2806 8000
rect 2846 7960 2855 8000
rect 2797 7959 2855 7960
rect 3130 8000 3188 8001
rect 3130 7960 3139 8000
rect 3179 7960 3188 8000
rect 3130 7959 3188 7960
rect 3243 8000 3285 8009
rect 4491 8000 4533 8009
rect 3243 7960 3244 8000
rect 3284 7960 3285 8000
rect 3243 7951 3285 7960
rect 3714 7991 3760 8000
rect 3714 7951 3715 7991
rect 3755 7951 3760 7991
rect 4491 7960 4492 8000
rect 4532 7960 4533 8000
rect 3714 7942 3760 7951
rect 4282 7958 4340 7959
rect 747 7916 789 7925
rect 4282 7918 4291 7958
rect 4331 7918 4340 7958
rect 4491 7951 4533 7960
rect 4603 8000 4661 8001
rect 5835 8000 5877 8009
rect 4603 7960 4612 8000
rect 4652 7960 4661 8000
rect 4603 7959 4661 7960
rect 5355 7991 5397 8000
rect 5355 7951 5356 7991
rect 5396 7951 5397 7991
rect 5835 7960 5836 8000
rect 5876 7960 5877 8000
rect 5835 7951 5877 7960
rect 6123 8000 6165 8009
rect 6123 7960 6124 8000
rect 6164 7960 6165 8000
rect 6123 7951 6165 7960
rect 6315 8000 6357 8009
rect 6315 7960 6316 8000
rect 6356 7960 6357 8000
rect 6315 7951 6357 7960
rect 6603 8000 6645 8009
rect 6603 7960 6604 8000
rect 6644 7960 6645 8000
rect 6603 7951 6645 7960
rect 7354 8000 7412 8001
rect 7354 7960 7363 8000
rect 7403 7960 7412 8000
rect 7354 7959 7412 7960
rect 8314 8000 8372 8001
rect 8314 7960 8323 8000
rect 8363 7960 8372 8000
rect 8314 7959 8372 7960
rect 8427 8000 8469 8009
rect 8427 7960 8428 8000
rect 8468 7960 8469 8000
rect 8427 7951 8469 7960
rect 9082 8000 9140 8001
rect 9082 7960 9091 8000
rect 9131 7960 9140 8000
rect 9082 7959 9140 7960
rect 9195 8000 9237 8009
rect 9195 7960 9196 8000
rect 9236 7960 9237 8000
rect 9195 7951 9237 7960
rect 9963 8000 10005 8009
rect 9963 7960 9964 8000
rect 10004 7960 10005 8000
rect 9963 7951 10005 7960
rect 10251 8000 10293 8009
rect 10870 8000 10912 8009
rect 10251 7960 10252 8000
rect 10292 7960 10293 8000
rect 10251 7951 10293 7960
rect 10731 7991 10773 8000
rect 10731 7951 10732 7991
rect 10772 7951 10773 7991
rect 10870 7960 10871 8000
rect 10911 7960 10912 8000
rect 10870 7951 10912 7960
rect 11115 8000 11157 8009
rect 11115 7960 11116 8000
rect 11156 7960 11157 8000
rect 11115 7951 11157 7960
rect 11580 8000 11622 8009
rect 11580 7960 11581 8000
rect 11621 7960 11622 8000
rect 11580 7951 11622 7960
rect 11691 8000 11733 8009
rect 11691 7960 11692 8000
rect 11732 7960 11733 8000
rect 11691 7951 11733 7960
rect 12250 8000 12308 8001
rect 13131 8000 13173 8009
rect 12250 7960 12259 8000
rect 12299 7960 12308 8000
rect 12250 7959 12308 7960
rect 12363 7991 12405 8000
rect 12363 7951 12364 7991
rect 12404 7951 12405 7991
rect 13131 7960 13132 8000
rect 13172 7960 13173 8000
rect 13131 7951 13173 7960
rect 13419 8000 13461 8009
rect 13419 7960 13420 8000
rect 13460 7960 13461 8000
rect 13419 7951 13461 7960
rect 14283 8000 14325 8009
rect 14283 7960 14284 8000
rect 14324 7960 14325 8000
rect 14283 7951 14325 7960
rect 14514 8000 14556 8009
rect 14514 7960 14515 8000
rect 14555 7960 14556 8000
rect 14514 7951 14556 7960
rect 14656 8000 14698 8009
rect 15472 8000 15530 8001
rect 14656 7960 14657 8000
rect 14697 7960 14698 8000
rect 14656 7951 14698 7960
rect 14955 7991 14997 8000
rect 14955 7951 14956 7991
rect 14996 7951 14997 7991
rect 15378 7991 15424 8000
rect 5355 7942 5397 7951
rect 10731 7942 10773 7951
rect 12363 7942 12405 7951
rect 14955 7942 14997 7951
rect 15243 7958 15285 7967
rect 4282 7917 4340 7918
rect 747 7876 748 7916
rect 788 7876 789 7916
rect 11002 7916 11060 7917
rect 747 7867 789 7876
rect 7306 7888 7364 7889
rect 7306 7848 7315 7888
rect 7355 7848 7364 7888
rect 11002 7876 11011 7916
rect 11051 7876 11060 7916
rect 11002 7875 11060 7876
rect 11211 7916 11253 7925
rect 15243 7918 15244 7958
rect 15284 7918 15285 7958
rect 15378 7951 15379 7991
rect 15419 7951 15424 7991
rect 15472 7960 15481 8000
rect 15521 7960 15530 8000
rect 15472 7959 15530 7960
rect 15994 8000 16052 8001
rect 15994 7960 16003 8000
rect 16043 7960 16052 8000
rect 15994 7959 16052 7960
rect 16107 8000 16149 8009
rect 16107 7960 16108 8000
rect 16148 7960 16149 8000
rect 16107 7951 16149 7960
rect 16875 8000 16917 8009
rect 16875 7960 16876 8000
rect 16916 7960 16917 8000
rect 16875 7951 16917 7960
rect 17163 8000 17205 8009
rect 17163 7960 17164 8000
rect 17204 7960 17205 8000
rect 17163 7951 17205 7960
rect 17739 8000 17781 8009
rect 17739 7960 17740 8000
rect 17780 7960 17781 8000
rect 17739 7951 17781 7960
rect 18123 8000 18165 8009
rect 18123 7960 18124 8000
rect 18164 7960 18165 8000
rect 18123 7951 18165 7960
rect 18490 8000 18548 8001
rect 18490 7960 18499 8000
rect 18539 7960 18548 8000
rect 18490 7959 18548 7960
rect 18603 8000 18645 8009
rect 18603 7960 18604 8000
rect 18644 7960 18645 8000
rect 18603 7951 18645 7960
rect 19083 8000 19125 8009
rect 19083 7960 19084 8000
rect 19124 7960 19125 8000
rect 19083 7951 19125 7960
rect 19258 8000 19316 8001
rect 19258 7960 19267 8000
rect 19307 7960 19316 8000
rect 19258 7959 19316 7960
rect 19759 8000 19817 8001
rect 19759 7960 19768 8000
rect 19808 7960 19817 8000
rect 19759 7959 19817 7960
rect 20314 8000 20372 8001
rect 20314 7960 20323 8000
rect 20363 7960 20372 8000
rect 20314 7959 20372 7960
rect 20427 8000 20469 8009
rect 20427 7960 20428 8000
rect 20468 7960 20469 8000
rect 20427 7951 20469 7960
rect 20907 8000 20949 8009
rect 20907 7960 20908 8000
rect 20948 7960 20949 8000
rect 21723 8000 21765 8009
rect 20907 7951 20949 7960
rect 21035 7976 21077 7985
rect 15378 7942 15424 7951
rect 21035 7936 21036 7976
rect 21076 7936 21077 7976
rect 21723 7960 21724 8000
rect 21764 7960 21765 8000
rect 21723 7951 21765 7960
rect 21867 8000 21909 8009
rect 21867 7960 21868 8000
rect 21908 7960 21909 8000
rect 21867 7951 21909 7960
rect 22347 8000 22389 8009
rect 22347 7960 22348 8000
rect 22388 7960 22389 8000
rect 22347 7951 22389 7960
rect 22491 8000 22533 8009
rect 22491 7960 22492 8000
rect 22532 7960 22533 8000
rect 22491 7951 22533 7960
rect 22635 8000 22677 8009
rect 22635 7960 22636 8000
rect 22676 7960 22677 8000
rect 22635 7951 22677 7960
rect 23403 8000 23445 8009
rect 23787 8000 23829 8009
rect 23403 7960 23404 8000
rect 23444 7960 23445 8000
rect 23403 7951 23445 7960
rect 23499 7991 23541 8000
rect 23499 7951 23500 7991
rect 23540 7951 23541 7991
rect 23787 7960 23788 8000
rect 23828 7960 23829 8000
rect 23787 7951 23829 7960
rect 24016 8000 24074 8001
rect 24016 7960 24025 8000
rect 24065 7960 24074 8000
rect 24016 7959 24074 7960
rect 24132 8000 24174 8009
rect 24132 7960 24133 8000
rect 24173 7960 24174 8000
rect 24132 7951 24174 7960
rect 24363 8000 24405 8009
rect 24363 7960 24364 8000
rect 24404 7960 24405 8000
rect 24363 7951 24405 7960
rect 24843 8000 24885 8009
rect 24843 7960 24844 8000
rect 24884 7960 24885 8000
rect 24843 7951 24885 7960
rect 25693 8000 25735 8009
rect 26176 8000 26218 8009
rect 26614 8000 26656 8009
rect 25693 7960 25694 8000
rect 25734 7960 25735 8000
rect 25693 7951 25735 7960
rect 25995 7991 26037 8000
rect 25995 7951 25996 7991
rect 26036 7951 26037 7991
rect 26176 7960 26177 8000
rect 26217 7960 26218 8000
rect 26176 7951 26218 7960
rect 26477 7991 26519 8000
rect 26477 7951 26478 7991
rect 26518 7951 26519 7991
rect 26614 7960 26615 8000
rect 26655 7960 26656 8000
rect 26614 7951 26656 7960
rect 26859 8000 26901 8009
rect 26859 7960 26860 8000
rect 26900 7960 26901 8000
rect 26859 7951 26901 7960
rect 23499 7942 23541 7951
rect 25995 7942 26037 7951
rect 26477 7942 26519 7951
rect 21035 7927 21077 7936
rect 11211 7876 11212 7916
rect 11252 7876 11253 7916
rect 11211 7867 11253 7876
rect 14418 7907 14464 7916
rect 15243 7909 15285 7918
rect 19594 7916 19652 7917
rect 14418 7867 14419 7907
rect 14459 7867 14464 7907
rect 19594 7876 19603 7916
rect 19643 7876 19652 7916
rect 19594 7875 19652 7876
rect 23906 7916 23948 7925
rect 23906 7876 23907 7916
rect 23947 7876 23948 7916
rect 23906 7867 23948 7876
rect 24250 7916 24308 7917
rect 24250 7876 24259 7916
rect 24299 7876 24308 7916
rect 24250 7875 24308 7876
rect 24459 7916 24501 7925
rect 24459 7876 24460 7916
rect 24500 7876 24501 7916
rect 24459 7867 24501 7876
rect 26746 7916 26804 7917
rect 26746 7876 26755 7916
rect 26795 7876 26804 7916
rect 26746 7875 26804 7876
rect 26955 7916 26997 7925
rect 26955 7876 26956 7916
rect 26996 7876 26997 7916
rect 26955 7867 26997 7876
rect 14418 7858 14464 7867
rect 7306 7847 7364 7848
rect 27147 7832 27189 7841
rect 27147 7792 27148 7832
rect 27188 7792 27189 7832
rect 27147 7783 27189 7792
rect 1515 7748 1557 7757
rect 1515 7708 1516 7748
rect 1556 7708 1557 7748
rect 1515 7699 1557 7708
rect 2187 7748 2229 7757
rect 2187 7708 2188 7748
rect 2228 7708 2229 7748
rect 2187 7699 2229 7708
rect 4779 7748 4821 7757
rect 4779 7708 4780 7748
rect 4820 7708 4821 7748
rect 4779 7699 4821 7708
rect 5050 7748 5108 7749
rect 5050 7708 5059 7748
rect 5099 7708 5108 7748
rect 5050 7707 5108 7708
rect 7546 7748 7604 7749
rect 7546 7708 7555 7748
rect 7595 7708 7604 7748
rect 7546 7707 7604 7708
rect 10426 7748 10484 7749
rect 10426 7708 10435 7748
rect 10475 7708 10484 7748
rect 10426 7707 10484 7708
rect 11499 7748 11541 7757
rect 11499 7708 11500 7748
rect 11540 7708 11541 7748
rect 11499 7699 11541 7708
rect 12651 7748 12693 7757
rect 12651 7708 12652 7748
rect 12692 7708 12693 7748
rect 12651 7699 12693 7708
rect 14650 7748 14708 7749
rect 14650 7708 14659 7748
rect 14699 7708 14708 7748
rect 14650 7707 14708 7708
rect 19258 7748 19316 7749
rect 19258 7708 19267 7748
rect 19307 7708 19316 7748
rect 19258 7707 19316 7708
rect 20523 7748 20565 7757
rect 20523 7708 20524 7748
rect 20564 7708 20565 7748
rect 20523 7699 20565 7708
rect 21754 7748 21812 7749
rect 21754 7708 21763 7748
rect 21803 7708 21812 7748
rect 21754 7707 21812 7708
rect 22827 7748 22869 7757
rect 22827 7708 22828 7748
rect 22868 7708 22869 7748
rect 22827 7699 22869 7708
rect 25515 7748 25557 7757
rect 25515 7708 25516 7748
rect 25556 7708 25557 7748
rect 25515 7699 25557 7708
rect 576 7580 31392 7604
rect 576 7540 3112 7580
rect 3480 7540 10886 7580
rect 11254 7540 18660 7580
rect 19028 7540 26434 7580
rect 26802 7540 31392 7580
rect 576 7516 31392 7540
rect 747 7412 789 7421
rect 747 7372 748 7412
rect 788 7372 789 7412
rect 747 7363 789 7372
rect 3243 7412 3285 7421
rect 3243 7372 3244 7412
rect 3284 7372 3285 7412
rect 3243 7363 3285 7372
rect 5338 7412 5396 7413
rect 5338 7372 5347 7412
rect 5387 7372 5396 7412
rect 5338 7371 5396 7372
rect 8763 7412 8805 7421
rect 8763 7372 8764 7412
rect 8804 7372 8805 7412
rect 8763 7363 8805 7372
rect 9579 7412 9621 7421
rect 9579 7372 9580 7412
rect 9620 7372 9621 7412
rect 9579 7363 9621 7372
rect 12699 7412 12741 7421
rect 12699 7372 12700 7412
rect 12740 7372 12741 7412
rect 12699 7363 12741 7372
rect 13978 7412 14036 7413
rect 13978 7372 13987 7412
rect 14027 7372 14036 7412
rect 13978 7371 14036 7372
rect 14554 7412 14612 7413
rect 14554 7372 14563 7412
rect 14603 7372 14612 7412
rect 14554 7371 14612 7372
rect 16587 7412 16629 7421
rect 16587 7372 16588 7412
rect 16628 7372 16629 7412
rect 16587 7363 16629 7372
rect 17979 7412 18021 7421
rect 17979 7372 17980 7412
rect 18020 7372 18021 7412
rect 17979 7363 18021 7372
rect 18747 7412 18789 7421
rect 18747 7372 18748 7412
rect 18788 7372 18789 7412
rect 18747 7363 18789 7372
rect 20523 7412 20565 7421
rect 20523 7372 20524 7412
rect 20564 7372 20565 7412
rect 20523 7363 20565 7372
rect 22827 7412 22869 7421
rect 22827 7372 22828 7412
rect 22868 7372 22869 7412
rect 22827 7363 22869 7372
rect 26091 7412 26133 7421
rect 26091 7372 26092 7412
rect 26132 7372 26133 7412
rect 26091 7363 26133 7372
rect 1035 7328 1077 7337
rect 1035 7288 1036 7328
rect 1076 7288 1077 7328
rect 1035 7279 1077 7288
rect 4491 7328 4533 7337
rect 4491 7288 4492 7328
rect 4532 7288 4533 7328
rect 4491 7279 4533 7288
rect 16347 7328 16389 7337
rect 16347 7288 16348 7328
rect 16388 7288 16389 7328
rect 16347 7279 16389 7288
rect 21483 7328 21525 7337
rect 21483 7288 21484 7328
rect 21524 7288 21525 7328
rect 21483 7279 21525 7288
rect 6315 7244 6357 7253
rect 5979 7202 6021 7211
rect 2959 7193 3001 7202
rect 651 7160 693 7169
rect 651 7120 652 7160
rect 692 7120 693 7160
rect 651 7111 693 7120
rect 848 7160 890 7169
rect 848 7120 849 7160
rect 889 7120 890 7160
rect 848 7111 890 7120
rect 1035 7160 1077 7169
rect 1035 7120 1036 7160
rect 1076 7120 1077 7160
rect 1035 7111 1077 7120
rect 1225 7160 1267 7169
rect 1225 7120 1226 7160
rect 1266 7120 1267 7160
rect 1225 7111 1267 7120
rect 1419 7160 1461 7169
rect 1419 7120 1420 7160
rect 1460 7120 1461 7160
rect 1419 7111 1461 7120
rect 1611 7160 1653 7169
rect 1611 7120 1612 7160
rect 1652 7120 1653 7160
rect 1611 7111 1653 7120
rect 1899 7160 1941 7169
rect 1899 7120 1900 7160
rect 1940 7120 1941 7160
rect 1899 7111 1941 7120
rect 2283 7160 2325 7169
rect 2283 7120 2284 7160
rect 2324 7120 2325 7160
rect 2283 7111 2325 7120
rect 2417 7160 2475 7161
rect 2417 7120 2426 7160
rect 2466 7120 2475 7160
rect 2417 7119 2475 7120
rect 2842 7160 2900 7161
rect 2842 7120 2851 7160
rect 2891 7120 2900 7160
rect 2959 7153 2960 7193
rect 3000 7153 3001 7193
rect 2959 7144 3001 7153
rect 3478 7160 3520 7169
rect 2842 7119 2900 7120
rect 3478 7120 3479 7160
rect 3519 7120 3520 7160
rect 3478 7111 3520 7120
rect 3610 7160 3668 7161
rect 3610 7120 3619 7160
rect 3659 7120 3668 7160
rect 3610 7119 3668 7120
rect 3723 7160 3765 7169
rect 3723 7120 3724 7160
rect 3764 7120 3765 7160
rect 3723 7111 3765 7120
rect 4107 7160 4149 7169
rect 4107 7120 4108 7160
rect 4148 7120 4149 7160
rect 4107 7111 4149 7120
rect 5050 7160 5108 7161
rect 5050 7120 5059 7160
rect 5099 7120 5108 7160
rect 5050 7119 5108 7120
rect 5163 7160 5205 7169
rect 5163 7120 5164 7160
rect 5204 7120 5205 7160
rect 5163 7111 5205 7120
rect 5643 7160 5685 7169
rect 5643 7120 5644 7160
rect 5684 7120 5685 7160
rect 5643 7111 5685 7120
rect 5835 7160 5877 7169
rect 5835 7120 5836 7160
rect 5876 7120 5877 7160
rect 5979 7162 5980 7202
rect 6020 7162 6021 7202
rect 6315 7204 6316 7244
rect 6356 7204 6357 7244
rect 6315 7195 6357 7204
rect 7546 7244 7604 7245
rect 7546 7204 7555 7244
rect 7595 7204 7604 7244
rect 7546 7203 7604 7204
rect 7755 7244 7797 7253
rect 7755 7204 7756 7244
rect 7796 7204 7797 7244
rect 7755 7195 7797 7204
rect 9003 7244 9045 7253
rect 9003 7204 9004 7244
rect 9044 7204 9045 7244
rect 9003 7195 9045 7204
rect 11595 7244 11637 7253
rect 11595 7204 11596 7244
rect 11636 7204 11637 7244
rect 11595 7195 11637 7204
rect 19732 7244 19774 7253
rect 19732 7204 19733 7244
rect 19773 7204 19774 7244
rect 19732 7195 19774 7204
rect 21003 7244 21045 7253
rect 21003 7204 21004 7244
rect 21044 7204 21045 7244
rect 21003 7195 21045 7204
rect 23133 7202 23191 7203
rect 5979 7153 6021 7162
rect 6106 7160 6164 7161
rect 5835 7111 5877 7120
rect 6106 7120 6115 7160
rect 6155 7120 6164 7160
rect 6106 7119 6164 7120
rect 6219 7160 6261 7169
rect 6219 7120 6220 7160
rect 6260 7120 6261 7160
rect 6219 7111 6261 7120
rect 6603 7160 6645 7169
rect 6603 7120 6604 7160
rect 6644 7120 6645 7160
rect 6603 7111 6645 7120
rect 7414 7160 7456 7169
rect 7414 7120 7415 7160
rect 7455 7120 7456 7160
rect 7414 7111 7456 7120
rect 7659 7160 7701 7169
rect 7659 7120 7660 7160
rect 7700 7120 7701 7160
rect 7659 7111 7701 7120
rect 8139 7160 8181 7169
rect 8139 7120 8140 7160
rect 8180 7120 8181 7160
rect 8139 7111 8181 7120
rect 8427 7160 8469 7169
rect 8427 7120 8428 7160
rect 8468 7120 8469 7160
rect 8427 7111 8469 7120
rect 9099 7160 9141 7169
rect 9099 7120 9100 7160
rect 9140 7120 9141 7160
rect 9099 7111 9141 7120
rect 9218 7160 9260 7169
rect 9218 7120 9219 7160
rect 9259 7120 9260 7160
rect 9218 7111 9260 7120
rect 9328 7160 9386 7161
rect 9328 7120 9337 7160
rect 9377 7120 9386 7160
rect 9328 7119 9386 7120
rect 9627 7160 9669 7169
rect 9627 7120 9628 7160
rect 9668 7120 9669 7160
rect 9627 7111 9669 7120
rect 9771 7160 9813 7169
rect 9771 7120 9772 7160
rect 9812 7120 9813 7160
rect 9771 7111 9813 7120
rect 10443 7160 10485 7169
rect 10443 7120 10444 7160
rect 10484 7120 10485 7160
rect 10443 7111 10485 7120
rect 11002 7160 11060 7161
rect 11002 7120 11011 7160
rect 11051 7120 11060 7160
rect 11002 7119 11060 7120
rect 11115 7160 11157 7169
rect 11115 7120 11116 7160
rect 11156 7120 11157 7160
rect 11115 7111 11157 7120
rect 11691 7160 11733 7169
rect 11691 7120 11692 7160
rect 11732 7120 11733 7160
rect 11691 7111 11733 7120
rect 11810 7160 11852 7169
rect 11810 7120 11811 7160
rect 11851 7120 11852 7160
rect 11810 7111 11852 7120
rect 11920 7160 11978 7161
rect 11920 7120 11929 7160
rect 11969 7120 11978 7160
rect 11920 7119 11978 7120
rect 12075 7160 12117 7169
rect 12075 7120 12076 7160
rect 12116 7120 12117 7160
rect 12075 7111 12117 7120
rect 12363 7160 12405 7169
rect 12363 7120 12364 7160
rect 12404 7120 12405 7160
rect 12363 7111 12405 7120
rect 13210 7160 13268 7161
rect 13210 7120 13219 7160
rect 13259 7120 13268 7160
rect 13210 7119 13268 7120
rect 13323 7160 13365 7169
rect 13323 7120 13324 7160
rect 13364 7120 13365 7160
rect 13323 7111 13365 7120
rect 13947 7160 13989 7169
rect 13947 7120 13948 7160
rect 13988 7120 13989 7160
rect 13947 7111 13989 7120
rect 14091 7160 14133 7169
rect 14091 7120 14092 7160
rect 14132 7120 14133 7160
rect 14091 7111 14133 7120
rect 14853 7160 14911 7161
rect 14853 7120 14862 7160
rect 14902 7120 14911 7160
rect 14853 7119 14911 7120
rect 15435 7160 15477 7169
rect 15435 7120 15436 7160
rect 15476 7120 15477 7160
rect 15435 7111 15477 7120
rect 15523 7160 15581 7161
rect 15523 7120 15532 7160
rect 15572 7120 15581 7160
rect 15523 7119 15581 7120
rect 15723 7160 15765 7169
rect 15723 7120 15724 7160
rect 15764 7120 15765 7160
rect 15723 7111 15765 7120
rect 16011 7160 16053 7169
rect 16011 7120 16012 7160
rect 16052 7120 16053 7160
rect 16011 7111 16053 7120
rect 16635 7160 16677 7169
rect 16635 7120 16636 7160
rect 16676 7120 16677 7160
rect 16635 7111 16677 7120
rect 16779 7160 16821 7169
rect 16779 7120 16780 7160
rect 16820 7120 16821 7160
rect 16779 7111 16821 7120
rect 17355 7160 17397 7169
rect 17355 7120 17356 7160
rect 17396 7120 17397 7160
rect 17355 7111 17397 7120
rect 17739 7160 17781 7169
rect 17739 7120 17740 7160
rect 17780 7120 17781 7160
rect 17739 7111 17781 7120
rect 18123 7160 18165 7169
rect 18123 7120 18124 7160
rect 18164 7120 18165 7160
rect 18123 7111 18165 7120
rect 18507 7160 18549 7169
rect 18507 7120 18508 7160
rect 18548 7120 18549 7160
rect 18507 7111 18549 7120
rect 18874 7160 18932 7161
rect 18874 7120 18883 7160
rect 18923 7120 18932 7160
rect 18874 7119 18932 7120
rect 18992 7160 19050 7161
rect 18992 7120 19001 7160
rect 19041 7120 19050 7160
rect 18992 7119 19050 7120
rect 19158 7160 19216 7161
rect 19158 7120 19167 7160
rect 19207 7120 19216 7160
rect 19158 7119 19216 7120
rect 19270 7160 19312 7169
rect 19270 7120 19271 7160
rect 19311 7120 19312 7160
rect 19270 7111 19312 7120
rect 19392 7160 19450 7161
rect 19392 7120 19401 7160
rect 19441 7120 19450 7160
rect 19392 7119 19450 7120
rect 19611 7160 19653 7169
rect 19611 7120 19612 7160
rect 19652 7120 19653 7160
rect 19611 7111 19653 7120
rect 19851 7160 19893 7169
rect 19851 7120 19852 7160
rect 19892 7120 19893 7160
rect 19851 7111 19893 7120
rect 20235 7160 20277 7169
rect 20235 7120 20236 7160
rect 20276 7120 20277 7160
rect 20235 7111 20277 7120
rect 20410 7160 20468 7161
rect 20410 7120 20419 7160
rect 20459 7120 20468 7160
rect 20410 7119 20468 7120
rect 20523 7160 20565 7169
rect 20523 7120 20524 7160
rect 20564 7120 20565 7160
rect 20523 7111 20565 7120
rect 20662 7160 20704 7169
rect 20662 7120 20663 7160
rect 20703 7120 20704 7160
rect 20662 7111 20704 7120
rect 20794 7160 20852 7161
rect 20794 7120 20803 7160
rect 20843 7120 20852 7160
rect 20794 7119 20852 7120
rect 20907 7160 20949 7169
rect 20907 7120 20908 7160
rect 20948 7120 20949 7160
rect 20907 7111 20949 7120
rect 21195 7160 21237 7169
rect 21195 7120 21196 7160
rect 21236 7120 21237 7160
rect 21195 7111 21237 7120
rect 21309 7160 21367 7161
rect 21309 7120 21318 7160
rect 21358 7120 21367 7160
rect 21309 7119 21367 7120
rect 21435 7160 21493 7161
rect 21435 7120 21444 7160
rect 21484 7120 21493 7160
rect 21435 7119 21493 7120
rect 22299 7160 22341 7169
rect 22299 7120 22300 7160
rect 22340 7120 22341 7160
rect 22299 7111 22341 7120
rect 22522 7160 22580 7161
rect 22522 7120 22531 7160
rect 22571 7120 22580 7160
rect 22522 7119 22580 7120
rect 22827 7160 22869 7169
rect 22827 7120 22828 7160
rect 22868 7120 22869 7160
rect 22827 7111 22869 7120
rect 23016 7160 23058 7169
rect 23133 7162 23142 7202
rect 23182 7162 23191 7202
rect 23133 7161 23191 7162
rect 23276 7193 23318 7202
rect 23016 7120 23017 7160
rect 23057 7120 23058 7160
rect 23276 7153 23277 7193
rect 23317 7153 23318 7193
rect 23276 7144 23318 7153
rect 24154 7160 24212 7161
rect 23016 7111 23058 7120
rect 24154 7120 24163 7160
rect 24203 7120 24212 7160
rect 24154 7119 24212 7120
rect 26955 7160 26997 7169
rect 26955 7120 26956 7160
rect 26996 7120 26997 7160
rect 26955 7111 26997 7120
rect 3802 7076 3860 7077
rect 3802 7036 3811 7076
rect 3851 7036 3860 7076
rect 3802 7035 3860 7036
rect 14560 7076 14602 7085
rect 14560 7036 14561 7076
rect 14601 7036 14602 7076
rect 14560 7027 14602 7036
rect 15229 7076 15271 7085
rect 15229 7036 15230 7076
rect 15270 7036 15271 7076
rect 15229 7027 15271 7036
rect 23770 7076 23828 7077
rect 23770 7036 23779 7076
rect 23819 7036 23828 7076
rect 23770 7035 23828 7036
rect 26266 7076 26324 7077
rect 26266 7036 26275 7076
rect 26315 7036 26324 7076
rect 26266 7035 26324 7036
rect 1594 6992 1652 6993
rect 1594 6952 1603 6992
rect 1643 6952 1652 6992
rect 1594 6951 1652 6952
rect 1786 6992 1844 6993
rect 1786 6952 1795 6992
rect 1835 6952 1844 6992
rect 1786 6951 1844 6952
rect 2091 6992 2133 7001
rect 2091 6952 2092 6992
rect 2132 6952 2133 6992
rect 2091 6943 2133 6952
rect 2571 6992 2613 7001
rect 2571 6952 2572 6992
rect 2612 6952 2613 6992
rect 2571 6943 2613 6952
rect 2698 6992 2756 6993
rect 2698 6952 2707 6992
rect 2747 6952 2756 6992
rect 2698 6951 2756 6952
rect 3994 6992 4052 6993
rect 3994 6952 4003 6992
rect 4043 6952 4052 6992
rect 3994 6951 4052 6952
rect 4299 6992 4341 7001
rect 4299 6952 4300 6992
rect 4340 6952 4341 6992
rect 4299 6943 4341 6952
rect 5739 6992 5781 7001
rect 5739 6952 5740 6992
rect 5780 6952 5781 6992
rect 5739 6943 5781 6952
rect 7275 6992 7317 7001
rect 7275 6952 7276 6992
rect 7316 6952 7317 6992
rect 7275 6943 7317 6952
rect 10330 6992 10388 6993
rect 10330 6952 10339 6992
rect 10379 6952 10388 6992
rect 10330 6951 10388 6952
rect 10635 6992 10677 7001
rect 10635 6952 10636 6992
rect 10676 6952 10677 6992
rect 10635 6943 10677 6952
rect 11403 6992 11445 7001
rect 11403 6952 11404 6992
rect 11444 6952 11445 6992
rect 11403 6943 11445 6952
rect 13611 6992 13653 7001
rect 13611 6952 13612 6992
rect 13652 6952 13653 6992
rect 13611 6943 13653 6952
rect 14763 6992 14805 7001
rect 14763 6952 14764 6992
rect 14804 6952 14805 6992
rect 14763 6943 14805 6952
rect 15322 6992 15380 6993
rect 15322 6952 15331 6992
rect 15371 6952 15380 6992
rect 15322 6951 15380 6952
rect 15435 6992 15477 7001
rect 15435 6952 15436 6992
rect 15476 6952 15477 6992
rect 15435 6943 15477 6952
rect 19354 6992 19412 6993
rect 19354 6952 19363 6992
rect 19403 6952 19412 6992
rect 19354 6951 19412 6952
rect 19930 6992 19988 6993
rect 19930 6952 19939 6992
rect 19979 6952 19988 6992
rect 19930 6951 19988 6952
rect 21675 6992 21717 7001
rect 21675 6952 21676 6992
rect 21716 6952 21717 6992
rect 21675 6943 21717 6952
rect 22731 6992 22773 7001
rect 22731 6952 22732 6992
rect 22772 6952 22773 6992
rect 22731 6943 22773 6952
rect 23307 6992 23349 7001
rect 23307 6952 23308 6992
rect 23348 6952 23349 6992
rect 23307 6943 23349 6952
rect 26091 6992 26133 7001
rect 26091 6952 26092 6992
rect 26132 6952 26133 6992
rect 26091 6943 26133 6952
rect 576 6824 31392 6848
rect 576 6784 4352 6824
rect 4720 6784 12126 6824
rect 12494 6784 19900 6824
rect 20268 6784 27674 6824
rect 28042 6784 31392 6824
rect 576 6760 31392 6784
rect 1227 6656 1269 6665
rect 1227 6616 1228 6656
rect 1268 6616 1269 6656
rect 1227 6607 1269 6616
rect 2283 6656 2325 6665
rect 2283 6616 2284 6656
rect 2324 6616 2325 6656
rect 2283 6607 2325 6616
rect 3435 6656 3477 6665
rect 3435 6616 3436 6656
rect 3476 6616 3477 6656
rect 3435 6607 3477 6616
rect 6027 6656 6069 6665
rect 6027 6616 6028 6656
rect 6068 6616 6069 6656
rect 6027 6607 6069 6616
rect 6874 6656 6932 6657
rect 6874 6616 6883 6656
rect 6923 6616 6932 6656
rect 6874 6615 6932 6616
rect 7851 6656 7893 6665
rect 7851 6616 7852 6656
rect 7892 6616 7893 6656
rect 7851 6607 7893 6616
rect 8314 6656 8372 6657
rect 8314 6616 8323 6656
rect 8363 6616 8372 6656
rect 8314 6615 8372 6616
rect 8667 6656 8709 6665
rect 8667 6616 8668 6656
rect 8708 6616 8709 6656
rect 8667 6607 8709 6616
rect 9147 6656 9189 6665
rect 9147 6616 9148 6656
rect 9188 6616 9189 6656
rect 9147 6607 9189 6616
rect 9466 6656 9524 6657
rect 9466 6616 9475 6656
rect 9515 6616 9524 6656
rect 9466 6615 9524 6616
rect 10234 6656 10292 6657
rect 10234 6616 10243 6656
rect 10283 6616 10292 6656
rect 10234 6615 10292 6616
rect 10539 6656 10581 6665
rect 10539 6616 10540 6656
rect 10580 6616 10581 6656
rect 10539 6607 10581 6616
rect 11979 6656 12021 6665
rect 11979 6616 11980 6656
rect 12020 6616 12021 6656
rect 11979 6607 12021 6616
rect 12442 6656 12500 6657
rect 12442 6616 12451 6656
rect 12491 6616 12500 6656
rect 12442 6615 12500 6616
rect 13018 6656 13076 6657
rect 13018 6616 13027 6656
rect 13067 6616 13076 6656
rect 13018 6615 13076 6616
rect 13131 6656 13173 6665
rect 13131 6616 13132 6656
rect 13172 6616 13173 6656
rect 13131 6607 13173 6616
rect 13498 6656 13556 6657
rect 13498 6616 13507 6656
rect 13547 6616 13556 6656
rect 13498 6615 13556 6616
rect 14667 6656 14709 6665
rect 14667 6616 14668 6656
rect 14708 6616 14709 6656
rect 14667 6607 14709 6616
rect 15147 6656 15189 6665
rect 15147 6616 15148 6656
rect 15188 6616 15189 6656
rect 15147 6607 15189 6616
rect 16107 6656 16149 6665
rect 16107 6616 16108 6656
rect 16148 6616 16149 6656
rect 16107 6607 16149 6616
rect 16666 6656 16724 6657
rect 16666 6616 16675 6656
rect 16715 6616 16724 6656
rect 16666 6615 16724 6616
rect 17434 6656 17492 6657
rect 17434 6616 17443 6656
rect 17483 6616 17492 6656
rect 17434 6615 17492 6616
rect 18202 6656 18260 6657
rect 18202 6616 18211 6656
rect 18251 6616 18260 6656
rect 18202 6615 18260 6616
rect 18507 6656 18549 6665
rect 18507 6616 18508 6656
rect 18548 6616 18549 6656
rect 18507 6607 18549 6616
rect 18778 6656 18836 6657
rect 18778 6616 18787 6656
rect 18827 6616 18836 6656
rect 18778 6615 18836 6616
rect 18891 6656 18933 6665
rect 18891 6616 18892 6656
rect 18932 6616 18933 6656
rect 18891 6607 18933 6616
rect 19371 6656 19413 6665
rect 19371 6616 19372 6656
rect 19412 6616 19413 6656
rect 19371 6607 19413 6616
rect 22635 6656 22677 6665
rect 22635 6616 22636 6656
rect 22676 6616 22677 6656
rect 22635 6607 22677 6616
rect 23194 6656 23252 6657
rect 23194 6616 23203 6656
rect 23243 6616 23252 6656
rect 23194 6615 23252 6616
rect 24267 6656 24309 6665
rect 24267 6616 24268 6656
rect 24308 6616 24309 6656
rect 24267 6607 24309 6616
rect 1611 6572 1653 6581
rect 1611 6532 1612 6572
rect 1652 6532 1653 6572
rect 1611 6523 1653 6532
rect 8427 6572 8469 6581
rect 8427 6532 8428 6572
rect 8468 6532 8469 6572
rect 8427 6523 8469 6532
rect 18685 6572 18727 6581
rect 18685 6532 18686 6572
rect 18726 6532 18727 6572
rect 18685 6523 18727 6532
rect 20043 6572 20085 6581
rect 20043 6532 20044 6572
rect 20084 6532 20085 6572
rect 20043 6523 20085 6532
rect 20314 6572 20372 6573
rect 20314 6532 20323 6572
rect 20363 6532 20372 6572
rect 20314 6531 20372 6532
rect 16961 6498 17019 6499
rect 1131 6488 1173 6497
rect 1131 6448 1132 6488
rect 1172 6448 1173 6488
rect 1131 6439 1173 6448
rect 1306 6488 1364 6489
rect 1306 6448 1315 6488
rect 1355 6448 1364 6488
rect 1306 6447 1364 6448
rect 1522 6488 1564 6497
rect 1522 6448 1523 6488
rect 1563 6448 1564 6488
rect 1522 6439 1564 6448
rect 1690 6488 1748 6489
rect 1690 6448 1699 6488
rect 1739 6448 1748 6488
rect 1690 6447 1748 6448
rect 2187 6488 2229 6497
rect 2187 6448 2188 6488
rect 2228 6448 2229 6488
rect 2187 6439 2229 6448
rect 2362 6488 2420 6489
rect 2362 6448 2371 6488
rect 2411 6448 2420 6488
rect 2362 6447 2420 6448
rect 2955 6488 2997 6497
rect 2955 6448 2956 6488
rect 2996 6448 2997 6488
rect 2955 6439 2997 6448
rect 3339 6488 3381 6497
rect 3339 6448 3340 6488
rect 3380 6448 3381 6488
rect 3339 6439 3381 6448
rect 4090 6488 4148 6489
rect 4090 6448 4099 6488
rect 4139 6448 4148 6488
rect 4090 6447 4148 6448
rect 6538 6488 6596 6489
rect 6538 6448 6547 6488
rect 6587 6448 6596 6488
rect 6538 6447 6596 6448
rect 6733 6488 6791 6489
rect 6733 6448 6742 6488
rect 6782 6448 6791 6488
rect 6733 6447 6791 6448
rect 6987 6488 7029 6497
rect 6987 6448 6988 6488
rect 7028 6448 7029 6488
rect 6987 6439 7029 6448
rect 7371 6488 7413 6497
rect 7371 6448 7372 6488
rect 7412 6448 7413 6488
rect 7371 6439 7413 6448
rect 7659 6488 7701 6497
rect 7659 6448 7660 6488
rect 7700 6448 7701 6488
rect 7659 6439 7701 6448
rect 8218 6488 8276 6489
rect 8218 6448 8227 6488
rect 8267 6448 8276 6488
rect 8218 6447 8276 6448
rect 8534 6488 8576 6497
rect 8534 6448 8535 6488
rect 8575 6448 8576 6488
rect 8534 6439 8576 6448
rect 8811 6488 8853 6497
rect 9627 6488 9669 6497
rect 8811 6448 8812 6488
rect 8852 6448 8853 6488
rect 8811 6439 8853 6448
rect 8994 6479 9040 6488
rect 8994 6439 8995 6479
rect 9035 6439 9040 6479
rect 9627 6448 9628 6488
rect 9668 6448 9669 6488
rect 9627 6439 9669 6448
rect 9771 6488 9813 6497
rect 9771 6448 9772 6488
rect 9812 6448 9813 6488
rect 9771 6439 9813 6448
rect 10347 6488 10389 6497
rect 10347 6448 10348 6488
rect 10388 6448 10389 6488
rect 10347 6439 10389 6448
rect 10875 6488 10917 6497
rect 10875 6448 10876 6488
rect 10916 6448 10917 6488
rect 10875 6439 10917 6448
rect 11019 6488 11061 6497
rect 11019 6448 11020 6488
rect 11060 6448 11061 6488
rect 11019 6439 11061 6448
rect 11499 6488 11541 6497
rect 11499 6448 11500 6488
rect 11540 6448 11541 6488
rect 11499 6439 11541 6448
rect 11787 6488 11829 6497
rect 11787 6448 11788 6488
rect 11828 6448 11829 6488
rect 11787 6439 11829 6448
rect 12555 6488 12597 6497
rect 12555 6448 12556 6488
rect 12596 6448 12597 6488
rect 12555 6439 12597 6448
rect 12928 6488 12970 6497
rect 13707 6488 13749 6497
rect 12928 6448 12929 6488
rect 12969 6448 12970 6488
rect 12928 6439 12970 6448
rect 13227 6479 13269 6488
rect 13227 6439 13228 6479
rect 13268 6439 13269 6479
rect 13707 6448 13708 6488
rect 13748 6448 13749 6488
rect 13707 6439 13749 6448
rect 13995 6488 14037 6497
rect 13995 6448 13996 6488
rect 14036 6448 14037 6488
rect 13995 6439 14037 6448
rect 14187 6488 14229 6497
rect 14187 6448 14188 6488
rect 14228 6448 14229 6488
rect 14187 6439 14229 6448
rect 14475 6488 14517 6497
rect 14475 6448 14476 6488
rect 14516 6448 14517 6488
rect 14475 6439 14517 6448
rect 14938 6488 14996 6489
rect 14938 6448 14947 6488
rect 14987 6448 14996 6488
rect 14938 6447 14996 6448
rect 15243 6488 15285 6497
rect 15243 6448 15244 6488
rect 15284 6448 15285 6488
rect 15243 6439 15285 6448
rect 15627 6488 15669 6497
rect 15627 6448 15628 6488
rect 15668 6448 15669 6488
rect 15627 6439 15669 6448
rect 16011 6488 16053 6497
rect 16011 6448 16012 6488
rect 16052 6448 16053 6488
rect 16011 6439 16053 6448
rect 16827 6488 16869 6497
rect 16827 6448 16828 6488
rect 16868 6448 16869 6488
rect 16961 6458 16970 6498
rect 17010 6458 17019 6498
rect 16961 6457 17019 6458
rect 17739 6488 17781 6497
rect 16827 6439 16869 6448
rect 17739 6448 17740 6488
rect 17780 6448 17781 6488
rect 17739 6439 17781 6448
rect 18315 6488 18357 6497
rect 19275 6488 19317 6497
rect 18315 6448 18316 6488
rect 18356 6448 18357 6488
rect 18315 6439 18357 6448
rect 18987 6479 19029 6488
rect 18987 6439 18988 6479
rect 19028 6439 19029 6479
rect 19275 6448 19276 6488
rect 19316 6448 19317 6488
rect 19275 6439 19317 6448
rect 19450 6488 19508 6489
rect 19450 6448 19459 6488
rect 19499 6448 19508 6488
rect 19450 6447 19508 6448
rect 19834 6488 19892 6489
rect 19834 6448 19843 6488
rect 19883 6448 19892 6488
rect 19834 6447 19892 6448
rect 20139 6488 20181 6497
rect 20139 6448 20140 6488
rect 20180 6448 20181 6488
rect 20139 6439 20181 6448
rect 20698 6488 20756 6489
rect 20698 6448 20707 6488
rect 20747 6448 20756 6488
rect 20698 6447 20756 6448
rect 23307 6488 23349 6497
rect 23307 6448 23308 6488
rect 23348 6448 23349 6488
rect 23307 6439 23349 6448
rect 23643 6488 23685 6497
rect 23643 6448 23644 6488
rect 23684 6448 23685 6488
rect 23643 6439 23685 6448
rect 23883 6488 23925 6497
rect 23883 6448 23884 6488
rect 23924 6448 23925 6488
rect 23883 6439 23925 6448
rect 24075 6488 24117 6497
rect 24075 6448 24076 6488
rect 24116 6448 24117 6488
rect 24075 6439 24117 6448
rect 24939 6488 24981 6497
rect 24939 6448 24940 6488
rect 24980 6448 24981 6488
rect 24939 6439 24981 6448
rect 25803 6488 25845 6497
rect 25803 6448 25804 6488
rect 25844 6448 25845 6488
rect 25803 6439 25845 6448
rect 8994 6430 9040 6439
rect 13227 6430 13269 6439
rect 18987 6430 19029 6439
rect 3723 6404 3765 6413
rect 3723 6364 3724 6404
rect 3764 6364 3765 6404
rect 3723 6355 3765 6364
rect 17649 6404 17691 6413
rect 17649 6364 17650 6404
rect 17690 6364 17691 6404
rect 17649 6355 17691 6364
rect 22251 6404 22293 6413
rect 22251 6364 22252 6404
rect 22292 6364 22293 6404
rect 22251 6355 22293 6364
rect 25114 6404 25172 6405
rect 25114 6364 25123 6404
rect 25163 6364 25172 6404
rect 25114 6363 25172 6364
rect 2571 6320 2613 6329
rect 2571 6280 2572 6320
rect 2612 6280 2613 6320
rect 2571 6271 2613 6280
rect 7179 6320 7221 6329
rect 7179 6280 7180 6320
rect 7220 6280 7221 6320
rect 7179 6271 7221 6280
rect 12747 6320 12789 6329
rect 12747 6280 12748 6320
rect 12788 6280 12789 6320
rect 12747 6271 12789 6280
rect 25995 6320 26037 6329
rect 25995 6280 25996 6320
rect 26036 6280 26037 6320
rect 25995 6271 26037 6280
rect 5643 6236 5685 6245
rect 5643 6196 5644 6236
rect 5684 6196 5685 6236
rect 5643 6187 5685 6196
rect 6027 6236 6069 6245
rect 6027 6196 6028 6236
rect 6068 6196 6069 6236
rect 6027 6187 6069 6196
rect 10827 6236 10869 6245
rect 10827 6196 10828 6236
rect 10868 6196 10869 6236
rect 10827 6187 10869 6196
rect 22635 6236 22677 6245
rect 22635 6196 22636 6236
rect 22676 6196 22677 6236
rect 22635 6187 22677 6196
rect 23883 6236 23925 6245
rect 23883 6196 23884 6236
rect 23924 6196 23925 6236
rect 23883 6187 23925 6196
rect 576 6068 31392 6092
rect 576 6028 3112 6068
rect 3480 6028 10886 6068
rect 11254 6028 18660 6068
rect 19028 6028 26434 6068
rect 26802 6028 31392 6068
rect 576 6004 31392 6028
rect 3531 5900 3573 5909
rect 3531 5860 3532 5900
rect 3572 5860 3573 5900
rect 3531 5851 3573 5860
rect 8427 5900 8469 5909
rect 8427 5860 8428 5900
rect 8468 5860 8469 5900
rect 8427 5851 8469 5860
rect 8811 5900 8853 5909
rect 8811 5860 8812 5900
rect 8852 5860 8853 5900
rect 8811 5851 8853 5860
rect 12171 5900 12213 5909
rect 12171 5860 12172 5900
rect 12212 5860 12213 5900
rect 12171 5851 12213 5860
rect 15723 5900 15765 5909
rect 15723 5860 15724 5900
rect 15764 5860 15765 5900
rect 15723 5851 15765 5860
rect 16971 5900 17013 5909
rect 16971 5860 16972 5900
rect 17012 5860 17013 5900
rect 16971 5851 17013 5860
rect 20331 5900 20373 5909
rect 20331 5860 20332 5900
rect 20372 5860 20373 5900
rect 20331 5851 20373 5860
rect 21483 5900 21525 5909
rect 21483 5860 21484 5900
rect 21524 5860 21525 5900
rect 21483 5851 21525 5860
rect 24267 5900 24309 5909
rect 24267 5860 24268 5900
rect 24308 5860 24309 5900
rect 24267 5851 24309 5860
rect 25131 5900 25173 5909
rect 25131 5860 25132 5900
rect 25172 5860 25173 5900
rect 25131 5851 25173 5860
rect 3915 5816 3957 5825
rect 4683 5816 4725 5825
rect 3915 5776 3916 5816
rect 3956 5776 3957 5816
rect 3915 5767 3957 5776
rect 4155 5807 4197 5816
rect 4155 5767 4156 5807
rect 4196 5767 4197 5807
rect 4683 5776 4684 5816
rect 4724 5776 4725 5816
rect 4683 5767 4725 5776
rect 12555 5816 12597 5825
rect 12555 5776 12556 5816
rect 12596 5776 12597 5816
rect 12555 5767 12597 5776
rect 17355 5816 17397 5825
rect 17355 5776 17356 5816
rect 17396 5776 17397 5816
rect 17355 5767 17397 5776
rect 21867 5816 21909 5825
rect 21867 5776 21868 5816
rect 21908 5776 21909 5816
rect 21867 5767 21909 5776
rect 24651 5816 24693 5825
rect 24651 5776 24652 5816
rect 24692 5776 24693 5816
rect 24651 5767 24693 5776
rect 4155 5758 4197 5767
rect 5355 5732 5397 5741
rect 5355 5692 5356 5732
rect 5396 5692 5397 5732
rect 5355 5683 5397 5692
rect 16426 5732 16484 5733
rect 16426 5692 16435 5732
rect 16475 5692 16484 5732
rect 16426 5691 16484 5692
rect 3531 5648 3573 5657
rect 3531 5608 3532 5648
rect 3572 5608 3573 5648
rect 3531 5599 3573 5608
rect 3723 5648 3765 5657
rect 3723 5608 3724 5648
rect 3764 5608 3765 5648
rect 3723 5599 3765 5608
rect 4090 5648 4148 5649
rect 4090 5608 4099 5648
rect 4139 5608 4148 5648
rect 4090 5607 4148 5608
rect 5026 5648 5084 5649
rect 5026 5608 5035 5648
rect 5075 5608 5084 5648
rect 5026 5607 5084 5608
rect 5146 5648 5204 5649
rect 5146 5608 5155 5648
rect 5195 5608 5204 5648
rect 5146 5607 5204 5608
rect 5259 5648 5301 5657
rect 5259 5608 5260 5648
rect 5300 5608 5301 5648
rect 5259 5599 5301 5608
rect 5827 5648 5885 5649
rect 5827 5608 5836 5648
rect 5876 5608 5885 5648
rect 5827 5607 5885 5608
rect 6007 5648 6065 5649
rect 6007 5608 6016 5648
rect 6056 5608 6065 5648
rect 6007 5607 6065 5608
rect 6874 5648 6932 5649
rect 6874 5608 6883 5648
rect 6923 5608 6932 5648
rect 6874 5607 6932 5608
rect 9195 5648 9237 5657
rect 9195 5608 9196 5648
rect 9236 5608 9237 5648
rect 9195 5599 9237 5608
rect 10618 5648 10676 5649
rect 10618 5608 10627 5648
rect 10667 5608 10676 5648
rect 10618 5607 10676 5608
rect 13035 5648 13077 5657
rect 13035 5608 13036 5648
rect 13076 5608 13077 5648
rect 13035 5599 13077 5608
rect 13179 5648 13221 5657
rect 13179 5608 13180 5648
rect 13220 5608 13221 5648
rect 13179 5599 13221 5608
rect 14170 5648 14228 5649
rect 14170 5608 14179 5648
rect 14219 5608 14228 5648
rect 14170 5607 14228 5608
rect 16621 5648 16679 5649
rect 16621 5608 16630 5648
rect 16670 5608 16679 5648
rect 16621 5607 16679 5608
rect 18874 5648 18932 5649
rect 18874 5608 18883 5648
rect 18923 5608 18932 5648
rect 18874 5607 18932 5608
rect 19467 5648 19509 5657
rect 19467 5608 19468 5648
rect 19508 5608 19509 5648
rect 19467 5599 19509 5608
rect 21003 5648 21045 5657
rect 21003 5608 21004 5648
rect 21044 5608 21045 5648
rect 21003 5599 21045 5608
rect 21178 5648 21236 5649
rect 21178 5608 21187 5648
rect 21227 5608 21236 5648
rect 21178 5607 21236 5608
rect 21291 5648 21333 5657
rect 21291 5608 21292 5648
rect 21332 5608 21333 5648
rect 21291 5599 21333 5608
rect 22714 5648 22772 5649
rect 22714 5608 22723 5648
rect 22763 5608 22772 5648
rect 22714 5607 22772 5608
rect 24826 5648 24884 5649
rect 24826 5608 24835 5648
rect 24875 5608 24884 5648
rect 24826 5607 24884 5608
rect 25131 5648 25173 5657
rect 25131 5608 25132 5648
rect 25172 5608 25173 5648
rect 25131 5599 25173 5608
rect 5533 5564 5575 5573
rect 5533 5524 5534 5564
rect 5574 5524 5575 5564
rect 5533 5515 5575 5524
rect 5626 5564 5684 5565
rect 5626 5524 5635 5564
rect 5675 5524 5684 5564
rect 5626 5523 5684 5524
rect 6490 5564 6548 5565
rect 6490 5524 6499 5564
rect 6539 5524 6548 5564
rect 6490 5523 6548 5524
rect 10234 5564 10292 5565
rect 10234 5524 10243 5564
rect 10283 5524 10292 5564
rect 10234 5523 10292 5524
rect 12826 5564 12884 5565
rect 12826 5524 12835 5564
rect 12875 5524 12884 5564
rect 12826 5523 12884 5524
rect 13786 5564 13844 5565
rect 13786 5524 13795 5564
rect 13835 5524 13844 5564
rect 13786 5523 13844 5524
rect 19258 5564 19316 5565
rect 19258 5524 19267 5564
rect 19307 5524 19316 5564
rect 19258 5523 19316 5524
rect 20139 5564 20181 5573
rect 20139 5524 20140 5564
rect 20180 5524 20181 5564
rect 20139 5515 20181 5524
rect 21494 5564 21536 5573
rect 21494 5524 21495 5564
rect 21535 5524 21536 5564
rect 21494 5515 21536 5524
rect 22330 5564 22388 5565
rect 22330 5524 22339 5564
rect 22379 5524 22388 5564
rect 22330 5523 22388 5524
rect 5739 5480 5781 5489
rect 5739 5440 5740 5480
rect 5780 5440 5781 5480
rect 5739 5431 5781 5440
rect 6171 5480 6213 5489
rect 6171 5440 6172 5480
rect 6212 5440 6213 5480
rect 6171 5431 6213 5440
rect 9867 5480 9909 5489
rect 9867 5440 9868 5480
rect 9908 5440 9909 5480
rect 9867 5431 9909 5440
rect 13131 5480 13173 5489
rect 13131 5440 13132 5480
rect 13172 5440 13173 5480
rect 13131 5431 13173 5440
rect 16107 5480 16149 5489
rect 16107 5440 16108 5480
rect 16148 5440 16149 5480
rect 16107 5431 16149 5440
rect 576 5312 31392 5336
rect 576 5272 4352 5312
rect 4720 5272 12126 5312
rect 12494 5272 19900 5312
rect 20268 5272 27674 5312
rect 28042 5272 31392 5312
rect 576 5248 31392 5272
rect 6363 5144 6405 5153
rect 6363 5104 6364 5144
rect 6404 5104 6405 5144
rect 6363 5095 6405 5104
rect 9130 5144 9188 5145
rect 9130 5104 9139 5144
rect 9179 5104 9188 5144
rect 9130 5103 9188 5104
rect 10059 5144 10101 5153
rect 10059 5104 10060 5144
rect 10100 5104 10101 5144
rect 10059 5095 10101 5104
rect 10827 5144 10869 5153
rect 10827 5104 10828 5144
rect 10868 5104 10869 5144
rect 10827 5095 10869 5104
rect 11770 5144 11828 5145
rect 11770 5104 11779 5144
rect 11819 5104 11828 5144
rect 11770 5103 11828 5104
rect 13786 5144 13844 5145
rect 13786 5104 13795 5144
rect 13835 5104 13844 5144
rect 13786 5103 13844 5104
rect 16971 5144 17013 5153
rect 16971 5104 16972 5144
rect 17012 5104 17013 5144
rect 16971 5095 17013 5104
rect 20715 5144 20757 5153
rect 20715 5104 20716 5144
rect 20756 5104 20757 5144
rect 20715 5095 20757 5104
rect 21195 5144 21237 5153
rect 21195 5104 21196 5144
rect 21236 5104 21237 5144
rect 21195 5095 21237 5104
rect 23595 5144 23637 5153
rect 23595 5104 23596 5144
rect 23636 5104 23637 5144
rect 23595 5095 23637 5104
rect 23962 5144 24020 5145
rect 23962 5104 23971 5144
rect 24011 5104 24020 5144
rect 23962 5103 24020 5104
rect 12075 5060 12117 5069
rect 12075 5020 12076 5060
rect 12116 5020 12117 5060
rect 12075 5011 12117 5020
rect 13899 5060 13941 5069
rect 13899 5020 13900 5060
rect 13940 5020 13941 5060
rect 13899 5011 13941 5020
rect 16011 5060 16053 5069
rect 16011 5020 16012 5060
rect 16052 5020 16053 5060
rect 16011 5011 16053 5020
rect 23869 5060 23911 5069
rect 23869 5020 23870 5060
rect 23910 5020 23911 5060
rect 23869 5011 23911 5020
rect 24075 5060 24117 5069
rect 24075 5020 24076 5060
rect 24116 5020 24117 5060
rect 24075 5011 24117 5020
rect 6219 4976 6261 4985
rect 6219 4936 6220 4976
rect 6260 4936 6261 4976
rect 6219 4927 6261 4936
rect 9325 4976 9383 4977
rect 9325 4936 9334 4976
rect 9374 4936 9383 4976
rect 9325 4935 9383 4936
rect 9658 4976 9716 4977
rect 9658 4936 9667 4976
rect 9707 4936 9716 4976
rect 9658 4935 9716 4936
rect 9771 4976 9813 4985
rect 9771 4936 9772 4976
rect 9812 4936 9813 4976
rect 9771 4927 9813 4936
rect 10539 4976 10581 4985
rect 10539 4936 10540 4976
rect 10580 4936 10581 4976
rect 10539 4927 10581 4936
rect 10731 4976 10773 4985
rect 10731 4936 10732 4976
rect 10772 4936 10773 4976
rect 10731 4927 10773 4936
rect 10923 4976 10965 4985
rect 10923 4936 10924 4976
rect 10964 4936 10965 4976
rect 10923 4927 10965 4936
rect 11446 4976 11488 4985
rect 11446 4936 11447 4976
rect 11487 4936 11488 4976
rect 11446 4927 11488 4936
rect 11691 4976 11733 4985
rect 11691 4936 11692 4976
rect 11732 4936 11733 4976
rect 11691 4927 11733 4936
rect 11979 4976 12021 4985
rect 11979 4936 11980 4976
rect 12020 4936 12021 4976
rect 11979 4927 12021 4936
rect 12171 4976 12213 4985
rect 12171 4936 12172 4976
rect 12212 4936 12213 4976
rect 12171 4927 12213 4936
rect 12747 4976 12789 4985
rect 12747 4936 12748 4976
rect 12788 4936 12789 4976
rect 12747 4927 12789 4936
rect 12922 4976 12980 4977
rect 12922 4936 12931 4976
rect 12971 4936 12980 4976
rect 12922 4935 12980 4936
rect 13035 4976 13077 4985
rect 13035 4936 13036 4976
rect 13076 4936 13077 4976
rect 13035 4927 13077 4936
rect 13227 4976 13269 4985
rect 13227 4936 13228 4976
rect 13268 4936 13269 4976
rect 13227 4927 13269 4936
rect 13341 4976 13399 4977
rect 13341 4936 13350 4976
rect 13390 4936 13399 4976
rect 13341 4935 13399 4936
rect 13468 4976 13526 4977
rect 13468 4936 13477 4976
rect 13517 4936 13526 4976
rect 13468 4935 13526 4936
rect 13690 4976 13748 4977
rect 13690 4936 13699 4976
rect 13739 4936 13748 4976
rect 13690 4935 13748 4936
rect 14006 4976 14048 4985
rect 14006 4936 14007 4976
rect 14047 4936 14048 4976
rect 14006 4927 14048 4936
rect 14235 4976 14277 4985
rect 14235 4936 14236 4976
rect 14276 4936 14277 4976
rect 14235 4927 14277 4936
rect 14859 4976 14901 4985
rect 14859 4936 14860 4976
rect 14900 4936 14901 4976
rect 14859 4927 14901 4936
rect 15610 4976 15668 4977
rect 15610 4936 15619 4976
rect 15659 4936 15668 4976
rect 15610 4935 15668 4936
rect 16299 4976 16341 4985
rect 16299 4936 16300 4976
rect 16340 4936 16341 4976
rect 16299 4927 16341 4936
rect 19083 4976 19125 4985
rect 19083 4936 19084 4976
rect 19124 4936 19125 4976
rect 19083 4927 19125 4936
rect 19258 4976 19316 4977
rect 19258 4936 19267 4976
rect 19307 4936 19316 4976
rect 19258 4935 19316 4936
rect 19642 4976 19700 4977
rect 19642 4936 19651 4976
rect 19691 4936 19700 4976
rect 19642 4935 19700 4936
rect 19755 4976 19797 4985
rect 19755 4936 19756 4976
rect 19796 4936 19797 4976
rect 19755 4927 19797 4936
rect 20235 4976 20277 4985
rect 20235 4936 20236 4976
rect 20276 4936 20277 4976
rect 20235 4927 20277 4936
rect 20404 4976 20446 4985
rect 20404 4936 20405 4976
rect 20445 4936 20446 4976
rect 20404 4927 20446 4936
rect 20523 4976 20565 4985
rect 20523 4936 20524 4976
rect 20564 4936 20565 4976
rect 20523 4927 20565 4936
rect 21003 4976 21045 4985
rect 21003 4936 21004 4976
rect 21044 4936 21045 4976
rect 21003 4927 21045 4936
rect 21195 4976 21237 4985
rect 21195 4936 21196 4976
rect 21236 4936 21237 4976
rect 21195 4927 21237 4936
rect 21387 4976 21429 4985
rect 21387 4936 21388 4976
rect 21428 4936 21429 4976
rect 21387 4927 21429 4936
rect 22635 4976 22677 4985
rect 22635 4936 22636 4976
rect 22676 4936 22677 4976
rect 22635 4927 22677 4936
rect 22810 4976 22868 4977
rect 22810 4936 22819 4976
rect 22859 4936 22868 4976
rect 22810 4935 22868 4936
rect 23019 4976 23061 4985
rect 23019 4936 23020 4976
rect 23060 4936 23061 4976
rect 23019 4927 23061 4936
rect 23194 4976 23252 4977
rect 23194 4936 23203 4976
rect 23243 4936 23252 4976
rect 23194 4935 23252 4936
rect 23305 4976 23363 4977
rect 23305 4936 23314 4976
rect 23354 4936 23363 4976
rect 23305 4935 23363 4936
rect 23506 4976 23564 4977
rect 23506 4936 23515 4976
rect 23555 4936 23564 4976
rect 23506 4935 23564 4936
rect 23691 4976 23733 4985
rect 23691 4936 23692 4976
rect 23732 4936 23733 4976
rect 23691 4927 23733 4936
rect 24171 4967 24213 4976
rect 24171 4927 24172 4967
rect 24212 4927 24213 4967
rect 24171 4918 24213 4927
rect 10443 4892 10485 4901
rect 10443 4852 10444 4892
rect 10484 4852 10485 4892
rect 10443 4843 10485 4852
rect 11578 4892 11636 4893
rect 11578 4852 11587 4892
rect 11627 4852 11636 4892
rect 11578 4851 11636 4852
rect 20859 4892 20901 4901
rect 20859 4852 20860 4892
rect 20900 4852 20901 4892
rect 20859 4843 20901 4852
rect 7563 4808 7605 4817
rect 7563 4768 7564 4808
rect 7604 4768 7605 4808
rect 7563 4759 7605 4768
rect 11122 4808 11164 4817
rect 11122 4768 11123 4808
rect 11163 4768 11164 4808
rect 11122 4759 11164 4768
rect 13035 4808 13077 4817
rect 13035 4768 13036 4808
rect 13076 4768 13077 4808
rect 13035 4759 13077 4768
rect 13515 4808 13557 4817
rect 13515 4768 13516 4808
rect 13556 4768 13557 4808
rect 13515 4759 13557 4768
rect 15051 4808 15093 4817
rect 15051 4768 15052 4808
rect 15092 4768 15093 4808
rect 15051 4759 15093 4768
rect 18219 4808 18261 4817
rect 18219 4768 18220 4808
rect 18260 4768 18261 4808
rect 18219 4759 18261 4768
rect 19258 4808 19316 4809
rect 19258 4768 19267 4808
rect 19307 4768 19316 4808
rect 19258 4767 19316 4768
rect 21579 4808 21621 4817
rect 21579 4768 21580 4808
rect 21620 4768 21621 4808
rect 21579 4759 21621 4768
rect 22810 4808 22868 4809
rect 22810 4768 22819 4808
rect 22859 4768 22868 4808
rect 22810 4767 22868 4768
rect 15819 4724 15861 4733
rect 15819 4684 15820 4724
rect 15860 4684 15861 4724
rect 15819 4675 15861 4684
rect 19851 4724 19893 4733
rect 19851 4684 19852 4724
rect 19892 4684 19893 4724
rect 19851 4675 19893 4684
rect 23307 4724 23349 4733
rect 23307 4684 23308 4724
rect 23348 4684 23349 4724
rect 23307 4675 23349 4684
rect 576 4556 31392 4580
rect 576 4516 3112 4556
rect 3480 4516 10886 4556
rect 11254 4516 18660 4556
rect 19028 4516 26434 4556
rect 26802 4516 31392 4556
rect 576 4492 31392 4516
rect 19834 4388 19892 4389
rect 19834 4348 19843 4388
rect 19883 4348 19892 4388
rect 19834 4347 19892 4348
rect 20331 4388 20373 4397
rect 20331 4348 20332 4388
rect 20372 4348 20373 4388
rect 20331 4339 20373 4348
rect 20667 4388 20709 4397
rect 20667 4348 20668 4388
rect 20708 4348 20709 4388
rect 20667 4339 20709 4348
rect 10059 4304 10101 4313
rect 10059 4264 10060 4304
rect 10100 4264 10101 4304
rect 10059 4255 10101 4264
rect 9963 4136 10005 4145
rect 9963 4096 9964 4136
rect 10004 4096 10005 4136
rect 9963 4087 10005 4096
rect 10155 4136 10197 4145
rect 10155 4096 10156 4136
rect 10196 4096 10197 4136
rect 10155 4087 10197 4096
rect 19659 4136 19701 4145
rect 19659 4096 19660 4136
rect 19700 4096 19701 4136
rect 19659 4087 19701 4096
rect 19834 4136 19892 4137
rect 19834 4096 19843 4136
rect 19883 4096 19892 4136
rect 19834 4095 19892 4096
rect 20331 4136 20373 4145
rect 20331 4096 20332 4136
rect 20372 4096 20373 4136
rect 20331 4087 20373 4096
rect 20523 4136 20565 4145
rect 20523 4096 20524 4136
rect 20564 4096 20565 4136
rect 20523 4087 20565 4096
rect 20811 4136 20853 4145
rect 20811 4096 20812 4136
rect 20852 4096 20853 4136
rect 20811 4087 20853 4096
rect 576 3800 31392 3824
rect 576 3760 4352 3800
rect 4720 3760 12126 3800
rect 12494 3760 19900 3800
rect 20268 3760 27674 3800
rect 28042 3760 31392 3800
rect 576 3736 31392 3760
rect 576 3044 31392 3068
rect 576 3004 3112 3044
rect 3480 3004 10886 3044
rect 11254 3004 18660 3044
rect 19028 3004 26434 3044
rect 26802 3004 31392 3044
rect 576 2980 31392 3004
rect 576 2288 31392 2312
rect 576 2248 4352 2288
rect 4720 2248 12126 2288
rect 12494 2248 19900 2288
rect 20268 2248 27674 2288
rect 28042 2248 31392 2288
rect 576 2224 31392 2248
rect 576 1532 31392 1556
rect 576 1492 3112 1532
rect 3480 1492 10886 1532
rect 11254 1492 18660 1532
rect 19028 1492 26434 1532
rect 26802 1492 31392 1532
rect 576 1468 31392 1492
rect 576 776 31392 800
rect 576 736 4352 776
rect 4720 736 12126 776
rect 12494 736 19900 776
rect 20268 736 27674 776
rect 28042 736 31392 776
rect 576 712 31392 736
<< via1 >>
rect 4352 27952 4720 27992
rect 12126 27952 12494 27992
rect 19900 27952 20268 27992
rect 27674 27952 28042 27992
rect 2092 27784 2132 27824
rect 2476 27784 2516 27824
rect 2947 27784 2987 27824
rect 4099 27784 4139 27824
rect 5164 27784 5204 27824
rect 13036 27784 13076 27824
rect 13516 27784 13556 27824
rect 19468 27784 19508 27824
rect 19747 27784 19787 27824
rect 22444 27784 22484 27824
rect 27868 27784 27908 27824
rect 6067 27700 6107 27740
rect 6604 27700 6644 27740
rect 6883 27700 6923 27740
rect 9955 27700 9995 27740
rect 12259 27700 12299 27740
rect 13795 27700 13835 27740
rect 13900 27700 13940 27740
rect 19939 27700 19979 27740
rect 844 27616 884 27656
rect 1036 27616 1076 27656
rect 1612 27616 1652 27656
rect 1802 27616 1842 27656
rect 2003 27616 2043 27656
rect 2179 27616 2219 27656
rect 2375 27616 2415 27656
rect 2566 27616 2606 27656
rect 2764 27616 2804 27656
rect 2955 27616 2995 27656
rect 3155 27616 3195 27656
rect 3331 27616 3371 27656
rect 3916 27616 3956 27656
rect 4112 27611 4152 27651
rect 4295 27635 4335 27675
rect 4492 27616 4532 27656
rect 5068 27616 5108 27656
rect 5251 27616 5291 27656
rect 5752 27616 5792 27656
rect 6232 27616 6272 27656
rect 6401 27616 6441 27656
rect 6700 27607 6740 27647
rect 7267 27616 7307 27656
rect 9688 27616 9728 27656
rect 11875 27616 11915 27656
rect 12643 27616 12683 27656
rect 12748 27616 12788 27656
rect 13228 27616 13268 27656
rect 13370 27584 13410 27624
rect 13694 27616 13734 27656
rect 13996 27607 14036 27647
rect 16291 27616 16331 27656
rect 16675 27616 16715 27656
rect 17251 27616 17291 27656
rect 19660 27616 19700 27656
rect 21859 27616 21899 27656
rect 24355 27616 24395 27656
rect 24940 27616 24980 27656
rect 25790 27616 25830 27656
rect 25900 27616 25940 27656
rect 26092 27616 26132 27656
rect 26275 27607 26315 27647
rect 26755 27607 26795 27647
rect 27235 27607 27275 27647
rect 27715 27607 27755 27647
rect 28195 27607 28235 27647
rect 28675 27607 28715 27647
rect 29155 27607 29195 27647
rect 30883 27607 30923 27647
rect 5587 27532 5627 27572
rect 9523 27532 9563 27572
rect 16876 27532 16916 27572
rect 22243 27532 22283 27572
rect 24739 27532 24779 27572
rect 26428 27532 26468 27572
rect 26908 27532 26948 27572
rect 27388 27532 27428 27572
rect 28348 27532 28388 27572
rect 28828 27532 28868 27572
rect 29308 27532 29348 27572
rect 31036 27532 31076 27572
rect 1420 27448 1460 27488
rect 1612 27448 1652 27488
rect 3724 27448 3764 27488
rect 4396 27448 4436 27488
rect 4876 27448 4916 27488
rect 19180 27448 19220 27488
rect 25612 27448 25652 27488
rect 29644 27448 29684 27488
rect 30028 27448 30068 27488
rect 30412 27448 30452 27488
rect 844 27364 884 27404
rect 3331 27364 3371 27404
rect 6403 27364 6443 27404
rect 9196 27364 9236 27404
rect 14380 27364 14420 27404
rect 19468 27364 19508 27404
rect 22828 27364 22868 27404
rect 25804 27364 25844 27404
rect 3112 27196 3480 27236
rect 10886 27196 11254 27236
rect 18660 27196 19028 27236
rect 26434 27196 26802 27236
rect 892 27028 932 27068
rect 1987 27028 2027 27068
rect 2371 27028 2411 27068
rect 9676 27028 9716 27068
rect 12172 27028 12212 27068
rect 17356 27028 17396 27068
rect 20524 27028 20564 27068
rect 21676 27028 21716 27068
rect 23500 27028 23540 27068
rect 29116 27028 29156 27068
rect 29644 27028 29684 27068
rect 3532 26944 3572 26984
rect 3916 26944 3956 26984
rect 15436 26944 15476 26984
rect 19372 26944 19412 26984
rect 21484 26944 21524 26984
rect 27148 26944 27188 26984
rect 27724 26944 27764 26984
rect 28780 26944 28820 26984
rect 31084 26944 31124 26984
rect 652 26860 692 26900
rect 1420 26860 1460 26900
rect 1660 26860 1700 26900
rect 13228 26860 13268 26900
rect 13459 26851 13499 26891
rect 29356 26860 29396 26900
rect 1036 26776 1076 26816
rect 1219 26776 1259 26816
rect 1804 26776 1844 26816
rect 1987 26776 2027 26816
rect 2195 26776 2235 26816
rect 2371 26776 2411 26816
rect 2572 26776 2612 26816
rect 2764 26776 2804 26816
rect 2956 26776 2996 26816
rect 3148 26776 3188 26816
rect 4780 26776 4820 26816
rect 5347 26776 5387 26816
rect 7468 26776 7508 26816
rect 8524 26776 8564 26816
rect 8668 26776 8708 26816
rect 9004 26776 9044 26816
rect 9868 26776 9908 26816
rect 10243 26776 10283 26816
rect 13036 26776 13076 26816
rect 13324 26776 13364 26816
rect 13561 26776 13601 26816
rect 13708 26776 13748 26816
rect 13830 26776 13870 26816
rect 13945 26776 13985 26816
rect 14041 26809 14081 26849
rect 14323 26776 14363 26816
rect 14572 26776 14612 26816
rect 14763 26776 14803 26816
rect 15100 26776 15140 26816
rect 15243 26776 15283 26816
rect 15724 26776 15764 26816
rect 15916 26776 15956 26816
rect 16876 26776 16916 26816
rect 17382 26818 17422 26858
rect 30412 26860 30452 26900
rect 30892 26860 30932 26900
rect 17260 26776 17300 26816
rect 17509 26776 17549 26816
rect 18040 26776 18080 26816
rect 18217 26776 18257 26816
rect 18342 26776 18382 26816
rect 18457 26809 18497 26849
rect 18556 26776 18596 26816
rect 18805 26776 18845 26816
rect 18940 26776 18980 26816
rect 19075 26776 19115 26816
rect 19180 26776 19220 26816
rect 19564 26776 19604 26816
rect 20428 26776 20468 26816
rect 20620 26776 20660 26816
rect 20812 26776 20852 26816
rect 22300 26776 22340 26816
rect 23308 26776 23348 26816
rect 24172 26776 24212 26816
rect 26371 26776 26411 26816
rect 26942 26776 26982 26816
rect 27052 26776 27092 26816
rect 27254 26776 27294 26816
rect 27427 26776 27467 26816
rect 27724 26776 27764 26816
rect 27904 26776 27944 26816
rect 28385 26776 28425 26816
rect 28588 26776 28628 26816
rect 29548 26776 29588 26816
rect 29733 26773 29773 26813
rect 29921 26776 29961 26816
rect 30124 26776 30164 26816
rect 30316 26776 30356 26816
rect 30508 26776 30548 26816
rect 4963 26692 5003 26732
rect 8323 26692 8363 26732
rect 15580 26692 15620 26732
rect 24451 26692 24491 26732
rect 26755 26692 26795 26732
rect 28060 26692 28100 26732
rect 1132 26608 1172 26648
rect 2755 26608 2795 26648
rect 3139 26608 3179 26648
rect 4108 26608 4148 26648
rect 7276 26608 7316 26648
rect 8140 26608 8180 26648
rect 8620 26608 8660 26648
rect 12364 26608 12404 26648
rect 13228 26608 13268 26648
rect 14092 26608 14132 26648
rect 14668 26608 14708 26648
rect 15148 26608 15188 26648
rect 16588 26608 16628 26648
rect 16771 26608 16811 26648
rect 17068 26608 17108 26648
rect 17875 26608 17915 26648
rect 18604 26608 18644 26648
rect 20236 26608 20276 26648
rect 22636 26608 22676 26648
rect 28396 26608 28436 26648
rect 29932 26608 29972 26648
rect 30652 26608 30692 26648
rect 4352 26440 4720 26480
rect 12126 26440 12494 26480
rect 19900 26440 20268 26480
rect 27674 26440 28042 26480
rect 5164 26272 5204 26312
rect 11212 26272 11252 26312
rect 11779 26272 11819 26312
rect 12163 26272 12203 26312
rect 14947 26272 14987 26312
rect 15997 26272 16037 26312
rect 17539 26272 17579 26312
rect 19276 26272 19316 26312
rect 21100 26272 21140 26312
rect 24652 26272 24692 26312
rect 30316 26272 30356 26312
rect 30604 26272 30644 26312
rect 30988 26272 31028 26312
rect 2188 26188 2228 26228
rect 12787 26188 12827 26228
rect 15162 26188 15202 26228
rect 17164 26188 17204 26228
rect 23011 26188 23051 26228
rect 27806 26188 27846 26228
rect 28012 26188 28052 26228
rect 652 26104 692 26144
rect 835 26104 875 26144
rect 1366 26104 1406 26144
rect 1987 26104 2027 26144
rect 2284 26104 2324 26144
rect 2471 26104 2511 26144
rect 2667 26104 2707 26144
rect 3235 26104 3275 26144
rect 5782 26104 5822 26144
rect 5932 26104 5972 26144
rect 6115 26104 6155 26144
rect 6220 26104 6260 26144
rect 7084 26104 7124 26144
rect 7948 26104 7988 26144
rect 8284 26104 8324 26144
rect 8428 26104 8468 26144
rect 9388 26104 9428 26144
rect 9859 26104 9899 26144
rect 10540 26104 10580 26144
rect 11062 26104 11102 26144
rect 11308 26104 11348 26144
rect 11545 26104 11585 26144
rect 11683 26104 11723 26144
rect 11994 26104 12034 26144
rect 12268 26104 12308 26144
rect 12952 26104 12992 26144
rect 1171 26020 1211 26060
rect 2860 26020 2900 26060
rect 5587 26020 5627 26060
rect 13084 26062 13124 26102
rect 13399 26104 13439 26144
rect 13555 26104 13595 26144
rect 13852 26095 13892 26135
rect 13965 26104 14005 26144
rect 14188 26104 14228 26144
rect 14380 26104 14420 26144
rect 14629 26104 14669 26144
rect 14851 26104 14891 26144
rect 15340 26104 15380 26144
rect 9298 26020 9338 26060
rect 10867 26020 10907 26060
rect 14519 26062 14559 26102
rect 15532 26104 15572 26144
rect 15763 26104 15803 26144
rect 16099 26104 16139 26144
rect 16204 26095 16244 26135
rect 16867 26104 16907 26144
rect 17468 26093 17508 26133
rect 17649 26104 17689 26144
rect 17752 26104 17792 26144
rect 17884 26095 17924 26135
rect 18019 26104 18059 26144
rect 18412 26104 18452 26144
rect 18547 26104 18587 26144
rect 18661 26104 18701 26144
rect 18988 26104 19028 26144
rect 19310 26104 19350 26144
rect 20140 26104 20180 26144
rect 20428 26104 20468 26144
rect 21259 26104 21299 26144
rect 21699 26104 21739 26144
rect 22254 26106 22294 26146
rect 11443 26011 11483 26051
rect 13228 26020 13268 26060
rect 16684 26020 16724 26060
rect 21571 26062 21611 26102
rect 22387 26104 22427 26144
rect 22684 26062 22724 26102
rect 22925 26104 22965 26144
rect 23395 26104 23435 26144
rect 23500 26104 23540 26144
rect 23980 26104 24020 26144
rect 26755 26104 26795 26144
rect 27304 26104 27344 26144
rect 27427 26104 27467 26144
rect 27532 26104 27572 26144
rect 28108 26095 28148 26135
rect 28300 26104 28340 26144
rect 28492 26104 28532 26144
rect 28684 26104 28724 26144
rect 28876 26104 28916 26144
rect 29069 26104 29109 26144
rect 29260 26104 29300 26144
rect 29452 26104 29492 26144
rect 29642 26104 29682 26144
rect 30220 26104 30260 26144
rect 30412 26104 30452 26144
rect 17260 26020 17300 26060
rect 19219 26011 19259 26051
rect 21388 26020 21428 26060
rect 22819 26020 22859 26060
rect 24835 26020 24875 26060
rect 27139 26020 27179 26060
rect 27628 26020 27668 26060
rect 30028 26020 30068 26060
rect 835 25936 875 25976
rect 1804 25936 1844 25976
rect 2659 25936 2699 25976
rect 12460 25936 12500 25976
rect 13324 25936 13364 25976
rect 16492 25936 16532 25976
rect 19084 25936 19124 25976
rect 21484 25936 21524 25976
rect 23683 25936 23723 25976
rect 28300 25936 28340 25976
rect 29788 25936 29828 25976
rect 6220 25852 6260 25892
rect 6412 25852 6452 25892
rect 7276 25852 7316 25892
rect 8323 25852 8363 25892
rect 9196 25852 9236 25892
rect 11980 25852 12020 25892
rect 13804 25852 13844 25892
rect 14092 25852 14132 25892
rect 14476 25852 14516 25892
rect 15148 25852 15188 25892
rect 15436 25852 15476 25892
rect 15868 25852 15908 25892
rect 18508 25852 18548 25892
rect 19747 25852 19787 25892
rect 22435 25852 22475 25892
rect 27811 25852 27851 25892
rect 28684 25852 28724 25892
rect 29164 25852 29204 25892
rect 29452 25852 29492 25892
rect 3112 25684 3480 25724
rect 10886 25684 11254 25724
rect 18660 25684 19028 25724
rect 26434 25684 26802 25724
rect 2476 25516 2516 25556
rect 3436 25516 3476 25556
rect 4684 25516 4724 25556
rect 9100 25516 9140 25556
rect 10924 25516 10964 25556
rect 13315 25516 13355 25556
rect 14092 25516 14132 25556
rect 14572 25516 14612 25556
rect 20995 25516 21035 25556
rect 23020 25516 23060 25556
rect 24748 25516 24788 25556
rect 29740 25516 29780 25556
rect 4876 25432 4916 25472
rect 12940 25432 12980 25472
rect 15907 25432 15947 25472
rect 19852 25432 19892 25472
rect 21292 25432 21332 25472
rect 30028 25432 30068 25472
rect 30412 25432 30452 25472
rect 30796 25432 30836 25472
rect 9859 25348 9899 25388
rect 10396 25348 10436 25388
rect 13036 25348 13076 25388
rect 16876 25348 16916 25388
rect 17347 25348 17387 25388
rect 19363 25348 19403 25388
rect 25411 25348 25451 25388
rect 844 25264 884 25304
rect 1027 25264 1067 25304
rect 1132 25264 1172 25304
rect 1996 25264 2036 25304
rect 2188 25264 2228 25304
rect 2860 25255 2900 25295
rect 3148 25264 3188 25304
rect 4108 25264 4148 25304
rect 4387 25264 4427 25304
rect 4492 25264 4532 25304
rect 6787 25264 6827 25304
rect 7372 25264 7412 25304
rect 7756 25264 7796 25304
rect 8812 25264 8852 25304
rect 9148 25264 9188 25304
rect 9292 25264 9332 25304
rect 9719 25264 9759 25304
rect 9964 25264 10004 25304
rect 10195 25264 10235 25304
rect 10828 25264 10868 25304
rect 11029 25264 11069 25304
rect 11404 25264 11444 25304
rect 11788 25264 11828 25304
rect 12163 25264 12203 25304
rect 12268 25264 12308 25304
rect 12717 25264 12757 25304
rect 12879 25264 12919 25304
rect 13157 25264 13197 25304
rect 13310 25264 13350 25304
rect 13612 25264 13652 25304
rect 13804 25264 13844 25304
rect 13987 25264 14027 25304
rect 14092 25264 14132 25304
rect 14284 25264 14324 25304
rect 14406 25264 14446 25304
rect 14524 25297 14564 25337
rect 14755 25264 14795 25304
rect 15063 25264 15103 25304
rect 15619 25264 15659 25304
rect 15724 25264 15764 25304
rect 16396 25264 16436 25304
rect 16492 25264 16532 25304
rect 16780 25264 16820 25304
rect 17083 25264 17123 25304
rect 17227 25264 17267 25304
rect 17452 25264 17492 25304
rect 17971 25264 18011 25304
rect 18211 25264 18251 25304
rect 18625 25264 18665 25304
rect 18892 25264 18932 25304
rect 19223 25264 19263 25304
rect 19466 25264 19506 25304
rect 19756 25297 19796 25337
rect 19891 25264 19931 25304
rect 20013 25297 20053 25337
rect 20332 25264 20372 25304
rect 20707 25264 20747 25304
rect 20812 25264 20852 25304
rect 21292 25264 21332 25304
rect 21484 25264 21524 25304
rect 22348 25264 22388 25304
rect 22723 25264 22763 25304
rect 22827 25264 22867 25304
rect 23212 25264 23252 25304
rect 24076 25264 24116 25304
rect 24940 25264 24980 25304
rect 25228 25264 25268 25304
rect 27331 25264 27371 25304
rect 29260 25306 29300 25346
rect 28588 25264 28628 25304
rect 29070 25264 29110 25304
rect 29452 25264 29492 25304
rect 29645 25264 29685 25304
rect 29836 25264 29876 25304
rect 931 25180 971 25220
rect 2764 25180 2804 25220
rect 4698 25180 4738 25220
rect 7171 25180 7211 25220
rect 8131 25180 8171 25220
rect 16193 25180 16233 25220
rect 19555 25180 19595 25220
rect 23884 25180 23924 25220
rect 27715 25180 27755 25220
rect 27907 25180 27947 25220
rect 28766 25180 28806 25220
rect 28867 25180 28907 25220
rect 1324 25096 1364 25136
rect 2332 25096 2372 25136
rect 7852 25096 7892 25136
rect 10051 25096 10091 25136
rect 10828 25096 10868 25136
rect 11299 25096 11339 25136
rect 12556 25096 12596 25136
rect 13516 25096 13556 25136
rect 14851 25096 14891 25136
rect 14956 25096 14996 25136
rect 16291 25096 16331 25136
rect 17539 25096 17579 25136
rect 18019 25096 18059 25136
rect 18787 25096 18827 25136
rect 19084 25096 19124 25136
rect 20188 25096 20228 25136
rect 21676 25096 21716 25136
rect 22732 25096 22772 25136
rect 25027 25096 25067 25136
rect 28972 25096 29012 25136
rect 29356 25096 29396 25136
rect 4352 24928 4720 24968
rect 12126 24928 12494 24968
rect 19900 24928 20268 24968
rect 27674 24928 28042 24968
rect 2956 24760 2996 24800
rect 4492 24760 4532 24800
rect 7468 24760 7508 24800
rect 8140 24760 8180 24800
rect 8524 24760 8564 24800
rect 8899 24760 8939 24800
rect 13411 24760 13451 24800
rect 14764 24760 14804 24800
rect 15187 24760 15227 24800
rect 17548 24760 17588 24800
rect 18787 24760 18827 24800
rect 22588 24760 22628 24800
rect 23011 24760 23051 24800
rect 643 24676 683 24716
rect 4876 24676 4916 24716
rect 5155 24676 5195 24716
rect 8801 24676 8841 24716
rect 17827 24676 17867 24716
rect 18220 24676 18260 24716
rect 19939 24676 19979 24716
rect 22243 24676 22283 24716
rect 25507 24676 25547 24716
rect 26083 24676 26123 24716
rect 1027 24592 1067 24632
rect 3820 24592 3860 24632
rect 4012 24592 4052 24632
rect 4396 24592 4436 24632
rect 4972 24592 5012 24632
rect 5539 24592 5579 24632
rect 7660 24592 7700 24632
rect 8044 24592 8084 24632
rect 8428 24592 8468 24632
rect 9004 24592 9044 24632
rect 8611 24550 8651 24590
rect 9100 24583 9140 24623
rect 11395 24592 11435 24632
rect 11980 24592 12020 24632
rect 12844 24592 12884 24632
rect 12959 24592 12999 24632
rect 13132 24592 13172 24632
rect 13516 24592 13556 24632
rect 13900 24592 13940 24632
rect 14092 24592 14132 24632
rect 15382 24592 15422 24632
rect 16396 24592 16436 24632
rect 16579 24583 16619 24623
rect 17155 24592 17195 24632
rect 17740 24592 17780 24632
rect 17923 24592 17963 24632
rect 18028 24592 18068 24632
rect 18403 24592 18443 24632
rect 18739 24592 18779 24632
rect 19027 24592 19067 24632
rect 19267 24592 19307 24632
rect 19459 24592 19499 24632
rect 21859 24592 21899 24632
rect 22444 24592 22484 24632
rect 22924 24592 22964 24632
rect 25123 24592 25163 24632
rect 25708 24592 25748 24632
rect 25900 24592 25940 24632
rect 26467 24592 26507 24632
rect 28918 24592 28958 24632
rect 29068 24592 29108 24632
rect 29260 24592 29300 24632
rect 29836 24592 29876 24632
rect 30028 24592 30068 24632
rect 9475 24508 9515 24548
rect 11779 24508 11819 24548
rect 16732 24508 16772 24548
rect 28723 24508 28763 24548
rect 2572 24424 2612 24464
rect 12844 24424 12884 24464
rect 17251 24424 17291 24464
rect 18448 24424 18488 24464
rect 23212 24424 23252 24464
rect 29452 24424 29492 24464
rect 30220 24424 30260 24464
rect 30604 24424 30644 24464
rect 30988 24424 31028 24464
rect 3148 24340 3188 24380
rect 12652 24340 12692 24380
rect 15724 24340 15764 24380
rect 20332 24340 20372 24380
rect 22732 24340 22772 24380
rect 25708 24340 25748 24380
rect 28396 24340 28436 24380
rect 29164 24340 29204 24380
rect 29836 24340 29876 24380
rect 3112 24172 3480 24212
rect 10886 24172 11254 24212
rect 18660 24172 19028 24212
rect 26434 24172 26802 24212
rect 1123 24004 1163 24044
rect 6787 24004 6827 24044
rect 12700 24004 12740 24044
rect 16588 24004 16628 24044
rect 19267 24004 19307 24044
rect 21955 24004 21995 24044
rect 23788 24004 23828 24044
rect 25891 24004 25931 24044
rect 27436 24004 27476 24044
rect 28588 24004 28628 24044
rect 29836 24004 29876 24044
rect 652 23920 692 23960
rect 3340 23920 3380 23960
rect 12844 23920 12884 23960
rect 15628 23920 15668 23960
rect 20332 23920 20372 23960
rect 30307 23920 30347 23960
rect 3532 23836 3572 23876
rect 652 23752 692 23792
rect 777 23752 817 23792
rect 940 23752 980 23792
rect 1420 23752 1460 23792
rect 2284 23752 2324 23792
rect 2668 23752 2708 23792
rect 2947 23752 2987 23792
rect 3907 23752 3947 23792
rect 6124 23752 6164 23792
rect 6430 23794 6470 23834
rect 8242 23836 8282 23876
rect 9772 23836 9812 23876
rect 15139 23836 15179 23876
rect 15724 23836 15764 23876
rect 20563 23864 20603 23904
rect 21292 23836 21332 23876
rect 21523 23827 21563 23867
rect 21970 23836 22010 23876
rect 22627 23836 22667 23876
rect 28924 23836 28964 23876
rect 6782 23752 6822 23792
rect 7084 23752 7124 23792
rect 7795 23752 7835 23792
rect 8332 23752 8372 23792
rect 9004 23752 9044 23792
rect 9196 23752 9236 23792
rect 9859 23752 9899 23792
rect 10531 23752 10571 23792
rect 11164 23752 11204 23792
rect 11308 23752 11348 23792
rect 12268 23752 12308 23792
rect 12556 23752 12596 23792
rect 14755 23752 14795 23792
rect 15388 23752 15428 23792
rect 15567 23752 15607 23792
rect 15859 23752 15899 23792
rect 16079 23752 16119 23792
rect 16209 23752 16249 23792
rect 16312 23752 16352 23792
rect 16444 23752 16484 23792
rect 16579 23752 16619 23792
rect 16876 23752 16916 23792
rect 17251 23752 17291 23792
rect 17644 23752 17684 23792
rect 18211 23752 18251 23792
rect 18316 23752 18356 23792
rect 18979 23752 19019 23792
rect 19084 23752 19124 23792
rect 19741 23752 19781 23792
rect 19852 23752 19892 23792
rect 20515 23752 20555 23792
rect 21004 23752 21044 23792
rect 21388 23752 21428 23792
rect 21625 23752 21665 23792
rect 22060 23752 22100 23792
rect 22507 23752 22547 23792
rect 22732 23752 22772 23792
rect 23116 23752 23156 23792
rect 23980 23752 24020 23792
rect 24940 23752 24980 23792
rect 25156 23752 25196 23792
rect 25315 23752 25355 23792
rect 25459 23752 25499 23792
rect 25603 23752 25643 23792
rect 25725 23752 25765 23792
rect 25889 23752 25929 23792
rect 26188 23752 26228 23792
rect 27244 23752 27284 23792
rect 28108 23752 28148 23792
rect 28396 23752 28436 23792
rect 28768 23752 28808 23792
rect 29356 23752 29396 23792
rect 29740 23752 29780 23792
rect 29932 23752 29972 23792
rect 30124 23752 30164 23792
rect 30315 23752 30355 23792
rect 30508 23794 30548 23834
rect 30693 23752 30733 23792
rect 30892 23752 30932 23792
rect 31084 23752 31124 23792
rect 1121 23668 1161 23708
rect 3052 23668 3092 23708
rect 6220 23668 6260 23708
rect 6988 23668 7028 23708
rect 10348 23668 10388 23708
rect 11875 23668 11915 23708
rect 17164 23668 17204 23708
rect 24259 23668 24299 23708
rect 30604 23668 30644 23708
rect 1324 23584 1364 23624
rect 1612 23584 1652 23624
rect 5836 23584 5876 23624
rect 6316 23584 6356 23624
rect 6604 23584 6644 23624
rect 7564 23584 7604 23624
rect 8035 23584 8075 23624
rect 9196 23584 9236 23624
rect 9475 23584 9515 23624
rect 10147 23584 10187 23624
rect 11011 23584 11051 23624
rect 16732 23584 16772 23624
rect 18604 23584 18644 23624
rect 19555 23584 19595 23624
rect 20812 23584 20852 23624
rect 21091 23584 21131 23624
rect 22819 23584 22859 23624
rect 25507 23584 25547 23624
rect 26092 23584 26132 23624
rect 26572 23584 26612 23624
rect 28291 23584 28331 23624
rect 29251 23584 29291 23624
rect 29548 23584 29588 23624
rect 30988 23584 31028 23624
rect 4352 23416 4720 23456
rect 12126 23416 12494 23456
rect 19900 23416 20268 23456
rect 27674 23416 28042 23456
rect 2956 23248 2996 23288
rect 3916 23248 3956 23288
rect 4492 23248 4532 23288
rect 5443 23248 5483 23288
rect 6796 23248 6836 23288
rect 7267 23248 7307 23288
rect 7900 23248 7940 23288
rect 11788 23248 11828 23288
rect 13891 23248 13931 23288
rect 15244 23248 15284 23288
rect 16444 23248 16484 23288
rect 19747 23248 19787 23288
rect 20707 23248 20747 23288
rect 26764 23248 26804 23288
rect 30028 23248 30068 23288
rect 643 23164 683 23204
rect 6268 23164 6308 23204
rect 7747 23164 7787 23204
rect 16972 23164 17012 23204
rect 20092 23164 20132 23204
rect 20606 23164 20646 23204
rect 20812 23164 20852 23204
rect 24259 23164 24299 23204
rect 1027 23080 1067 23120
rect 3436 23080 3476 23120
rect 3820 23080 3860 23120
rect 4300 23080 4340 23120
rect 5164 23080 5204 23120
rect 5731 23080 5771 23120
rect 6115 23071 6155 23111
rect 6892 23080 6932 23120
rect 7084 23080 7124 23120
rect 7280 23075 7320 23115
rect 7420 23038 7460 23078
rect 7660 23080 7700 23120
rect 8092 23080 8132 23120
rect 8236 23080 8276 23120
rect 8419 23080 8459 23120
rect 8951 23080 8991 23120
rect 9196 23080 9236 23120
rect 9859 23080 9899 23120
rect 11980 23080 12020 23120
rect 12652 23080 12692 23120
rect 13324 23080 13364 23120
rect 13820 23069 13860 23109
rect 14001 23080 14041 23120
rect 14104 23080 14144 23120
rect 14243 23080 14283 23120
rect 14371 23080 14411 23120
rect 14572 23080 14612 23120
rect 15556 23080 15596 23120
rect 15715 23080 15755 23120
rect 15832 23080 15872 23120
rect 16003 23080 16043 23120
rect 16105 23080 16145 23120
rect 16243 23080 16283 23120
rect 17068 23080 17108 23120
rect 17305 23080 17345 23120
rect 17452 23080 17492 23120
rect 17635 23080 17675 23120
rect 17932 23080 17972 23120
rect 18124 23080 18164 23120
rect 18316 23080 18356 23120
rect 18565 23080 18605 23120
rect 19468 23080 19508 23120
rect 5347 22996 5387 23036
rect 5923 22996 5963 23036
rect 7555 22996 7595 23036
rect 9091 22996 9131 23036
rect 9292 22996 9332 23036
rect 9484 22996 9524 23036
rect 18439 23038 18479 23078
rect 19651 23080 19691 23120
rect 19962 23080 20002 23120
rect 20908 23071 20948 23111
rect 21091 23080 21131 23120
rect 21772 23080 21812 23120
rect 22732 23080 22772 23120
rect 23596 23080 23636 23120
rect 23831 23080 23871 23120
rect 23971 23071 24011 23111
rect 24076 23080 24116 23120
rect 26179 23080 26219 23120
rect 28675 23080 28715 23120
rect 29059 23080 29099 23120
rect 30028 23080 30068 23120
rect 30220 23080 30260 23120
rect 31180 23080 31220 23120
rect 17187 22996 17227 23036
rect 20332 22996 20372 23036
rect 26563 22996 26603 23036
rect 8812 22912 8852 22952
rect 11404 22912 11444 22952
rect 18028 22912 18068 22952
rect 18604 22912 18644 22952
rect 22924 22912 22964 22952
rect 23788 22912 23828 22952
rect 29260 22912 29300 22952
rect 29644 22912 29684 22952
rect 30412 22912 30452 22952
rect 30796 22912 30836 22952
rect 2572 22828 2612 22868
rect 8419 22828 8459 22868
rect 12931 22828 12971 22868
rect 16108 22828 16148 22868
rect 17635 22828 17675 22868
rect 18796 22828 18836 22868
rect 19948 22828 19988 22868
rect 22060 22828 22100 22868
rect 3112 22660 3480 22700
rect 10886 22660 11254 22700
rect 18660 22660 19028 22700
rect 26434 22660 26802 22700
rect 6403 22492 6443 22532
rect 10732 22492 10772 22532
rect 16300 22492 16340 22532
rect 21100 22492 21140 22532
rect 21724 22492 21764 22532
rect 24364 22492 24404 22532
rect 25219 22492 25259 22532
rect 26572 22492 26612 22532
rect 27052 22492 27092 22532
rect 8227 22408 8267 22448
rect 10348 22408 10388 22448
rect 12844 22408 12884 22448
rect 17452 22408 17492 22448
rect 30604 22408 30644 22448
rect 30988 22408 31028 22448
rect 748 22324 788 22364
rect 4579 22324 4619 22364
rect 5155 22324 5195 22364
rect 5356 22324 5396 22364
rect 1459 22282 1499 22322
rect 5571 22324 5611 22364
rect 5836 22324 5876 22364
rect 6067 22315 6107 22355
rect 7180 22324 7220 22364
rect 7372 22324 7412 22364
rect 7948 22324 7988 22364
rect 8131 22324 8171 22364
rect 8707 22324 8747 22364
rect 12643 22324 12683 22364
rect 14908 22324 14948 22364
rect 16579 22324 16619 22364
rect 16972 22324 17012 22364
rect 17548 22324 17588 22364
rect 21379 22324 21419 22364
rect 22060 22324 22100 22364
rect 1804 22240 1844 22280
rect 1948 22240 1988 22280
rect 2572 22240 2612 22280
rect 2956 22240 2996 22280
rect 3523 22240 3563 22280
rect 3628 22240 3668 22280
rect 4055 22240 4095 22280
rect 4195 22240 4235 22280
rect 4300 22240 4340 22280
rect 4963 22240 5003 22280
rect 5452 22240 5492 22280
rect 5669 22240 5709 22280
rect 5932 22240 5972 22280
rect 6169 22240 6209 22280
rect 6401 22240 6441 22280
rect 6698 22273 6738 22313
rect 6839 22240 6879 22280
rect 6979 22240 7019 22280
rect 7084 22240 7124 22280
rect 7555 22240 7595 22280
rect 8515 22240 8555 22280
rect 8947 22240 8987 22280
rect 9868 22240 9908 22280
rect 12259 22240 12299 22280
rect 13242 22240 13282 22280
rect 13516 22240 13556 22280
rect 13987 22240 14027 22280
rect 14707 22240 14747 22280
rect 15244 22240 15284 22280
rect 15388 22240 15428 22280
rect 15532 22240 15572 22280
rect 15715 22240 15755 22280
rect 15820 22240 15860 22280
rect 16012 22240 16052 22280
rect 16151 22240 16191 22280
rect 16261 22240 16301 22280
rect 16459 22240 16499 22280
rect 16684 22240 16724 22280
rect 17155 22240 17195 22280
rect 18028 22240 18068 22280
rect 18616 22240 18656 22280
rect 19171 22240 19211 22280
rect 21239 22240 21279 22280
rect 21484 22240 21524 22280
rect 21868 22240 21908 22280
rect 22435 22240 22475 22280
rect 24940 22240 24980 22280
rect 25504 22273 25544 22313
rect 25603 22240 25643 22280
rect 25900 22240 25940 22280
rect 26764 22240 26804 22280
rect 26899 22240 26939 22280
rect 27004 22240 27044 22280
rect 29155 22240 29195 22280
rect 29726 22240 29766 22280
rect 30028 22240 30068 22280
rect 30220 22240 30260 22280
rect 30403 22240 30443 22280
rect 1603 22156 1643 22196
rect 4387 22156 4427 22196
rect 7852 22156 7892 22196
rect 13132 22156 13172 22196
rect 14380 22156 14420 22196
rect 15619 22156 15659 22196
rect 18787 22156 18827 22196
rect 27235 22156 27275 22196
rect 29539 22156 29579 22196
rect 988 22072 1028 22112
rect 1267 22072 1307 22112
rect 1900 22072 1940 22112
rect 3052 22072 3092 22112
rect 3916 22072 3956 22112
rect 4675 22072 4715 22112
rect 6604 22072 6644 22112
rect 9148 22072 9188 22112
rect 9676 22072 9716 22112
rect 9955 22072 9995 22112
rect 16771 22072 16811 22112
rect 17836 22072 17876 22112
rect 18115 22072 18155 22112
rect 18451 22072 18491 22112
rect 21571 22072 21611 22112
rect 24748 22072 24788 22112
rect 25027 22072 25067 22112
rect 25747 22072 25787 22112
rect 29827 22072 29867 22112
rect 29932 22072 29972 22112
rect 30316 22072 30356 22112
rect 4352 21904 4720 21944
rect 12126 21904 12494 21944
rect 19900 21904 20268 21944
rect 27674 21904 28042 21944
rect 883 21736 923 21776
rect 5443 21736 5483 21776
rect 5548 21736 5588 21776
rect 6115 21736 6155 21776
rect 6595 21736 6635 21776
rect 6988 21736 7028 21776
rect 7660 21736 7700 21776
rect 9532 21736 9572 21776
rect 11443 21736 11483 21776
rect 13324 21736 13364 21776
rect 15043 21736 15083 21776
rect 18076 21736 18116 21776
rect 18787 21736 18827 21776
rect 24700 21736 24740 21776
rect 25516 21736 25556 21776
rect 28012 21736 28052 21776
rect 5176 21652 5216 21692
rect 5656 21652 5696 21692
rect 6807 21652 6847 21692
rect 8227 21652 8267 21692
rect 9043 21652 9083 21692
rect 10963 21652 11003 21692
rect 16204 21652 16244 21692
rect 16972 21652 17012 21692
rect 17731 21652 17771 21692
rect 20620 21652 20660 21692
rect 25324 21652 25364 21692
rect 1075 21568 1115 21608
rect 1315 21568 1355 21608
rect 1420 21568 1460 21608
rect 1180 21526 1220 21566
rect 1795 21568 1835 21608
rect 2572 21568 2612 21608
rect 2809 21568 2849 21608
rect 2956 21568 2996 21608
rect 3139 21568 3179 21608
rect 3523 21568 3563 21608
rect 3638 21568 3678 21608
rect 4363 21568 4403 21608
rect 4588 21568 4628 21608
rect 4865 21568 4905 21608
rect 4972 21568 5012 21608
rect 5347 21568 5387 21608
rect 5803 21568 5843 21608
rect 6499 21568 6539 21608
rect 7084 21568 7124 21608
rect 1516 21484 1556 21524
rect 2476 21484 2516 21524
rect 2691 21484 2731 21524
rect 4483 21484 4523 21524
rect 4684 21484 4724 21524
rect 5909 21484 5949 21524
rect 6028 21526 6068 21566
rect 7301 21568 7341 21608
rect 7454 21568 7494 21608
rect 7756 21559 7796 21599
rect 7203 21484 7243 21524
rect 7900 21526 7940 21566
rect 8140 21568 8180 21608
rect 8728 21568 8768 21608
rect 9238 21568 9278 21608
rect 9379 21559 9419 21599
rect 9859 21559 9899 21599
rect 10339 21559 10379 21599
rect 11128 21568 11168 21608
rect 11608 21568 11648 21608
rect 11788 21568 11828 21608
rect 12844 21568 12884 21608
rect 13228 21568 13268 21608
rect 13655 21568 13695 21608
rect 13900 21568 13940 21608
rect 14371 21568 14411 21608
rect 15331 21568 15371 21608
rect 15724 21568 15764 21608
rect 15916 21568 15956 21608
rect 16108 21568 16148 21608
rect 16300 21568 16340 21608
rect 16588 21568 16628 21608
rect 16780 21568 16820 21608
rect 17068 21568 17108 21608
rect 17305 21568 17345 21608
rect 17419 21568 17459 21608
rect 17644 21568 17684 21608
rect 17923 21559 17963 21599
rect 18892 21568 18932 21608
rect 19852 21568 19892 21608
rect 20236 21568 20276 21608
rect 20515 21568 20555 21608
rect 21100 21568 21140 21608
rect 21475 21568 21515 21608
rect 23971 21610 24011 21650
rect 23596 21568 23636 21608
rect 23779 21568 23819 21608
rect 24097 21568 24137 21608
rect 24403 21568 24443 21608
rect 24547 21559 24587 21599
rect 25123 21568 25163 21608
rect 27427 21568 27467 21608
rect 27811 21568 27851 21608
rect 29923 21568 29963 21608
rect 30307 21568 30347 21608
rect 8035 21484 8075 21524
rect 8563 21484 8603 21524
rect 10012 21484 10052 21524
rect 10492 21484 10532 21524
rect 13795 21484 13835 21524
rect 13996 21484 14036 21524
rect 14188 21484 14228 21524
rect 14764 21484 14804 21524
rect 14947 21484 14987 21524
rect 15523 21484 15563 21524
rect 17187 21484 17227 21524
rect 17539 21484 17579 21524
rect 18604 21484 18644 21524
rect 19459 21484 19499 21524
rect 24268 21484 24308 21524
rect 14668 21400 14708 21440
rect 23404 21400 23444 21440
rect 24172 21400 24212 21440
rect 25095 21400 25135 21440
rect 30508 21400 30548 21440
rect 30892 21400 30932 21440
rect 2188 21316 2228 21356
rect 3139 21316 3179 21356
rect 3811 21316 3851 21356
rect 5164 21316 5204 21356
rect 6796 21316 6836 21356
rect 7459 21316 7499 21356
rect 12460 21316 12500 21356
rect 15724 21316 15764 21356
rect 16588 21316 16628 21356
rect 18364 21316 18404 21356
rect 19084 21316 19124 21356
rect 20908 21316 20948 21356
rect 23779 21316 23819 21356
rect 3112 21148 3480 21188
rect 10886 21148 11254 21188
rect 18660 21148 19028 21188
rect 26434 21148 26802 21188
rect 6316 20980 6356 21020
rect 7939 20980 7979 21020
rect 9004 20980 9044 21020
rect 10348 20980 10388 21020
rect 24556 20980 24596 21020
rect 25228 20980 25268 21020
rect 29740 20980 29780 21020
rect 30076 20980 30116 21020
rect 30508 20980 30548 21020
rect 1804 20896 1844 20936
rect 2179 20896 2219 20936
rect 5068 20896 5108 20936
rect 9772 20896 9812 20936
rect 14764 20896 14804 20936
rect 20803 20896 20843 20936
rect 27244 20896 27284 20936
rect 30892 20896 30932 20936
rect 844 20812 884 20852
rect 1075 20803 1115 20843
rect 1324 20812 1364 20852
rect 1900 20812 1940 20852
rect 2083 20812 2123 20852
rect 2659 20812 2699 20852
rect 3667 20803 3707 20843
rect 5395 20812 5435 20852
rect 7276 20812 7316 20852
rect 9388 20812 9428 20852
rect 940 20728 980 20768
rect 1177 20728 1217 20768
rect 1507 20728 1547 20768
rect 2467 20728 2507 20768
rect 3190 20728 3230 20768
rect 3532 20728 3572 20768
rect 3769 20728 3809 20768
rect 4099 20728 4139 20768
rect 4204 20728 4244 20768
rect 5590 20728 5630 20768
rect 5836 20728 5876 20768
rect 6019 20728 6059 20768
rect 6219 20728 6259 20768
rect 6412 20728 6452 20768
rect 6604 20728 6644 20768
rect 6787 20728 6827 20768
rect 6955 20728 6995 20768
rect 7075 20728 7115 20768
rect 7180 20728 7220 20768
rect 7612 20728 7652 20768
rect 7756 20728 7796 20768
rect 7939 20728 7979 20768
rect 8044 20739 8084 20779
rect 8189 20728 8229 20768
rect 8323 20728 8363 20768
rect 8500 20728 8540 20768
rect 8707 20728 8747 20768
rect 9676 20728 9716 20768
rect 9868 20728 9908 20768
rect 10156 20728 10196 20768
rect 12796 20770 12836 20810
rect 13397 20812 13437 20852
rect 14092 20812 14132 20852
rect 14284 20812 14324 20852
rect 14860 20812 14900 20852
rect 15139 20812 15179 20852
rect 15340 20812 15380 20852
rect 17068 20812 17108 20852
rect 17251 20812 17291 20852
rect 17827 20812 17867 20852
rect 18019 20812 18059 20852
rect 18595 20812 18635 20852
rect 23203 20812 23243 20852
rect 30316 20812 30356 20852
rect 11020 20728 11060 20768
rect 11704 20728 11744 20768
rect 11872 20728 11912 20768
rect 12322 20728 12362 20768
rect 12931 20728 12971 20768
rect 13036 20728 13076 20768
rect 13291 20728 13331 20768
rect 13514 20728 13554 20768
rect 13751 20728 13791 20768
rect 13891 20728 13931 20768
rect 13996 20728 14036 20768
rect 14467 20728 14507 20768
rect 14999 20728 15039 20768
rect 15244 20728 15284 20768
rect 16120 20728 16160 20768
rect 16295 20728 16335 20768
rect 16483 20728 16523 20768
rect 16727 20728 16767 20768
rect 16867 20728 16907 20768
rect 16972 20728 17012 20768
rect 17635 20728 17675 20768
rect 18403 20728 18443 20768
rect 18739 20728 18779 20768
rect 19267 20761 19307 20801
rect 20033 20728 20073 20768
rect 20332 20728 20372 20768
rect 20620 20728 20660 20768
rect 21088 20761 21128 20801
rect 21187 20728 21227 20768
rect 21661 20728 21701 20768
rect 21772 20728 21812 20768
rect 22348 20728 22388 20768
rect 22467 20728 22507 20768
rect 22585 20728 22625 20768
rect 23404 20728 23444 20768
rect 23635 20728 23675 20768
rect 23836 20728 23876 20768
rect 24259 20728 24299 20768
rect 24931 20728 24971 20768
rect 25242 20728 25282 20768
rect 26092 20728 26132 20768
rect 26380 20728 26420 20768
rect 29155 20728 29195 20768
rect 29740 20728 29780 20768
rect 29932 20728 29972 20768
rect 30508 20728 30548 20768
rect 30700 20728 30740 20768
rect 9015 20644 9055 20684
rect 13123 20644 13163 20684
rect 15955 20644 15995 20684
rect 19420 20644 19460 20684
rect 24364 20644 24404 20684
rect 24570 20644 24610 20684
rect 27052 20644 27092 20684
rect 29539 20644 29579 20684
rect 2995 20560 3035 20600
rect 3436 20560 3476 20600
rect 4492 20560 4532 20600
rect 5932 20560 5972 20600
rect 6700 20560 6740 20600
rect 7459 20560 7499 20600
rect 8803 20560 8843 20600
rect 9148 20560 9188 20600
rect 10003 20560 10043 20600
rect 10915 20560 10955 20600
rect 11212 20560 11252 20600
rect 11539 20560 11579 20600
rect 12028 20560 12068 20600
rect 12508 20560 12548 20600
rect 13603 20560 13643 20600
rect 16396 20560 16436 20600
rect 17347 20560 17387 20600
rect 18115 20560 18155 20600
rect 18940 20560 18980 20600
rect 20131 20560 20171 20600
rect 20236 20560 20276 20600
rect 20476 20560 20516 20600
rect 21307 20560 21347 20600
rect 21475 20560 21515 20600
rect 22252 20560 22292 20600
rect 25027 20560 25067 20600
rect 25420 20560 25460 20600
rect 4352 20392 4720 20432
rect 12126 20392 12494 20432
rect 19900 20392 20268 20432
rect 27674 20392 28042 20432
rect 1132 20224 1172 20264
rect 2371 20224 2411 20264
rect 3628 20224 3668 20264
rect 4060 20224 4100 20264
rect 5443 20224 5483 20264
rect 9571 20224 9611 20264
rect 10444 20224 10484 20264
rect 1603 20140 1643 20180
rect 3425 20140 3465 20180
rect 6616 20182 6656 20222
rect 13804 20224 13844 20264
rect 14083 20224 14123 20264
rect 14563 20224 14603 20264
rect 16483 20224 16523 20264
rect 18691 20224 18731 20264
rect 19852 20224 19892 20264
rect 21580 20224 21620 20264
rect 23980 20224 24020 20264
rect 28876 20224 28916 20264
rect 7267 20140 7307 20180
rect 8044 20140 8084 20180
rect 844 20056 884 20096
rect 986 20053 1026 20093
rect 1291 20056 1331 20096
rect 1517 20056 1557 20096
rect 1771 20056 1811 20096
rect 1996 20056 2036 20096
rect 2275 20056 2315 20096
rect 2583 20056 2623 20096
rect 3052 20056 3092 20096
rect 3289 20056 3329 20096
rect 3724 20047 3764 20087
rect 3916 20056 3956 20096
rect 4204 20056 4244 20096
rect 4387 20056 4427 20096
rect 4535 20056 4575 20096
rect 4780 20056 4820 20096
rect 5092 20056 5132 20096
rect 5251 20056 5291 20096
rect 5827 20098 5867 20138
rect 6403 20098 6443 20138
rect 6835 20098 6875 20138
rect 9148 20140 9188 20180
rect 9783 20140 9823 20180
rect 10924 20140 10964 20180
rect 12460 20140 12500 20180
rect 12979 20140 13019 20180
rect 14188 20140 14228 20180
rect 15134 20140 15174 20180
rect 16972 20140 17012 20180
rect 19555 20140 19595 20180
rect 22147 20140 22187 20180
rect 25132 20140 25172 20180
rect 29212 20140 29252 20180
rect 30268 20140 30308 20180
rect 5368 20056 5408 20096
rect 5539 20056 5579 20096
rect 5661 20056 5701 20096
rect 1411 19972 1451 20012
rect 1891 19972 1931 20012
rect 2092 19972 2132 20012
rect 2956 19972 2996 20012
rect 3187 19963 3227 20003
rect 4675 19972 4715 20012
rect 4876 19972 4916 20012
rect 5932 20014 5972 20054
rect 6259 20014 6299 20054
rect 6536 20014 6576 20054
rect 6940 20056 6980 20096
rect 7180 20056 7220 20096
rect 7564 20056 7604 20096
rect 7683 20056 7723 20096
rect 7801 20056 7841 20096
rect 7948 20056 7988 20096
rect 8140 20056 8180 20096
rect 8279 20056 8319 20096
rect 8524 20056 8564 20096
rect 8812 20056 8852 20096
rect 9004 20056 9044 20096
rect 9292 20056 9332 20096
rect 9475 20056 9515 20096
rect 6124 19972 6164 20012
rect 6693 19972 6733 20012
rect 7075 19972 7115 20012
rect 7468 19972 7508 20012
rect 8419 19972 8459 20012
rect 8620 19972 8660 20012
rect 9916 20014 9956 20054
rect 10156 20056 10196 20096
rect 10539 20056 10579 20096
rect 10659 20056 10699 20096
rect 10777 20056 10817 20096
rect 11020 20056 11060 20096
rect 11139 20056 11179 20096
rect 11257 20056 11297 20096
rect 11980 20056 12020 20096
rect 12355 20056 12395 20096
rect 12666 20056 12706 20096
rect 13174 20056 13214 20096
rect 13372 20056 13412 20096
rect 13493 20056 13533 20096
rect 13612 20056 13652 20096
rect 13982 20056 14022 20096
rect 14284 20047 14324 20087
rect 14465 20056 14505 20096
rect 14668 20056 14708 20096
rect 14764 20047 14804 20087
rect 15340 20056 15380 20096
rect 15436 20047 15476 20087
rect 15883 20056 15923 20096
rect 16106 20056 16146 20096
rect 16387 20056 16427 20096
rect 16695 20056 16735 20096
rect 16877 20061 16917 20101
rect 17178 20056 17218 20096
rect 17452 20056 17492 20096
rect 17827 20056 17867 20096
rect 18115 20056 18155 20096
rect 18359 20056 18399 20096
rect 18604 20056 18644 20096
rect 19084 20056 19124 20096
rect 19267 20056 19307 20096
rect 19372 20056 19412 20096
rect 19756 20056 19796 20096
rect 19900 20056 19940 20096
rect 20428 20056 20468 20096
rect 20812 20056 20852 20096
rect 21571 20056 21611 20096
rect 21676 20056 21716 20096
rect 22435 20056 22475 20096
rect 23116 20056 23156 20096
rect 23692 20056 23732 20096
rect 23940 20056 23980 20096
rect 24119 20056 24159 20096
rect 10051 19972 10091 20012
rect 10252 19972 10292 20012
rect 16003 19972 16043 20012
rect 16204 19972 16244 20012
rect 17644 19972 17684 20012
rect 18220 19972 18260 20012
rect 18499 19972 18539 20012
rect 22051 19972 22091 20012
rect 22627 19972 22667 20012
rect 23815 20014 23855 20054
rect 24364 20056 24404 20096
rect 24748 20056 24788 20096
rect 25027 20056 25067 20096
rect 27619 20056 27659 20096
rect 28204 20056 28244 20096
rect 29059 20047 29099 20087
rect 30412 20056 30452 20096
rect 23026 19972 23066 20012
rect 24259 19972 24299 20012
rect 24460 19972 24500 20012
rect 28003 19972 28043 20012
rect 6028 19888 6068 19928
rect 17308 19888 17348 19928
rect 19276 19888 19316 19928
rect 21004 19888 21044 19928
rect 21868 19888 21908 19928
rect 25420 19888 25460 19928
rect 29548 19888 29588 19928
rect 29932 19888 29972 19928
rect 2572 19804 2612 19844
rect 3427 19804 3467 19844
rect 4387 19804 4427 19844
rect 8812 19804 8852 19844
rect 9772 19804 9812 19844
rect 11587 19804 11627 19844
rect 12652 19804 12692 19844
rect 15139 19804 15179 19844
rect 16684 19804 16724 19844
rect 17164 19804 17204 19844
rect 20188 19804 20228 19844
rect 22924 19804 22964 19844
rect 25708 19804 25748 19844
rect 3112 19636 3480 19676
rect 10886 19636 11254 19676
rect 18660 19636 19028 19676
rect 26434 19636 26802 19676
rect 3139 19468 3179 19508
rect 3619 19468 3659 19508
rect 7747 19468 7787 19508
rect 9955 19468 9995 19508
rect 11203 19468 11243 19508
rect 13036 19468 13076 19508
rect 14275 19468 14315 19508
rect 15235 19468 15275 19508
rect 16195 19468 16235 19508
rect 16675 19468 16715 19508
rect 17452 19468 17492 19508
rect 20716 19468 20756 19508
rect 22684 19468 22724 19508
rect 28108 19468 28148 19508
rect 9724 19375 9764 19415
rect 12460 19384 12500 19424
rect 18604 19384 18644 19424
rect 22348 19384 22388 19424
rect 28780 19384 28820 19424
rect 1027 19300 1067 19340
rect 1228 19300 1268 19340
rect 1420 19300 1460 19340
rect 1996 19300 2036 19340
rect 2188 19300 2228 19340
rect 4204 19300 4244 19340
rect 5932 19300 5972 19340
rect 6163 19291 6203 19331
rect 6723 19300 6763 19340
rect 8707 19300 8747 19340
rect 8908 19300 8948 19340
rect 17731 19300 17771 19340
rect 17932 19300 17972 19340
rect 23251 19291 23291 19331
rect 25132 19300 25172 19340
rect 26284 19300 26324 19340
rect 27676 19300 27716 19340
rect 887 19216 927 19256
rect 1132 19216 1172 19256
rect 1603 19216 1643 19256
rect 2284 19216 2324 19256
rect 2403 19216 2443 19256
rect 2521 19216 2561 19256
rect 2764 19216 2804 19256
rect 2883 19216 2923 19256
rect 2995 19216 3035 19256
rect 3436 19216 3476 19256
rect 3916 19216 3956 19256
rect 4300 19216 4340 19256
rect 4419 19216 4459 19256
rect 4537 19216 4577 19256
rect 4780 19216 4820 19256
rect 4899 19216 4939 19256
rect 5017 19216 5057 19256
rect 5260 19216 5300 19256
rect 5587 19216 5627 19256
rect 6028 19216 6068 19256
rect 6265 19216 6305 19256
rect 6604 19216 6644 19256
rect 6841 19216 6881 19256
rect 6990 19216 7030 19256
rect 7097 19216 7137 19256
rect 7229 19216 7269 19256
rect 7363 19216 7403 19256
rect 7539 19216 7579 19256
rect 7759 19227 7799 19267
rect 7891 19216 7931 19256
rect 7997 19216 8037 19256
rect 8131 19216 8171 19256
rect 8308 19216 8348 19256
rect 8587 19216 8627 19256
rect 8812 19216 8852 19256
rect 9196 19216 9236 19256
rect 9388 19216 9428 19256
rect 9763 19216 9803 19256
rect 10241 19216 10281 19256
rect 10540 19216 10580 19256
rect 10828 19216 10868 19256
rect 11201 19216 11241 19256
rect 11500 19216 11540 19256
rect 11635 19216 11675 19256
rect 11836 19216 11876 19256
rect 12652 19216 12692 19256
rect 13036 19216 13076 19256
rect 13228 19216 13268 19256
rect 13516 19216 13556 19256
rect 13996 19216 14036 19256
rect 14270 19216 14310 19256
rect 14574 19216 14614 19256
rect 14725 19216 14765 19256
rect 14851 19216 14891 19256
rect 14956 19216 14996 19256
rect 15532 19216 15572 19256
rect 16054 19216 16094 19256
rect 16492 19216 16532 19256
rect 16972 19216 17012 19256
rect 17155 19216 17195 19256
rect 17463 19216 17503 19256
rect 17611 19216 17651 19256
rect 17836 19216 17876 19256
rect 18124 19216 18164 19256
rect 18316 19216 18356 19256
rect 18988 19207 19028 19247
rect 19276 19216 19316 19256
rect 20236 19216 20276 19256
rect 20524 19216 20564 19256
rect 20851 19216 20891 19256
rect 21004 19216 21044 19256
rect 21763 19216 21803 19256
rect 21868 19216 21908 19256
rect 22348 19216 22388 19256
rect 22540 19216 22580 19256
rect 22780 19216 22820 19256
rect 23116 19216 23156 19256
rect 23353 19216 23393 19256
rect 23500 19216 23540 19256
rect 23692 19216 23732 19256
rect 24076 19216 24116 19256
rect 24195 19216 24235 19256
rect 24313 19216 24353 19256
rect 24460 19216 24500 19256
rect 25324 19216 25364 19256
rect 26177 19216 26217 19256
rect 26380 19216 26420 19256
rect 26668 19216 26708 19256
rect 27475 19216 27515 19256
rect 28010 19221 28050 19261
rect 28204 19216 28244 19256
rect 28396 19216 28436 19256
rect 28588 19216 28628 19256
rect 1900 19132 1940 19172
rect 3137 19132 3177 19172
rect 3614 19132 3654 19172
rect 5452 19132 5492 19172
rect 6508 19132 6548 19172
rect 9484 19132 9524 19172
rect 10339 19132 10379 19172
rect 13708 19132 13748 19172
rect 15233 19132 15273 19172
rect 16190 19132 16230 19172
rect 16673 19132 16713 19172
rect 17260 19132 17300 19172
rect 18892 19132 18932 19172
rect 27340 19132 27380 19172
rect 2668 19048 2708 19088
rect 3340 19048 3380 19088
rect 3820 19048 3860 19088
rect 4684 19048 4724 19088
rect 6979 19048 7019 19088
rect 9955 19048 9995 19088
rect 10444 19048 10484 19088
rect 10723 19048 10763 19088
rect 11020 19048 11060 19088
rect 11404 19048 11444 19088
rect 12739 19048 12779 19088
rect 13411 19048 13451 19088
rect 14476 19048 14516 19088
rect 15043 19048 15083 19088
rect 15436 19048 15476 19088
rect 15859 19048 15899 19088
rect 16396 19048 16436 19088
rect 16876 19048 16916 19088
rect 18220 19048 18260 19088
rect 19564 19048 19604 19088
rect 21100 19048 21140 19088
rect 22156 19048 22196 19088
rect 23020 19048 23060 19088
rect 23500 19048 23540 19088
rect 23980 19048 24020 19088
rect 25996 19048 26036 19088
rect 28396 19048 28436 19088
rect 29164 19048 29204 19088
rect 29548 19048 29588 19088
rect 4352 18880 4720 18920
rect 12126 18880 12494 18920
rect 19900 18880 20268 18920
rect 27674 18880 28042 18920
rect 3235 18712 3275 18752
rect 3340 18712 3380 18752
rect 3724 18712 3764 18752
rect 6499 18754 6539 18794
rect 4780 18712 4820 18752
rect 5059 18712 5099 18752
rect 10732 18712 10772 18752
rect 12691 18712 12731 18752
rect 16099 18712 16139 18752
rect 17251 18712 17291 18752
rect 18307 18712 18347 18752
rect 22540 18712 22580 18752
rect 787 18628 827 18668
rect 1612 18628 1652 18668
rect 3134 18628 3174 18668
rect 4204 18628 4244 18668
rect 6616 18670 6656 18710
rect 25132 18712 25172 18752
rect 27916 18712 27956 18752
rect 14558 18628 14598 18668
rect 982 18544 1022 18584
rect 1099 18544 1139 18584
rect 1324 18544 1364 18584
rect 1708 18544 1748 18584
rect 1925 18544 1965 18584
rect 2284 18544 2324 18584
rect 2403 18544 2443 18584
rect 2524 18544 2564 18584
rect 2773 18544 2813 18584
rect 2981 18544 3021 18584
rect 3436 18535 3476 18575
rect 3628 18544 3668 18584
rect 3811 18544 3851 18584
rect 4108 18544 4148 18584
rect 4291 18544 4331 18584
rect 4972 18544 5012 18584
rect 5356 18544 5396 18584
rect 5644 18544 5684 18584
rect 5861 18544 5901 18584
rect 6028 18544 6068 18584
rect 6219 18544 6259 18584
rect 6835 18586 6875 18626
rect 18019 18628 18059 18668
rect 18499 18628 18539 18668
rect 25315 18628 25355 18668
rect 6543 18544 6583 18584
rect 6980 18533 7020 18573
rect 7084 18535 7124 18575
rect 7267 18535 7307 18575
rect 7371 18544 7411 18584
rect 7489 18533 7529 18573
rect 7708 18544 7748 18584
rect 8023 18544 8063 18584
rect 8163 18544 8203 18584
rect 8428 18544 8468 18584
rect 8665 18544 8705 18584
rect 8908 18544 8948 18584
rect 9100 18544 9140 18584
rect 9688 18544 9728 18584
rect 9868 18544 9908 18584
rect 10060 18544 10100 18584
rect 10339 18544 10379 18584
rect 11107 18544 11147 18584
rect 11500 18544 11540 18584
rect 11793 18544 11833 18584
rect 12115 18544 12155 18584
rect 13132 18544 13172 18584
rect 1219 18460 1259 18500
rect 1420 18460 1460 18500
rect 1827 18460 1867 18500
rect 2188 18460 2228 18500
rect 2668 18460 2708 18500
rect 2883 18460 2923 18500
rect 5548 18460 5588 18500
rect 5779 18451 5819 18491
rect 6700 18460 6740 18500
rect 7852 18460 7892 18500
rect 12883 18502 12923 18542
rect 13507 18544 13547 18584
rect 13900 18544 13940 18584
rect 14039 18544 14079 18584
rect 14284 18544 14324 18584
rect 14764 18544 14804 18584
rect 14860 18535 14900 18575
rect 15139 18535 15179 18575
rect 15436 18544 15476 18584
rect 15767 18544 15807 18584
rect 16012 18544 16052 18584
rect 16324 18544 16364 18584
rect 16483 18544 16523 18584
rect 16600 18544 16640 18584
rect 16766 18544 16806 18584
rect 16867 18544 16907 18584
rect 17092 18544 17132 18584
rect 17251 18544 17291 18584
rect 17368 18544 17408 18584
rect 17535 18533 17575 18573
rect 17641 18544 17681 18584
rect 18220 18544 18260 18584
rect 18883 18544 18923 18584
rect 21091 18544 21131 18584
rect 22102 18544 22142 18584
rect 22336 18536 22376 18576
rect 22540 18544 22580 18584
rect 22828 18544 22868 18584
rect 23203 18544 23243 18584
rect 25699 18544 25739 18584
rect 27820 18544 27860 18584
rect 28003 18544 28043 18584
rect 28588 18544 28628 18584
rect 28780 18544 28820 18584
rect 29068 18544 29108 18584
rect 8332 18460 8372 18500
rect 8563 18451 8603 18491
rect 9523 18460 9563 18500
rect 13420 18460 13460 18500
rect 14179 18460 14219 18500
rect 14380 18460 14420 18500
rect 15331 18460 15371 18500
rect 15907 18460 15947 18500
rect 21907 18460 21947 18500
rect 24748 18460 24788 18500
rect 27244 18460 27284 18500
rect 6211 18376 6251 18416
rect 7948 18376 7988 18416
rect 9100 18376 9140 18416
rect 10435 18376 10475 18416
rect 20428 18376 20468 18416
rect 20812 18376 20852 18416
rect 28204 18376 28244 18416
rect 28684 18376 28724 18416
rect 5212 18292 5252 18332
rect 6979 18292 7019 18332
rect 9964 18292 10004 18332
rect 11020 18292 11060 18332
rect 11980 18292 12020 18332
rect 12988 18292 13028 18332
rect 14563 18292 14603 18332
rect 16876 18292 16916 18332
rect 21292 18292 21332 18332
rect 27628 18292 27668 18332
rect 28924 18292 28964 18332
rect 3112 18124 3480 18164
rect 10886 18124 11254 18164
rect 18660 18124 19028 18164
rect 26434 18124 26802 18164
rect 739 17956 779 17996
rect 1996 17956 2036 17996
rect 3331 17956 3371 17996
rect 3811 17956 3851 17996
rect 5443 17956 5483 17996
rect 11587 17956 11627 17996
rect 15916 17956 15956 17996
rect 23587 17956 23627 17996
rect 1708 17872 1748 17912
rect 5068 17872 5108 17912
rect 6412 17872 6452 17912
rect 7020 17863 7060 17903
rect 9676 17872 9716 17912
rect 17932 17872 17972 17912
rect 21196 17872 21236 17912
rect 24268 17872 24308 17912
rect 25132 17872 25172 17912
rect 26860 17872 26900 17912
rect 27628 17872 27668 17912
rect 28012 17872 28052 17912
rect 1228 17788 1268 17828
rect 1804 17788 1844 17828
rect 2595 17788 2635 17828
rect 3075 17788 3115 17828
rect 940 17704 980 17744
rect 1036 17704 1076 17744
rect 1411 17704 1451 17744
rect 1996 17704 2036 17744
rect 2188 17704 2228 17744
rect 2476 17704 2516 17744
rect 2713 17704 2753 17744
rect 4972 17746 5012 17786
rect 5164 17788 5204 17828
rect 6508 17788 6548 17828
rect 12291 17788 12331 17828
rect 13155 17788 13195 17828
rect 13507 17788 13547 17828
rect 14668 17788 14708 17828
rect 18892 17788 18932 17828
rect 20812 17788 20852 17828
rect 22243 17788 22283 17828
rect 23788 17788 23828 17828
rect 24364 17788 24404 17828
rect 2956 17704 2996 17744
rect 3193 17704 3233 17744
rect 3628 17704 3668 17744
rect 4108 17704 4148 17744
rect 4723 17704 4763 17744
rect 4845 17704 4885 17744
rect 5299 17704 5339 17744
rect 5443 17704 5483 17744
rect 5548 17715 5588 17755
rect 5835 17704 5875 17744
rect 5971 17704 6011 17744
rect 6189 17704 6229 17744
rect 6351 17704 6391 17744
rect 6643 17704 6683 17744
rect 6979 17704 7019 17744
rect 7300 17704 7340 17744
rect 7459 17704 7499 17744
rect 7576 17704 7616 17744
rect 7715 17704 7755 17744
rect 7843 17704 7883 17744
rect 8224 17704 8264 17744
rect 9016 17704 9056 17744
rect 9196 17704 9236 17744
rect 9571 17704 9611 17744
rect 9955 17704 9995 17744
rect 10252 17704 10292 17744
rect 10540 17704 10580 17744
rect 10732 17704 10772 17744
rect 11104 17704 11144 17744
rect 11788 17704 11828 17744
rect 11884 17704 11924 17744
rect 12172 17704 12212 17744
rect 12412 17704 12452 17744
rect 12556 17704 12596 17744
rect 12748 17704 12788 17744
rect 13036 17704 13076 17744
rect 13273 17704 13313 17744
rect 13381 17704 13421 17744
rect 13612 17704 13652 17744
rect 13891 17704 13931 17744
rect 13996 17715 14036 17755
rect 14149 17704 14189 17744
rect 14270 17704 14310 17744
rect 14452 17704 14492 17744
rect 14773 17704 14813 17744
rect 14899 17695 14939 17735
rect 15004 17704 15044 17744
rect 15364 17704 15404 17744
rect 15523 17704 15563 17744
rect 15640 17704 15680 17744
rect 15811 17704 15851 17744
rect 15933 17704 15973 17744
rect 16103 17704 16143 17744
rect 16291 17704 16331 17744
rect 16588 17704 16628 17744
rect 16771 17704 16811 17744
rect 17272 17704 17312 17744
rect 17410 17704 17450 17744
rect 17933 17704 17973 17744
rect 18124 17704 18164 17744
rect 18403 17704 18443 17744
rect 18508 17704 18548 17744
rect 18988 17704 19028 17744
rect 19468 17704 19508 17744
rect 19987 17704 20027 17744
rect 20332 17704 20372 17744
rect 21580 17695 21620 17735
rect 21868 17704 21908 17744
rect 22103 17704 22143 17744
rect 22348 17704 22388 17744
rect 23224 17704 23264 17744
rect 23399 17704 23439 17744
rect 23587 17704 23627 17744
rect 23971 17704 24011 17744
rect 24739 17704 24779 17744
rect 25720 17704 25760 17744
rect 25996 17704 26036 17744
rect 26668 17704 26708 17744
rect 27244 17704 27284 17744
rect 27436 17704 27476 17744
rect 737 17620 777 17660
rect 3329 17620 3369 17660
rect 3809 17620 3849 17660
rect 5731 17653 5771 17693
rect 6796 17620 6836 17660
rect 11582 17620 11622 17660
rect 13699 17620 13739 17660
rect 16684 17620 16724 17660
rect 17596 17620 17636 17660
rect 20476 17620 20516 17660
rect 21484 17620 21524 17660
rect 2380 17536 2420 17576
rect 2860 17536 2900 17576
rect 3532 17536 3572 17576
rect 4012 17536 4052 17576
rect 4531 17536 4571 17576
rect 7363 17536 7403 17576
rect 8380 17536 8420 17576
rect 8851 17536 8891 17576
rect 10156 17536 10196 17576
rect 10636 17536 10676 17576
rect 11260 17536 11300 17576
rect 12076 17536 12116 17576
rect 12556 17536 12596 17576
rect 12940 17536 12980 17576
rect 14275 17536 14315 17576
rect 16204 17536 16244 17576
rect 17107 17536 17147 17576
rect 20140 17536 20180 17576
rect 20572 17536 20612 17576
rect 22435 17536 22475 17576
rect 23059 17536 23099 17576
rect 24940 17536 24980 17576
rect 25555 17536 25595 17576
rect 27340 17536 27380 17576
rect 4352 17368 4720 17408
rect 12126 17368 12494 17408
rect 19900 17368 20268 17408
rect 27674 17368 28042 17408
rect 1612 17200 1652 17240
rect 3148 17200 3188 17240
rect 3532 17200 3572 17240
rect 4876 17200 4916 17240
rect 6307 17200 6347 17240
rect 10924 17200 10964 17240
rect 929 17116 969 17156
rect 1722 17116 1762 17156
rect 1900 17116 1940 17156
rect 4204 17116 4244 17156
rect 5368 17158 5408 17198
rect 11683 17200 11723 17240
rect 11971 17200 12011 17240
rect 12835 17200 12875 17240
rect 14083 17200 14123 17240
rect 15427 17200 15467 17240
rect 17068 17200 17108 17240
rect 18316 17200 18356 17240
rect 8044 17116 8084 17156
rect 12259 17107 12299 17147
rect 13047 17116 13087 17156
rect 17491 17116 17531 17156
rect 21004 17116 21044 17156
rect 1132 17032 1172 17072
rect 1228 17023 1268 17063
rect 1411 17032 1451 17072
rect 1516 17032 1556 17072
rect 1996 17032 2036 17072
rect 2131 17023 2171 17063
rect 2236 17032 2276 17072
rect 2347 17032 2387 17072
rect 2572 17032 2612 17072
rect 3052 17032 3092 17072
rect 3235 17032 3275 17072
rect 3436 17032 3476 17072
rect 3628 17032 3668 17072
rect 3916 17032 3956 17072
rect 4103 17032 4143 17072
rect 4291 17032 4331 17072
rect 4775 17032 4815 17072
rect 4963 17032 5003 17072
rect 5116 17032 5156 17072
rect 5707 17032 5747 17072
rect 6147 17032 6187 17072
rect 2453 16948 2493 16988
rect 2668 16948 2708 16988
rect 5288 16990 5328 17030
rect 5587 16990 5627 17030
rect 5462 16948 5502 16988
rect 6019 16990 6059 17030
rect 6460 17032 6500 17072
rect 6604 17032 6644 17072
rect 7180 17032 7220 17072
rect 7315 17023 7355 17063
rect 5836 16948 5876 16988
rect 7084 16948 7124 16988
rect 7420 16990 7460 17030
rect 7852 17032 7892 17072
rect 8179 17032 8219 17072
rect 8380 17032 8420 17072
rect 8695 17032 8735 17072
rect 8845 17032 8885 17072
rect 8971 17032 9011 17072
rect 9257 17032 9297 17072
rect 9427 17032 9467 17072
rect 9672 17032 9712 17072
rect 9868 17032 9908 17072
rect 10648 17032 10688 17072
rect 11020 17032 11060 17072
rect 11257 17032 11297 17072
rect 11371 17032 11411 17072
rect 11596 17032 11636 17072
rect 11971 17032 12011 17072
rect 12076 17023 12116 17063
rect 12355 17032 12395 17072
rect 12532 17021 12572 17061
rect 12739 17032 12779 17072
rect 13324 17032 13364 17072
rect 13651 17065 13691 17105
rect 13996 17032 14036 17072
rect 14755 17074 14795 17114
rect 21964 17116 22004 17156
rect 28099 17116 28139 17156
rect 14284 17032 14324 17072
rect 14467 17032 14507 17072
rect 14881 17032 14921 17072
rect 15187 17032 15227 17072
rect 15356 17021 15396 17061
rect 15537 17032 15577 17072
rect 15667 17032 15707 17072
rect 15811 17032 15851 17072
rect 15916 17021 15956 17061
rect 16438 17032 16478 17072
rect 16588 17032 16628 17072
rect 16780 17032 16820 17072
rect 16973 17032 17013 17072
rect 17157 17032 17197 17072
rect 17686 17032 17726 17072
rect 17932 17032 17972 17072
rect 18124 17032 18164 17072
rect 18499 17032 18539 17072
rect 18988 17023 19028 17063
rect 19468 17032 19508 17072
rect 19948 17032 19988 17072
rect 20066 17032 20106 17072
rect 20620 17032 20660 17072
rect 20899 17032 20939 17072
rect 22093 17032 22133 17072
rect 22348 17032 22388 17072
rect 23020 17032 23060 17072
rect 23130 17065 23170 17105
rect 23404 17032 23444 17072
rect 23971 17032 24011 17072
rect 24460 17023 24500 17063
rect 24940 17032 24980 17072
rect 25420 17032 25460 17072
rect 25521 17032 25561 17072
rect 27715 17032 27755 17072
rect 8524 16948 8564 16988
rect 9100 16948 9140 16988
rect 10483 16948 10523 16988
rect 11155 16939 11195 16979
rect 11491 16948 11531 16988
rect 13420 16948 13460 16988
rect 15052 16948 15092 16988
rect 16243 16948 16283 16988
rect 19564 16948 19604 16988
rect 25036 16948 25076 16988
rect 931 16780 971 16820
rect 3772 16780 3812 16820
rect 5932 16822 5972 16862
rect 8620 16864 8660 16904
rect 9196 16864 9236 16904
rect 9868 16864 9908 16904
rect 14956 16864 14996 16904
rect 16588 16864 16628 16904
rect 21292 16864 21332 16904
rect 22732 16864 22772 16904
rect 13036 16780 13076 16820
rect 13804 16780 13844 16820
rect 14467 16780 14507 16820
rect 17932 16780 17972 16820
rect 21676 16780 21716 16820
rect 23740 16780 23780 16820
rect 25804 16780 25844 16820
rect 26188 16780 26228 16820
rect 3112 16612 3480 16652
rect 10886 16612 11254 16652
rect 18660 16612 19028 16652
rect 26434 16612 26802 16652
rect 2563 16444 2603 16484
rect 10819 16444 10859 16484
rect 15436 16444 15476 16484
rect 15619 16444 15659 16484
rect 21580 16444 21620 16484
rect 22444 16444 22484 16484
rect 23884 16444 23924 16484
rect 5644 16360 5684 16400
rect 6796 16360 6836 16400
rect 8135 16360 8175 16400
rect 8803 16360 8843 16400
rect 10604 16351 10644 16391
rect 11212 16360 11252 16400
rect 13036 16360 13076 16400
rect 17356 16360 17396 16400
rect 20428 16360 20468 16400
rect 21763 16360 21803 16400
rect 24268 16360 24308 16400
rect 29068 16360 29108 16400
rect 796 16234 836 16274
rect 1132 16276 1172 16316
rect 1315 16276 1355 16316
rect 1891 16276 1931 16316
rect 3619 16276 3659 16316
rect 3820 16276 3860 16316
rect 4707 16276 4747 16316
rect 4972 16276 5012 16316
rect 5187 16276 5227 16316
rect 5740 16276 5780 16316
rect 6339 16276 6379 16316
rect 6892 16276 6932 16316
rect 8236 16276 8276 16316
rect 931 16192 971 16232
rect 1036 16192 1076 16232
rect 1699 16192 1739 16232
rect 2081 16192 2121 16232
rect 2378 16192 2418 16232
rect 2860 16192 2900 16232
rect 3352 16192 3392 16232
rect 3484 16192 3524 16232
rect 3724 16192 3764 16232
rect 4108 16192 4148 16232
rect 4227 16192 4267 16232
rect 4345 16192 4385 16232
rect 4588 16192 4628 16232
rect 4825 16192 4865 16232
rect 5077 16192 5117 16232
rect 5299 16192 5339 16232
rect 5583 16192 5623 16232
rect 5875 16192 5915 16232
rect 6220 16192 6260 16232
rect 6457 16192 6497 16232
rect 7027 16234 7067 16274
rect 9004 16276 9044 16316
rect 10291 16267 10331 16307
rect 11308 16276 11348 16316
rect 11884 16276 11924 16316
rect 6735 16192 6775 16232
rect 7204 16192 7244 16232
rect 7363 16192 7403 16232
rect 7480 16192 7520 16232
rect 7612 16192 7652 16232
rect 7754 16192 7794 16232
rect 7917 16192 7957 16232
rect 8079 16192 8119 16232
rect 8371 16192 8411 16232
rect 8620 16192 8660 16232
rect 8803 16192 8843 16232
rect 9331 16192 9371 16232
rect 10156 16192 10196 16232
rect 10393 16192 10433 16232
rect 10627 16192 10667 16232
rect 10972 16192 11012 16232
rect 11443 16234 11483 16274
rect 12595 16267 12635 16307
rect 12940 16276 12980 16316
rect 17260 16276 17300 16316
rect 11151 16192 11191 16232
rect 11548 16192 11588 16232
rect 11727 16192 11767 16232
rect 12005 16192 12045 16232
rect 12460 16192 12500 16232
rect 13123 16234 13163 16274
rect 17827 16276 17867 16316
rect 18028 16276 18068 16316
rect 19372 16276 19412 16316
rect 12700 16192 12740 16232
rect 12811 16192 12851 16232
rect 13269 16192 13309 16232
rect 13411 16165 13451 16205
rect 13615 16192 13655 16232
rect 13795 16192 13835 16232
rect 13900 16203 13940 16243
rect 14045 16192 14085 16232
rect 14179 16192 14219 16232
rect 14356 16192 14396 16232
rect 14884 16192 14924 16232
rect 15043 16192 15083 16232
rect 15160 16192 15200 16232
rect 15292 16203 15332 16243
rect 15427 16192 15467 16232
rect 15631 16192 15671 16232
rect 15737 16192 15777 16232
rect 15903 16192 15943 16232
rect 16011 16192 16051 16232
rect 16137 16192 16177 16232
rect 16387 16192 16427 16232
rect 16505 16192 16545 16232
rect 16665 16192 16705 16232
rect 16771 16192 16811 16232
rect 16905 16192 16945 16232
rect 17116 16192 17156 16232
rect 17431 16192 17471 16232
rect 17587 16192 17627 16232
rect 17692 16192 17732 16232
rect 19027 16234 19067 16274
rect 26860 16276 26900 16316
rect 17932 16192 17972 16232
rect 18520 16192 18560 16232
rect 19564 16192 19604 16232
rect 19843 16183 19883 16223
rect 20140 16192 20180 16232
rect 20908 16192 20948 16232
rect 21187 16192 21227 16232
rect 21964 16192 22004 16232
rect 22085 16192 22125 16232
rect 22487 16192 22527 16232
rect 22627 16183 22667 16223
rect 22732 16192 22772 16232
rect 23212 16192 23252 16232
rect 23491 16192 23531 16232
rect 24119 16192 24159 16232
rect 24259 16183 24299 16223
rect 24364 16192 24404 16232
rect 24556 16192 24596 16232
rect 26092 16192 26132 16232
rect 26371 16192 26411 16232
rect 26476 16192 26516 16232
rect 26956 16192 26996 16232
rect 27436 16192 27476 16232
rect 27955 16192 27995 16232
rect 28300 16192 28340 16232
rect 28492 16192 28532 16232
rect 28684 16234 28724 16274
rect 28876 16192 28916 16232
rect 2561 16108 2601 16148
rect 4492 16108 4532 16148
rect 6124 16108 6164 16148
rect 9532 16108 9572 16148
rect 1411 16024 1451 16064
rect 2179 16024 2219 16064
rect 2284 16024 2324 16064
rect 2764 16024 2804 16064
rect 3187 16024 3227 16064
rect 4012 16024 4052 16064
rect 7267 16024 7307 16064
rect 9244 16024 9284 16064
rect 5539 15982 5579 16022
rect 6691 15982 6731 16022
rect 10060 16024 10100 16064
rect 11800 16066 11840 16106
rect 19132 16108 19172 16148
rect 19948 16108 19988 16148
rect 21292 16108 21332 16148
rect 23596 16108 23636 16148
rect 25228 16108 25268 16148
rect 12364 16024 12404 16064
rect 13603 16024 13643 16064
rect 14275 16024 14315 16064
rect 16867 16024 16907 16064
rect 18355 16024 18395 16064
rect 18835 16024 18875 16064
rect 19708 16024 19748 16064
rect 22060 16024 22100 16064
rect 25420 16024 25460 16064
rect 28108 16024 28148 16064
rect 28396 16024 28436 16064
rect 28780 16024 28820 16064
rect 4352 15856 4720 15896
rect 12126 15856 12494 15896
rect 19900 15856 20268 15896
rect 27674 15856 28042 15896
rect 1507 15688 1547 15728
rect 1612 15688 1652 15728
rect 1987 15688 2027 15728
rect 2956 15688 2996 15728
rect 3436 15688 3476 15728
rect 4003 15688 4043 15728
rect 4483 15688 4523 15728
rect 4876 15688 4916 15728
rect 5740 15688 5780 15728
rect 6307 15688 6347 15728
rect 7756 15688 7796 15728
rect 8140 15688 8180 15728
rect 10732 15688 10772 15728
rect 12028 15688 12068 15728
rect 13804 15688 13844 15728
rect 14860 15688 14900 15728
rect 16012 15688 16052 15728
rect 16867 15688 16907 15728
rect 17827 15688 17867 15728
rect 17932 15688 17972 15728
rect 21772 15688 21812 15728
rect 22339 15688 22379 15728
rect 23788 15688 23828 15728
rect 24940 15688 24980 15728
rect 25219 15688 25259 15728
rect 25900 15688 25940 15728
rect 28972 15688 29012 15728
rect 3233 15604 3273 15644
rect 3715 15604 3755 15644
rect 7180 15604 7220 15644
rect 8995 15604 9035 15644
rect 10819 15595 10859 15635
rect 12353 15604 12393 15644
rect 15628 15604 15668 15644
rect 931 15520 971 15560
rect 1228 15520 1268 15560
rect 1409 15520 1449 15560
rect 1708 15511 1748 15551
rect 1900 15520 1940 15560
rect 2188 15520 2228 15560
rect 2327 15520 2367 15560
rect 2467 15520 2507 15560
rect 2572 15520 2612 15560
rect 2860 15520 2900 15560
rect 3052 15520 3092 15560
rect 3532 15511 3572 15551
rect 3916 15520 3956 15560
rect 4151 15520 4191 15560
rect 4396 15520 4436 15560
rect 4972 15520 5012 15560
rect 5203 15520 5243 15560
rect 5356 15520 5396 15560
rect 5548 15520 5588 15560
rect 5836 15520 5876 15560
rect 6067 15520 6107 15560
rect 6211 15520 6251 15560
rect 6519 15520 6559 15560
rect 6796 15520 6836 15560
rect 6979 15520 7019 15560
rect 7276 15520 7316 15560
rect 7493 15520 7533 15560
rect 7660 15520 7700 15560
rect 7843 15520 7883 15560
rect 8044 15520 8084 15560
rect 2668 15436 2708 15476
rect 4291 15436 4331 15476
rect 5091 15436 5131 15476
rect 5955 15436 5995 15476
rect 7395 15436 7435 15476
rect 8236 15478 8276 15518
rect 8428 15520 8468 15560
rect 8683 15520 8723 15560
rect 8908 15520 8948 15560
rect 9283 15520 9323 15560
rect 9571 15520 9611 15560
rect 10060 15520 10100 15560
rect 10277 15520 10317 15560
rect 10523 15520 10563 15560
rect 10687 15520 10727 15560
rect 10911 15520 10951 15560
rect 11092 15520 11132 15560
rect 11452 15520 11492 15560
rect 11907 15520 11947 15560
rect 8803 15436 8843 15476
rect 9187 15436 9227 15476
rect 9724 15436 9764 15476
rect 9964 15436 10004 15476
rect 10179 15436 10219 15476
rect 11779 15478 11819 15518
rect 12172 15520 12212 15560
rect 13219 15562 13259 15602
rect 17249 15604 17289 15644
rect 17726 15604 17766 15644
rect 21004 15604 21044 15644
rect 21114 15604 21154 15644
rect 22842 15604 22882 15644
rect 23203 15604 23243 15644
rect 12556 15520 12596 15560
rect 12652 15511 12692 15551
rect 13420 15520 13460 15560
rect 12796 15478 12836 15518
rect 11596 15436 11636 15476
rect 13123 15478 13163 15518
rect 13612 15520 13652 15560
rect 13900 15520 13940 15560
rect 14137 15520 14177 15560
rect 14253 15520 14293 15560
rect 14401 15520 14441 15560
rect 14693 15520 14733 15560
rect 15043 15520 15083 15560
rect 15532 15520 15572 15560
rect 15724 15520 15764 15560
rect 15916 15520 15956 15560
rect 16108 15520 16148 15560
rect 16675 15520 16715 15560
rect 17452 15520 17492 15560
rect 17548 15511 17588 15551
rect 18028 15511 18068 15551
rect 18223 15520 18263 15560
rect 18345 15520 18385 15560
rect 18508 15520 18548 15560
rect 18743 15520 18783 15560
rect 18988 15520 19028 15560
rect 19243 15520 19283 15560
rect 19468 15520 19508 15560
rect 19708 15520 19748 15560
rect 19887 15520 19927 15560
rect 20428 15520 20468 15560
rect 12938 15436 12978 15476
rect 14019 15436 14059 15476
rect 14572 15436 14612 15476
rect 15091 15408 15131 15448
rect 18883 15436 18923 15476
rect 19084 15436 19124 15476
rect 19363 15436 19403 15476
rect 19564 15436 19604 15476
rect 20179 15478 20219 15518
rect 20668 15520 20708 15560
rect 20803 15520 20843 15560
rect 20908 15520 20948 15560
rect 21484 15520 21524 15560
rect 21823 15520 21863 15560
rect 22027 15520 22067 15560
rect 22252 15520 22292 15560
rect 22531 15520 22571 15560
rect 22636 15520 22676 15560
rect 23301 15531 23341 15571
rect 23500 15520 23540 15560
rect 23831 15520 23871 15560
rect 23971 15511 24011 15551
rect 24076 15520 24116 15560
rect 24547 15520 24587 15560
rect 24652 15520 24692 15560
rect 25420 15520 25460 15560
rect 25708 15520 25748 15560
rect 27811 15520 27851 15560
rect 28195 15520 28235 15560
rect 28387 15511 28427 15551
rect 28876 15520 28916 15560
rect 29068 15520 29108 15560
rect 29260 15520 29300 15560
rect 20044 15436 20084 15476
rect 20332 15436 20372 15476
rect 20547 15436 20587 15476
rect 21706 15436 21746 15476
rect 22147 15436 22187 15476
rect 26275 15436 26315 15476
rect 28540 15436 28580 15476
rect 1228 15352 1268 15392
rect 11692 15352 11732 15392
rect 13036 15352 13076 15392
rect 13516 15352 13556 15392
rect 14476 15352 14516 15392
rect 16647 15352 16687 15392
rect 19948 15352 19988 15392
rect 21580 15352 21620 15392
rect 3235 15268 3275 15308
rect 5452 15268 5492 15308
rect 6508 15268 6548 15308
rect 6979 15268 7019 15308
rect 8572 15268 8612 15308
rect 10531 15268 10571 15308
rect 12355 15268 12395 15308
rect 17251 15268 17291 15308
rect 18220 15268 18260 15308
rect 22828 15268 22868 15308
rect 23980 15268 24020 15308
rect 3112 15100 3480 15140
rect 10886 15100 11254 15140
rect 18660 15100 19028 15140
rect 26434 15100 26802 15140
rect 4675 14932 4715 14972
rect 5068 14932 5108 14972
rect 9964 14932 10004 14972
rect 12844 14932 12884 14972
rect 13612 14932 13652 14972
rect 14956 14932 14996 14972
rect 17443 14932 17483 14972
rect 17932 14932 17972 14972
rect 18604 14932 18644 14972
rect 19084 14932 19124 14972
rect 20524 14932 20564 14972
rect 21964 14932 22004 14972
rect 23500 14932 23540 14972
rect 28012 14932 28052 14972
rect 28972 14932 29012 14972
rect 3148 14848 3188 14888
rect 4003 14848 4043 14888
rect 8947 14848 8987 14888
rect 11020 14848 11060 14888
rect 15427 14848 15467 14888
rect 19468 14848 19508 14888
rect 20812 14848 20852 14888
rect 23980 14848 24020 14888
rect 26956 14848 26996 14888
rect 29836 14848 29876 14888
rect 1027 14764 1067 14804
rect 2947 14764 2987 14804
rect 5980 14764 6020 14804
rect 6403 14764 6443 14804
rect 6604 14764 6644 14804
rect 7651 14764 7691 14804
rect 7852 14764 7892 14804
rect 9571 14764 9611 14804
rect 9772 14764 9812 14804
rect 10563 14764 10603 14804
rect 2563 14680 2603 14720
rect 3148 14680 3188 14720
rect 3273 14680 3313 14720
rect 3436 14680 3476 14720
rect 3820 14680 3860 14720
rect 4003 14680 4043 14720
rect 4481 14680 4521 14720
rect 4588 14680 4628 14720
rect 4972 14680 5012 14720
rect 5164 14680 5204 14720
rect 5303 14680 5343 14720
rect 5443 14680 5483 14720
rect 5548 14680 5588 14720
rect 5824 14680 5864 14720
rect 6263 14680 6303 14720
rect 6508 14680 6548 14720
rect 6973 14680 7013 14720
rect 7084 14680 7124 14720
rect 7511 14680 7551 14720
rect 7756 14680 7796 14720
rect 8032 14680 8072 14720
rect 8854 14680 8894 14720
rect 9148 14713 9188 14753
rect 9244 14680 9284 14720
rect 9448 14680 9488 14720
rect 9676 14680 9716 14720
rect 9964 14680 10004 14720
rect 10156 14680 10196 14720
rect 10444 14680 10484 14720
rect 10952 14722 10992 14762
rect 11116 14764 11156 14804
rect 11788 14764 11828 14804
rect 12652 14764 12692 14804
rect 14563 14764 14603 14804
rect 22371 14764 22411 14804
rect 10661 14680 10701 14720
rect 10797 14680 10837 14720
rect 11452 14680 11492 14720
rect 11251 14638 11291 14678
rect 11587 14680 11627 14720
rect 11692 14680 11732 14720
rect 11980 14680 12020 14720
rect 12172 14680 12212 14720
rect 12887 14680 12927 14720
rect 13027 14671 13067 14711
rect 13132 14680 13172 14720
rect 13315 14680 13355 14720
rect 13420 14680 13460 14720
rect 13900 14680 13940 14720
rect 14019 14680 14059 14720
rect 14137 14680 14177 14720
rect 14371 14671 14411 14711
rect 14668 14680 14708 14720
rect 14956 14680 14996 14720
rect 15148 14680 15188 14720
rect 15712 14713 15752 14753
rect 15811 14680 15851 14720
rect 16097 14680 16137 14720
rect 16396 14680 16436 14720
rect 16588 14680 16628 14720
rect 16780 14680 16820 14720
rect 17260 14680 17300 14720
rect 17443 14680 17483 14720
rect 17932 14680 17972 14720
rect 18124 14680 18164 14720
rect 18412 14680 18452 14720
rect 18647 14680 18687 14720
rect 18787 14713 18827 14753
rect 23020 14764 23060 14804
rect 23154 14764 23194 14804
rect 26572 14764 26612 14804
rect 18887 14680 18927 14720
rect 19084 14680 19124 14720
rect 19276 14680 19316 14720
rect 20227 14680 20267 14720
rect 20535 14680 20575 14720
rect 20716 14680 20756 14720
rect 20851 14680 20891 14720
rect 20965 14680 21005 14720
rect 21340 14713 21380 14753
rect 21436 14680 21476 14720
rect 21676 14680 21716 14720
rect 21816 14680 21856 14720
rect 21925 14680 21965 14720
rect 22252 14680 22292 14720
rect 22469 14680 22509 14720
rect 22675 14680 22715 14720
rect 22924 14680 22964 14720
rect 23263 14680 23303 14720
rect 23543 14713 23583 14753
rect 23683 14671 23723 14711
rect 23788 14680 23828 14720
rect 24141 14680 24181 14720
rect 24257 14680 24297 14720
rect 24369 14680 24409 14720
rect 25027 14680 25067 14720
rect 27340 14680 27380 14720
rect 28147 14680 28187 14720
rect 29644 14680 29684 14720
rect 5635 14596 5675 14636
rect 12076 14596 12116 14636
rect 13623 14596 13663 14636
rect 20332 14596 20372 14636
rect 24643 14596 24683 14636
rect 28348 14596 28388 14636
rect 652 14512 692 14552
rect 6787 14512 6827 14552
rect 8188 14512 8228 14552
rect 8659 14512 8699 14552
rect 10348 14512 10388 14552
rect 12412 14512 12452 14552
rect 13804 14512 13844 14552
rect 15955 14512 15995 14552
rect 16195 14512 16235 14552
rect 16300 14512 16340 14552
rect 16684 14512 16724 14552
rect 18268 14512 18308 14552
rect 19852 14512 19892 14552
rect 21187 14512 21227 14552
rect 22156 14512 22196 14552
rect 22780 14512 22820 14552
rect 23020 14512 23060 14552
rect 4352 14344 4720 14384
rect 12126 14344 12494 14384
rect 19900 14344 20268 14384
rect 27674 14344 28042 14384
rect 739 14176 779 14216
rect 1228 14176 1268 14216
rect 3052 14176 3092 14216
rect 3724 14176 3764 14216
rect 4195 14176 4235 14216
rect 4972 14176 5012 14216
rect 5827 14176 5867 14216
rect 6124 14176 6164 14216
rect 7180 14176 7220 14216
rect 7372 14176 7412 14216
rect 8035 14176 8075 14216
rect 9331 14176 9371 14216
rect 9763 14176 9803 14216
rect 10540 14176 10580 14216
rect 12595 14176 12635 14216
rect 13987 14176 14027 14216
rect 15235 14176 15275 14216
rect 16003 14176 16043 14216
rect 16579 14176 16619 14216
rect 18892 14176 18932 14216
rect 19372 14176 19412 14216
rect 21955 14176 21995 14216
rect 22252 14176 22292 14216
rect 24163 14176 24203 14216
rect 24748 14176 24788 14216
rect 29452 14176 29492 14216
rect 5059 14083 5099 14123
rect 10263 14092 10303 14132
rect 12508 14092 12548 14132
rect 15902 14092 15942 14132
rect 19948 14092 19988 14132
rect 21379 14092 21419 14132
rect 22540 14092 22580 14132
rect 24643 14092 24683 14132
rect 844 14008 884 14048
rect 1900 14008 1940 14048
rect 2753 14008 2793 14048
rect 2860 14008 2900 14048
rect 3244 14008 3284 14048
rect 3532 14008 3572 14048
rect 4028 13997 4068 14037
rect 4227 14008 4267 14048
rect 4339 14008 4379 14048
rect 4483 14008 4523 14048
rect 4605 14008 4645 14048
rect 4771 14008 4811 14048
rect 4876 13999 4916 14039
rect 5155 14008 5195 14048
rect 5332 14008 5372 14048
rect 5495 14008 5535 14048
rect 5740 14008 5780 14048
rect 6028 14008 6068 14048
rect 6220 14008 6260 14048
rect 6379 14008 6419 14048
rect 6499 14008 6539 14048
rect 6604 14008 6644 14048
rect 6892 14008 6932 14048
rect 7141 14008 7181 14048
rect 5635 13924 5675 13964
rect 7014 13966 7054 14006
rect 7533 13999 7573 14039
rect 7651 13999 7691 14039
rect 7760 14008 7800 14048
rect 8188 14008 8228 14048
rect 8332 14008 8372 14048
rect 9088 13999 9128 14039
rect 9187 14008 9227 14048
rect 9431 14008 9471 14048
rect 9676 14008 9716 14048
rect 9955 14008 9995 14048
rect 10060 14008 10100 14048
rect 10444 14008 10484 14048
rect 10634 14008 10674 14048
rect 10819 13999 10859 14039
rect 10972 14008 11012 14048
rect 11404 14008 11444 14048
rect 11519 14008 11559 14048
rect 11692 14008 11732 14048
rect 11884 14008 11924 14048
rect 12268 14008 12308 14048
rect 12739 14008 12779 14048
rect 12844 13999 12884 14039
rect 13324 14008 13364 14048
rect 13507 14008 13547 14048
rect 13893 14008 13933 14048
rect 13660 13966 13700 14006
rect 14179 13999 14219 14039
rect 14476 14008 14516 14048
rect 14903 14008 14943 14048
rect 15148 14008 15188 14048
rect 15532 14008 15572 14048
rect 15769 14008 15809 14048
rect 16108 14008 16148 14048
rect 16204 13999 16244 14039
rect 16876 14008 16916 14048
rect 17644 14008 17684 14048
rect 18268 14008 18308 14048
rect 18569 14008 18609 14048
rect 18739 14008 18779 14048
rect 18988 14008 19028 14048
rect 19225 14008 19265 14048
rect 19705 14008 19745 14048
rect 19852 14008 19892 14048
rect 6700 13924 6740 13964
rect 9571 13924 9611 13964
rect 13795 13924 13835 13964
rect 15043 13924 15083 13964
rect 15436 13924 15476 13964
rect 15651 13924 15691 13964
rect 16786 13924 16826 13964
rect 17554 13924 17594 13964
rect 18412 13924 18452 13964
rect 19107 13924 19147 13964
rect 19468 13966 19508 14006
rect 20140 14008 20180 14048
rect 20332 14008 20372 14048
rect 20515 14008 20555 14048
rect 20620 14008 20660 14048
rect 20812 14008 20852 14048
rect 21151 14008 21191 14048
rect 21433 13999 21473 14039
rect 21531 14008 21571 14048
rect 21667 13999 21707 14039
rect 21772 14008 21812 14048
rect 22060 14008 22100 14048
rect 22444 14008 22484 14048
rect 22636 14008 22676 14048
rect 22797 14008 22837 14048
rect 23404 14008 23444 14048
rect 22924 13966 22964 14006
rect 19587 13924 19627 13964
rect 23251 13966 23291 14006
rect 23743 14008 23783 14048
rect 24076 14008 24116 14048
rect 24364 14008 24404 14048
rect 24545 14008 24585 14048
rect 24844 13999 24884 14039
rect 25708 14008 25748 14048
rect 26572 14008 26612 14048
rect 26764 14008 26804 14048
rect 26956 14008 26996 14048
rect 27523 14008 27563 14048
rect 21043 13915 21083 13955
rect 23119 13924 23159 13964
rect 23635 13915 23675 13955
rect 27148 13924 27188 13964
rect 1036 13840 1076 13880
rect 2092 13840 2132 13880
rect 11404 13840 11444 13880
rect 13132 13840 13172 13880
rect 13507 13840 13547 13880
rect 14476 13840 14516 13880
rect 18508 13840 18548 13880
rect 21196 13840 21236 13880
rect 23020 13840 23060 13880
rect 23788 13840 23828 13880
rect 26764 13840 26804 13880
rect 29644 13840 29684 13880
rect 8140 13756 8180 13796
rect 8803 13756 8843 13796
rect 10252 13756 10292 13796
rect 12508 13756 12548 13796
rect 14275 13756 14315 13796
rect 17452 13756 17492 13796
rect 20620 13756 20660 13796
rect 20908 13756 20948 13796
rect 23500 13756 23540 13796
rect 25036 13756 25076 13796
rect 25900 13756 25940 13796
rect 29068 13756 29108 13796
rect 3112 13588 3480 13628
rect 10886 13588 11254 13628
rect 18660 13588 19028 13628
rect 26434 13588 26802 13628
rect 2563 13420 2603 13460
rect 3820 13420 3860 13460
rect 9139 13420 9179 13460
rect 12355 13420 12395 13460
rect 15724 13420 15764 13460
rect 18403 13420 18443 13460
rect 19084 13420 19124 13460
rect 19468 13420 19508 13460
rect 20236 13420 20276 13460
rect 20899 13420 20939 13460
rect 21763 13420 21803 13460
rect 22828 13420 22868 13460
rect 23404 13420 23444 13460
rect 24028 13420 24068 13460
rect 24652 13420 24692 13460
rect 28780 13420 28820 13460
rect 4771 13336 4811 13376
rect 9379 13336 9419 13376
rect 18124 13336 18164 13376
rect 19852 13336 19892 13376
rect 21196 13336 21236 13376
rect 22348 13336 22388 13376
rect 5347 13252 5387 13292
rect 5548 13252 5588 13292
rect 5827 13252 5867 13292
rect 6307 13252 6347 13292
rect 6508 13252 6548 13292
rect 940 13168 980 13208
rect 2275 13168 2315 13208
rect 2380 13168 2420 13208
rect 2947 13168 2987 13208
rect 3244 13168 3284 13208
rect 3523 13168 3563 13208
rect 3628 13168 3668 13208
rect 4483 13168 4523 13208
rect 4588 13168 4628 13208
rect 5227 13168 5267 13208
rect 5452 13168 5492 13208
rect 5692 13210 5732 13250
rect 7852 13252 7892 13292
rect 10258 13252 10298 13292
rect 10915 13252 10955 13292
rect 13084 13252 13124 13292
rect 13635 13252 13675 13292
rect 17187 13252 17227 13292
rect 25987 13252 26027 13292
rect 5930 13168 5970 13208
rect 6167 13168 6207 13208
rect 6412 13168 6452 13208
rect 6691 13168 6731 13208
rect 6796 13168 6836 13208
rect 7342 13168 7382 13208
rect 7459 13140 7499 13180
rect 7948 13168 7988 13208
rect 8428 13168 8468 13208
rect 8916 13168 8956 13208
rect 9664 13201 9704 13241
rect 9763 13168 9803 13208
rect 10351 13168 10391 13208
rect 10775 13168 10815 13208
rect 11020 13168 11060 13208
rect 11704 13168 11744 13208
rect 12214 13168 12254 13208
rect 12652 13168 12692 13208
rect 12928 13168 12968 13208
rect 13516 13168 13556 13208
rect 13753 13168 13793 13208
rect 14188 13168 14228 13208
rect 14307 13168 14347 13208
rect 14425 13168 14465 13208
rect 14711 13168 14751 13208
rect 14851 13168 14891 13208
rect 14956 13168 14996 13208
rect 15235 13168 15275 13208
rect 15546 13168 15586 13208
rect 16108 13159 16148 13199
rect 16396 13168 16436 13208
rect 17068 13168 17108 13208
rect 17305 13168 17345 13208
rect 17740 13168 17780 13208
rect 17851 13201 17891 13241
rect 17954 13210 17994 13250
rect 18796 13168 18836 13208
rect 19084 13168 19124 13208
rect 19276 13168 19316 13208
rect 19468 13168 19508 13208
rect 19660 13168 19700 13208
rect 19852 13168 19892 13208
rect 20044 13168 20084 13208
rect 20236 13168 20276 13208
rect 20524 13168 20564 13208
rect 20716 13168 20756 13208
rect 20907 13168 20947 13208
rect 21090 13201 21130 13241
rect 21272 13168 21312 13208
rect 21388 13168 21428 13208
rect 21575 13168 21615 13208
rect 21771 13168 21811 13208
rect 22003 13168 22043 13208
rect 22252 13168 22292 13208
rect 22387 13168 22427 13208
rect 22501 13168 22541 13208
rect 22732 13168 22772 13208
rect 22917 13165 22957 13205
rect 23107 13168 23147 13208
rect 23596 13168 23636 13208
rect 23740 13201 23780 13241
rect 24172 13168 24212 13208
rect 24364 13168 24404 13208
rect 24547 13168 24587 13208
rect 24652 13168 24692 13208
rect 25027 13168 25067 13208
rect 28627 13210 28667 13250
rect 25132 13168 25172 13208
rect 27523 13168 27563 13208
rect 28780 13168 28820 13208
rect 28972 13168 29012 13208
rect 3148 13084 3188 13124
rect 3831 13084 3871 13124
rect 7002 13084 7042 13124
rect 11107 13084 11147 13124
rect 11539 13084 11579 13124
rect 12353 13084 12393 13124
rect 13420 13084 13460 13124
rect 15043 13084 15083 13124
rect 16012 13084 16052 13124
rect 16972 13084 17012 13124
rect 23212 13084 23252 13124
rect 23418 13084 23458 13124
rect 23932 13084 23972 13124
rect 25603 13084 25643 13124
rect 27907 13084 27947 13124
rect 1612 13000 1652 13040
rect 6019 13000 6059 13040
rect 6892 13000 6932 13040
rect 10051 13000 10091 13040
rect 12019 13000 12059 13040
rect 12556 13000 12596 13040
rect 9907 12958 9947 12998
rect 14092 13000 14132 13040
rect 15331 13000 15371 13040
rect 15436 13000 15476 13040
rect 22108 13000 22148 13040
rect 25420 13000 25460 13040
rect 28435 13000 28475 13040
rect 4352 12832 4720 12872
rect 12126 12832 12494 12872
rect 19900 12832 20268 12872
rect 27674 12832 28042 12872
rect 835 12664 875 12704
rect 1804 12664 1844 12704
rect 2035 12664 2075 12704
rect 3043 12664 3083 12704
rect 3571 12664 3611 12704
rect 4588 12664 4628 12704
rect 6028 12664 6068 12704
rect 6307 12664 6347 12704
rect 6412 12664 6452 12704
rect 9283 12664 9323 12704
rect 9763 12664 9803 12704
rect 10867 12664 10907 12704
rect 11404 12664 11444 12704
rect 13420 12664 13460 12704
rect 15091 12664 15131 12704
rect 16012 12664 16052 12704
rect 16291 12664 16331 12704
rect 16876 12664 16916 12704
rect 17644 12664 17684 12704
rect 18211 12664 18251 12704
rect 19075 12664 19115 12704
rect 20611 12664 20651 12704
rect 21100 12664 21140 12704
rect 23788 12664 23828 12704
rect 24940 12664 24980 12704
rect 25507 12664 25547 12704
rect 26860 12664 26900 12704
rect 28204 12664 28244 12704
rect 6689 12580 6729 12620
rect 8332 12580 8372 12620
rect 8716 12580 8756 12620
rect 11201 12580 11241 12620
rect 11971 12580 12011 12620
rect 14179 12571 14219 12611
rect 16190 12580 16230 12620
rect 16396 12580 16436 12620
rect 17438 12580 17478 12620
rect 21475 12580 21515 12620
rect 26967 12580 27007 12620
rect 27614 12580 27654 12620
rect 940 12496 980 12536
rect 1324 12496 1364 12536
rect 1708 12496 1748 12536
rect 2179 12496 2219 12536
rect 2284 12487 2324 12527
rect 2731 12496 2771 12536
rect 2956 12496 2996 12536
rect 3766 12496 3806 12536
rect 4195 12496 4235 12536
rect 4300 12496 4340 12536
rect 4747 12496 4787 12536
rect 4972 12496 5012 12536
rect 5635 12496 5675 12536
rect 5740 12496 5780 12536
rect 6209 12496 6249 12536
rect 6508 12487 6548 12527
rect 6892 12496 6932 12536
rect 6988 12487 7028 12527
rect 7180 12496 7220 12536
rect 7375 12496 7415 12536
rect 7852 12496 7892 12536
rect 8042 12496 8082 12536
rect 8236 12496 8276 12536
rect 8428 12496 8468 12536
rect 8609 12496 8649 12536
rect 8812 12496 8852 12536
rect 9004 12496 9044 12536
rect 9444 12496 9484 12536
rect 9580 12496 9620 12536
rect 9916 12496 9956 12536
rect 10060 12496 10100 12536
rect 11062 12496 11102 12536
rect 11500 12487 11540 12527
rect 12172 12496 12212 12536
rect 12739 12496 12779 12536
rect 12846 12496 12886 12536
rect 13516 12496 13556 12536
rect 13753 12496 13793 12536
rect 13891 12496 13931 12536
rect 13996 12487 14036 12527
rect 14275 12496 14315 12536
rect 14452 12485 14492 12525
rect 15286 12496 15326 12536
rect 15619 12496 15659 12536
rect 15724 12496 15764 12536
rect 16492 12487 16532 12527
rect 16972 12496 17012 12536
rect 17209 12496 17249 12536
rect 17740 12487 17780 12527
rect 18508 12496 18548 12536
rect 19276 12496 19316 12536
rect 19564 12496 19604 12536
rect 19756 12496 19796 12536
rect 20140 12496 20180 12536
rect 20332 12496 20372 12536
rect 20716 12496 20756 12536
rect 21100 12496 21140 12536
rect 21292 12496 21332 12536
rect 21859 12496 21899 12536
rect 24652 12496 24692 12536
rect 24940 12496 24980 12536
rect 25130 12496 25170 12536
rect 25411 12496 25451 12536
rect 25719 12496 25759 12536
rect 25891 12487 25931 12527
rect 26044 12496 26084 12536
rect 26659 12496 26699 12536
rect 26764 12496 26804 12536
rect 27095 12496 27135 12536
rect 27340 12496 27380 12536
rect 27820 12496 27860 12536
rect 27916 12487 27956 12527
rect 28108 12496 28148 12536
rect 28281 12496 28321 12536
rect 2851 12412 2891 12452
rect 4867 12412 4907 12452
rect 5068 12412 5108 12452
rect 13651 12403 13691 12443
rect 17091 12412 17131 12452
rect 18418 12412 18458 12452
rect 23404 12412 23444 12452
rect 27221 12412 27261 12452
rect 27436 12412 27476 12452
rect 1132 12328 1172 12368
rect 2572 12328 2612 12368
rect 7276 12328 7316 12368
rect 21196 12328 21236 12368
rect 28492 12328 28532 12368
rect 28876 12328 28916 12368
rect 6691 12244 6731 12284
rect 7852 12244 7892 12284
rect 9148 12244 9188 12284
rect 11203 12244 11243 12284
rect 13027 12244 13067 12284
rect 13891 12244 13931 12284
rect 17443 12244 17483 12284
rect 19852 12244 19892 12284
rect 20140 12244 20180 12284
rect 20908 12244 20948 12284
rect 23980 12244 24020 12284
rect 25708 12244 25748 12284
rect 27619 12244 27659 12284
rect 3112 12076 3480 12116
rect 10886 12076 11254 12116
rect 18660 12076 19028 12116
rect 26434 12076 26802 12116
rect 3340 11908 3380 11948
rect 6883 11908 6923 11948
rect 8332 11908 8372 11948
rect 10444 11908 10484 11948
rect 12748 11908 12788 11948
rect 13996 11908 14036 11948
rect 14764 11908 14804 11948
rect 15724 11908 15764 11948
rect 17443 11908 17483 11948
rect 19372 11908 19412 11948
rect 22732 11908 22772 11948
rect 24076 11908 24116 11948
rect 25516 11908 25556 11948
rect 16460 11815 16500 11855
rect 27628 11824 27668 11864
rect 28108 11824 28148 11864
rect 979 11740 1019 11780
rect 2380 11740 2420 11780
rect 3619 11740 3659 11780
rect 3820 11740 3860 11780
rect 1174 11656 1214 11696
rect 1507 11656 1547 11696
rect 1612 11656 1652 11696
rect 2039 11656 2079 11696
rect 2179 11656 2219 11696
rect 2899 11698 2939 11738
rect 6220 11740 6260 11780
rect 6451 11731 6491 11771
rect 6898 11740 6938 11780
rect 11218 11740 11258 11780
rect 11731 11740 11771 11780
rect 13635 11740 13675 11780
rect 15436 11740 15476 11780
rect 15826 11740 15866 11780
rect 16972 11740 17012 11780
rect 18883 11740 18923 11780
rect 23443 11740 23483 11780
rect 27427 11740 27467 11780
rect 2284 11656 2324 11696
rect 3041 11656 3081 11696
rect 3351 11656 3391 11696
rect 3484 11656 3524 11696
rect 3724 11656 3764 11696
rect 4300 11656 4340 11696
rect 4972 11656 5012 11696
rect 5107 11656 5147 11696
rect 5495 11656 5535 11696
rect 5635 11656 5675 11696
rect 5740 11656 5780 11696
rect 6316 11656 6356 11696
rect 6553 11656 6593 11696
rect 6988 11656 7028 11696
rect 7756 11656 7796 11696
rect 8044 11656 8084 11696
rect 8413 11656 8453 11696
rect 8524 11656 8564 11696
rect 9004 11656 9044 11696
rect 9388 11656 9428 11696
rect 9772 11656 9812 11696
rect 9955 11656 9995 11696
rect 10150 11656 10190 11696
rect 10455 11656 10495 11696
rect 10636 11656 10676 11696
rect 10828 11656 10868 11696
rect 11308 11656 11348 11696
rect 11980 11656 12020 11696
rect 12364 11656 12404 11696
rect 12796 11656 12836 11696
rect 12940 11656 12980 11696
rect 13516 11656 13556 11696
rect 13733 11656 13773 11696
rect 13900 11656 13940 11696
rect 14092 11656 14132 11696
rect 14275 11656 14315 11696
rect 14380 11656 14420 11696
rect 14764 11656 14804 11696
rect 14956 11656 14996 11696
rect 15095 11656 15135 11696
rect 15235 11656 15275 11696
rect 15341 11656 15381 11696
rect 15916 11656 15956 11696
rect 16483 11656 16523 11696
rect 16684 11656 16724 11696
rect 17068 11656 17108 11696
rect 17187 11656 17227 11696
rect 17305 11656 17345 11696
rect 17441 11656 17481 11696
rect 17740 11656 17780 11696
rect 18508 11656 18548 11696
rect 18743 11656 18783 11696
rect 18988 11656 19028 11696
rect 19468 11656 19508 11696
rect 20035 11656 20075 11696
rect 20140 11656 20180 11696
rect 21187 11656 21227 11696
rect 23608 11656 23648 11696
rect 23788 11656 23828 11696
rect 23910 11656 23950 11696
rect 24037 11689 24077 11729
rect 24268 11656 24308 11696
rect 27043 11656 27083 11696
rect 27628 11689 27668 11729
rect 27726 11656 27766 11696
rect 27916 11689 27956 11729
rect 5827 11572 5867 11612
rect 9868 11572 9908 11612
rect 10252 11572 10292 11612
rect 10732 11572 10772 11612
rect 14476 11572 14516 11612
rect 14583 11572 14623 11612
rect 17644 11572 17684 11612
rect 18115 11572 18155 11612
rect 20803 11572 20843 11612
rect 25123 11572 25163 11612
rect 1900 11488 1940 11528
rect 2707 11488 2747 11528
rect 3139 11488 3179 11528
rect 4195 11488 4235 11528
rect 4492 11488 4532 11528
rect 5260 11488 5300 11528
rect 7555 11488 7595 11528
rect 9484 11488 9524 11528
rect 11011 11488 11051 11528
rect 13420 11488 13460 11528
rect 14371 11488 14411 11528
rect 19075 11488 19115 11528
rect 20428 11488 20468 11528
rect 23116 11488 23156 11528
rect 24940 11488 24980 11528
rect 4352 11320 4720 11360
rect 12126 11320 12494 11360
rect 19900 11320 20268 11360
rect 27674 11320 28042 11360
rect 748 11152 788 11192
rect 1612 11152 1652 11192
rect 2380 11152 2420 11192
rect 2764 11152 2804 11192
rect 3235 11152 3275 11192
rect 4195 11152 4235 11192
rect 4483 11152 4523 11192
rect 5452 11152 5492 11192
rect 6499 11152 6539 11192
rect 7324 11152 7364 11192
rect 7555 11152 7595 11192
rect 8524 11152 8564 11192
rect 9100 11152 9140 11192
rect 9868 11152 9908 11192
rect 10147 11152 10187 11192
rect 12355 11152 12395 11192
rect 12931 11152 12971 11192
rect 13219 11152 13259 11192
rect 13987 11152 14027 11192
rect 14755 11152 14795 11192
rect 16483 11152 16523 11192
rect 17740 11152 17780 11192
rect 18019 11152 18059 11192
rect 18499 11152 18539 11192
rect 20035 11152 20075 11192
rect 21772 11152 21812 11192
rect 23356 11152 23396 11192
rect 23980 11152 24020 11192
rect 24604 11152 24644 11192
rect 27715 11152 27755 11192
rect 4588 11068 4628 11108
rect 7770 11068 7810 11108
rect 8428 11068 8468 11108
rect 9571 11068 9611 11108
rect 10348 11068 10388 11108
rect 19708 11068 19748 11108
rect 652 10984 692 11024
rect 835 10984 875 11024
rect 1324 10984 1364 11024
rect 1459 10984 1499 11024
rect 1987 10984 2027 11024
rect 2092 10984 2132 11024
rect 2764 10984 2804 11024
rect 2956 10984 2996 11024
rect 3340 10984 3380 11024
rect 3724 10984 3764 11024
rect 3863 10984 3903 11024
rect 4108 10984 4148 11024
rect 4387 10984 4427 11024
rect 4695 10984 4735 11024
rect 5059 10984 5099 11024
rect 5164 10984 5204 11024
rect 5596 10984 5636 11024
rect 5897 10984 5937 11024
rect 6051 10984 6091 11024
rect 6604 10984 6644 11024
rect 6988 10984 7028 11024
rect 7180 10984 7220 11024
rect 7459 10984 7499 11024
rect 7948 10984 7988 11024
rect 8140 10984 8180 11024
rect 8323 10984 8363 11024
rect 8631 10984 8671 11024
rect 8812 10984 8852 11024
rect 8954 10984 8994 11024
rect 9239 10984 9279 11024
rect 9484 10984 9524 11024
rect 10060 10984 10100 11024
rect 10531 10984 10571 11024
rect 11128 10984 11168 11024
rect 11692 10984 11732 11024
rect 11875 10984 11915 11024
rect 4003 10900 4043 10940
rect 5740 10900 5780 10940
rect 9379 10900 9419 10940
rect 10963 10900 11003 10940
rect 11308 10900 11348 10940
rect 12028 10942 12068 10982
rect 12269 10984 12309 11024
rect 12604 10984 12644 11024
rect 12844 10984 12884 11024
rect 13420 10984 13460 11024
rect 13708 10984 13748 11024
rect 14092 10984 14132 11024
rect 14476 10984 14516 11024
rect 14956 10984 14996 11024
rect 15244 10984 15284 11024
rect 16012 10984 16052 11024
rect 16147 10984 16187 11024
rect 16780 10984 16820 11024
rect 17251 10984 17291 11024
rect 17548 10984 17588 11024
rect 17932 10984 17972 11024
rect 18167 10984 18207 11024
rect 18412 10984 18452 11024
rect 19030 10984 19070 11024
rect 19555 10975 19595 11015
rect 20332 10984 20372 11024
rect 20908 10984 20948 11024
rect 22444 10984 22484 11024
rect 22732 10984 22772 11024
rect 22924 10984 22964 11024
rect 23203 10975 23243 11015
rect 24172 10984 24212 11024
rect 24451 10975 24491 11015
rect 26947 10984 26987 11024
rect 27532 10984 27572 11024
rect 27724 10984 27764 11024
rect 5836 10816 5876 10856
rect 10572 10858 10612 10898
rect 12163 10900 12203 10940
rect 12739 10900 12779 10940
rect 16690 10900 16730 10940
rect 18307 10900 18347 10940
rect 18835 10900 18875 10940
rect 20242 10900 20282 10940
rect 25411 10900 25451 10940
rect 27331 10900 27371 10940
rect 11875 10816 11915 10856
rect 16195 10816 16235 10856
rect 17548 10816 17588 10856
rect 19372 10816 19412 10856
rect 22723 10816 22763 10856
rect 7756 10732 7796 10772
rect 8044 10732 8084 10772
rect 11548 10732 11588 10772
rect 21580 10732 21620 10772
rect 25036 10732 25076 10772
rect 3112 10564 3480 10604
rect 10886 10564 11254 10604
rect 18660 10564 19028 10604
rect 26434 10564 26802 10604
rect 1756 10396 1796 10436
rect 3139 10396 3179 10436
rect 3532 10396 3572 10436
rect 4483 10396 4523 10436
rect 6595 10396 6635 10436
rect 8716 10396 8756 10436
rect 9196 10396 9236 10436
rect 12067 10396 12107 10436
rect 13699 10396 13739 10436
rect 14188 10396 14228 10436
rect 16195 10396 16235 10436
rect 16588 10396 16628 10436
rect 21484 10396 21524 10436
rect 24076 10396 24116 10436
rect 931 10312 971 10352
rect 2524 10312 2564 10352
rect 4012 10312 4052 10352
rect 5356 10312 5396 10352
rect 8035 10312 8075 10352
rect 15532 10312 15572 10352
rect 17740 10312 17780 10352
rect 21868 10312 21908 10352
rect 23683 10312 23723 10352
rect 27148 10312 27188 10352
rect 1987 10228 2027 10268
rect 2188 10228 2228 10268
rect 4771 10228 4811 10268
rect 4972 10228 5012 10268
rect 5260 10228 5300 10268
rect 7276 10228 7316 10268
rect 11683 10228 11723 10268
rect 12643 10228 12683 10268
rect 12844 10228 12884 10268
rect 13228 10228 13268 10268
rect 13459 10219 13499 10259
rect 748 10144 788 10184
rect 931 10144 971 10184
rect 1132 10144 1172 10184
rect 1516 10144 1556 10184
rect 1847 10144 1887 10184
rect 2092 10144 2132 10184
rect 2380 10144 2420 10184
rect 2851 10144 2891 10184
rect 2956 10144 2996 10184
rect 3436 10144 3476 10184
rect 3628 10144 3668 10184
rect 3916 10144 3956 10184
rect 4108 10144 4148 10184
rect 4300 10144 4340 10184
rect 4491 10144 4531 10184
rect 4631 10144 4671 10184
rect 4876 10144 4916 10184
rect 5131 10144 5171 10184
rect 5417 10144 5457 10184
rect 5587 10144 5627 10184
rect 5740 10144 5780 10184
rect 5937 10144 5977 10184
rect 6307 10144 6347 10184
rect 6412 10144 6452 10184
rect 6957 10144 6997 10184
rect 7105 10144 7145 10184
rect 7397 10144 7437 10184
rect 7747 10144 7787 10184
rect 7852 10144 7892 10184
rect 8515 10144 8555 10184
rect 8620 10144 8660 10184
rect 9244 10144 9284 10184
rect 9388 10144 9428 10184
rect 10045 10144 10085 10184
rect 10156 10144 10196 10184
rect 10636 10144 10676 10184
rect 10775 10144 10815 10184
rect 11107 10177 11147 10217
rect 11543 10144 11583 10184
rect 11788 10144 11828 10184
rect 12062 10144 12102 10184
rect 12364 10144 12404 10184
rect 12523 10144 12563 10184
rect 12748 10144 12788 10184
rect 14188 10186 14228 10226
rect 13324 10144 13364 10184
rect 13561 10144 13601 10184
rect 13996 10144 14036 10184
rect 16690 10228 16730 10268
rect 14380 10186 14420 10226
rect 19564 10228 19604 10268
rect 24178 10228 24218 10268
rect 24883 10228 24923 10268
rect 14611 10144 14651 10184
rect 14713 10144 14753 10184
rect 15139 10144 15179 10184
rect 15256 10177 15296 10217
rect 16012 10144 16052 10184
rect 16147 10144 16187 10184
rect 16780 10144 16820 10184
rect 17260 10144 17300 10184
rect 17402 10144 17442 10184
rect 17932 10144 17972 10184
rect 18220 10144 18260 10184
rect 18403 10144 18443 10184
rect 18891 10144 18931 10184
rect 19027 10144 19067 10184
rect 19939 10144 19979 10184
rect 22060 10144 22100 10184
rect 23020 10144 23060 10184
rect 23395 10144 23435 10184
rect 23500 10144 23540 10184
rect 24268 10144 24308 10184
rect 25048 10144 25088 10184
rect 25420 10144 25460 10184
rect 26956 10144 26996 10184
rect 5740 9976 5780 10016
rect 7194 10018 7234 10058
rect 10972 10060 11012 10100
rect 13694 10060 13734 10100
rect 14908 10060 14948 10100
rect 17596 10060 17636 10100
rect 18316 10060 18356 10100
rect 9859 9976 9899 10016
rect 11260 9976 11300 10016
rect 11875 9976 11915 10016
rect 12268 9976 12308 10016
rect 13900 9976 13940 10016
rect 15043 9967 15083 10007
rect 18019 9976 18059 10016
rect 19180 9976 19220 10016
rect 22348 9976 22388 10016
rect 26092 9976 26132 10016
rect 26284 9976 26324 10016
rect 4352 9808 4720 9848
rect 12126 9808 12494 9848
rect 19900 9808 20268 9848
rect 27674 9808 28042 9848
rect 1123 9640 1163 9680
rect 1507 9640 1547 9680
rect 4780 9640 4820 9680
rect 4963 9640 5003 9680
rect 6316 9640 6356 9680
rect 7180 9640 7220 9680
rect 7564 9640 7604 9680
rect 8323 9640 8363 9680
rect 9475 9640 9515 9680
rect 11500 9640 11540 9680
rect 12364 9640 12404 9680
rect 13123 9640 13163 9680
rect 13795 9640 13835 9680
rect 13900 9640 13940 9680
rect 14275 9640 14315 9680
rect 15043 9640 15083 9680
rect 16291 9640 16331 9680
rect 18412 9640 18452 9680
rect 18787 9640 18827 9680
rect 19555 9640 19595 9680
rect 21091 9640 21131 9680
rect 22819 9640 22859 9680
rect 24172 9640 24212 9680
rect 25036 9640 25076 9680
rect 26188 9640 26228 9680
rect 1722 9556 1762 9596
rect 2179 9556 2219 9596
rect 7468 9556 7508 9596
rect 8812 9556 8852 9596
rect 10636 9556 10676 9596
rect 22147 9556 22187 9596
rect 652 9472 692 9512
rect 940 9472 980 9512
rect 1132 9472 1172 9512
rect 1411 9472 1451 9512
rect 1516 9472 1556 9512
rect 1847 9472 1887 9512
rect 2092 9472 2132 9512
rect 3052 9472 3092 9512
rect 3436 9472 3476 9512
rect 3724 9472 3764 9512
rect 4387 9472 4427 9512
rect 4492 9472 4532 9512
rect 5260 9472 5300 9512
rect 5836 9472 5876 9512
rect 6220 9472 6260 9512
rect 6787 9472 6827 9512
rect 6892 9472 6932 9512
rect 7363 9472 7403 9512
rect 7671 9472 7711 9512
rect 8236 9472 8276 9512
rect 8707 9472 8747 9512
rect 9015 9472 9055 9512
rect 9143 9472 9183 9512
rect 9388 9472 9428 9512
rect 9739 9472 9779 9512
rect 9964 9472 10004 9512
rect 10435 9472 10475 9512
rect 10732 9472 10772 9512
rect 11020 9472 11060 9512
rect 11404 9472 11444 9512
rect 11971 9472 12011 9512
rect 12076 9472 12116 9512
rect 12508 9472 12548 9512
rect 1987 9388 2027 9428
rect 5170 9388 5210 9428
rect 9283 9388 9323 9428
rect 9859 9388 9899 9428
rect 10060 9388 10100 9428
rect 12652 9388 12692 9428
rect 12816 9430 12856 9470
rect 12963 9472 13003 9512
rect 13276 9472 13316 9512
rect 13420 9472 13460 9512
rect 13694 9472 13734 9512
rect 13996 9463 14036 9503
rect 14476 9472 14516 9512
rect 14764 9472 14804 9512
rect 15244 9472 15284 9512
rect 15532 9472 15572 9512
rect 15767 9472 15807 9512
rect 16012 9472 16052 9512
rect 16444 9472 16484 9512
rect 16588 9472 16628 9512
rect 17212 9472 17252 9512
rect 17356 9472 17396 9512
rect 17548 9472 17588 9512
rect 17731 9472 17771 9512
rect 17932 9472 17972 9512
rect 18316 9472 18356 9512
rect 18973 9472 19013 9512
rect 19084 9472 19124 9512
rect 19708 9472 19748 9512
rect 19852 9472 19892 9512
rect 20620 9472 20660 9512
rect 21388 9472 21428 9512
rect 22540 9472 22580 9512
rect 23119 9472 23159 9512
rect 23779 9472 23819 9512
rect 23884 9472 23924 9512
rect 24643 9472 24683 9512
rect 24748 9472 24788 9512
rect 25411 9472 25451 9512
rect 26092 9472 26132 9512
rect 26275 9472 26315 9512
rect 15907 9388 15947 9428
rect 16108 9388 16148 9428
rect 20530 9388 20570 9428
rect 21298 9388 21338 9428
rect 23026 9388 23066 9428
rect 26476 9388 26516 9428
rect 4675 9304 4715 9344
rect 12748 9304 12788 9344
rect 17011 9304 17051 9344
rect 26716 9304 26756 9344
rect 796 9220 836 9260
rect 1708 9220 1748 9260
rect 2380 9220 2420 9260
rect 4060 9220 4100 9260
rect 7075 9220 7115 9260
rect 8044 9220 8084 9260
rect 9004 9220 9044 9260
rect 17731 9220 17771 9260
rect 20428 9220 20468 9260
rect 25612 9220 25652 9260
rect 3112 9052 3480 9092
rect 10886 9052 11254 9092
rect 18660 9052 19028 9092
rect 26434 9052 26802 9092
rect 2860 8884 2900 8924
rect 3619 8884 3659 8924
rect 5548 8884 5588 8924
rect 6028 8884 6068 8924
rect 7948 8884 7988 8924
rect 12652 8884 12692 8924
rect 16291 8884 16331 8924
rect 17539 8884 17579 8924
rect 18595 8884 18635 8924
rect 20131 8884 20171 8924
rect 21244 8884 21284 8924
rect 21868 8884 21908 8924
rect 23404 8884 23444 8924
rect 25708 8884 25748 8924
rect 5116 8800 5156 8840
rect 6268 8791 6308 8831
rect 6499 8800 6539 8840
rect 9859 8800 9899 8840
rect 13315 8800 13355 8840
rect 14092 8800 14132 8840
rect 24547 8800 24587 8840
rect 26860 8800 26900 8840
rect 940 8716 980 8756
rect 7267 8716 7307 8756
rect 8338 8716 8378 8756
rect 9139 8707 9179 8747
rect 10156 8716 10196 8756
rect 10732 8716 10772 8756
rect 13612 8716 13652 8756
rect 14188 8716 14228 8756
rect 15538 8716 15578 8756
rect 16963 8716 17003 8756
rect 18883 8716 18923 8756
rect 19459 8716 19499 8756
rect 23506 8716 23546 8756
rect 1315 8632 1355 8672
rect 3580 8632 3620 8672
rect 3724 8632 3764 8672
rect 4492 8632 4532 8672
rect 4780 8632 4820 8672
rect 5251 8632 5291 8672
rect 5356 8632 5396 8672
rect 5731 8632 5771 8672
rect 6307 8632 6347 8672
rect 6647 8632 6687 8672
rect 6787 8632 6827 8672
rect 6892 8632 6932 8672
rect 7127 8632 7167 8672
rect 7372 8632 7412 8672
rect 7651 8632 7691 8672
rect 7962 8632 8002 8672
rect 8428 8632 8468 8672
rect 9004 8632 9044 8672
rect 9241 8632 9281 8672
rect 9571 8632 9611 8672
rect 9676 8632 9716 8672
rect 10339 8632 10379 8672
rect 10924 8632 10964 8672
rect 11116 8632 11156 8672
rect 11308 8632 11348 8672
rect 11596 8632 11636 8672
rect 12460 8632 12500 8672
rect 13138 8632 13178 8672
rect 13267 8632 13307 8672
rect 13795 8632 13835 8672
rect 14524 8632 14564 8672
rect 14668 8632 14708 8672
rect 15628 8632 15668 8672
rect 16252 8632 16292 8672
rect 16396 8632 16436 8672
rect 16823 8632 16863 8672
rect 17061 8632 17101 8672
rect 17356 8632 17396 8672
rect 17539 8632 17579 8672
rect 17932 8632 17972 8672
rect 18412 8665 18452 8705
rect 25042 8716 25082 8756
rect 26595 8716 26635 8756
rect 18508 8632 18548 8672
rect 19267 8632 19307 8672
rect 19948 8632 19988 8672
rect 20083 8632 20123 8672
rect 20620 8632 20660 8672
rect 21004 8632 21044 8672
rect 21678 8632 21718 8672
rect 21868 8632 21908 8672
rect 22041 8632 22081 8672
rect 22243 8665 22283 8705
rect 22684 8632 22724 8672
rect 22874 8632 22914 8672
rect 23596 8632 23636 8672
rect 24370 8632 24410 8672
rect 24499 8632 24539 8672
rect 25132 8632 25172 8672
rect 25756 8632 25796 8672
rect 25900 8632 25940 8672
rect 26476 8632 26516 8672
rect 26716 8674 26756 8714
rect 26860 8632 26900 8672
rect 27052 8632 27092 8672
rect 27244 8632 27284 8672
rect 27436 8632 27476 8672
rect 5562 8548 5602 8588
rect 6039 8548 6079 8588
rect 7459 8548 7499 8588
rect 10636 8548 10676 8588
rect 17155 8548 17195 8588
rect 18979 8548 19019 8588
rect 21374 8548 21414 8588
rect 21475 8548 21515 8588
rect 26380 8548 26420 8588
rect 3244 8464 3284 8504
rect 5827 8464 5867 8504
rect 6979 8464 7019 8504
rect 7747 8464 7787 8504
rect 8131 8464 8171 8504
rect 8908 8464 8948 8504
rect 9964 8464 10004 8504
rect 11107 8464 11147 8504
rect 11788 8464 11828 8504
rect 12355 8464 12395 8504
rect 14371 8464 14411 8504
rect 15331 8464 15371 8504
rect 17788 8464 17828 8504
rect 21580 8464 21620 8504
rect 22396 8464 22436 8504
rect 23020 8464 23060 8504
rect 24835 8464 24875 8504
rect 27244 8464 27284 8504
rect 4352 8296 4720 8336
rect 12126 8296 12494 8336
rect 19900 8296 20268 8336
rect 27674 8296 28042 8336
rect 1219 8128 1259 8168
rect 3532 8128 3572 8168
rect 3868 8128 3908 8168
rect 4396 8128 4436 8168
rect 5260 8128 5300 8168
rect 5635 8128 5675 8168
rect 6796 8128 6836 8168
rect 7756 8128 7796 8168
rect 8716 8128 8756 8168
rect 9484 8128 9524 8168
rect 9763 8128 9803 8168
rect 10636 8128 10676 8168
rect 11395 8128 11435 8168
rect 12115 8128 12155 8168
rect 13612 8128 13652 8168
rect 14188 8128 14228 8168
rect 14860 8128 14900 8168
rect 16396 8128 16436 8168
rect 16675 8128 16715 8168
rect 17635 8128 17675 8168
rect 18892 8128 18932 8168
rect 21196 8128 21236 8168
rect 21571 8128 21611 8168
rect 23299 8128 23339 8168
rect 25795 8128 25835 8168
rect 25900 8128 25940 8168
rect 26275 8128 26315 8168
rect 5057 8044 5097 8084
rect 10433 8044 10473 8084
rect 15148 8044 15188 8084
rect 23201 8044 23241 8084
rect 23692 8044 23732 8084
rect 26380 8044 26420 8084
rect 652 7960 692 8000
rect 844 7960 884 8000
rect 1036 7960 1076 8000
rect 1227 7960 1267 8000
rect 1403 7960 1443 8000
rect 1612 7960 1652 8000
rect 2092 7960 2132 8000
rect 2284 7960 2324 8000
rect 2611 7960 2651 8000
rect 2806 7960 2846 8000
rect 3139 7960 3179 8000
rect 3244 7960 3284 8000
rect 3715 7951 3755 7991
rect 4492 7960 4532 8000
rect 4291 7918 4331 7958
rect 4612 7960 4652 8000
rect 5356 7951 5396 7991
rect 5836 7960 5876 8000
rect 6124 7960 6164 8000
rect 6316 7960 6356 8000
rect 6604 7960 6644 8000
rect 7363 7960 7403 8000
rect 8323 7960 8363 8000
rect 8428 7960 8468 8000
rect 9091 7960 9131 8000
rect 9196 7960 9236 8000
rect 9964 7960 10004 8000
rect 10252 7960 10292 8000
rect 10732 7951 10772 7991
rect 10871 7960 10911 8000
rect 11116 7960 11156 8000
rect 11581 7960 11621 8000
rect 11692 7960 11732 8000
rect 12259 7960 12299 8000
rect 12364 7951 12404 7991
rect 13132 7960 13172 8000
rect 13420 7960 13460 8000
rect 14284 7960 14324 8000
rect 14515 7960 14555 8000
rect 14657 7960 14697 8000
rect 14956 7951 14996 7991
rect 748 7876 788 7916
rect 7315 7848 7355 7888
rect 11011 7876 11051 7916
rect 15244 7918 15284 7958
rect 15379 7951 15419 7991
rect 15481 7960 15521 8000
rect 16003 7960 16043 8000
rect 16108 7960 16148 8000
rect 16876 7960 16916 8000
rect 17164 7960 17204 8000
rect 17740 7960 17780 8000
rect 18124 7960 18164 8000
rect 18499 7960 18539 8000
rect 18604 7960 18644 8000
rect 19084 7960 19124 8000
rect 19267 7960 19307 8000
rect 19768 7960 19808 8000
rect 20323 7960 20363 8000
rect 20428 7960 20468 8000
rect 20908 7960 20948 8000
rect 21036 7936 21076 7976
rect 21724 7960 21764 8000
rect 21868 7960 21908 8000
rect 22348 7960 22388 8000
rect 22492 7960 22532 8000
rect 22636 7960 22676 8000
rect 23404 7960 23444 8000
rect 23500 7951 23540 7991
rect 23788 7960 23828 8000
rect 24025 7960 24065 8000
rect 24133 7960 24173 8000
rect 24364 7960 24404 8000
rect 24844 7960 24884 8000
rect 25694 7960 25734 8000
rect 25996 7951 26036 7991
rect 26177 7960 26217 8000
rect 26478 7951 26518 7991
rect 26615 7960 26655 8000
rect 26860 7960 26900 8000
rect 11212 7876 11252 7916
rect 14419 7867 14459 7907
rect 19603 7876 19643 7916
rect 23907 7876 23947 7916
rect 24259 7876 24299 7916
rect 24460 7876 24500 7916
rect 26755 7876 26795 7916
rect 26956 7876 26996 7916
rect 27148 7792 27188 7832
rect 1516 7708 1556 7748
rect 2188 7708 2228 7748
rect 4780 7708 4820 7748
rect 5059 7708 5099 7748
rect 7555 7708 7595 7748
rect 10435 7708 10475 7748
rect 11500 7708 11540 7748
rect 12652 7708 12692 7748
rect 14659 7708 14699 7748
rect 19267 7708 19307 7748
rect 20524 7708 20564 7748
rect 21763 7708 21803 7748
rect 22828 7708 22868 7748
rect 25516 7708 25556 7748
rect 3112 7540 3480 7580
rect 10886 7540 11254 7580
rect 18660 7540 19028 7580
rect 26434 7540 26802 7580
rect 748 7372 788 7412
rect 3244 7372 3284 7412
rect 5347 7372 5387 7412
rect 8764 7372 8804 7412
rect 9580 7372 9620 7412
rect 12700 7372 12740 7412
rect 13987 7372 14027 7412
rect 14563 7372 14603 7412
rect 16588 7372 16628 7412
rect 17980 7372 18020 7412
rect 18748 7372 18788 7412
rect 20524 7372 20564 7412
rect 22828 7372 22868 7412
rect 26092 7372 26132 7412
rect 1036 7288 1076 7328
rect 4492 7288 4532 7328
rect 16348 7288 16388 7328
rect 21484 7288 21524 7328
rect 652 7120 692 7160
rect 849 7120 889 7160
rect 1036 7120 1076 7160
rect 1226 7120 1266 7160
rect 1420 7120 1460 7160
rect 1612 7120 1652 7160
rect 1900 7120 1940 7160
rect 2284 7120 2324 7160
rect 2426 7120 2466 7160
rect 2851 7120 2891 7160
rect 2960 7153 3000 7193
rect 3479 7120 3519 7160
rect 3619 7120 3659 7160
rect 3724 7120 3764 7160
rect 4108 7120 4148 7160
rect 5059 7120 5099 7160
rect 5164 7120 5204 7160
rect 5644 7120 5684 7160
rect 5836 7120 5876 7160
rect 5980 7162 6020 7202
rect 6316 7204 6356 7244
rect 7555 7204 7595 7244
rect 7756 7204 7796 7244
rect 9004 7204 9044 7244
rect 11596 7204 11636 7244
rect 19733 7204 19773 7244
rect 21004 7204 21044 7244
rect 6115 7120 6155 7160
rect 6220 7120 6260 7160
rect 6604 7120 6644 7160
rect 7415 7120 7455 7160
rect 7660 7120 7700 7160
rect 8140 7120 8180 7160
rect 8428 7120 8468 7160
rect 9100 7120 9140 7160
rect 9219 7120 9259 7160
rect 9337 7120 9377 7160
rect 9628 7120 9668 7160
rect 9772 7120 9812 7160
rect 10444 7120 10484 7160
rect 11011 7120 11051 7160
rect 11116 7120 11156 7160
rect 11692 7120 11732 7160
rect 11811 7120 11851 7160
rect 11929 7120 11969 7160
rect 12076 7120 12116 7160
rect 12364 7120 12404 7160
rect 13219 7120 13259 7160
rect 13324 7120 13364 7160
rect 13948 7120 13988 7160
rect 14092 7120 14132 7160
rect 14862 7120 14902 7160
rect 15436 7120 15476 7160
rect 15532 7120 15572 7160
rect 15724 7120 15764 7160
rect 16012 7120 16052 7160
rect 16636 7120 16676 7160
rect 16780 7120 16820 7160
rect 17356 7120 17396 7160
rect 17740 7120 17780 7160
rect 18124 7120 18164 7160
rect 18508 7120 18548 7160
rect 18883 7120 18923 7160
rect 19001 7120 19041 7160
rect 19167 7120 19207 7160
rect 19271 7120 19311 7160
rect 19401 7120 19441 7160
rect 19612 7120 19652 7160
rect 19852 7120 19892 7160
rect 20236 7120 20276 7160
rect 20419 7120 20459 7160
rect 20524 7120 20564 7160
rect 20663 7120 20703 7160
rect 20803 7120 20843 7160
rect 20908 7120 20948 7160
rect 21196 7120 21236 7160
rect 21318 7120 21358 7160
rect 21444 7120 21484 7160
rect 22300 7120 22340 7160
rect 22531 7120 22571 7160
rect 22828 7120 22868 7160
rect 23142 7162 23182 7202
rect 23017 7120 23057 7160
rect 23277 7153 23317 7193
rect 24163 7120 24203 7160
rect 26956 7120 26996 7160
rect 3811 7036 3851 7076
rect 14561 7036 14601 7076
rect 15230 7036 15270 7076
rect 23779 7036 23819 7076
rect 26275 7036 26315 7076
rect 1603 6952 1643 6992
rect 1795 6952 1835 6992
rect 2092 6952 2132 6992
rect 2572 6952 2612 6992
rect 2707 6952 2747 6992
rect 4003 6952 4043 6992
rect 4300 6952 4340 6992
rect 5740 6952 5780 6992
rect 7276 6952 7316 6992
rect 10339 6952 10379 6992
rect 10636 6952 10676 6992
rect 11404 6952 11444 6992
rect 13612 6952 13652 6992
rect 14764 6952 14804 6992
rect 15331 6952 15371 6992
rect 15436 6952 15476 6992
rect 19363 6952 19403 6992
rect 19939 6952 19979 6992
rect 21676 6952 21716 6992
rect 22732 6952 22772 6992
rect 23308 6952 23348 6992
rect 26092 6952 26132 6992
rect 4352 6784 4720 6824
rect 12126 6784 12494 6824
rect 19900 6784 20268 6824
rect 27674 6784 28042 6824
rect 1228 6616 1268 6656
rect 2284 6616 2324 6656
rect 3436 6616 3476 6656
rect 6028 6616 6068 6656
rect 6883 6616 6923 6656
rect 7852 6616 7892 6656
rect 8323 6616 8363 6656
rect 8668 6616 8708 6656
rect 9148 6616 9188 6656
rect 9475 6616 9515 6656
rect 10243 6616 10283 6656
rect 10540 6616 10580 6656
rect 11980 6616 12020 6656
rect 12451 6616 12491 6656
rect 13027 6616 13067 6656
rect 13132 6616 13172 6656
rect 13507 6616 13547 6656
rect 14668 6616 14708 6656
rect 15148 6616 15188 6656
rect 16108 6616 16148 6656
rect 16675 6616 16715 6656
rect 17443 6616 17483 6656
rect 18211 6616 18251 6656
rect 18508 6616 18548 6656
rect 18787 6616 18827 6656
rect 18892 6616 18932 6656
rect 19372 6616 19412 6656
rect 22636 6616 22676 6656
rect 23203 6616 23243 6656
rect 24268 6616 24308 6656
rect 1612 6532 1652 6572
rect 8428 6532 8468 6572
rect 18686 6532 18726 6572
rect 20044 6532 20084 6572
rect 20323 6532 20363 6572
rect 1132 6448 1172 6488
rect 1315 6448 1355 6488
rect 1523 6448 1563 6488
rect 1699 6448 1739 6488
rect 2188 6448 2228 6488
rect 2371 6448 2411 6488
rect 2956 6448 2996 6488
rect 3340 6448 3380 6488
rect 4099 6448 4139 6488
rect 6547 6448 6587 6488
rect 6742 6448 6782 6488
rect 6988 6448 7028 6488
rect 7372 6448 7412 6488
rect 7660 6448 7700 6488
rect 8227 6448 8267 6488
rect 8535 6448 8575 6488
rect 8812 6448 8852 6488
rect 8995 6439 9035 6479
rect 9628 6448 9668 6488
rect 9772 6448 9812 6488
rect 10348 6448 10388 6488
rect 10876 6448 10916 6488
rect 11020 6448 11060 6488
rect 11500 6448 11540 6488
rect 11788 6448 11828 6488
rect 12556 6448 12596 6488
rect 12929 6448 12969 6488
rect 13228 6439 13268 6479
rect 13708 6448 13748 6488
rect 13996 6448 14036 6488
rect 14188 6448 14228 6488
rect 14476 6448 14516 6488
rect 14947 6448 14987 6488
rect 15244 6448 15284 6488
rect 15628 6448 15668 6488
rect 16012 6448 16052 6488
rect 16828 6448 16868 6488
rect 16970 6458 17010 6498
rect 17740 6448 17780 6488
rect 18316 6448 18356 6488
rect 18988 6439 19028 6479
rect 19276 6448 19316 6488
rect 19459 6448 19499 6488
rect 19843 6448 19883 6488
rect 20140 6448 20180 6488
rect 20707 6448 20747 6488
rect 23308 6448 23348 6488
rect 23644 6448 23684 6488
rect 23884 6448 23924 6488
rect 24076 6448 24116 6488
rect 24940 6448 24980 6488
rect 25804 6448 25844 6488
rect 3724 6364 3764 6404
rect 17650 6364 17690 6404
rect 22252 6364 22292 6404
rect 25123 6364 25163 6404
rect 2572 6280 2612 6320
rect 7180 6280 7220 6320
rect 12748 6280 12788 6320
rect 25996 6280 26036 6320
rect 5644 6196 5684 6236
rect 6028 6196 6068 6236
rect 10828 6196 10868 6236
rect 22636 6196 22676 6236
rect 23884 6196 23924 6236
rect 3112 6028 3480 6068
rect 10886 6028 11254 6068
rect 18660 6028 19028 6068
rect 26434 6028 26802 6068
rect 3532 5860 3572 5900
rect 8428 5860 8468 5900
rect 8812 5860 8852 5900
rect 12172 5860 12212 5900
rect 15724 5860 15764 5900
rect 16972 5860 17012 5900
rect 20332 5860 20372 5900
rect 21484 5860 21524 5900
rect 24268 5860 24308 5900
rect 25132 5860 25172 5900
rect 3916 5776 3956 5816
rect 4156 5767 4196 5807
rect 4684 5776 4724 5816
rect 12556 5776 12596 5816
rect 17356 5776 17396 5816
rect 21868 5776 21908 5816
rect 24652 5776 24692 5816
rect 5356 5692 5396 5732
rect 16435 5692 16475 5732
rect 3532 5608 3572 5648
rect 3724 5608 3764 5648
rect 4099 5608 4139 5648
rect 5035 5608 5075 5648
rect 5155 5608 5195 5648
rect 5260 5608 5300 5648
rect 5836 5608 5876 5648
rect 6016 5608 6056 5648
rect 6883 5608 6923 5648
rect 9196 5608 9236 5648
rect 10627 5608 10667 5648
rect 13036 5608 13076 5648
rect 13180 5608 13220 5648
rect 14179 5608 14219 5648
rect 16630 5608 16670 5648
rect 18883 5608 18923 5648
rect 19468 5608 19508 5648
rect 21004 5608 21044 5648
rect 21187 5608 21227 5648
rect 21292 5608 21332 5648
rect 22723 5608 22763 5648
rect 24835 5608 24875 5648
rect 25132 5608 25172 5648
rect 5534 5524 5574 5564
rect 5635 5524 5675 5564
rect 6499 5524 6539 5564
rect 10243 5524 10283 5564
rect 12835 5524 12875 5564
rect 13795 5524 13835 5564
rect 19267 5524 19307 5564
rect 20140 5524 20180 5564
rect 21495 5524 21535 5564
rect 22339 5524 22379 5564
rect 5740 5440 5780 5480
rect 6172 5440 6212 5480
rect 9868 5440 9908 5480
rect 13132 5440 13172 5480
rect 16108 5440 16148 5480
rect 4352 5272 4720 5312
rect 12126 5272 12494 5312
rect 19900 5272 20268 5312
rect 27674 5272 28042 5312
rect 6364 5104 6404 5144
rect 9139 5104 9179 5144
rect 10060 5104 10100 5144
rect 10828 5104 10868 5144
rect 11779 5104 11819 5144
rect 13795 5104 13835 5144
rect 16972 5104 17012 5144
rect 20716 5104 20756 5144
rect 21196 5104 21236 5144
rect 23596 5104 23636 5144
rect 23971 5104 24011 5144
rect 12076 5020 12116 5060
rect 13900 5020 13940 5060
rect 16012 5020 16052 5060
rect 23870 5020 23910 5060
rect 24076 5020 24116 5060
rect 6220 4936 6260 4976
rect 9334 4936 9374 4976
rect 9667 4936 9707 4976
rect 9772 4936 9812 4976
rect 10540 4936 10580 4976
rect 10732 4936 10772 4976
rect 10924 4936 10964 4976
rect 11447 4936 11487 4976
rect 11692 4936 11732 4976
rect 11980 4936 12020 4976
rect 12172 4936 12212 4976
rect 12748 4936 12788 4976
rect 12931 4936 12971 4976
rect 13036 4936 13076 4976
rect 13228 4936 13268 4976
rect 13350 4936 13390 4976
rect 13477 4936 13517 4976
rect 13699 4936 13739 4976
rect 14007 4936 14047 4976
rect 14236 4936 14276 4976
rect 14860 4936 14900 4976
rect 15619 4936 15659 4976
rect 16300 4936 16340 4976
rect 19084 4936 19124 4976
rect 19267 4936 19307 4976
rect 19651 4936 19691 4976
rect 19756 4936 19796 4976
rect 20236 4936 20276 4976
rect 20405 4936 20445 4976
rect 20524 4936 20564 4976
rect 21004 4936 21044 4976
rect 21196 4936 21236 4976
rect 21388 4936 21428 4976
rect 22636 4936 22676 4976
rect 22819 4936 22859 4976
rect 23020 4936 23060 4976
rect 23203 4936 23243 4976
rect 23314 4936 23354 4976
rect 23515 4936 23555 4976
rect 23692 4936 23732 4976
rect 24172 4927 24212 4967
rect 10444 4852 10484 4892
rect 11587 4852 11627 4892
rect 20860 4852 20900 4892
rect 7564 4768 7604 4808
rect 11123 4768 11163 4808
rect 13036 4768 13076 4808
rect 13516 4768 13556 4808
rect 15052 4768 15092 4808
rect 18220 4768 18260 4808
rect 19267 4768 19307 4808
rect 21580 4768 21620 4808
rect 22819 4768 22859 4808
rect 15820 4684 15860 4724
rect 19852 4684 19892 4724
rect 23308 4684 23348 4724
rect 3112 4516 3480 4556
rect 10886 4516 11254 4556
rect 18660 4516 19028 4556
rect 26434 4516 26802 4556
rect 19843 4348 19883 4388
rect 20332 4348 20372 4388
rect 20668 4348 20708 4388
rect 10060 4264 10100 4304
rect 9964 4096 10004 4136
rect 10156 4096 10196 4136
rect 19660 4096 19700 4136
rect 19843 4096 19883 4136
rect 20332 4096 20372 4136
rect 20524 4096 20564 4136
rect 20812 4096 20852 4136
rect 4352 3760 4720 3800
rect 12126 3760 12494 3800
rect 19900 3760 20268 3800
rect 27674 3760 28042 3800
rect 3112 3004 3480 3044
rect 10886 3004 11254 3044
rect 18660 3004 19028 3044
rect 26434 3004 26802 3044
rect 4352 2248 4720 2288
rect 12126 2248 12494 2288
rect 19900 2248 20268 2288
rect 27674 2248 28042 2288
rect 3112 1492 3480 1532
rect 10886 1492 11254 1532
rect 18660 1492 19028 1532
rect 26434 1492 26802 1532
rect 4352 736 4720 776
rect 12126 736 12494 776
rect 19900 736 20268 776
rect 27674 736 28042 776
<< metal2 >>
rect 2083 28876 2092 28916
rect 2132 28876 13516 28916
rect 13556 28876 13565 28916
rect 5635 28624 5644 28664
rect 5684 28624 12652 28664
rect 12692 28624 12701 28664
rect 4867 28540 4876 28580
rect 4916 28540 14092 28580
rect 14132 28540 14141 28580
rect 16483 28540 16492 28580
rect 16532 28540 30028 28580
rect 30068 28540 30077 28580
rect 2371 28456 2380 28496
rect 2420 28456 2900 28496
rect 4099 28456 4108 28496
rect 4148 28456 12980 28496
rect 24643 28456 24652 28496
rect 24692 28456 27244 28496
rect 27284 28456 27293 28496
rect 2860 28412 2900 28456
rect 12940 28412 12980 28456
rect 2860 28372 9196 28412
rect 9236 28372 9245 28412
rect 12940 28372 13708 28412
rect 13748 28372 13757 28412
rect 19459 28372 19468 28412
rect 19508 28372 28972 28412
rect 29012 28372 29021 28412
rect 2467 28288 2476 28328
rect 2516 28288 12556 28328
rect 12596 28288 12605 28328
rect 23875 28288 23884 28328
rect 23924 28288 26764 28328
rect 26804 28288 26813 28328
rect 23107 28204 23116 28244
rect 23156 28204 30028 28244
rect 30068 28204 30077 28244
rect 23779 28120 23788 28160
rect 23828 28120 28876 28160
rect 28916 28120 28925 28160
rect 2083 28036 2092 28076
rect 2132 28036 2141 28076
rect 2188 28036 13804 28076
rect 13844 28036 13853 28076
rect 24556 28036 29684 28076
rect 1036 27868 1900 27908
rect 1940 27868 1949 27908
rect 1036 27656 1076 27868
rect 2092 27824 2132 28036
rect 2083 27784 2092 27824
rect 2132 27784 2141 27824
rect 1891 27700 1900 27740
rect 1940 27700 1949 27740
rect 1997 27700 2092 27740
rect 2132 27700 2141 27740
rect 1900 27656 1940 27700
rect 1997 27656 2037 27700
rect 2188 27656 2228 28036
rect 13132 27992 13172 28036
rect 4343 27952 4352 27992
rect 4720 27952 4729 27992
rect 5347 27952 5356 27992
rect 5396 27952 11308 27992
rect 11348 27952 11357 27992
rect 12117 27952 12126 27992
rect 12494 27952 12503 27992
rect 13123 27952 13132 27992
rect 13172 27952 13248 27992
rect 19891 27952 19900 27992
rect 20268 27952 20277 27992
rect 24556 27908 24596 28036
rect 27665 27952 27674 27992
rect 28042 27952 28051 27992
rect 2275 27868 2284 27908
rect 2324 27868 3052 27908
rect 3092 27868 4972 27908
rect 5012 27868 5021 27908
rect 5164 27868 8620 27908
rect 8660 27868 8669 27908
rect 13036 27868 13900 27908
rect 13940 27868 13949 27908
rect 20044 27868 24596 27908
rect 25324 27868 26380 27908
rect 26420 27868 26429 27908
rect 27043 27868 27052 27908
rect 27092 27868 27908 27908
rect 5164 27824 5204 27868
rect 13036 27824 13076 27868
rect 2345 27784 2476 27824
rect 2516 27784 2525 27824
rect 2938 27784 2947 27824
rect 2996 27784 3127 27824
rect 3977 27784 4099 27824
rect 4148 27784 4157 27824
rect 4204 27784 5108 27824
rect 5155 27784 5164 27824
rect 5204 27784 5213 27824
rect 5539 27784 5548 27824
rect 5588 27784 7316 27824
rect 9283 27784 9292 27824
rect 9332 27784 10732 27824
rect 10772 27784 10781 27824
rect 13027 27784 13036 27824
rect 13076 27784 13085 27824
rect 13507 27784 13516 27824
rect 13556 27784 14228 27824
rect 19337 27784 19468 27824
rect 19508 27784 19517 27824
rect 19738 27784 19747 27824
rect 19787 27784 19872 27824
rect 4204 27740 4244 27784
rect 835 27616 844 27656
rect 884 27616 893 27656
rect 1027 27616 1036 27656
rect 1076 27616 1085 27656
rect 1132 27616 1516 27656
rect 1556 27616 1612 27656
rect 1652 27616 1687 27656
rect 1793 27616 1802 27656
rect 1842 27616 1940 27656
rect 1994 27616 2003 27656
rect 2043 27616 2052 27656
rect 2170 27616 2179 27656
rect 2219 27616 2228 27656
rect 2284 27700 2380 27740
rect 2420 27700 2429 27740
rect 2851 27700 2860 27740
rect 2900 27700 3188 27740
rect 2284 27656 2324 27700
rect 3148 27656 3188 27700
rect 3916 27700 4244 27740
rect 5068 27740 5108 27784
rect 5068 27700 6067 27740
rect 6107 27700 6604 27740
rect 6644 27700 6653 27740
rect 6874 27700 6883 27740
rect 6932 27700 7063 27740
rect 3916 27656 3956 27700
rect 2284 27616 2375 27656
rect 2415 27616 2424 27656
rect 2557 27616 2566 27656
rect 2606 27616 2615 27656
rect 2755 27616 2764 27656
rect 2804 27616 2851 27656
rect 2946 27616 2955 27656
rect 2995 27616 3092 27656
rect 3146 27616 3155 27656
rect 3195 27616 3204 27656
rect 3322 27616 3331 27656
rect 3380 27616 3511 27656
rect 3907 27616 3916 27656
rect 3956 27616 3965 27656
rect 844 27572 884 27616
rect 1132 27572 1172 27616
rect 2572 27572 2612 27616
rect 2764 27572 2804 27616
rect 3052 27572 3092 27616
rect 4103 27611 4112 27651
rect 4152 27611 4161 27651
rect 844 27532 1172 27572
rect 1420 27532 2380 27572
rect 2420 27532 2429 27572
rect 2563 27532 2572 27572
rect 2612 27532 2653 27572
rect 2755 27532 2764 27572
rect 2804 27532 2813 27572
rect 3043 27532 3052 27572
rect 3092 27532 3101 27572
rect 3244 27532 3724 27572
rect 3764 27532 3773 27572
rect 1420 27488 1460 27532
rect 3244 27488 3284 27532
rect 1411 27448 1420 27488
rect 1460 27448 1469 27488
rect 1603 27448 1612 27488
rect 1652 27448 3284 27488
rect 3593 27448 3628 27488
rect 3668 27448 3724 27488
rect 3764 27448 3773 27488
rect 4108 27404 4148 27611
rect 4204 27572 4244 27700
rect 4286 27635 4295 27675
rect 4335 27635 4344 27675
rect 7276 27656 7316 27784
rect 9946 27700 9955 27740
rect 9995 27700 10540 27740
rect 10580 27700 12116 27740
rect 12250 27700 12259 27740
rect 12299 27700 13795 27740
rect 13835 27700 13844 27740
rect 13891 27700 13900 27740
rect 13940 27700 14071 27740
rect 12076 27667 12116 27700
rect 12076 27656 12212 27667
rect 14188 27656 14228 27784
rect 19756 27740 19796 27784
rect 16300 27700 17300 27740
rect 18019 27700 18028 27740
rect 18068 27700 19939 27740
rect 19979 27700 19988 27740
rect 16300 27656 16340 27700
rect 17260 27656 17300 27700
rect 4300 27572 4340 27635
rect 4483 27616 4492 27656
rect 4532 27616 4663 27656
rect 4937 27616 5068 27656
rect 5108 27616 5117 27656
rect 5242 27616 5251 27656
rect 5300 27616 5431 27656
rect 5731 27616 5740 27656
rect 5792 27616 5911 27656
rect 6110 27616 6220 27656
rect 6272 27616 6290 27656
rect 6392 27616 6401 27656
rect 6441 27616 6452 27656
rect 6691 27616 6700 27656
rect 6740 27616 6871 27656
rect 7258 27616 7267 27656
rect 7307 27616 7316 27656
rect 9566 27616 9676 27656
rect 9728 27616 9746 27656
rect 11491 27616 11500 27656
rect 11540 27616 11875 27656
rect 11915 27616 11924 27656
rect 12076 27627 12643 27656
rect 12172 27616 12643 27627
rect 12683 27616 12692 27656
rect 12739 27616 12748 27656
rect 12788 27616 12797 27656
rect 13097 27616 13228 27656
rect 13268 27616 13277 27656
rect 6412 27572 6452 27616
rect 6700 27598 6740 27607
rect 12748 27572 12788 27616
rect 13361 27584 13370 27624
rect 13410 27584 13419 27624
rect 13507 27616 13516 27656
rect 13556 27616 13694 27656
rect 13734 27616 13743 27656
rect 13996 27647 14228 27656
rect 14036 27616 14228 27647
rect 14275 27616 14284 27656
rect 14324 27616 16291 27656
rect 16331 27616 16340 27656
rect 16666 27616 16675 27656
rect 16724 27616 16855 27656
rect 17242 27616 17251 27656
rect 17291 27616 17300 27656
rect 19529 27616 19660 27656
rect 19700 27616 19709 27656
rect 13996 27598 14036 27607
rect 4195 27532 4204 27572
rect 4244 27532 4253 27572
rect 4300 27532 5356 27572
rect 5396 27532 5405 27572
rect 5539 27532 5548 27572
rect 5627 27532 5719 27572
rect 6307 27532 6316 27572
rect 6356 27532 6452 27572
rect 8419 27532 8428 27572
rect 8468 27532 8477 27572
rect 9475 27532 9484 27572
rect 9563 27532 9655 27572
rect 10636 27563 10676 27572
rect 12355 27532 12364 27572
rect 12404 27532 12788 27572
rect 13379 27572 13419 27584
rect 20044 27572 20084 27868
rect 25324 27824 25364 27868
rect 27868 27824 27908 27868
rect 22435 27784 22444 27824
rect 22484 27784 25364 27824
rect 25411 27784 25420 27824
rect 25460 27784 27724 27824
rect 27764 27784 27773 27824
rect 27859 27784 27868 27824
rect 27908 27784 27917 27824
rect 22060 27700 23788 27740
rect 23828 27700 23837 27740
rect 24163 27700 24172 27740
rect 24212 27700 25804 27740
rect 25844 27700 25853 27740
rect 26179 27700 26188 27740
rect 26228 27700 27860 27740
rect 28483 27700 28492 27740
rect 28532 27700 29204 27740
rect 21737 27616 21859 27656
rect 21908 27616 21917 27656
rect 13379 27532 13804 27572
rect 13844 27532 13853 27572
rect 14083 27532 14092 27572
rect 14132 27532 15072 27572
rect 16745 27532 16876 27572
rect 16916 27532 16925 27572
rect 18528 27532 20084 27572
rect 22060 27552 22100 27700
rect 25790 27656 25830 27700
rect 27820 27656 27860 27700
rect 29164 27656 29204 27700
rect 24233 27616 24355 27656
rect 24404 27616 24413 27656
rect 24931 27616 24940 27656
rect 24980 27616 25228 27656
rect 25268 27616 25277 27656
rect 25781 27616 25790 27656
rect 25830 27616 25839 27656
rect 25889 27616 25900 27656
rect 25940 27616 25949 27656
rect 26083 27616 26092 27656
rect 26132 27616 26141 27656
rect 26266 27647 26380 27656
rect 25889 27572 25929 27616
rect 26092 27572 26132 27616
rect 26266 27607 26275 27647
rect 26315 27616 26380 27647
rect 26420 27616 26455 27656
rect 26633 27647 26764 27656
rect 26633 27616 26755 27647
rect 26804 27616 26813 27656
rect 27113 27647 27244 27656
rect 27113 27616 27235 27647
rect 27284 27616 27293 27656
rect 27593 27647 27724 27656
rect 27593 27616 27715 27647
rect 27764 27616 27773 27656
rect 27820 27647 28244 27656
rect 27820 27616 28195 27647
rect 26315 27607 26324 27616
rect 26266 27606 26324 27607
rect 26746 27607 26755 27616
rect 26795 27607 26804 27616
rect 26746 27606 26804 27607
rect 27226 27607 27235 27616
rect 27275 27607 27284 27616
rect 27226 27606 27284 27607
rect 27706 27607 27715 27616
rect 27755 27607 27764 27616
rect 27706 27606 27764 27607
rect 28186 27607 28195 27616
rect 28235 27607 28244 27647
rect 28553 27647 28684 27656
rect 28553 27616 28675 27647
rect 28724 27616 28733 27656
rect 29146 27647 29204 27656
rect 28186 27606 28244 27607
rect 28666 27607 28675 27616
rect 28715 27607 28724 27616
rect 28666 27606 28724 27607
rect 29146 27607 29155 27647
rect 29195 27607 29204 27647
rect 29146 27606 29204 27607
rect 22234 27532 22243 27572
rect 22292 27532 22423 27572
rect 24547 27532 24556 27572
rect 24596 27532 24605 27572
rect 24730 27532 24739 27572
rect 24788 27532 24919 27572
rect 25889 27532 25900 27572
rect 25940 27532 25965 27572
rect 26092 27532 26188 27572
rect 26228 27532 26237 27572
rect 26419 27532 26428 27572
rect 26468 27532 26476 27572
rect 26516 27532 26599 27572
rect 26851 27532 26860 27572
rect 26900 27532 26908 27572
rect 26948 27532 27031 27572
rect 27379 27532 27388 27572
rect 27428 27532 27436 27572
rect 27476 27532 27559 27572
rect 28339 27532 28348 27572
rect 28388 27532 28492 27572
rect 28532 27532 28541 27572
rect 28771 27532 28780 27572
rect 28820 27532 28828 27572
rect 28868 27532 28951 27572
rect 29251 27532 29260 27572
rect 29300 27532 29308 27572
rect 29348 27532 29431 27572
rect 10636 27514 10676 27523
rect 29644 27488 29684 28036
rect 30787 27616 30796 27656
rect 30836 27647 30967 27656
rect 30836 27616 30883 27647
rect 30874 27607 30883 27616
rect 30923 27616 30967 27647
rect 30923 27607 30932 27616
rect 30874 27606 30932 27607
rect 30979 27532 30988 27572
rect 31028 27532 31036 27572
rect 31076 27532 31159 27572
rect 4265 27448 4396 27488
rect 4436 27448 4445 27488
rect 4745 27448 4876 27488
rect 4916 27448 4925 27488
rect 8620 27448 10580 27488
rect 643 27364 652 27404
rect 692 27364 844 27404
rect 884 27364 893 27404
rect 3322 27364 3331 27404
rect 3371 27364 4052 27404
rect 4108 27364 6218 27404
rect 6281 27364 6403 27404
rect 6452 27364 6461 27404
rect 4012 27320 4052 27364
rect 6178 27320 6218 27364
rect 8620 27320 8660 27448
rect 10540 27404 10580 27448
rect 11596 27448 11980 27488
rect 12020 27448 12029 27488
rect 19171 27448 19180 27488
rect 19220 27448 19564 27488
rect 19604 27448 19613 27488
rect 25603 27448 25612 27488
rect 25652 27448 27532 27488
rect 27572 27448 27581 27488
rect 29635 27448 29644 27488
rect 29684 27448 29693 27488
rect 29897 27448 29932 27488
rect 29972 27448 30028 27488
rect 30068 27448 30077 27488
rect 30211 27448 30220 27488
rect 30260 27448 30412 27488
rect 30452 27448 30461 27488
rect 11596 27404 11636 27448
rect 9065 27364 9196 27404
rect 9236 27364 9245 27404
rect 10540 27364 11636 27404
rect 14371 27364 14380 27404
rect 14420 27364 14429 27404
rect 18307 27364 18316 27404
rect 18356 27364 19468 27404
rect 19508 27364 19517 27404
rect 22819 27364 22828 27404
rect 22868 27364 23692 27404
rect 23732 27364 23741 27404
rect 25795 27364 25804 27404
rect 25844 27364 25975 27404
rect 26371 27364 26380 27404
rect 26420 27364 30260 27404
rect 2179 27280 2188 27320
rect 2228 27280 3956 27320
rect 4003 27280 4012 27320
rect 4052 27280 4061 27320
rect 4108 27280 4972 27320
rect 5012 27280 5021 27320
rect 6178 27280 8660 27320
rect 2188 27236 2228 27280
rect 3916 27236 3956 27280
rect 4108 27236 4148 27280
rect 1804 27196 2228 27236
rect 3103 27196 3112 27236
rect 3480 27196 3489 27236
rect 3916 27196 4148 27236
rect 4579 27196 4588 27236
rect 4628 27196 6316 27236
rect 6356 27196 8332 27236
rect 8372 27196 9484 27236
rect 9524 27196 9533 27236
rect 10877 27196 10886 27236
rect 11254 27196 11263 27236
rect 1804 27068 1844 27196
rect 1996 27112 9868 27152
rect 9908 27112 9917 27152
rect 1996 27068 2036 27112
rect 14380 27068 14420 27364
rect 30220 27320 30260 27364
rect 16003 27280 16012 27320
rect 16052 27280 23116 27320
rect 23156 27280 23165 27320
rect 30220 27280 30932 27320
rect 18651 27196 18660 27236
rect 19028 27196 19037 27236
rect 23395 27196 23404 27236
rect 23444 27196 25996 27236
rect 26036 27196 26045 27236
rect 26425 27196 26434 27236
rect 26802 27196 26811 27236
rect 26947 27196 26956 27236
rect 26996 27196 30644 27236
rect 15235 27112 15244 27152
rect 15284 27112 19276 27152
rect 19316 27112 19325 27152
rect 19747 27112 19756 27152
rect 19796 27112 29156 27152
rect 17356 27068 17396 27112
rect 29116 27068 29156 27112
rect 883 27028 892 27068
rect 932 27028 1844 27068
rect 1978 27028 1987 27068
rect 2027 27028 2036 27068
rect 2362 27028 2371 27068
rect 2411 27028 3340 27068
rect 3380 27028 3389 27068
rect 9545 27028 9676 27068
rect 9716 27028 9725 27068
rect 9772 27028 10348 27068
rect 10388 27028 10397 27068
rect 11971 27028 11980 27068
rect 12020 27028 12172 27068
rect 12212 27028 12221 27068
rect 14179 27028 14188 27068
rect 14228 27028 15764 27068
rect 17347 27028 17356 27068
rect 17396 27028 17405 27068
rect 18403 27028 18412 27068
rect 18452 27028 20524 27068
rect 20564 27028 20573 27068
rect 21667 27028 21676 27068
rect 21716 27028 22252 27068
rect 22292 27028 22301 27068
rect 22435 27028 22444 27068
rect 22484 27028 23500 27068
rect 23540 27028 23596 27068
rect 23636 27028 23700 27068
rect 25036 27028 28108 27068
rect 28148 27028 28157 27068
rect 29107 27028 29116 27068
rect 29156 27028 29165 27068
rect 29513 27028 29644 27068
rect 29684 27028 29693 27068
rect 9772 26984 9812 27028
rect 3523 26944 3532 26984
rect 3572 26944 3628 26984
rect 3668 26944 3703 26984
rect 3907 26944 3916 26984
rect 3956 26944 5108 26984
rect 643 26860 652 26900
rect 692 26860 1036 26900
rect 1076 26860 1085 26900
rect 1385 26860 1420 26900
rect 1460 26860 1516 26900
rect 1556 26860 1565 26900
rect 1651 26860 1660 26900
rect 1700 26860 2380 26900
rect 2420 26860 2429 26900
rect 2476 26860 2764 26900
rect 2804 26860 2813 26900
rect 2956 26860 3148 26900
rect 3188 26860 3197 26900
rect 3331 26860 3340 26900
rect 3380 26860 4780 26900
rect 4820 26860 4829 26900
rect 2476 26816 2516 26860
rect 2956 26816 2996 26860
rect 643 26776 652 26816
rect 692 26776 1036 26816
rect 1076 26776 1085 26816
rect 1210 26776 1219 26816
rect 1268 26776 1399 26816
rect 1673 26776 1804 26816
rect 1844 26776 1853 26816
rect 1961 26776 1987 26816
rect 2027 26776 2092 26816
rect 2132 26776 2141 26816
rect 2186 26776 2195 26816
rect 2235 26776 2275 26816
rect 2332 26776 2371 26816
rect 2411 26776 2516 26816
rect 2563 26776 2572 26816
rect 2612 26776 2708 26816
rect 2755 26776 2764 26816
rect 2804 26776 2900 26816
rect 2947 26776 2956 26816
rect 2996 26776 3005 26816
rect 3139 26776 3148 26816
rect 3188 26776 4588 26816
rect 4628 26776 4637 26816
rect 4771 26776 4780 26816
rect 4820 26776 4876 26816
rect 4916 26776 4951 26816
rect 2188 26732 2228 26776
rect 2179 26692 2188 26732
rect 2228 26692 2237 26732
rect 2332 26648 2372 26776
rect 2668 26732 2708 26776
rect 2659 26692 2668 26732
rect 2708 26692 2717 26732
rect 1123 26608 1132 26648
rect 1172 26608 1303 26648
rect 1987 26608 1996 26648
rect 2036 26608 2372 26648
rect 2633 26608 2755 26648
rect 2804 26608 2813 26648
rect 2860 26396 2900 26776
rect 5068 26732 5108 26944
rect 6700 26944 9812 26984
rect 6307 26860 6316 26900
rect 6356 26860 6365 26900
rect 5338 26776 5347 26816
rect 5387 26776 5548 26816
rect 5588 26776 5597 26816
rect 6700 26732 6740 26944
rect 2947 26692 2956 26732
rect 2996 26692 4244 26732
rect 4841 26692 4963 26732
rect 5012 26692 5021 26732
rect 5068 26692 6740 26732
rect 6796 26860 8468 26900
rect 4204 26648 4244 26692
rect 6796 26648 6836 26860
rect 7276 26776 7468 26816
rect 7508 26776 7517 26816
rect 7276 26648 7316 26776
rect 8428 26732 8468 26860
rect 8524 26860 8908 26900
rect 8948 26860 8957 26900
rect 10051 26860 10060 26900
rect 10100 26860 10109 26900
rect 8524 26816 8564 26860
rect 12172 26816 12212 27028
rect 12259 26944 12268 26984
rect 12308 26944 13748 26984
rect 13097 26860 13228 26900
rect 13268 26860 13277 26900
rect 13450 26891 13516 26900
rect 13450 26851 13459 26891
rect 13499 26860 13516 26891
rect 13556 26860 13639 26900
rect 13499 26851 13508 26860
rect 13450 26850 13508 26851
rect 13708 26816 13748 26944
rect 13804 26944 13900 26984
rect 13940 26944 13949 26984
rect 15305 26944 15436 26984
rect 15476 26944 15485 26984
rect 13804 26816 13844 26944
rect 15724 26900 15764 27028
rect 25036 26984 25076 27028
rect 15811 26944 15820 26984
rect 15860 26944 17431 26984
rect 19363 26944 19372 26984
rect 19412 26944 19421 26984
rect 21475 26944 21484 26984
rect 21524 26944 25076 26984
rect 26755 26944 26764 26984
rect 26804 26944 26813 26984
rect 27017 26944 27148 26984
rect 27188 26944 27197 26984
rect 27244 26944 27724 26984
rect 27764 26944 27773 26984
rect 28649 26944 28780 26984
rect 28820 26944 28829 26984
rect 29251 26944 29260 26984
rect 29300 26944 30164 26984
rect 15724 26860 17260 26900
rect 17300 26860 17309 26900
rect 14041 26849 14081 26858
rect 8515 26776 8524 26816
rect 8564 26776 8573 26816
rect 8659 26776 8668 26816
rect 8708 26776 8812 26816
rect 8852 26776 8861 26816
rect 8995 26776 9004 26816
rect 9044 26776 9196 26816
rect 9236 26776 9245 26816
rect 9737 26776 9868 26816
rect 9908 26776 9917 26816
rect 10234 26776 10243 26816
rect 10292 26776 10423 26816
rect 12172 26776 13036 26816
rect 13076 26776 13085 26816
rect 13193 26776 13324 26816
rect 13364 26776 13373 26816
rect 13552 26776 13561 26816
rect 13601 26776 13610 26816
rect 13699 26776 13708 26816
rect 13748 26776 13757 26816
rect 13804 26776 13830 26816
rect 13870 26776 13879 26816
rect 13936 26776 13945 26816
rect 13985 26776 13994 26816
rect 15916 26816 15956 26860
rect 17391 26858 17431 26944
rect 19372 26900 19412 26944
rect 26764 26900 26804 26944
rect 27244 26900 27284 26944
rect 18211 26860 18220 26900
rect 18260 26860 18269 26900
rect 18460 26860 18796 26900
rect 18836 26860 18845 26900
rect 19363 26860 19372 26900
rect 19412 26860 19459 26900
rect 19651 26860 19660 26900
rect 19700 26860 20756 26900
rect 17373 26818 17382 26858
rect 17422 26818 17431 26858
rect 18220 26816 18260 26860
rect 18460 26858 18500 26860
rect 18457 26849 18500 26858
rect 13570 26732 13610 26776
rect 13948 26732 13988 26776
rect 14041 26774 14081 26809
rect 14314 26776 14323 26816
rect 14363 26776 14420 26816
rect 14563 26776 14572 26816
rect 14612 26776 14621 26816
rect 14754 26776 14763 26816
rect 14803 26776 14812 26816
rect 14969 26776 15052 26816
rect 15092 26776 15100 26816
rect 15140 26776 15149 26816
rect 15234 26776 15243 26816
rect 15283 26776 15340 26816
rect 15380 26776 15423 26816
rect 15715 26776 15724 26816
rect 15764 26776 15773 26816
rect 15907 26776 15916 26816
rect 15956 26776 15965 26816
rect 16771 26776 16780 26816
rect 16820 26776 16876 26816
rect 16916 26776 17260 26816
rect 17300 26776 17309 26816
rect 17500 26776 17509 26816
rect 17588 26776 17689 26816
rect 17918 26776 18028 26816
rect 18080 26776 18098 26816
rect 18173 26776 18217 26816
rect 18257 26776 18266 26816
rect 18333 26776 18342 26816
rect 18382 26776 18391 26816
rect 18497 26818 18500 26849
rect 18796 26816 18836 26860
rect 18940 26816 18980 26825
rect 19180 26816 19220 26825
rect 18457 26800 18497 26809
rect 18547 26776 18556 26816
rect 18596 26776 18644 26816
rect 18796 26776 18805 26816
rect 18845 26776 18883 26816
rect 19066 26776 19075 26816
rect 19115 26776 19124 26816
rect 14041 26734 14092 26774
rect 14132 26734 14141 26774
rect 14380 26732 14420 26776
rect 7948 26692 8140 26732
rect 8180 26692 8323 26732
rect 8363 26692 8372 26732
rect 8428 26692 12980 26732
rect 13507 26692 13516 26732
rect 13556 26692 13610 26732
rect 13891 26692 13900 26732
rect 13940 26692 13988 26732
rect 14220 26692 14284 26732
rect 14324 26692 14420 26732
rect 14572 26732 14612 26776
rect 14572 26692 14668 26732
rect 14708 26692 14717 26732
rect 3130 26608 3139 26648
rect 3179 26608 3188 26648
rect 3977 26608 4108 26648
rect 4148 26608 4157 26648
rect 4204 26608 6836 26648
rect 7267 26608 7276 26648
rect 7316 26608 7325 26648
rect 3148 26564 3188 26608
rect 7948 26564 7988 26692
rect 12940 26648 12980 26692
rect 8035 26608 8044 26648
rect 8084 26608 8140 26648
rect 8180 26608 8215 26648
rect 8323 26608 8332 26648
rect 8372 26608 8620 26648
rect 8660 26608 8669 26648
rect 8716 26608 12172 26648
rect 12212 26608 12221 26648
rect 12355 26608 12364 26648
rect 12404 26608 12413 26648
rect 12940 26608 13228 26648
rect 13268 26608 13277 26648
rect 13411 26608 13420 26648
rect 13460 26608 13804 26648
rect 13844 26608 14092 26648
rect 14132 26608 14141 26648
rect 8716 26564 8756 26608
rect 12364 26564 12404 26608
rect 14380 26564 14420 26692
rect 14537 26608 14572 26648
rect 14612 26608 14668 26648
rect 14708 26608 14717 26648
rect 3148 26524 6700 26564
rect 6740 26524 6749 26564
rect 6796 26524 7988 26564
rect 8611 26524 8620 26564
rect 8660 26524 8756 26564
rect 11107 26524 11116 26564
rect 11156 26524 12404 26564
rect 12931 26524 12940 26564
rect 12980 26524 14420 26564
rect 6796 26480 6836 26524
rect 14764 26480 14804 26776
rect 15724 26732 15764 26776
rect 18351 26732 18391 26776
rect 18604 26732 18644 26776
rect 18940 26732 18980 26776
rect 14851 26692 14860 26732
rect 14900 26692 15580 26732
rect 15620 26692 15629 26732
rect 15724 26692 17644 26732
rect 17684 26692 17693 26732
rect 18304 26692 18316 26732
rect 18356 26692 18391 26732
rect 18595 26692 18604 26732
rect 18644 26692 18980 26732
rect 15724 26648 15764 26692
rect 19084 26648 19124 26776
rect 15134 26608 15148 26648
rect 15188 26608 15197 26648
rect 15427 26608 15436 26648
rect 15476 26608 15764 26648
rect 16457 26608 16588 26648
rect 16628 26608 16637 26648
rect 16762 26608 16771 26648
rect 16811 26608 16820 26648
rect 17059 26608 17068 26648
rect 17108 26608 17356 26648
rect 17396 26608 17405 26648
rect 17866 26608 17875 26648
rect 17915 26608 17924 26648
rect 18595 26608 18604 26648
rect 18644 26608 18653 26648
rect 18883 26608 18892 26648
rect 18932 26608 19124 26648
rect 19433 26776 19564 26816
rect 19604 26776 19613 26816
rect 20227 26776 20236 26816
rect 20276 26776 20428 26816
rect 20468 26776 20477 26816
rect 20611 26776 20620 26816
rect 20660 26776 20669 26816
rect 4343 26440 4352 26480
rect 4720 26440 4729 26480
rect 6787 26440 6796 26480
rect 6836 26440 6845 26480
rect 7171 26440 7180 26480
rect 7220 26440 9484 26480
rect 9524 26440 9533 26480
rect 9667 26440 9676 26480
rect 9716 26440 9964 26480
rect 10004 26440 10100 26480
rect 12117 26440 12126 26480
rect 12494 26440 12503 26480
rect 14755 26440 14764 26480
rect 14804 26440 14813 26480
rect 10060 26396 10100 26440
rect 15134 26396 15174 26608
rect 16780 26564 16820 26608
rect 16106 26524 16820 26564
rect 16106 26396 16146 26524
rect 17884 26480 17924 26608
rect 18604 26564 18644 26608
rect 19180 26564 19220 26776
rect 20620 26732 20660 26776
rect 20419 26692 20428 26732
rect 20468 26692 20660 26732
rect 20716 26732 20756 26860
rect 22263 26860 23020 26900
rect 23060 26860 23069 26900
rect 23308 26860 23692 26900
rect 23732 26860 24940 26900
rect 24980 26860 24989 26900
rect 26275 26860 26284 26900
rect 26324 26860 26333 26900
rect 26764 26860 27284 26900
rect 28387 26860 28396 26900
rect 28436 26860 28472 26900
rect 29225 26860 29356 26900
rect 29396 26860 29405 26900
rect 29539 26860 29548 26900
rect 29588 26860 29684 26900
rect 29923 26860 29932 26900
rect 29972 26860 30008 26900
rect 22263 26816 22303 26860
rect 23308 26816 23348 26860
rect 26942 26816 26982 26860
rect 28396 26816 28436 26860
rect 29644 26816 29684 26860
rect 29932 26816 29972 26860
rect 30124 26816 30164 26944
rect 30281 26860 30316 26900
rect 30356 26860 30412 26900
rect 30452 26860 30461 26900
rect 30604 26816 30644 27196
rect 30892 26900 30932 27280
rect 31075 26944 31084 26984
rect 31124 26944 31133 26984
rect 30883 26860 30892 26900
rect 30932 26860 30941 26900
rect 31084 26816 31124 26944
rect 20803 26776 20812 26816
rect 20852 26776 20983 26816
rect 22263 26776 22300 26816
rect 22340 26776 22349 26816
rect 23299 26776 23308 26816
rect 23348 26776 23357 26816
rect 24163 26776 24172 26816
rect 24212 26776 24221 26816
rect 26284 26776 26371 26816
rect 26411 26776 26420 26816
rect 26933 26776 26942 26816
rect 26982 26776 26991 26816
rect 27043 26776 27052 26816
rect 27092 26776 27101 26816
rect 27245 26776 27254 26816
rect 27294 26776 27356 26816
rect 27418 26776 27427 26816
rect 27467 26776 27476 26816
rect 27593 26776 27724 26816
rect 27764 26776 27773 26816
rect 27895 26776 27904 26816
rect 27956 26776 28084 26816
rect 28376 26776 28385 26816
rect 28425 26776 28436 26816
rect 28492 26776 28588 26816
rect 28628 26776 28637 26816
rect 28963 26776 28972 26816
rect 29012 26776 29548 26816
rect 29588 26776 29597 26816
rect 29644 26813 29780 26816
rect 29644 26776 29733 26813
rect 24172 26732 24212 26776
rect 20716 26692 21964 26732
rect 22004 26692 24451 26732
rect 24491 26692 24500 26732
rect 26284 26648 26324 26776
rect 26371 26692 26380 26732
rect 26420 26692 26755 26732
rect 26795 26692 26804 26732
rect 20227 26608 20236 26648
rect 20276 26608 20407 26648
rect 21091 26608 21100 26648
rect 21140 26608 22444 26648
rect 22484 26608 22493 26648
rect 22627 26608 22636 26648
rect 22676 26608 22807 26648
rect 26284 26608 26764 26648
rect 26804 26608 26813 26648
rect 18604 26524 19084 26564
rect 19124 26524 19133 26564
rect 19180 26524 20372 26564
rect 19180 26480 19220 26524
rect 20332 26480 20372 26524
rect 27052 26480 27092 26776
rect 27316 26732 27356 26776
rect 27235 26692 27244 26732
rect 27284 26692 27356 26732
rect 27436 26732 27476 26776
rect 27436 26692 27628 26732
rect 27668 26692 27956 26732
rect 28051 26692 28060 26732
rect 28100 26692 28300 26732
rect 28340 26692 28349 26732
rect 27916 26648 27956 26692
rect 28492 26648 28532 26776
rect 29724 26773 29733 26776
rect 29773 26773 29782 26813
rect 29912 26776 29921 26816
rect 29961 26776 29972 26816
rect 30115 26776 30124 26816
rect 30164 26776 30173 26816
rect 30307 26776 30316 26816
rect 30356 26776 30365 26816
rect 30412 26776 30508 26816
rect 30548 26776 30557 26816
rect 30604 26776 31124 26816
rect 30316 26732 30356 26776
rect 29836 26692 30356 26732
rect 29836 26648 29876 26692
rect 30412 26648 30452 26776
rect 27916 26608 28204 26648
rect 28244 26608 28253 26648
rect 28387 26608 28396 26648
rect 28436 26608 28445 26648
rect 28492 26608 29876 26648
rect 29923 26608 29932 26648
rect 29972 26608 29981 26648
rect 30115 26608 30124 26648
rect 30164 26608 30652 26648
rect 30692 26608 30701 26648
rect 28396 26480 28436 26608
rect 17884 26440 18988 26480
rect 19028 26440 19220 26480
rect 19891 26440 19900 26480
rect 20268 26440 20277 26480
rect 20332 26440 20524 26480
rect 20564 26440 21676 26480
rect 21716 26440 21725 26480
rect 24652 26440 27092 26480
rect 27427 26440 27436 26480
rect 27476 26440 27572 26480
rect 27665 26440 27674 26480
rect 28042 26440 28051 26480
rect 28387 26440 28396 26480
rect 28436 26440 28445 26480
rect 2860 26356 5644 26396
rect 5684 26356 5693 26396
rect 10060 26356 11828 26396
rect 11788 26312 11828 26356
rect 13612 26356 14476 26396
rect 14516 26356 14525 26396
rect 14638 26356 15174 26396
rect 15331 26356 15340 26396
rect 15380 26356 16146 26396
rect 16387 26356 16396 26396
rect 16436 26356 22924 26396
rect 22964 26356 22973 26396
rect 2860 26272 3532 26312
rect 3572 26272 3581 26312
rect 4867 26272 4876 26312
rect 4916 26272 5164 26312
rect 5204 26272 5213 26312
rect 6211 26272 6220 26312
rect 6260 26272 6892 26312
rect 6932 26272 6941 26312
rect 7363 26272 7372 26312
rect 7412 26272 11212 26312
rect 11252 26272 11261 26312
rect 11770 26272 11779 26312
rect 11819 26272 11828 26312
rect 11875 26272 11884 26312
rect 11924 26272 12163 26312
rect 12203 26272 13516 26312
rect 13556 26272 13565 26312
rect 2860 26228 2900 26272
rect 1123 26188 1132 26228
rect 1172 26188 2188 26228
rect 2228 26188 2237 26228
rect 2284 26188 2900 26228
rect 3427 26188 3436 26228
rect 3476 26188 6028 26228
rect 6068 26188 6077 26228
rect 6124 26188 6412 26228
rect 6452 26188 6461 26228
rect 7171 26188 7180 26228
rect 7220 26188 12787 26228
rect 12827 26188 12940 26228
rect 12980 26188 12996 26228
rect 13108 26188 13132 26228
rect 13172 26188 13181 26228
rect 2284 26144 2324 26188
rect 5932 26144 5972 26188
rect 6124 26144 6164 26188
rect 521 26104 652 26144
rect 692 26104 701 26144
rect 826 26104 835 26144
rect 884 26104 1015 26144
rect 1357 26104 1366 26144
rect 1406 26104 1420 26144
rect 1460 26104 1546 26144
rect 1795 26104 1804 26144
rect 1844 26104 1987 26144
rect 2027 26104 2036 26144
rect 2275 26104 2284 26144
rect 2324 26104 2333 26144
rect 2380 26104 2471 26144
rect 2511 26104 2520 26144
rect 2658 26104 2667 26144
rect 2707 26104 2860 26144
rect 2900 26104 2909 26144
rect 3226 26104 3235 26144
rect 3275 26104 4204 26144
rect 4244 26104 4628 26144
rect 5631 26104 5740 26144
rect 5780 26104 5782 26144
rect 5822 26104 5876 26144
rect 5923 26104 5932 26144
rect 5972 26104 5981 26144
rect 6106 26104 6115 26144
rect 6155 26104 6164 26144
rect 6211 26104 6220 26144
rect 6260 26104 6796 26144
rect 6836 26104 6845 26144
rect 7075 26104 7084 26144
rect 7124 26104 7604 26144
rect 7747 26104 7756 26144
rect 7796 26104 7948 26144
rect 7988 26104 7997 26144
rect 8044 26104 8236 26144
rect 8276 26104 8284 26144
rect 8324 26104 8333 26144
rect 8419 26104 8428 26144
rect 8468 26104 8524 26144
rect 8564 26104 8599 26144
rect 9283 26104 9292 26144
rect 9332 26104 9388 26144
rect 9428 26104 9524 26144
rect 9763 26104 9772 26144
rect 9812 26104 9859 26144
rect 9899 26104 9943 26144
rect 10409 26104 10540 26144
rect 10580 26104 10589 26144
rect 10985 26104 11062 26144
rect 11102 26104 11116 26144
rect 11156 26104 11165 26144
rect 11273 26104 11308 26144
rect 11348 26104 11404 26144
rect 11444 26104 11453 26144
rect 11536 26104 11545 26144
rect 11585 26104 11594 26144
rect 11674 26104 11683 26144
rect 11732 26104 11863 26144
rect 11985 26104 11994 26144
rect 12034 26104 12212 26144
rect 12259 26104 12268 26144
rect 12308 26104 12439 26144
rect 12835 26104 12844 26144
rect 12884 26104 12952 26144
rect 12992 26104 13015 26144
rect 2380 26060 2420 26104
rect 4588 26060 4628 26104
rect 931 26020 940 26060
rect 980 26020 1171 26060
rect 1211 26020 1996 26060
rect 2036 26020 2045 26060
rect 2380 26020 2476 26060
rect 2516 26020 2525 26060
rect 2851 26020 2860 26060
rect 2900 26020 2909 26060
rect 3619 26020 3628 26060
rect 3668 26020 3677 26060
rect 4588 26020 5587 26060
rect 5627 26020 5636 26060
rect 2860 25976 2900 26020
rect 826 25936 835 25976
rect 875 25936 1612 25976
rect 1652 25936 1661 25976
rect 1795 25936 1804 25976
rect 1844 25936 2284 25976
rect 2324 25936 2333 25976
rect 2537 25936 2659 25976
rect 2708 25936 2717 25976
rect 2764 25936 2900 25976
rect 5836 25976 5876 26104
rect 7084 26060 7124 26104
rect 6403 26020 6412 26060
rect 6452 26020 7124 26060
rect 7564 26060 7604 26104
rect 8044 26060 8084 26104
rect 9484 26060 9524 26104
rect 11554 26060 11594 26104
rect 7564 26020 8084 26060
rect 8131 26020 8140 26060
rect 8180 26020 9298 26060
rect 9338 26020 9347 26060
rect 9484 26020 10867 26060
rect 10907 26020 11348 26060
rect 5836 25936 11212 25976
rect 11252 25936 11261 25976
rect 2764 25892 2804 25936
rect 11308 25892 11348 26020
rect 11434 26051 11492 26060
rect 11434 26011 11443 26051
rect 11483 26011 11492 26051
rect 11554 26020 11788 26060
rect 11828 26020 11837 26060
rect 11434 26010 11492 26011
rect 11452 25976 11492 26010
rect 12172 25976 12212 26104
rect 13108 26102 13148 26188
rect 13612 26144 13652 26356
rect 14638 26312 14678 26356
rect 14179 26272 14188 26312
rect 14228 26272 14678 26312
rect 14825 26272 14947 26312
rect 14996 26272 15997 26312
rect 16052 26272 16061 26312
rect 13891 26188 13900 26228
rect 13940 26188 13998 26228
rect 13958 26144 13998 26188
rect 14380 26188 14476 26228
rect 14516 26188 14525 26228
rect 14380 26144 14420 26188
rect 14638 26144 14678 26272
rect 15153 26188 15162 26228
rect 15202 26188 15532 26228
rect 15572 26188 15581 26228
rect 15715 26188 15724 26228
rect 15764 26188 15860 26228
rect 15820 26144 15860 26188
rect 16106 26144 16146 26356
rect 24652 26312 24692 26440
rect 27532 26396 27572 26440
rect 28492 26396 28532 26608
rect 29932 26564 29972 26608
rect 29347 26524 29356 26564
rect 29396 26524 29972 26564
rect 29155 26440 29164 26480
rect 29204 26440 30316 26480
rect 30356 26440 30365 26480
rect 25123 26356 25132 26396
rect 25172 26356 27476 26396
rect 27532 26356 28532 26396
rect 17530 26272 17539 26312
rect 17579 26272 17588 26312
rect 18473 26272 18604 26312
rect 18644 26272 19084 26312
rect 19124 26272 19133 26312
rect 19267 26272 19276 26312
rect 19316 26272 19948 26312
rect 19988 26272 19997 26312
rect 21091 26272 21100 26312
rect 21140 26272 24460 26312
rect 24500 26272 24509 26312
rect 24643 26272 24652 26312
rect 24692 26272 24701 26312
rect 17548 26228 17588 26272
rect 17033 26188 17164 26228
rect 17204 26188 17213 26228
rect 17260 26188 17588 26228
rect 17705 26188 17740 26228
rect 17780 26188 17789 26228
rect 17884 26188 18316 26228
rect 18356 26188 18452 26228
rect 13289 26104 13399 26144
rect 13460 26104 13469 26144
rect 13546 26104 13555 26144
rect 13595 26104 13652 26144
rect 13721 26104 13804 26144
rect 13844 26135 13892 26144
rect 13844 26104 13852 26135
rect 13075 26062 13084 26102
rect 13124 26062 13148 26102
rect 13956 26104 13965 26144
rect 14005 26104 14014 26144
rect 14083 26104 14092 26144
rect 14132 26104 14188 26144
rect 14228 26104 14263 26144
rect 14371 26104 14380 26144
rect 14420 26104 14429 26144
rect 14620 26104 14629 26144
rect 14669 26104 14678 26144
rect 14842 26104 14851 26144
rect 14900 26104 15031 26144
rect 15209 26104 15340 26144
rect 15380 26104 15389 26144
rect 15497 26104 15532 26144
rect 15572 26104 15628 26144
rect 15668 26104 15677 26144
rect 15754 26104 15763 26144
rect 15803 26104 15860 26144
rect 16090 26104 16099 26144
rect 16139 26104 16148 26144
rect 16195 26104 16204 26144
rect 16244 26104 16375 26144
rect 16745 26104 16867 26144
rect 16916 26104 16925 26144
rect 13852 26086 13892 26095
rect 14510 26062 14519 26102
rect 14559 26062 14569 26102
rect 16204 26086 16244 26095
rect 14529 26060 14569 26062
rect 13219 26020 13228 26060
rect 13268 26020 13791 26060
rect 14529 26020 15436 26060
rect 15476 26020 15485 26060
rect 16675 26020 16684 26060
rect 16724 26020 16733 26060
rect 13751 25976 13791 26020
rect 16684 25976 16724 26020
rect 11452 25936 12076 25976
rect 12116 25936 12125 25976
rect 12172 25936 12460 25976
rect 12500 25936 13076 25976
rect 13219 25936 13228 25976
rect 13268 25936 13324 25976
rect 13364 25936 13399 25976
rect 13751 25936 15188 25976
rect 16483 25936 16492 25976
rect 16532 25936 16724 25976
rect 16876 25976 16916 26104
rect 17260 26060 17300 26188
rect 17740 26144 17780 26188
rect 17347 26104 17356 26144
rect 17396 26104 17468 26144
rect 17428 26093 17468 26104
rect 17508 26093 17517 26133
rect 17640 26104 17649 26144
rect 17689 26104 17698 26144
rect 17740 26104 17752 26144
rect 17792 26104 17801 26144
rect 17884 26135 17924 26188
rect 18412 26144 18452 26188
rect 18556 26144 18596 26272
rect 18892 26188 22156 26228
rect 22196 26188 22205 26228
rect 22263 26188 22636 26228
rect 22676 26188 22685 26228
rect 22732 26188 22828 26228
rect 22868 26188 22877 26228
rect 23002 26188 23011 26228
rect 23051 26188 23308 26228
rect 23348 26188 23357 26228
rect 23404 26188 26476 26228
rect 26516 26188 26525 26228
rect 26659 26188 26668 26228
rect 26708 26188 27092 26228
rect 18892 26144 18932 26188
rect 22263 26146 22303 26188
rect 17649 26060 17689 26104
rect 18010 26104 18019 26144
rect 18068 26104 18199 26144
rect 18403 26104 18412 26144
rect 18452 26104 18461 26144
rect 18538 26104 18547 26144
rect 18587 26104 18596 26144
rect 18652 26104 18661 26144
rect 18701 26104 18932 26144
rect 18979 26104 18988 26144
rect 19028 26104 19159 26144
rect 19267 26104 19276 26144
rect 19350 26104 19447 26144
rect 20131 26104 20140 26144
rect 20180 26104 20236 26144
rect 20276 26104 20311 26144
rect 20419 26104 20428 26144
rect 20468 26104 20477 26144
rect 21161 26104 21259 26144
rect 21332 26104 21341 26144
rect 21667 26104 21676 26144
rect 21739 26104 21847 26144
rect 22245 26106 22254 26146
rect 22294 26106 22303 26146
rect 22732 26144 22772 26188
rect 23404 26144 23444 26188
rect 27052 26144 27092 26188
rect 27436 26144 27476 26356
rect 28492 26312 28532 26356
rect 28099 26272 28108 26312
rect 28148 26272 28436 26312
rect 28492 26272 29204 26312
rect 29731 26272 29740 26312
rect 29780 26272 30316 26312
rect 30356 26272 30365 26312
rect 30473 26272 30604 26312
rect 30644 26272 30653 26312
rect 30857 26272 30988 26312
rect 31028 26272 31037 26312
rect 28396 26228 28436 26272
rect 27523 26188 27532 26228
rect 27572 26188 27806 26228
rect 27846 26188 27855 26228
rect 27907 26188 27916 26228
rect 27956 26188 28012 26228
rect 28052 26188 28087 26228
rect 28396 26188 28724 26228
rect 28771 26188 28780 26228
rect 28820 26188 28829 26228
rect 28963 26188 28972 26228
rect 29012 26188 29021 26228
rect 28684 26144 28724 26188
rect 28780 26144 28820 26188
rect 28972 26144 29012 26188
rect 29164 26144 29204 26272
rect 22378 26104 22387 26144
rect 22427 26104 22444 26144
rect 22484 26104 22567 26144
rect 22708 26104 22772 26144
rect 22916 26104 22925 26144
rect 22965 26104 23020 26144
rect 23060 26104 23096 26144
rect 23386 26104 23395 26144
rect 23435 26104 23444 26144
rect 23491 26104 23500 26144
rect 23540 26104 23596 26144
rect 23636 26104 23671 26144
rect 23971 26104 23980 26144
rect 24020 26104 25460 26144
rect 26633 26104 26755 26144
rect 26804 26104 26813 26144
rect 27052 26104 27304 26144
rect 27344 26104 27353 26144
rect 27418 26104 27427 26144
rect 27467 26104 27476 26144
rect 27523 26104 27532 26144
rect 27572 26104 27628 26144
rect 27668 26104 27703 26144
rect 28108 26135 28148 26144
rect 17884 26060 17924 26095
rect 18700 26060 18740 26104
rect 20428 26060 20468 26104
rect 22708 26102 22748 26104
rect 21562 26062 21571 26102
rect 21611 26062 21620 26102
rect 22675 26062 22684 26102
rect 22724 26062 22748 26102
rect 17251 26020 17260 26060
rect 17300 26020 17309 26060
rect 17602 26020 17644 26060
rect 17684 26020 17693 26060
rect 17827 26020 17836 26060
rect 17876 26020 17924 26060
rect 18307 26020 18316 26060
rect 18356 26020 18740 26060
rect 18787 26020 18796 26060
rect 18836 26051 19359 26060
rect 18836 26020 19219 26051
rect 19210 26011 19219 26020
rect 19259 26020 19359 26051
rect 19747 26020 19756 26060
rect 19796 26020 20468 26060
rect 20707 26020 20716 26060
rect 20756 26020 21388 26060
rect 21428 26020 21437 26060
rect 19259 26011 19268 26020
rect 19210 26010 19268 26011
rect 19319 25976 19359 26020
rect 21580 25976 21620 26062
rect 22810 26020 22819 26060
rect 22859 26020 23156 26060
rect 24713 26020 24835 26060
rect 24884 26020 24893 26060
rect 23116 25976 23156 26020
rect 16876 25936 18644 25976
rect 18883 25936 18892 25976
rect 18932 25936 19084 25976
rect 19124 25936 19133 25976
rect 19319 25936 19660 25976
rect 19700 25936 20044 25976
rect 20084 25936 20093 25976
rect 21353 25936 21484 25976
rect 21524 25936 21533 25976
rect 21580 25936 21676 25976
rect 21716 25936 21725 25976
rect 23107 25936 23116 25976
rect 23156 25936 23165 25976
rect 23561 25936 23683 25976
rect 23732 25936 23741 25976
rect 2476 25852 2804 25892
rect 6089 25852 6220 25892
rect 6260 25852 6269 25892
rect 6403 25852 6412 25892
rect 6452 25852 6461 25892
rect 7145 25852 7276 25892
rect 7316 25852 7325 25892
rect 8314 25852 8323 25892
rect 8363 25852 8524 25892
rect 8564 25852 8573 25892
rect 9065 25852 9196 25892
rect 9236 25852 9245 25892
rect 11308 25852 11692 25892
rect 11732 25852 11741 25892
rect 11849 25852 11980 25892
rect 12020 25852 12029 25892
rect 2476 25556 2516 25852
rect 6412 25808 6452 25852
rect 13036 25808 13076 25936
rect 15148 25892 15188 25936
rect 18604 25892 18644 25936
rect 25420 25892 25460 26104
rect 28291 26104 28300 26144
rect 28340 26104 28349 26144
rect 28483 26104 28492 26144
rect 28532 26104 28541 26144
rect 28675 26104 28684 26144
rect 28724 26104 28733 26144
rect 28780 26104 28876 26144
rect 28916 26104 28925 26144
rect 28972 26104 29069 26144
rect 29109 26104 29118 26144
rect 29164 26104 29260 26144
rect 29300 26104 29309 26144
rect 29443 26104 29452 26144
rect 29492 26104 29501 26144
rect 29633 26104 29642 26144
rect 29684 26104 29813 26144
rect 30211 26104 30220 26144
rect 30260 26104 30269 26144
rect 30403 26104 30412 26144
rect 30452 26104 30583 26144
rect 28108 26060 28148 26095
rect 26947 26020 26956 26060
rect 26996 26020 27005 26060
rect 27130 26020 27139 26060
rect 27188 26020 27319 26060
rect 27619 26020 27628 26060
rect 27668 26020 27724 26060
rect 27764 26020 27799 26060
rect 28003 26020 28012 26060
rect 28052 26020 28148 26060
rect 28300 26060 28340 26104
rect 28492 26060 28532 26104
rect 29452 26060 29492 26104
rect 28300 26020 28436 26060
rect 28492 26020 28684 26060
rect 28724 26020 28733 26060
rect 29347 26020 29356 26060
rect 29396 26020 29492 26060
rect 29897 26020 30028 26060
rect 30068 26020 30077 26060
rect 27907 25936 27916 25976
rect 27956 25936 28300 25976
rect 28340 25936 28349 25976
rect 13795 25852 13804 25892
rect 13844 25852 13900 25892
rect 13940 25852 13975 25892
rect 14057 25852 14092 25892
rect 14132 25852 14188 25892
rect 14228 25852 14237 25892
rect 14467 25852 14476 25892
rect 14516 25852 14572 25892
rect 14612 25852 14647 25892
rect 15139 25852 15148 25892
rect 15188 25852 15197 25892
rect 15305 25852 15340 25892
rect 15380 25852 15436 25892
rect 15476 25852 15485 25892
rect 15859 25852 15868 25892
rect 15908 25852 16396 25892
rect 16436 25852 16445 25892
rect 18377 25852 18508 25892
rect 18548 25852 18557 25892
rect 18604 25852 19747 25892
rect 19787 25852 20620 25892
rect 20660 25852 20669 25892
rect 22426 25852 22435 25892
rect 22475 25852 25132 25892
rect 25172 25852 25181 25892
rect 25420 25852 27811 25892
rect 27851 25852 27860 25892
rect 28396 25808 28436 26020
rect 28579 25936 28588 25976
rect 28628 25936 28724 25976
rect 29443 25936 29452 25976
rect 29492 25936 29788 25976
rect 29828 25936 29837 25976
rect 28684 25892 28724 25936
rect 30220 25892 30260 26104
rect 28675 25852 28684 25892
rect 28724 25852 28733 25892
rect 28867 25852 28876 25892
rect 28916 25852 29164 25892
rect 29204 25852 29213 25892
rect 29417 25852 29452 25892
rect 29492 25852 29548 25892
rect 29588 25852 29597 25892
rect 30019 25852 30028 25892
rect 30068 25852 30260 25892
rect 2860 25768 6452 25808
rect 8803 25768 8812 25808
rect 8852 25768 12980 25808
rect 13036 25768 14860 25808
rect 14900 25768 14909 25808
rect 17731 25768 17740 25808
rect 17780 25768 24268 25808
rect 24308 25768 24317 25808
rect 24748 25768 27764 25808
rect 27907 25768 27916 25808
rect 27956 25768 28436 25808
rect 28579 25768 28588 25808
rect 28628 25768 30548 25808
rect 2467 25516 2476 25556
rect 2516 25516 2525 25556
rect 2860 25472 2900 25768
rect 3103 25684 3112 25724
rect 3480 25684 3489 25724
rect 6787 25684 6796 25724
rect 6836 25684 10100 25724
rect 10877 25684 10886 25724
rect 11254 25684 11263 25724
rect 6691 25600 6700 25640
rect 6740 25600 10004 25640
rect 3401 25516 3436 25556
rect 3476 25516 3532 25556
rect 3572 25516 3581 25556
rect 4675 25516 4684 25556
rect 4724 25516 4972 25556
rect 5012 25516 5021 25556
rect 5452 25516 6412 25556
rect 6452 25516 6461 25556
rect 7756 25516 9100 25556
rect 9140 25516 9908 25556
rect 5452 25472 5492 25516
rect 2188 25432 2900 25472
rect 2956 25432 4244 25472
rect 4867 25432 4876 25472
rect 4916 25432 5492 25472
rect 1027 25348 1036 25388
rect 1076 25348 1123 25388
rect 1036 25304 1076 25348
rect 2188 25304 2228 25432
rect 2956 25388 2996 25432
rect 4204 25388 4244 25432
rect 2668 25348 2996 25388
rect 3052 25348 4108 25388
rect 4148 25348 4157 25388
rect 4204 25348 5260 25388
rect 5300 25348 5309 25388
rect 6979 25348 6988 25388
rect 7028 25348 7037 25388
rect 713 25264 844 25304
rect 884 25264 893 25304
rect 1018 25264 1027 25304
rect 1067 25264 1076 25304
rect 1123 25264 1132 25304
rect 1172 25264 1303 25304
rect 1987 25264 1996 25304
rect 2036 25264 2045 25304
rect 2179 25264 2188 25304
rect 2228 25264 2237 25304
rect 1996 25220 2036 25264
rect 922 25180 931 25220
rect 971 25180 2036 25220
rect 2668 25220 2708 25348
rect 3052 25304 3092 25348
rect 7756 25304 7796 25516
rect 9868 25388 9908 25516
rect 9292 25348 9580 25388
rect 9620 25348 9629 25388
rect 9850 25348 9859 25388
rect 9899 25348 9908 25388
rect 9292 25304 9332 25348
rect 9964 25304 10004 25600
rect 10060 25388 10100 25684
rect 12940 25640 12980 25768
rect 18651 25684 18660 25724
rect 19028 25684 19037 25724
rect 20131 25684 20140 25724
rect 20180 25684 20908 25724
rect 20948 25684 20957 25724
rect 24748 25640 24788 25768
rect 26425 25684 26434 25724
rect 26802 25684 26811 25724
rect 12940 25600 14036 25640
rect 10915 25516 10924 25556
rect 10964 25516 11404 25556
rect 11444 25516 11453 25556
rect 13306 25516 13315 25556
rect 13355 25516 13364 25556
rect 11779 25432 11788 25472
rect 11828 25432 12940 25472
rect 12980 25432 12989 25472
rect 13324 25388 13364 25516
rect 13507 25432 13516 25472
rect 13556 25432 13940 25472
rect 13900 25388 13940 25432
rect 13996 25388 14036 25600
rect 20140 25600 24788 25640
rect 27724 25640 27764 25768
rect 27724 25600 29300 25640
rect 20140 25556 20180 25600
rect 14083 25516 14092 25556
rect 14132 25516 14380 25556
rect 14420 25516 14429 25556
rect 14563 25516 14572 25556
rect 14612 25516 14764 25556
rect 14804 25516 14813 25556
rect 17452 25516 19564 25556
rect 19604 25516 19613 25556
rect 19939 25516 19948 25556
rect 19988 25516 20180 25556
rect 20873 25516 20995 25556
rect 21044 25516 21053 25556
rect 23011 25516 23020 25556
rect 23060 25516 24172 25556
rect 24212 25516 24221 25556
rect 24617 25516 24748 25556
rect 24788 25516 24797 25556
rect 24844 25516 28876 25556
rect 28916 25516 28925 25556
rect 14083 25432 14092 25472
rect 14132 25432 14476 25472
rect 14516 25432 14564 25472
rect 10060 25348 10396 25388
rect 10436 25348 10445 25388
rect 11107 25348 11116 25388
rect 11156 25348 11165 25388
rect 13027 25348 13036 25388
rect 13076 25348 13364 25388
rect 13891 25348 13900 25388
rect 13940 25348 13949 25388
rect 13996 25348 14132 25388
rect 14371 25348 14380 25388
rect 14420 25348 14429 25388
rect 11116 25304 11156 25348
rect 13612 25304 13652 25313
rect 13900 25304 13940 25348
rect 14092 25304 14132 25348
rect 14380 25304 14420 25348
rect 14524 25337 14564 25432
rect 14764 25388 14804 25516
rect 14947 25432 14956 25472
rect 14996 25432 15724 25472
rect 15764 25432 15773 25472
rect 15898 25432 15907 25472
rect 15947 25432 17396 25472
rect 17356 25388 17396 25432
rect 14764 25348 15668 25388
rect 16867 25348 16876 25388
rect 16916 25348 17227 25388
rect 17338 25348 17347 25388
rect 17387 25348 17396 25388
rect 2860 25295 3092 25304
rect 2900 25264 3092 25295
rect 3139 25264 3148 25304
rect 3188 25264 3319 25304
rect 4099 25264 4108 25304
rect 4148 25264 4195 25304
rect 4378 25264 4387 25304
rect 4427 25264 4436 25304
rect 4483 25264 4492 25304
rect 4532 25264 6604 25304
rect 6644 25264 6653 25304
rect 6778 25264 6787 25304
rect 6827 25299 6932 25304
rect 7084 25299 7180 25304
rect 6827 25264 7180 25299
rect 7220 25264 7229 25304
rect 7363 25264 7372 25304
rect 7412 25264 7543 25304
rect 7747 25264 7756 25304
rect 7796 25264 7805 25304
rect 8803 25264 8812 25304
rect 8852 25264 8861 25304
rect 9017 25264 9100 25304
rect 9140 25264 9148 25304
rect 9188 25264 9197 25304
rect 9283 25264 9292 25304
rect 9332 25264 9341 25304
rect 9484 25264 9719 25304
rect 9759 25264 9768 25304
rect 9955 25264 9964 25304
rect 10004 25264 10013 25304
rect 10060 25264 10195 25304
rect 10235 25264 10244 25304
rect 10819 25264 10828 25304
rect 10868 25264 10877 25304
rect 11020 25264 11029 25304
rect 11069 25264 11156 25304
rect 11203 25264 11212 25304
rect 11252 25264 11404 25304
rect 11444 25264 11453 25304
rect 11683 25264 11692 25304
rect 11732 25264 11788 25304
rect 11828 25264 11863 25304
rect 11971 25264 11980 25304
rect 12020 25264 12163 25304
rect 12203 25264 12212 25304
rect 12259 25264 12268 25304
rect 12308 25264 12317 25304
rect 12617 25264 12717 25304
rect 12788 25264 12797 25304
rect 12870 25264 12879 25304
rect 12919 25264 12940 25304
rect 12980 25264 13050 25304
rect 13132 25264 13157 25304
rect 13197 25264 13310 25304
rect 13350 25264 13359 25304
rect 2860 25246 2900 25255
rect 4108 25220 4148 25264
rect 2668 25180 2764 25220
rect 2804 25180 2813 25220
rect 4099 25180 4108 25220
rect 4148 25180 4157 25220
rect 4396 25136 4436 25264
rect 6892 25259 7124 25264
rect 4689 25180 4698 25220
rect 4738 25180 6836 25220
rect 7162 25180 7171 25220
rect 7211 25180 8131 25220
rect 8171 25180 8180 25220
rect 6796 25136 6836 25180
rect 8812 25136 8852 25264
rect 9484 25220 9524 25264
rect 10060 25220 10100 25264
rect 8899 25180 8908 25220
rect 8948 25180 9524 25220
rect 9667 25180 9676 25220
rect 9716 25180 10100 25220
rect 10828 25220 10868 25264
rect 10828 25180 11404 25220
rect 11444 25180 11453 25220
rect 1315 25096 1324 25136
rect 1364 25096 1373 25136
rect 2323 25096 2332 25136
rect 2372 25096 2900 25136
rect 4396 25096 6412 25136
rect 6452 25096 6461 25136
rect 6796 25096 7084 25136
rect 7124 25096 7133 25136
rect 7721 25096 7852 25136
rect 7892 25096 7901 25136
rect 8812 25096 8948 25136
rect 9929 25096 9964 25136
rect 10004 25096 10051 25136
rect 10091 25096 10164 25136
rect 10697 25096 10828 25136
rect 10868 25096 10877 25136
rect 11177 25096 11299 25136
rect 11348 25096 11357 25136
rect 1324 24716 1364 25096
rect 2860 25052 2900 25096
rect 2860 25012 8140 25052
rect 8180 25012 8189 25052
rect 4343 24928 4352 24968
rect 4720 24928 4729 24968
rect 4108 24844 4876 24884
rect 4916 24844 4925 24884
rect 8380 24844 8716 24884
rect 8756 24844 8765 24884
rect 2083 24760 2092 24800
rect 2132 24760 2956 24800
rect 2996 24760 3340 24800
rect 3380 24760 3389 24800
rect 4108 24716 4148 24844
rect 4361 24760 4492 24800
rect 4532 24760 4541 24800
rect 7459 24760 7468 24800
rect 7508 24760 7756 24800
rect 7796 24760 7805 24800
rect 8009 24760 8140 24800
rect 8180 24760 8189 24800
rect 634 24676 643 24716
rect 683 24676 1364 24716
rect 4012 24676 4148 24716
rect 4841 24676 4876 24716
rect 4916 24676 4972 24716
rect 5012 24676 5021 24716
rect 5146 24676 5155 24716
rect 5195 24676 6796 24716
rect 6836 24676 6845 24716
rect 4012 24632 4052 24676
rect 8380 24632 8420 24844
rect 8908 24800 8948 25096
rect 12268 25052 12308 25264
rect 13132 25220 13172 25264
rect 13612 25220 13652 25264
rect 13708 25264 13804 25304
rect 13844 25264 13853 25304
rect 13900 25264 13987 25304
rect 14027 25264 14036 25304
rect 14083 25264 14092 25304
rect 14132 25301 14144 25304
rect 14275 25301 14284 25304
rect 14132 25264 14284 25301
rect 14324 25264 14333 25304
rect 14380 25264 14406 25304
rect 14446 25264 14467 25304
rect 15628 25304 15668 25348
rect 16492 25304 16532 25313
rect 14524 25288 14564 25297
rect 14746 25264 14755 25304
rect 14795 25264 14804 25304
rect 14851 25264 14860 25304
rect 14900 25264 15063 25304
rect 15103 25264 15112 25304
rect 15610 25264 15619 25304
rect 15659 25264 15668 25304
rect 15715 25264 15724 25304
rect 15764 25264 15773 25304
rect 15907 25264 15916 25304
rect 15956 25264 16396 25304
rect 16436 25264 16445 25304
rect 16649 25264 16780 25304
rect 16820 25264 16829 25304
rect 16952 25264 16972 25304
rect 17012 25264 17083 25304
rect 17123 25264 17132 25304
rect 17187 25264 17227 25348
rect 17452 25304 17492 25516
rect 24844 25472 24884 25516
rect 17836 25432 18988 25472
rect 19028 25432 19037 25472
rect 19084 25432 19852 25472
rect 19892 25432 19901 25472
rect 20131 25432 20140 25472
rect 20180 25432 20852 25472
rect 20899 25432 20908 25472
rect 20948 25432 21292 25472
rect 21332 25432 21341 25472
rect 23011 25432 23020 25472
rect 23060 25432 24884 25472
rect 24931 25432 24940 25472
rect 24980 25432 24989 25472
rect 28675 25432 28684 25472
rect 28724 25432 29204 25472
rect 17267 25264 17396 25304
rect 17443 25264 17452 25304
rect 17492 25264 17501 25304
rect 13708 25220 13748 25264
rect 14104 25261 14324 25264
rect 14764 25220 14804 25264
rect 15724 25220 15764 25264
rect 12835 25180 12844 25220
rect 12884 25180 13172 25220
rect 13315 25180 13324 25220
rect 13364 25180 13652 25220
rect 13699 25180 13708 25220
rect 13748 25180 13757 25220
rect 14371 25180 14380 25220
rect 14420 25180 14804 25220
rect 15427 25180 15436 25220
rect 15476 25180 15764 25220
rect 16073 25180 16193 25220
rect 16244 25180 16253 25220
rect 12425 25096 12556 25136
rect 12596 25096 12605 25136
rect 13132 25052 13172 25180
rect 13411 25096 13420 25136
rect 13460 25096 13516 25136
rect 13556 25096 13591 25136
rect 13891 25096 13900 25136
rect 13940 25096 14851 25136
rect 14891 25096 14900 25136
rect 14947 25096 14956 25136
rect 14996 25096 15724 25136
rect 15764 25096 15773 25136
rect 16099 25096 16108 25136
rect 16148 25096 16291 25136
rect 16331 25096 16340 25136
rect 16492 25052 16532 25264
rect 17356 25220 17396 25264
rect 17836 25220 17876 25432
rect 19084 25388 19124 25432
rect 20812 25388 20852 25432
rect 18220 25348 18604 25388
rect 18644 25348 18653 25388
rect 18892 25348 19124 25388
rect 19241 25348 19363 25388
rect 19412 25348 19421 25388
rect 19651 25348 19660 25388
rect 19700 25348 19781 25388
rect 19843 25348 19852 25388
rect 19892 25348 19901 25388
rect 20669 25348 20716 25388
rect 20756 25348 20765 25388
rect 20812 25348 21908 25388
rect 18220 25304 18260 25348
rect 18892 25304 18932 25348
rect 19741 25346 19781 25348
rect 19741 25337 19796 25346
rect 19741 25306 19756 25337
rect 17962 25264 17971 25304
rect 18011 25264 18020 25304
rect 18202 25264 18211 25304
rect 18251 25264 18260 25304
rect 18499 25264 18508 25304
rect 18548 25264 18625 25304
rect 18665 25264 18679 25304
rect 18883 25264 18892 25304
rect 18932 25264 18941 25304
rect 19092 25264 19180 25304
rect 19220 25264 19223 25304
rect 19263 25264 19272 25304
rect 19337 25264 19466 25304
rect 19508 25264 19517 25304
rect 19756 25288 19796 25297
rect 19852 25304 19892 25348
rect 20013 25337 20054 25346
rect 19852 25264 19891 25304
rect 19931 25264 19940 25304
rect 20053 25325 20054 25337
rect 20053 25297 20073 25325
rect 20716 25304 20756 25348
rect 20013 25288 20073 25297
rect 20014 25285 20073 25288
rect 17356 25180 17876 25220
rect 17980 25220 18020 25264
rect 19852 25261 19940 25264
rect 20033 25220 20073 25285
rect 20131 25264 20140 25304
rect 20180 25264 20189 25304
rect 20323 25264 20332 25304
rect 20372 25264 20381 25304
rect 20698 25264 20707 25304
rect 20747 25264 20756 25304
rect 20803 25264 20812 25304
rect 20852 25264 20908 25304
rect 20948 25264 20983 25304
rect 21161 25264 21292 25304
rect 21332 25264 21341 25304
rect 21449 25264 21484 25304
rect 21524 25264 21580 25304
rect 21620 25264 21629 25304
rect 20140 25220 20180 25264
rect 20332 25220 20372 25264
rect 17980 25180 18028 25220
rect 18068 25180 18077 25220
rect 18211 25180 18220 25220
rect 18260 25180 19220 25220
rect 19433 25180 19555 25220
rect 19604 25180 19613 25220
rect 20033 25180 20044 25220
rect 20084 25180 20093 25220
rect 20140 25180 20372 25220
rect 19180 25136 19220 25180
rect 16675 25096 16684 25136
rect 16724 25096 17539 25136
rect 17579 25096 17588 25136
rect 17635 25096 17644 25136
rect 17684 25096 18019 25136
rect 18059 25096 18068 25136
rect 18665 25096 18787 25136
rect 18836 25096 18845 25136
rect 19075 25096 19084 25136
rect 19124 25096 19133 25136
rect 19180 25096 20188 25136
rect 20228 25096 20237 25136
rect 21667 25096 21676 25136
rect 21716 25096 21725 25136
rect 12268 25012 12692 25052
rect 13132 25012 14476 25052
rect 14516 25012 15092 25052
rect 16492 25012 16724 25052
rect 12652 24968 12692 25012
rect 9091 24928 9100 24968
rect 9140 24928 11884 24968
rect 11924 24928 11933 24968
rect 12117 24928 12126 24968
rect 12494 24928 12503 24968
rect 12652 24928 13460 24968
rect 9283 24844 9292 24884
rect 9332 24844 10732 24884
rect 10772 24844 10781 24884
rect 11203 24844 11212 24884
rect 11252 24844 11980 24884
rect 12020 24844 12029 24884
rect 13420 24800 13460 24928
rect 15052 24800 15092 25012
rect 16684 24968 16724 25012
rect 16675 24928 16684 24968
rect 16724 24928 16733 24968
rect 17548 24800 17588 24809
rect 8489 24760 8524 24800
rect 8564 24760 8620 24800
rect 8660 24760 8669 24800
rect 8890 24760 8899 24800
rect 8939 24760 8948 24800
rect 9091 24760 9100 24800
rect 9140 24760 13228 24800
rect 13268 24760 13277 24800
rect 13402 24760 13411 24800
rect 13451 24760 13460 24800
rect 14755 24760 14764 24800
rect 14804 24760 14956 24800
rect 14996 24760 15005 24800
rect 15052 24760 15187 24800
rect 15227 24760 15236 24800
rect 16099 24760 16108 24800
rect 16148 24760 16157 24800
rect 17588 24760 18124 24800
rect 18164 24760 18173 24800
rect 18307 24760 18316 24800
rect 18356 24760 18508 24800
rect 18548 24760 18557 24800
rect 18665 24760 18787 24800
rect 18836 24760 18845 24800
rect 8681 24676 8801 24716
rect 8852 24676 8861 24716
rect 9100 24676 12844 24716
rect 12884 24676 12893 24716
rect 1018 24592 1027 24632
rect 1076 24592 1207 24632
rect 3628 24592 3820 24632
rect 3860 24592 3869 24632
rect 4003 24592 4012 24632
rect 4052 24592 4061 24632
rect 4265 24592 4396 24632
rect 4436 24592 4445 24632
rect 4937 24592 4972 24632
rect 5012 24592 5068 24632
rect 5108 24592 5117 24632
rect 5530 24592 5539 24632
rect 5588 24592 5719 24632
rect 6595 24592 6604 24632
rect 6644 24592 7660 24632
rect 7700 24592 7709 24632
rect 8035 24592 8044 24632
rect 8084 24592 8093 24632
rect 8380 24592 8428 24632
rect 8468 24592 8477 24632
rect 8873 24592 8908 24632
rect 8948 24592 9004 24632
rect 9044 24592 9053 24632
rect 9100 24623 9140 24676
rect 12940 24632 12980 24760
rect 16108 24716 16148 24760
rect 17548 24751 17588 24760
rect 17836 24716 17876 24760
rect 19084 24716 19124 25096
rect 19267 25012 19276 25052
rect 19316 25012 21388 25052
rect 21428 25012 21437 25052
rect 19891 24928 19900 24968
rect 20268 24928 20277 24968
rect 19267 24844 19276 24884
rect 19316 24844 21004 24884
rect 21044 24844 21053 24884
rect 19459 24760 19468 24800
rect 19508 24760 21292 24800
rect 21332 24760 21341 24800
rect 21676 24716 21716 25096
rect 21868 25052 21908 25348
rect 22348 25348 23308 25388
rect 23348 25348 23357 25388
rect 22348 25304 22388 25348
rect 24940 25304 24980 25432
rect 25289 25348 25411 25388
rect 25460 25348 25469 25388
rect 27552 25348 28588 25388
rect 28628 25348 28637 25388
rect 28867 25348 28876 25388
rect 28916 25348 29012 25388
rect 28972 25304 29012 25348
rect 29070 25304 29110 25313
rect 22339 25264 22348 25304
rect 22388 25264 22397 25304
rect 22714 25264 22723 25304
rect 22763 25264 22772 25304
rect 22818 25264 22827 25304
rect 22867 25264 22924 25304
rect 22964 25264 23007 25304
rect 23203 25264 23212 25304
rect 23252 25264 23383 25304
rect 23945 25264 24076 25304
rect 24116 25264 24125 25304
rect 24931 25264 24940 25304
rect 24980 25264 24989 25304
rect 25097 25264 25228 25304
rect 25268 25264 25277 25304
rect 27209 25264 27331 25304
rect 27380 25264 27389 25304
rect 28579 25264 28588 25304
rect 28628 25264 28916 25304
rect 28972 25264 29070 25304
rect 22732 25220 22772 25264
rect 28876 25220 28916 25264
rect 29070 25255 29110 25264
rect 22732 25180 23308 25220
rect 23348 25180 23357 25220
rect 23875 25180 23884 25220
rect 23924 25180 25996 25220
rect 26036 25180 26045 25220
rect 26092 25180 27572 25220
rect 27706 25180 27715 25220
rect 27755 25180 27907 25220
rect 27947 25180 27956 25220
rect 28099 25180 28108 25220
rect 28148 25180 28766 25220
rect 28806 25180 28815 25220
rect 28858 25180 28867 25220
rect 28907 25180 28916 25220
rect 29164 25220 29204 25432
rect 29260 25346 29300 25600
rect 29635 25516 29644 25556
rect 29684 25516 29740 25556
rect 29780 25516 29815 25556
rect 30508 25472 30548 25768
rect 29347 25432 29356 25472
rect 29396 25432 30028 25472
rect 30068 25432 30077 25472
rect 30403 25432 30412 25472
rect 30452 25432 30461 25472
rect 30508 25432 30796 25472
rect 30836 25432 30845 25472
rect 29443 25348 29452 25388
rect 29492 25348 29588 25388
rect 29251 25306 29260 25346
rect 29300 25306 29309 25346
rect 29548 25304 29588 25348
rect 29356 25264 29452 25304
rect 29492 25264 29501 25304
rect 29548 25264 29645 25304
rect 29685 25264 29694 25304
rect 29827 25264 29836 25304
rect 29876 25264 30260 25304
rect 29356 25220 29396 25264
rect 30220 25220 30260 25264
rect 29164 25180 29396 25220
rect 30211 25180 30220 25220
rect 30260 25180 30269 25220
rect 26092 25136 26132 25180
rect 22723 25096 22732 25136
rect 22772 25096 23212 25136
rect 23252 25096 23261 25136
rect 24259 25096 24268 25136
rect 24308 25096 25027 25136
rect 25067 25096 25076 25136
rect 25132 25096 26132 25136
rect 27532 25136 27572 25180
rect 30412 25136 30452 25432
rect 27532 25096 28396 25136
rect 28436 25096 28445 25136
rect 28963 25096 28972 25136
rect 29012 25096 29021 25136
rect 29347 25096 29356 25136
rect 29396 25096 29405 25136
rect 30220 25096 30452 25136
rect 25132 25052 25172 25096
rect 28972 25052 29012 25096
rect 29356 25052 29396 25096
rect 21868 25012 25172 25052
rect 28963 25012 28972 25052
rect 29012 25012 29059 25052
rect 29155 25012 29164 25052
rect 29204 25012 29396 25052
rect 30220 24968 30260 25096
rect 27665 24928 27674 24968
rect 28042 24928 28051 24968
rect 28108 24928 30260 24968
rect 28108 24884 28148 24928
rect 25315 24844 25324 24884
rect 25364 24844 28148 24884
rect 22505 24760 22588 24800
rect 22628 24760 22636 24800
rect 22676 24760 22685 24800
rect 22889 24760 23011 24800
rect 23060 24760 23069 24800
rect 25027 24760 25036 24800
rect 25076 24760 29108 24800
rect 13516 24676 14380 24716
rect 14420 24676 14429 24716
rect 14476 24676 16012 24716
rect 16052 24676 16061 24716
rect 16108 24676 16436 24716
rect 17818 24676 17827 24716
rect 17867 24676 17876 24716
rect 17932 24676 18220 24716
rect 18260 24676 19028 24716
rect 19084 24676 19508 24716
rect 19747 24676 19756 24716
rect 19796 24676 19939 24716
rect 19979 24676 19988 24716
rect 20131 24676 20140 24716
rect 20180 24676 21580 24716
rect 21620 24676 21629 24716
rect 21676 24676 22243 24716
rect 22283 24676 22292 24716
rect 22339 24676 22348 24716
rect 22388 24676 25364 24716
rect 25498 24676 25507 24716
rect 25547 24676 25804 24716
rect 25844 24676 25853 24716
rect 26074 24676 26083 24716
rect 26123 24676 27436 24716
rect 27476 24676 27485 24716
rect 13516 24632 13556 24676
rect 14092 24632 14132 24676
rect 3628 24548 3668 24592
rect 8044 24548 8084 24592
rect 8602 24550 8611 24590
rect 8651 24550 8660 24590
rect 9100 24574 9140 24583
rect 9484 24592 11212 24632
rect 11252 24592 11261 24632
rect 11369 24592 11395 24632
rect 11435 24592 11500 24632
rect 11540 24592 11549 24632
rect 11971 24592 11980 24632
rect 12020 24592 12151 24632
rect 12748 24592 12844 24632
rect 12884 24592 12893 24632
rect 12940 24592 12959 24632
rect 12999 24592 13008 24632
rect 13123 24592 13132 24632
rect 13172 24592 13324 24632
rect 13364 24592 13373 24632
rect 13507 24592 13516 24632
rect 13556 24592 13687 24632
rect 13769 24592 13900 24632
rect 13940 24592 13949 24632
rect 14083 24592 14092 24632
rect 14132 24592 14141 24632
rect 8620 24548 8660 24550
rect 9484 24548 9524 24592
rect 1699 24508 1708 24548
rect 1748 24508 1757 24548
rect 2476 24508 2900 24548
rect 3331 24508 3340 24548
rect 3380 24508 3668 24548
rect 3715 24508 3724 24548
rect 3764 24508 5376 24548
rect 8044 24508 8236 24548
rect 8276 24508 8428 24548
rect 8468 24508 8477 24548
rect 8620 24508 9058 24548
rect 9466 24508 9475 24548
rect 9515 24508 9524 24548
rect 10339 24508 10348 24548
rect 10388 24508 10397 24548
rect 11770 24508 11779 24548
rect 11828 24508 11959 24548
rect 2476 24380 2516 24508
rect 2860 24464 2900 24508
rect 9018 24464 9058 24508
rect 12748 24464 12788 24592
rect 14476 24548 14516 24676
rect 16396 24632 16436 24676
rect 17932 24632 17972 24676
rect 18988 24632 19028 24676
rect 19468 24632 19508 24676
rect 25324 24651 25364 24676
rect 25324 24632 25460 24651
rect 29068 24632 29108 24760
rect 29788 24676 29836 24716
rect 29876 24676 29885 24716
rect 29788 24632 29828 24676
rect 15373 24592 15382 24632
rect 15422 24592 16108 24632
rect 16148 24592 16157 24632
rect 16387 24592 16396 24632
rect 16436 24592 16445 24632
rect 16570 24623 16588 24632
rect 16570 24583 16579 24623
rect 16628 24592 16759 24632
rect 17033 24592 17155 24632
rect 17204 24592 17213 24632
rect 17609 24592 17740 24632
rect 17780 24592 17789 24632
rect 17914 24592 17923 24632
rect 17963 24592 17972 24632
rect 18019 24592 18028 24632
rect 18068 24592 18220 24632
rect 18260 24592 18269 24632
rect 18377 24592 18403 24632
rect 18443 24592 18508 24632
rect 18548 24592 18557 24632
rect 18617 24592 18700 24632
rect 18779 24592 18797 24632
rect 18905 24592 18988 24632
rect 19067 24592 19076 24632
rect 19145 24592 19267 24632
rect 19316 24592 19325 24632
rect 19450 24592 19459 24632
rect 19499 24592 19508 24632
rect 20524 24592 21859 24632
rect 21908 24592 21917 24632
rect 22435 24592 22444 24632
rect 22484 24592 22493 24632
rect 22793 24592 22924 24632
rect 22964 24592 22973 24632
rect 24355 24592 24364 24632
rect 24404 24592 25123 24632
rect 25163 24592 25172 24632
rect 25324 24611 25708 24632
rect 25420 24592 25708 24611
rect 25748 24592 25757 24632
rect 25891 24592 25900 24632
rect 25940 24592 25949 24632
rect 26458 24592 26467 24632
rect 26507 24592 27340 24632
rect 27380 24592 27389 24632
rect 28909 24592 28918 24632
rect 28958 24592 29012 24632
rect 29059 24592 29068 24632
rect 29108 24592 29117 24632
rect 29251 24592 29260 24632
rect 29300 24592 29644 24632
rect 29684 24592 29693 24632
rect 29788 24592 29836 24632
rect 29876 24592 29885 24632
rect 30019 24592 30028 24632
rect 30068 24592 30124 24632
rect 30164 24592 30199 24632
rect 16619 24583 16628 24592
rect 16570 24582 16628 24583
rect 20524 24548 20564 24592
rect 22444 24548 22484 24592
rect 25900 24548 25940 24592
rect 28972 24548 29012 24592
rect 12844 24508 14516 24548
rect 16723 24508 16732 24548
rect 16772 24508 20564 24548
rect 21571 24508 21580 24548
rect 21620 24508 21629 24548
rect 22444 24508 23788 24548
rect 23828 24508 23837 24548
rect 25315 24508 25324 24548
rect 25364 24508 25373 24548
rect 25420 24508 25940 24548
rect 27744 24508 28628 24548
rect 28714 24508 28723 24548
rect 28763 24508 28780 24548
rect 28820 24508 28903 24548
rect 28972 24508 29068 24548
rect 29108 24508 29117 24548
rect 29164 24508 30260 24548
rect 12844 24464 12884 24508
rect 2563 24424 2572 24464
rect 2612 24424 2743 24464
rect 2860 24424 4148 24464
rect 9018 24424 9580 24464
rect 9620 24424 9629 24464
rect 11971 24424 11980 24464
rect 12020 24424 12788 24464
rect 12835 24424 12844 24464
rect 12884 24424 12893 24464
rect 12940 24424 17108 24464
rect 17225 24424 17251 24464
rect 17291 24424 17356 24464
rect 17396 24424 17405 24464
rect 18377 24424 18448 24464
rect 18488 24424 18508 24464
rect 18548 24424 18557 24464
rect 18700 24424 19564 24464
rect 19604 24424 19613 24464
rect 22435 24424 22444 24464
rect 22484 24424 23212 24464
rect 23252 24424 23261 24464
rect 451 24340 460 24380
rect 500 24340 2516 24380
rect 3139 24340 3148 24380
rect 3188 24340 3532 24380
rect 3572 24340 3581 24380
rect 4108 24296 4148 24424
rect 12940 24380 12980 24424
rect 17068 24380 17108 24424
rect 18700 24380 18740 24424
rect 25420 24380 25460 24508
rect 28588 24464 28628 24508
rect 29164 24464 29204 24508
rect 30220 24464 30260 24508
rect 28588 24424 29204 24464
rect 29251 24424 29260 24464
rect 29300 24424 29452 24464
rect 29492 24424 29501 24464
rect 30211 24424 30220 24464
rect 30260 24424 30269 24464
rect 30595 24424 30604 24464
rect 30644 24424 30653 24464
rect 30857 24424 30988 24464
rect 31028 24424 31037 24464
rect 30604 24380 30644 24424
rect 4867 24340 4876 24380
rect 4916 24340 9196 24380
rect 9236 24340 9245 24380
rect 12521 24340 12556 24380
rect 12596 24340 12652 24380
rect 12692 24340 12701 24380
rect 12748 24340 12980 24380
rect 13036 24340 14860 24380
rect 14900 24340 14909 24380
rect 15139 24340 15148 24380
rect 15188 24340 15724 24380
rect 15764 24340 15773 24380
rect 17068 24340 18740 24380
rect 20201 24340 20332 24380
rect 20372 24340 20908 24380
rect 20948 24340 20957 24380
rect 21004 24340 22732 24380
rect 22772 24340 22781 24380
rect 24451 24340 24460 24380
rect 24500 24340 25460 24380
rect 25577 24340 25708 24380
rect 25748 24340 25757 24380
rect 28265 24340 28396 24380
rect 28436 24340 28445 24380
rect 28675 24340 28684 24380
rect 28724 24340 29164 24380
rect 29204 24340 29213 24380
rect 29443 24340 29452 24380
rect 29492 24340 29836 24380
rect 29876 24340 29885 24380
rect 30019 24340 30028 24380
rect 30068 24340 30644 24380
rect 12748 24296 12788 24340
rect 13036 24296 13076 24340
rect 21004 24296 21044 24340
rect 4108 24256 12788 24296
rect 12835 24256 12844 24296
rect 12884 24256 13076 24296
rect 14179 24256 14188 24296
rect 14228 24256 21044 24296
rect 22051 24256 22060 24296
rect 22100 24256 25516 24296
rect 25556 24256 25565 24296
rect 3103 24172 3112 24212
rect 3480 24172 3489 24212
rect 8995 24172 9004 24212
rect 9044 24172 10636 24212
rect 10676 24172 10685 24212
rect 10877 24172 10886 24212
rect 11254 24172 11263 24212
rect 11308 24172 14324 24212
rect 18651 24172 18660 24212
rect 19028 24172 19037 24212
rect 19276 24172 24460 24212
rect 24500 24172 24509 24212
rect 26425 24172 26434 24212
rect 26802 24172 26811 24212
rect 11308 24128 11348 24172
rect 10051 24088 10060 24128
rect 10100 24088 11348 24128
rect 14284 24044 14324 24172
rect 19276 24044 19316 24172
rect 23788 24088 29740 24128
rect 29780 24088 29789 24128
rect 23788 24044 23828 24088
rect 1114 24004 1123 24044
rect 1163 24004 1172 24044
rect 4771 24004 4780 24044
rect 4820 24004 6356 24044
rect 6665 24004 6787 24044
rect 6836 24004 6845 24044
rect 9955 24004 9964 24044
rect 10004 24004 10828 24044
rect 10868 24004 10877 24044
rect 12617 24004 12700 24044
rect 12740 24004 12748 24044
rect 12788 24004 12797 24044
rect 12844 24004 13516 24044
rect 13556 24004 13565 24044
rect 14284 24004 15820 24044
rect 15860 24004 15869 24044
rect 16195 24004 16204 24044
rect 16244 24004 16588 24044
rect 16628 24004 16637 24044
rect 19258 24004 19267 24044
rect 19307 24004 19316 24044
rect 19843 24004 19852 24044
rect 19892 24004 21955 24044
rect 21995 24004 22348 24044
rect 22388 24004 22397 24044
rect 23779 24004 23788 24044
rect 23828 24004 23837 24044
rect 25769 24004 25891 24044
rect 25940 24004 25949 24044
rect 27305 24004 27436 24044
rect 27476 24004 27485 24044
rect 28195 24004 28204 24044
rect 28244 24004 28532 24044
rect 28579 24004 28588 24044
rect 28628 24004 28876 24044
rect 28916 24004 28925 24044
rect 29635 24004 29644 24044
rect 29684 24004 29836 24044
rect 29876 24004 29885 24044
rect 1132 23960 1172 24004
rect 521 23920 556 23960
rect 596 23920 652 23960
rect 692 23920 701 23960
rect 1132 23920 2324 23960
rect 3331 23920 3340 23960
rect 3380 23920 3572 23960
rect 1420 23792 1460 23801
rect 2284 23792 2324 23920
rect 3532 23876 3572 23920
rect 3523 23836 3532 23876
rect 3572 23836 3581 23876
rect 5184 23836 5260 23876
rect 5300 23836 5309 23876
rect 355 23752 364 23792
rect 404 23752 652 23792
rect 692 23752 701 23792
rect 768 23752 777 23792
rect 817 23752 884 23792
rect 931 23752 940 23792
rect 980 23752 1111 23792
rect 1289 23752 1420 23792
rect 1460 23752 1469 23792
rect 2275 23752 2284 23792
rect 2324 23752 2333 23792
rect 2537 23752 2668 23792
rect 2708 23752 2717 23792
rect 2938 23752 2947 23792
rect 2987 23752 3691 23792
rect 3898 23752 3907 23792
rect 3947 23752 4204 23792
rect 4244 23752 4253 23792
rect 4867 23752 4876 23792
rect 4916 23752 6124 23792
rect 6164 23752 6173 23792
rect 652 23456 692 23752
rect 844 23540 884 23752
rect 1420 23743 1460 23752
rect 3651 23708 3691 23752
rect 6316 23708 6356 24004
rect 12844 23960 12884 24004
rect 6412 23920 12364 23960
rect 12404 23920 12413 23960
rect 12835 23920 12844 23960
rect 12884 23920 12893 23960
rect 15619 23920 15628 23960
rect 15668 23920 18316 23960
rect 18356 23920 18365 23960
rect 6412 23834 6452 23920
rect 19276 23876 19316 24004
rect 28492 23960 28532 24004
rect 19651 23920 19660 23960
rect 19700 23920 20332 23960
rect 20372 23920 20381 23960
rect 21970 23920 22772 23960
rect 24355 23920 24364 23960
rect 24404 23920 26324 23960
rect 7075 23836 7084 23876
rect 7124 23836 7200 23876
rect 7852 23836 8140 23876
rect 8180 23836 8242 23876
rect 8282 23836 8311 23876
rect 9004 23836 9524 23876
rect 9763 23836 9772 23876
rect 9812 23836 11308 23876
rect 11348 23836 11357 23876
rect 11491 23836 11500 23876
rect 11540 23836 12980 23876
rect 13507 23836 13516 23876
rect 13556 23836 13565 23876
rect 15130 23836 15139 23876
rect 15188 23836 15319 23876
rect 15593 23836 15724 23876
rect 15764 23836 15773 23876
rect 16204 23836 16300 23876
rect 16340 23836 16349 23876
rect 16588 23836 16684 23876
rect 16724 23836 18124 23876
rect 18164 23836 18173 23876
rect 18220 23836 19316 23876
rect 19372 23836 20180 23876
rect 20554 23864 20563 23904
rect 20603 23876 20612 23904
rect 21970 23876 22010 23920
rect 22732 23876 22772 23920
rect 26284 23876 26324 23920
rect 28108 23920 28436 23960
rect 28492 23920 30307 23960
rect 30347 23920 30356 23960
rect 30499 23920 30508 23960
rect 30548 23920 30557 23960
rect 28108 23876 28148 23920
rect 20603 23864 21044 23876
rect 20572 23836 21044 23864
rect 21161 23836 21292 23876
rect 21332 23836 21341 23876
rect 21514 23867 21970 23876
rect 6412 23794 6430 23834
rect 6470 23794 6479 23834
rect 7084 23792 7124 23836
rect 7852 23792 7892 23836
rect 9004 23792 9044 23836
rect 9484 23792 9524 23836
rect 12940 23792 12980 23836
rect 16204 23792 16244 23836
rect 16444 23792 16484 23801
rect 16588 23792 16628 23836
rect 18220 23792 18260 23836
rect 19372 23792 19412 23836
rect 20140 23792 20180 23836
rect 6604 23752 6782 23792
rect 6822 23752 6831 23792
rect 7786 23752 7795 23792
rect 7835 23752 7892 23792
rect 8323 23752 8332 23792
rect 8372 23752 8620 23792
rect 8660 23752 8669 23792
rect 8899 23752 8908 23792
rect 8948 23752 9004 23792
rect 9044 23752 9079 23792
rect 9187 23752 9196 23792
rect 9236 23752 9367 23792
rect 9484 23752 9859 23792
rect 9899 23752 9908 23792
rect 9955 23752 9964 23792
rect 10004 23752 10252 23792
rect 10292 23752 10301 23792
rect 10522 23752 10531 23792
rect 10571 23752 10580 23792
rect 11033 23752 11116 23792
rect 11156 23752 11164 23792
rect 11204 23752 11213 23792
rect 11299 23752 11308 23792
rect 11348 23752 11357 23792
rect 12259 23752 12268 23792
rect 12308 23752 12317 23792
rect 12425 23752 12556 23792
rect 12596 23752 12605 23792
rect 12940 23752 13036 23792
rect 13076 23752 14755 23792
rect 14795 23752 14804 23792
rect 15235 23752 15244 23792
rect 15284 23752 15388 23792
rect 15428 23752 15437 23792
rect 15497 23752 15567 23792
rect 15607 23752 15628 23792
rect 15668 23752 15677 23792
rect 15785 23752 15859 23792
rect 15899 23752 15916 23792
rect 15956 23752 15965 23792
rect 16070 23752 16079 23792
rect 16119 23752 16128 23792
rect 16200 23752 16209 23792
rect 16249 23752 16258 23792
rect 16303 23752 16312 23792
rect 16352 23752 16387 23792
rect 16570 23752 16579 23792
rect 16619 23752 16628 23792
rect 16745 23752 16876 23792
rect 16916 23752 16925 23792
rect 17068 23752 17251 23792
rect 17291 23752 17300 23792
rect 17347 23752 17356 23792
rect 17396 23752 17644 23792
rect 17684 23752 17693 23792
rect 18202 23752 18211 23792
rect 18251 23752 18260 23792
rect 18307 23752 18316 23792
rect 18356 23752 18487 23792
rect 18857 23752 18892 23792
rect 18932 23752 18979 23792
rect 19019 23752 19028 23792
rect 19075 23752 19084 23792
rect 19124 23752 19412 23792
rect 19732 23752 19741 23792
rect 19781 23752 19796 23792
rect 19843 23752 19852 23792
rect 19892 23752 20023 23792
rect 20140 23752 20236 23792
rect 20276 23752 20515 23792
rect 20555 23752 20564 23792
rect 6604 23708 6644 23752
rect 7084 23708 7124 23752
rect 9196 23708 9236 23752
rect 1112 23668 1121 23708
rect 1161 23668 1228 23708
rect 1268 23668 1292 23708
rect 1516 23668 2900 23708
rect 3043 23668 3052 23708
rect 3092 23668 3223 23708
rect 3651 23668 4780 23708
rect 4820 23668 4829 23708
rect 6089 23668 6220 23708
rect 6260 23668 6269 23708
rect 6316 23668 6644 23708
rect 6857 23668 6988 23708
rect 7028 23668 7037 23708
rect 7084 23668 9100 23708
rect 9140 23668 9149 23708
rect 9196 23668 9524 23708
rect 1516 23624 1556 23668
rect 2860 23624 2900 23668
rect 9484 23624 9524 23668
rect 1315 23584 1324 23624
rect 1364 23584 1556 23624
rect 1603 23584 1612 23624
rect 1652 23584 1661 23624
rect 2860 23584 3532 23624
rect 3572 23584 3581 23624
rect 5059 23584 5068 23624
rect 5108 23584 5836 23624
rect 5876 23584 5885 23624
rect 6281 23584 6316 23624
rect 6356 23584 6412 23624
rect 6452 23584 6461 23624
rect 6595 23584 6604 23624
rect 6644 23584 6653 23624
rect 7555 23584 7564 23624
rect 7604 23584 7660 23624
rect 7700 23584 7735 23624
rect 7913 23584 7948 23624
rect 7988 23584 8035 23624
rect 8075 23584 8093 23624
rect 9065 23584 9196 23624
rect 9236 23584 9245 23624
rect 9466 23584 9475 23624
rect 9515 23584 9524 23624
rect 9868 23624 9908 23752
rect 10217 23668 10348 23708
rect 10388 23668 10397 23708
rect 9868 23584 10147 23624
rect 10187 23584 10196 23624
rect 1612 23540 1652 23584
rect 6604 23540 6644 23584
rect 9196 23540 9236 23584
rect 844 23500 1652 23540
rect 2860 23500 6644 23540
rect 7171 23500 7180 23540
rect 7220 23500 9236 23540
rect 9484 23540 9524 23584
rect 10540 23540 10580 23752
rect 11308 23708 11348 23752
rect 12268 23708 12308 23752
rect 10819 23668 10828 23708
rect 10868 23668 11348 23708
rect 11395 23668 11404 23708
rect 11444 23668 11875 23708
rect 11915 23668 11924 23708
rect 12268 23668 12460 23708
rect 12500 23668 12509 23708
rect 10627 23584 10636 23624
rect 10676 23584 11011 23624
rect 11051 23584 11060 23624
rect 9484 23500 10580 23540
rect 16088 23540 16128 23752
rect 16312 23708 16352 23752
rect 16291 23668 16300 23708
rect 16340 23668 16352 23708
rect 16444 23708 16484 23752
rect 16444 23668 16972 23708
rect 17012 23668 17021 23708
rect 16195 23584 16204 23624
rect 16244 23584 16732 23624
rect 16772 23584 16781 23624
rect 17068 23540 17108 23752
rect 18988 23708 19028 23752
rect 19756 23708 19796 23752
rect 20606 23708 20646 23836
rect 21004 23792 21044 23836
rect 21514 23827 21523 23867
rect 21563 23836 21970 23867
rect 22010 23836 22019 23876
rect 22505 23836 22627 23876
rect 22676 23836 22685 23876
rect 22732 23836 23156 23876
rect 24067 23836 24076 23876
rect 24116 23836 25472 23876
rect 21563 23827 21572 23836
rect 21514 23826 21572 23827
rect 23116 23792 23156 23836
rect 25432 23792 25472 23836
rect 25756 23836 25804 23876
rect 25844 23836 25853 23876
rect 26284 23836 28148 23876
rect 28396 23876 28436 23920
rect 28396 23836 28924 23876
rect 28964 23836 28973 23876
rect 29155 23836 29164 23876
rect 29204 23836 29396 23876
rect 25756 23792 25796 23836
rect 26188 23792 26228 23801
rect 20873 23752 21004 23792
rect 21044 23752 21053 23792
rect 21379 23752 21388 23792
rect 21428 23752 21437 23792
rect 21616 23752 21625 23792
rect 21665 23752 21772 23792
rect 21812 23752 21821 23792
rect 21929 23752 22060 23792
rect 22100 23752 22109 23792
rect 22498 23752 22507 23792
rect 22547 23752 22676 23792
rect 22723 23752 22732 23792
rect 22772 23752 22781 23792
rect 22985 23752 23116 23792
rect 23156 23752 23165 23792
rect 23971 23752 23980 23792
rect 24020 23752 24364 23792
rect 24404 23752 24413 23792
rect 24809 23752 24940 23792
rect 24980 23752 24989 23792
rect 25034 23752 25132 23792
rect 25196 23752 25214 23792
rect 25306 23752 25315 23792
rect 25355 23752 25364 23792
rect 25432 23752 25459 23792
rect 25499 23752 25508 23792
rect 25594 23752 25603 23792
rect 25643 23752 25652 23792
rect 25716 23752 25725 23792
rect 25765 23752 25796 23792
rect 25865 23752 25889 23792
rect 25929 23752 25996 23792
rect 26036 23752 26045 23792
rect 26179 23752 26188 23792
rect 26228 23752 26359 23792
rect 27235 23752 27244 23792
rect 27284 23752 27415 23792
rect 28099 23752 28108 23792
rect 28148 23752 28204 23792
rect 28244 23752 28279 23792
rect 28387 23752 28396 23792
rect 28436 23752 28445 23792
rect 21388 23708 21428 23752
rect 17155 23668 17164 23708
rect 17204 23668 17452 23708
rect 17492 23668 17501 23708
rect 18988 23668 19700 23708
rect 19747 23668 19756 23708
rect 19796 23668 19828 23708
rect 20140 23668 20646 23708
rect 20812 23668 21428 23708
rect 19660 23624 19700 23668
rect 20140 23624 20180 23668
rect 20812 23624 20852 23668
rect 18473 23584 18508 23624
rect 18548 23584 18604 23624
rect 18644 23584 18653 23624
rect 19546 23584 19555 23624
rect 19595 23584 19604 23624
rect 19660 23584 20180 23624
rect 20606 23584 20812 23624
rect 20852 23584 20861 23624
rect 21082 23584 21091 23624
rect 21131 23584 21388 23624
rect 21428 23584 22444 23624
rect 22484 23584 22493 23624
rect 19564 23540 19604 23584
rect 16088 23500 16876 23540
rect 16916 23500 17108 23540
rect 19363 23500 19372 23540
rect 19412 23500 19604 23540
rect 2860 23456 2900 23500
rect 652 23416 2900 23456
rect 4343 23416 4352 23456
rect 4720 23416 4729 23456
rect 9379 23416 9388 23456
rect 9428 23416 11884 23456
rect 11924 23416 11933 23456
rect 12117 23416 12126 23456
rect 12494 23416 12503 23456
rect 15148 23416 15916 23456
rect 15956 23416 15965 23456
rect 16291 23416 16300 23456
rect 16340 23416 19796 23456
rect 19891 23416 19900 23456
rect 20268 23416 20277 23456
rect 748 23332 5492 23372
rect 521 23164 556 23204
rect 596 23164 643 23204
rect 683 23164 701 23204
rect 748 23120 788 23332
rect 5452 23288 5492 23332
rect 7276 23332 9004 23372
rect 9044 23332 9053 23372
rect 10723 23332 10732 23372
rect 10772 23332 12980 23372
rect 13411 23332 13420 23372
rect 13460 23332 14041 23372
rect 7276 23288 7316 23332
rect 12940 23288 12980 23332
rect 2563 23248 2572 23288
rect 2612 23248 2956 23288
rect 2996 23248 3005 23288
rect 3907 23248 3916 23288
rect 3956 23248 4300 23288
rect 4340 23248 4349 23288
rect 4483 23248 4492 23288
rect 4532 23248 4780 23288
rect 4820 23248 4829 23288
rect 5434 23248 5443 23288
rect 5483 23248 5492 23288
rect 5635 23248 5644 23288
rect 5684 23248 6796 23288
rect 6836 23248 6988 23288
rect 7028 23248 7037 23288
rect 7258 23248 7267 23288
rect 7307 23248 7316 23288
rect 7363 23248 7372 23288
rect 7412 23248 7900 23288
rect 7940 23248 7949 23288
rect 8140 23248 8236 23288
rect 8276 23248 8285 23288
rect 11683 23248 11692 23288
rect 11732 23248 11788 23288
rect 11828 23248 11863 23288
rect 12940 23248 13891 23288
rect 13931 23248 13940 23288
rect 4300 23164 5548 23204
rect 5588 23164 5597 23204
rect 6259 23164 6268 23204
rect 6308 23164 6604 23204
rect 6644 23164 6653 23204
rect 6892 23164 7084 23204
rect 7124 23164 7133 23204
rect 7444 23164 7468 23204
rect 7508 23164 7517 23204
rect 7625 23164 7747 23204
rect 7796 23164 7805 23204
rect 4300 23120 4340 23164
rect 6892 23120 6932 23164
rect 163 23080 172 23120
rect 212 23080 788 23120
rect 1018 23080 1027 23120
rect 1076 23080 1207 23120
rect 3305 23080 3340 23120
rect 3380 23080 3436 23120
rect 3476 23080 3485 23120
rect 3785 23080 3820 23120
rect 3860 23080 3916 23120
rect 3956 23080 3965 23120
rect 4291 23080 4300 23120
rect 4340 23080 4349 23120
rect 5059 23080 5068 23120
rect 5108 23080 5164 23120
rect 5204 23080 5239 23120
rect 5722 23080 5731 23120
rect 5771 23111 6412 23120
rect 5771 23080 6115 23111
rect 6106 23071 6115 23080
rect 6155 23080 6412 23111
rect 6452 23080 6461 23120
rect 6883 23080 6892 23120
rect 6932 23080 6941 23120
rect 7075 23080 7084 23120
rect 7124 23080 7133 23120
rect 6155 23071 6164 23080
rect 6106 23070 6164 23071
rect 7084 23036 7124 23080
rect 7271 23075 7280 23115
rect 7320 23075 7329 23115
rect 7444 23078 7484 23164
rect 8140 23120 8180 23248
rect 8236 23164 13228 23204
rect 13268 23164 13277 23204
rect 8236 23120 8276 23164
rect 14001 23120 14041 23332
rect 14188 23248 14668 23288
rect 14708 23248 14717 23288
rect 14188 23204 14228 23248
rect 14104 23164 14228 23204
rect 14467 23164 14476 23204
rect 14516 23164 14525 23204
rect 14104 23120 14144 23164
rect 14476 23120 14516 23164
rect 15148 23120 15188 23416
rect 19756 23372 19796 23416
rect 20606 23372 20646 23584
rect 22636 23540 22676 23752
rect 22732 23708 22772 23752
rect 25324 23708 25364 23752
rect 22732 23668 23732 23708
rect 23779 23668 23788 23708
rect 23828 23668 24259 23708
rect 24299 23668 24308 23708
rect 24547 23668 24556 23708
rect 24596 23668 25364 23708
rect 25612 23708 25652 23752
rect 26188 23743 26228 23752
rect 28396 23708 28436 23752
rect 25612 23668 25900 23708
rect 25940 23668 25949 23708
rect 26275 23668 26284 23708
rect 26324 23668 28436 23708
rect 23692 23624 23732 23668
rect 22810 23584 22819 23624
rect 22859 23584 23060 23624
rect 23692 23584 25324 23624
rect 25364 23584 25373 23624
rect 25498 23584 25507 23624
rect 25556 23584 25687 23624
rect 26083 23584 26092 23624
rect 26132 23584 26141 23624
rect 26563 23584 26572 23624
rect 26612 23584 26621 23624
rect 28282 23584 28291 23624
rect 28331 23584 28340 23624
rect 22636 23500 22732 23540
rect 22772 23500 22781 23540
rect 15244 23332 17452 23372
rect 17492 23332 17501 23372
rect 19756 23332 20180 23372
rect 15244 23288 15284 23332
rect 20140 23288 20180 23332
rect 20572 23332 20646 23372
rect 20572 23288 20612 23332
rect 15235 23248 15244 23288
rect 15284 23248 15293 23288
rect 15619 23248 15628 23288
rect 15668 23248 15872 23288
rect 16195 23248 16204 23288
rect 16244 23248 16253 23288
rect 16435 23248 16444 23288
rect 16484 23248 16684 23288
rect 16724 23248 16733 23288
rect 17068 23248 17356 23288
rect 17396 23248 17405 23288
rect 19459 23248 19468 23288
rect 19508 23248 19747 23288
rect 19787 23248 19796 23288
rect 20140 23248 20236 23288
rect 20276 23248 20285 23288
rect 20428 23248 20612 23288
rect 20698 23248 20707 23288
rect 20747 23248 20812 23288
rect 20852 23248 20887 23288
rect 21091 23248 21100 23288
rect 21140 23248 21149 23288
rect 15235 23164 15244 23204
rect 15284 23164 15764 23204
rect 15724 23120 15764 23164
rect 15832 23120 15872 23248
rect 16204 23204 16244 23248
rect 16108 23164 16244 23204
rect 16963 23164 16972 23204
rect 17012 23164 17021 23204
rect 16108 23120 16148 23164
rect 7651 23080 7660 23120
rect 7700 23080 7892 23120
rect 8083 23080 8092 23120
rect 8132 23080 8180 23120
rect 8227 23080 8236 23120
rect 8276 23080 8285 23120
rect 8410 23080 8419 23120
rect 8459 23080 8716 23120
rect 8756 23080 8765 23120
rect 8820 23080 8908 23120
rect 8948 23080 8951 23120
rect 8991 23080 9000 23120
rect 9187 23080 9196 23120
rect 9236 23080 9388 23120
rect 9428 23080 9437 23120
rect 9850 23080 9859 23120
rect 9908 23080 11788 23120
rect 11828 23080 11837 23120
rect 11971 23080 11980 23120
rect 12020 23080 12029 23120
rect 12643 23080 12652 23120
rect 12692 23080 13132 23120
rect 13172 23080 13181 23120
rect 13315 23080 13324 23120
rect 13364 23080 13516 23120
rect 13556 23080 13565 23120
rect 13612 23109 13860 23120
rect 13612 23080 13820 23109
rect 7276 23038 7320 23075
rect 7411 23038 7420 23078
rect 7460 23038 7484 23078
rect 1987 22996 1996 23036
rect 2036 22996 2045 23036
rect 4675 22996 4684 23036
rect 4724 22996 5347 23036
rect 5387 22996 5396 23036
rect 5635 22996 5644 23036
rect 5684 22996 5923 23036
rect 5963 22996 5972 23036
rect 6211 22996 6220 23036
rect 6260 22996 7180 23036
rect 7220 22996 7229 23036
rect 7276 22952 7316 23038
rect 7852 23036 7892 23080
rect 11980 23036 12020 23080
rect 13612 23036 13652 23080
rect 13811 23069 13820 23080
rect 13860 23069 13869 23109
rect 13992 23080 14001 23120
rect 14041 23080 14050 23120
rect 14095 23080 14104 23120
rect 14144 23080 14153 23120
rect 14234 23080 14243 23120
rect 14283 23080 14310 23120
rect 14362 23080 14371 23120
rect 14411 23080 14516 23120
rect 14563 23080 14572 23120
rect 14612 23080 14743 23120
rect 15148 23080 15556 23120
rect 15596 23080 15605 23120
rect 15706 23080 15715 23120
rect 15755 23080 15764 23120
rect 15823 23080 15832 23120
rect 15872 23080 15881 23120
rect 15994 23080 16003 23120
rect 16043 23080 16052 23120
rect 16096 23080 16105 23120
rect 16145 23080 16154 23120
rect 16204 23080 16243 23120
rect 16283 23080 16292 23120
rect 7546 22996 7555 23036
rect 7604 22996 7735 23036
rect 7843 22996 7852 23036
rect 7892 22996 7901 23036
rect 8969 22996 9091 23036
rect 9140 22996 9149 23036
rect 9283 22996 9292 23036
rect 9332 22996 9484 23036
rect 9524 22996 9533 23036
rect 10339 22996 10348 23036
rect 10388 22996 10397 23036
rect 11491 22996 11500 23036
rect 11540 22996 12844 23036
rect 12884 22996 12893 23036
rect 13411 22996 13420 23036
rect 13460 22996 13652 23036
rect 14001 23036 14041 23080
rect 14270 23036 14310 23080
rect 16012 23036 16052 23080
rect 16204 23036 16244 23080
rect 14001 22996 14081 23036
rect 14179 22996 14188 23036
rect 14228 22996 14310 23036
rect 15715 22996 15724 23036
rect 15764 22996 16052 23036
rect 16099 22996 16108 23036
rect 16148 22996 16244 23036
rect 16972 23036 17012 23164
rect 17068 23120 17108 23248
rect 17155 23164 17164 23204
rect 17204 23164 17684 23204
rect 17644 23120 17684 23164
rect 18124 23164 18892 23204
rect 18932 23164 18941 23204
rect 19555 23164 19564 23204
rect 19604 23164 20092 23204
rect 20132 23164 20141 23204
rect 18124 23120 18164 23164
rect 20428 23120 20468 23248
rect 21100 23204 21140 23248
rect 20515 23164 20524 23204
rect 20564 23164 20606 23204
rect 20646 23164 20695 23204
rect 20803 23164 20812 23204
rect 20852 23164 21140 23204
rect 21571 23164 21580 23204
rect 21620 23164 22484 23204
rect 17059 23080 17068 23120
rect 17108 23080 17117 23120
rect 17292 23080 17305 23120
rect 17345 23080 17452 23120
rect 17492 23080 17501 23120
rect 17626 23080 17635 23120
rect 17675 23080 17684 23120
rect 17827 23080 17836 23120
rect 17876 23080 17932 23120
rect 17972 23080 18007 23120
rect 18115 23080 18124 23120
rect 18164 23080 18173 23120
rect 18307 23080 18316 23120
rect 18356 23080 18365 23120
rect 18556 23080 18565 23120
rect 18644 23080 18745 23120
rect 19459 23080 19468 23120
rect 19508 23080 19517 23120
rect 19642 23080 19651 23120
rect 19700 23080 19831 23120
rect 19953 23080 19962 23120
rect 20002 23080 20468 23120
rect 20908 23111 20948 23120
rect 18316 23036 18356 23080
rect 18430 23038 18439 23078
rect 18479 23038 18488 23078
rect 16972 22996 17108 23036
rect 17155 22996 17164 23036
rect 17227 22996 17335 23036
rect 18278 22996 18316 23036
rect 18356 22996 18365 23036
rect 14041 22952 14081 22996
rect 7267 22912 7276 22952
rect 7316 22912 7325 22952
rect 8803 22912 8812 22952
rect 8852 22912 8861 22952
rect 11395 22912 11404 22952
rect 11444 22912 13076 22952
rect 14041 22912 16396 22952
rect 16436 22912 16445 22952
rect 8812 22868 8852 22912
rect 13036 22868 13076 22912
rect 2563 22828 2572 22868
rect 2612 22828 5836 22868
rect 5876 22828 5885 22868
rect 8410 22828 8419 22868
rect 8459 22828 8468 22868
rect 8812 22828 11212 22868
rect 11252 22828 11261 22868
rect 11875 22828 11884 22868
rect 11924 22828 12931 22868
rect 12971 22828 12980 22868
rect 13036 22828 14572 22868
rect 14612 22828 14621 22868
rect 16099 22828 16108 22868
rect 16148 22828 16300 22868
rect 16340 22828 16349 22868
rect 3103 22660 3112 22700
rect 3480 22660 3489 22700
rect 8428 22616 8468 22828
rect 17068 22784 17108 22996
rect 18448 22952 18488 23038
rect 19468 22952 19508 23080
rect 21082 23080 21091 23120
rect 21140 23080 21271 23120
rect 21379 23080 21388 23120
rect 21428 23080 21772 23120
rect 21812 23080 21821 23120
rect 20908 23060 20948 23071
rect 20908 23036 21024 23060
rect 19555 22996 19564 23036
rect 19604 22996 20332 23036
rect 20372 22996 20381 23036
rect 20899 22996 20908 23036
rect 20948 23020 21024 23036
rect 22444 23036 22484 23164
rect 23020 23120 23060 23584
rect 26092 23540 26132 23584
rect 23299 23500 23308 23540
rect 23348 23500 26132 23540
rect 26572 23456 26612 23584
rect 28300 23540 28340 23584
rect 28195 23500 28204 23540
rect 28244 23500 28340 23540
rect 28588 23456 28628 23836
rect 29356 23792 29396 23836
rect 29452 23836 30220 23876
rect 30260 23836 30269 23876
rect 28759 23752 28768 23792
rect 28808 23752 29068 23792
rect 29108 23752 29117 23792
rect 29347 23752 29356 23792
rect 29396 23752 29405 23792
rect 29452 23708 29492 23836
rect 29932 23792 29972 23836
rect 30508 23834 30548 23920
rect 30604 23836 31124 23876
rect 30499 23794 30508 23834
rect 30548 23794 30557 23834
rect 30604 23792 30644 23836
rect 31084 23792 31124 23836
rect 29609 23752 29644 23792
rect 29684 23752 29740 23792
rect 29780 23752 29789 23792
rect 29923 23752 29932 23792
rect 29972 23752 29981 23792
rect 30115 23752 30124 23792
rect 30164 23752 30173 23792
rect 30240 23752 30315 23792
rect 30355 23752 30364 23792
rect 30604 23752 30693 23792
rect 30733 23752 30742 23792
rect 30883 23752 30892 23792
rect 30932 23752 30941 23792
rect 31075 23752 31084 23792
rect 31124 23752 31133 23792
rect 30124 23708 30164 23752
rect 30316 23708 30356 23752
rect 30892 23708 30932 23752
rect 28963 23668 28972 23708
rect 29012 23668 29492 23708
rect 29644 23668 30164 23708
rect 30307 23668 30316 23708
rect 30356 23668 30604 23708
rect 30644 23668 30653 23708
rect 30700 23668 30932 23708
rect 29155 23584 29164 23624
rect 29204 23584 29251 23624
rect 29291 23584 29335 23624
rect 29417 23584 29548 23624
rect 29588 23584 29597 23624
rect 29644 23540 29684 23668
rect 30700 23624 30740 23668
rect 29827 23584 29836 23624
rect 29876 23584 30740 23624
rect 30857 23584 30988 23624
rect 31028 23584 31037 23624
rect 31084 23540 31124 23752
rect 28867 23500 28876 23540
rect 28916 23500 29684 23540
rect 30220 23500 31124 23540
rect 30220 23456 30260 23500
rect 23788 23416 26612 23456
rect 27665 23416 27674 23456
rect 28042 23416 28051 23456
rect 28579 23416 28588 23456
rect 28628 23416 28637 23456
rect 29539 23416 29548 23456
rect 29588 23416 30260 23456
rect 23788 23120 23828 23416
rect 25315 23332 25324 23372
rect 25364 23332 26572 23372
rect 26612 23332 26621 23372
rect 26755 23248 26764 23288
rect 26804 23248 27244 23288
rect 27284 23248 27293 23288
rect 28396 23248 30028 23288
rect 30068 23248 30077 23288
rect 24250 23164 24259 23204
rect 24299 23164 28204 23204
rect 28244 23164 28253 23204
rect 28396 23120 28436 23248
rect 29155 23164 29164 23204
rect 29204 23164 30260 23204
rect 30220 23120 30260 23164
rect 22601 23080 22732 23120
rect 22772 23080 22781 23120
rect 23020 23080 23596 23120
rect 23636 23080 23645 23120
rect 23788 23080 23831 23120
rect 23871 23080 23880 23120
rect 23962 23111 24020 23120
rect 23962 23071 23971 23111
rect 24011 23071 24020 23111
rect 24067 23080 24076 23120
rect 24116 23080 24247 23120
rect 26153 23080 26179 23120
rect 26219 23080 26284 23120
rect 26324 23080 26333 23120
rect 26563 23080 26572 23120
rect 26612 23080 28436 23120
rect 28579 23080 28588 23120
rect 28628 23080 28675 23120
rect 28715 23080 28759 23120
rect 28963 23080 28972 23120
rect 29012 23080 29059 23120
rect 29099 23080 29452 23120
rect 29492 23080 29501 23120
rect 29731 23080 29740 23120
rect 29780 23080 30028 23120
rect 30068 23080 30077 23120
rect 30211 23080 30220 23120
rect 30260 23080 30269 23120
rect 30316 23080 31180 23120
rect 31220 23080 31229 23120
rect 23962 23070 24020 23071
rect 20948 22996 20957 23020
rect 22444 22996 23060 23036
rect 23020 22952 23060 22996
rect 23980 22952 24020 23070
rect 30316 23036 30356 23080
rect 26371 22996 26380 23036
rect 26420 22996 26429 23036
rect 26554 22996 26563 23036
rect 26603 22996 26860 23036
rect 26900 22996 26909 23036
rect 28896 22996 30028 23036
rect 30068 22996 30077 23036
rect 30124 22996 30356 23036
rect 18019 22912 18028 22952
rect 18068 22912 18488 22952
rect 18595 22912 18604 22952
rect 18644 22912 19508 22952
rect 22051 22912 22060 22952
rect 22100 22912 22924 22952
rect 22964 22912 22973 22952
rect 23020 22912 23788 22952
rect 23828 22912 23837 22952
rect 23980 22912 24116 22952
rect 29155 22912 29164 22952
rect 29204 22912 29260 22952
rect 29300 22912 29335 22952
rect 29513 22912 29644 22952
rect 29684 22912 29693 22952
rect 24076 22868 24116 22912
rect 30124 22868 30164 22996
rect 30281 22912 30412 22952
rect 30452 22912 30461 22952
rect 30508 22912 30796 22952
rect 30836 22912 30845 22952
rect 17513 22828 17548 22868
rect 17588 22828 17635 22868
rect 17675 22828 17693 22868
rect 18787 22828 18796 22868
rect 18836 22828 19084 22868
rect 19124 22828 19133 22868
rect 19843 22828 19852 22868
rect 19892 22828 19948 22868
rect 19988 22828 20023 22868
rect 21571 22828 21580 22868
rect 21620 22828 22060 22868
rect 22100 22828 22109 22868
rect 24076 22828 24940 22868
rect 24980 22828 24989 22868
rect 28771 22828 28780 22868
rect 28820 22828 30164 22868
rect 24076 22784 24116 22828
rect 9283 22744 9292 22784
rect 9332 22744 11500 22784
rect 11540 22744 11549 22784
rect 17068 22744 19124 22784
rect 21475 22744 21484 22784
rect 21524 22744 24116 22784
rect 24748 22744 30124 22784
rect 30164 22744 30173 22784
rect 19084 22700 19124 22744
rect 24748 22700 24788 22744
rect 8803 22660 8812 22700
rect 8852 22660 9236 22700
rect 10877 22660 10886 22700
rect 11254 22660 11263 22700
rect 16209 22660 16300 22700
rect 16340 22660 16349 22700
rect 18651 22660 18660 22700
rect 19028 22660 19037 22700
rect 19084 22660 24788 22700
rect 26425 22660 26434 22700
rect 26802 22660 26811 22700
rect 9196 22616 9236 22660
rect 16209 22616 16249 22660
rect 30508 22616 30548 22912
rect 6702 22576 7276 22616
rect 7316 22576 7325 22616
rect 8428 22576 9100 22616
rect 9140 22576 9149 22616
rect 9196 22576 16249 22616
rect 16300 22576 18316 22616
rect 18356 22576 18365 22616
rect 23692 22576 30548 22616
rect 748 22492 6403 22532
rect 6443 22492 6452 22532
rect 748 22448 788 22492
rect 652 22408 788 22448
rect 1603 22408 1612 22448
rect 1652 22408 5492 22448
rect 5635 22408 5644 22448
rect 5684 22408 5876 22448
rect 0 22364 400 22384
rect 652 22364 692 22408
rect 5452 22364 5492 22408
rect 5836 22364 5876 22408
rect 0 22324 692 22364
rect 739 22324 748 22364
rect 788 22324 797 22364
rect 1516 22324 2612 22364
rect 0 22304 400 22324
rect 748 22280 788 22324
rect 1516 22322 1556 22324
rect 1450 22282 1459 22322
rect 1499 22282 1556 22322
rect 2572 22280 2612 22324
rect 2956 22324 4204 22364
rect 4244 22324 4253 22364
rect 4553 22324 4579 22364
rect 4619 22324 4684 22364
rect 4724 22324 4733 22364
rect 5146 22324 5155 22364
rect 5195 22324 5356 22364
rect 5396 22324 5405 22364
rect 5452 22324 5571 22364
rect 5611 22324 5620 22364
rect 5827 22324 5836 22364
rect 5876 22324 5885 22364
rect 6058 22355 6124 22364
rect 2956 22280 2996 22324
rect 6058 22315 6067 22355
rect 6107 22324 6124 22355
rect 6164 22324 6247 22364
rect 6401 22324 6508 22364
rect 6548 22324 6557 22364
rect 6107 22315 6116 22324
rect 6058 22314 6116 22315
rect 6401 22280 6441 22324
rect 6702 22313 6742 22576
rect 16300 22532 16340 22576
rect 6883 22492 6892 22532
rect 6932 22492 10484 22532
rect 10601 22492 10732 22532
rect 10772 22492 10781 22532
rect 11491 22492 11500 22532
rect 11540 22492 12980 22532
rect 16291 22492 16300 22532
rect 16340 22492 16349 22532
rect 16487 22492 19468 22532
rect 19508 22492 19517 22532
rect 20969 22492 21004 22532
rect 21044 22492 21100 22532
rect 21140 22492 21149 22532
rect 21667 22492 21676 22532
rect 21716 22492 21724 22532
rect 21764 22492 21847 22532
rect 10444 22448 10484 22492
rect 12940 22448 12980 22492
rect 16487 22448 16527 22492
rect 8105 22408 8227 22448
rect 8276 22408 8285 22448
rect 9763 22408 9772 22448
rect 9812 22408 10252 22448
rect 10292 22408 10348 22448
rect 10388 22408 10397 22448
rect 10444 22408 11060 22448
rect 7171 22324 7180 22364
rect 7220 22324 7372 22364
rect 7412 22324 7421 22364
rect 7747 22324 7756 22364
rect 7796 22324 7948 22364
rect 7988 22324 8131 22364
rect 8171 22324 8180 22364
rect 8242 22324 8707 22364
rect 8747 22324 8756 22364
rect 9091 22324 9100 22364
rect 9140 22324 10060 22364
rect 10100 22324 10109 22364
rect 11020 22344 11060 22408
rect 12652 22408 12844 22448
rect 12884 22408 12893 22448
rect 12940 22408 13940 22448
rect 14755 22408 14764 22448
rect 14804 22408 16527 22448
rect 17321 22408 17452 22448
rect 17492 22408 17501 22448
rect 12652 22364 12692 22408
rect 13900 22364 13940 22408
rect 12634 22324 12643 22364
rect 12683 22324 12692 22364
rect 13123 22324 13132 22364
rect 13172 22324 13181 22364
rect 13900 22324 14908 22364
rect 14948 22324 14957 22364
rect 547 22240 556 22280
rect 596 22240 788 22280
rect 1673 22240 1804 22280
rect 1844 22240 1853 22280
rect 1939 22240 1948 22280
rect 1988 22240 2092 22280
rect 2132 22240 2141 22280
rect 2563 22240 2572 22280
rect 2612 22240 2743 22280
rect 2947 22240 2956 22280
rect 2996 22240 3005 22280
rect 3052 22240 3523 22280
rect 3563 22240 3572 22280
rect 3619 22240 3628 22280
rect 3668 22240 3677 22280
rect 3907 22240 3916 22280
rect 3956 22240 4055 22280
rect 4095 22240 4104 22280
rect 4186 22240 4195 22280
rect 4235 22240 4244 22280
rect 4291 22240 4300 22280
rect 4340 22240 4894 22280
rect 4954 22240 4963 22280
rect 5012 22240 5143 22280
rect 5443 22240 5452 22280
rect 5492 22240 5501 22280
rect 5635 22240 5644 22280
rect 5709 22240 5815 22280
rect 5923 22240 5932 22280
rect 5972 22240 5981 22280
rect 6160 22240 6169 22280
rect 6209 22240 6260 22280
rect 6392 22240 6401 22280
rect 6441 22240 6450 22280
rect 6689 22273 6698 22313
rect 6738 22273 6747 22313
rect 8242 22280 8282 22324
rect 13132 22280 13172 22324
rect 15244 22280 15284 22408
rect 15677 22324 15724 22364
rect 15764 22324 15773 22364
rect 15820 22324 16012 22364
rect 16052 22324 16061 22364
rect 16291 22324 16300 22364
rect 16340 22324 16357 22364
rect 15724 22280 15764 22324
rect 15820 22280 15860 22324
rect 16300 22280 16340 22324
rect 16487 22280 16527 22408
rect 16570 22324 16579 22364
rect 16619 22324 16684 22364
rect 16724 22324 16759 22364
rect 16841 22324 16972 22364
rect 17012 22324 17021 22364
rect 17417 22324 17548 22364
rect 17588 22324 17597 22364
rect 20448 22324 20812 22364
rect 20852 22324 20861 22364
rect 21353 22324 21379 22364
rect 21419 22324 21484 22364
rect 21524 22324 21533 22364
rect 21763 22324 21772 22364
rect 21812 22324 21821 22364
rect 21929 22324 22060 22364
rect 22100 22324 22109 22364
rect 23692 22344 23732 22576
rect 24329 22492 24364 22532
rect 24404 22492 24460 22532
rect 24500 22492 24509 22532
rect 25210 22492 25219 22532
rect 25259 22492 26380 22532
rect 26420 22492 26429 22532
rect 26563 22492 26572 22532
rect 26612 22492 26860 22532
rect 26900 22492 26909 22532
rect 27043 22492 27052 22532
rect 27092 22492 27223 22532
rect 27820 22492 28972 22532
rect 29012 22492 29021 22532
rect 27820 22448 27860 22492
rect 25420 22408 27860 22448
rect 29726 22408 30316 22448
rect 30356 22408 30365 22448
rect 30473 22408 30604 22448
rect 30644 22408 30653 22448
rect 30787 22408 30796 22448
rect 30836 22408 30988 22448
rect 31028 22408 31037 22448
rect 21772 22280 21812 22324
rect 25420 22322 25460 22408
rect 25612 22324 25804 22364
rect 25844 22324 25853 22364
rect 27148 22324 27532 22364
rect 27572 22324 27581 22364
rect 29347 22324 29356 22364
rect 29396 22324 29405 22364
rect 25420 22313 25544 22322
rect 25420 22282 25504 22313
rect 6796 22240 6839 22280
rect 6879 22240 6888 22280
rect 6970 22240 6979 22280
rect 7019 22240 7028 22280
rect 7075 22240 7084 22280
rect 7124 22240 7255 22280
rect 7433 22240 7555 22280
rect 7604 22240 7613 22280
rect 8227 22240 8236 22280
rect 8276 22240 8285 22280
rect 8506 22240 8515 22280
rect 8555 22240 8612 22280
rect 8899 22240 8908 22280
rect 8987 22240 9079 22280
rect 9187 22240 9196 22280
rect 9236 22240 9868 22280
rect 9908 22240 9917 22280
rect 11779 22240 11788 22280
rect 11828 22240 12259 22280
rect 12299 22240 12308 22280
rect 13132 22240 13242 22280
rect 13282 22240 13291 22280
rect 13385 22240 13516 22280
rect 13556 22240 13565 22280
rect 13978 22240 13987 22280
rect 14027 22240 14036 22280
rect 14275 22240 14284 22280
rect 14324 22240 14707 22280
rect 14747 22240 14860 22280
rect 14900 22240 14916 22280
rect 15235 22240 15244 22280
rect 15284 22240 15293 22280
rect 15379 22240 15388 22280
rect 15428 22240 15532 22280
rect 15572 22240 15581 22280
rect 15706 22240 15715 22280
rect 15755 22240 15764 22280
rect 15811 22240 15820 22280
rect 15860 22240 15869 22280
rect 16003 22240 16012 22280
rect 16052 22240 16061 22280
rect 16142 22240 16151 22280
rect 16191 22240 16200 22280
rect 16252 22240 16261 22280
rect 16301 22240 16340 22280
rect 16450 22240 16459 22280
rect 16499 22240 16527 22280
rect 16588 22240 16684 22280
rect 16724 22240 16780 22280
rect 16820 22240 16884 22280
rect 17033 22240 17155 22280
rect 17204 22240 17213 22280
rect 17452 22240 18028 22280
rect 18068 22240 18077 22280
rect 18403 22240 18412 22280
rect 18452 22240 18616 22280
rect 18656 22240 18665 22280
rect 19162 22240 19171 22280
rect 19220 22240 19351 22280
rect 19555 22240 19564 22280
rect 19604 22240 21239 22280
rect 21279 22240 21288 22280
rect 21475 22240 21484 22280
rect 21524 22240 21812 22280
rect 21859 22240 21868 22280
rect 21908 22240 22156 22280
rect 22196 22240 22205 22280
rect 22426 22240 22435 22280
rect 22484 22240 22615 22280
rect 24809 22240 24940 22280
rect 24980 22240 24989 22280
rect 25612 22280 25652 22324
rect 27148 22287 27188 22324
rect 27021 22280 27188 22287
rect 29726 22280 29766 22408
rect 30115 22324 30124 22364
rect 30164 22324 30173 22364
rect 30028 22280 30068 22289
rect 30124 22280 30164 22324
rect 25504 22264 25544 22273
rect 25594 22240 25603 22280
rect 25643 22240 25652 22280
rect 25769 22240 25900 22280
rect 25940 22240 25949 22280
rect 26633 22240 26764 22280
rect 26804 22240 26813 22280
rect 26890 22240 26899 22280
rect 26939 22240 26948 22280
rect 26995 22240 27004 22280
rect 27044 22247 27188 22280
rect 27044 22240 27061 22247
rect 27331 22240 27340 22280
rect 27380 22240 28780 22280
rect 28820 22240 29155 22280
rect 29195 22240 29204 22280
rect 29445 22240 29726 22280
rect 29766 22240 29775 22280
rect 29897 22240 30028 22280
rect 30068 22240 30077 22280
rect 30124 22240 30220 22280
rect 30260 22240 30269 22280
rect 30394 22240 30403 22280
rect 30443 22240 30508 22280
rect 30548 22240 30700 22280
rect 30740 22240 30749 22280
rect 835 22156 844 22196
rect 884 22156 1603 22196
rect 1643 22156 1652 22196
rect 3052 22112 3092 22240
rect 3628 22196 3668 22240
rect 3628 22156 4108 22196
rect 4148 22156 4157 22196
rect 979 22072 988 22112
rect 1028 22072 1037 22112
rect 1219 22072 1228 22112
rect 1307 22072 1900 22112
rect 1940 22072 2860 22112
rect 2900 22072 2909 22112
rect 3043 22072 3052 22112
rect 3092 22072 3101 22112
rect 3811 22072 3820 22112
rect 3860 22072 3916 22112
rect 3956 22072 3991 22112
rect 988 22028 1028 22072
rect 4204 22028 4244 22240
rect 4854 22196 4894 22240
rect 5452 22196 5492 22240
rect 5932 22196 5972 22240
rect 6220 22196 6260 22240
rect 6796 22196 6836 22240
rect 4378 22156 4387 22196
rect 4436 22156 4567 22196
rect 4854 22156 6124 22196
rect 6164 22156 6173 22196
rect 6220 22156 6700 22196
rect 6740 22156 6836 22196
rect 6988 22196 7028 22240
rect 8572 22196 8612 22240
rect 6988 22156 7372 22196
rect 7412 22156 7421 22196
rect 7843 22156 7852 22196
rect 7892 22156 7901 22196
rect 8035 22156 8044 22196
rect 8084 22156 8612 22196
rect 13097 22156 13132 22196
rect 13172 22156 13228 22196
rect 13268 22156 13277 22196
rect 6220 22112 6260 22156
rect 4553 22072 4675 22112
rect 4724 22072 4733 22112
rect 6019 22072 6028 22112
rect 6068 22072 6260 22112
rect 6473 22072 6604 22112
rect 6644 22072 6653 22112
rect 7852 22028 7892 22156
rect 8572 22112 8612 22156
rect 13996 22112 14036 22240
rect 16012 22196 16052 22240
rect 16159 22196 16199 22240
rect 14249 22156 14380 22196
rect 14420 22156 14429 22196
rect 15610 22156 15619 22196
rect 15659 22156 16012 22196
rect 16052 22156 16061 22196
rect 16159 22156 16396 22196
rect 16436 22156 16445 22196
rect 8572 22072 9148 22112
rect 9188 22072 9197 22112
rect 9545 22072 9676 22112
rect 9716 22072 9725 22112
rect 9946 22072 9955 22112
rect 9995 22072 10252 22112
rect 10292 22072 10301 22112
rect 10636 22072 12940 22112
rect 12980 22072 14036 22112
rect 14380 22112 14420 22156
rect 16588 22112 16628 22240
rect 17452 22112 17492 22240
rect 26908 22196 26948 22240
rect 18778 22156 18787 22196
rect 18827 22156 19084 22196
rect 19124 22156 19133 22196
rect 26908 22156 26956 22196
rect 26996 22156 27005 22196
rect 27139 22156 27148 22196
rect 27188 22156 27235 22196
rect 27275 22156 27319 22196
rect 29445 22112 29485 22240
rect 30028 22231 30068 22240
rect 29530 22156 29539 22196
rect 29579 22156 29588 22196
rect 14380 22072 16628 22112
rect 16762 22072 16771 22112
rect 16811 22072 17492 22112
rect 17827 22072 17836 22112
rect 17876 22072 17885 22112
rect 18106 22072 18115 22112
rect 18155 22072 18164 22112
rect 18329 22072 18412 22112
rect 18491 22072 18509 22112
rect 21562 22072 21571 22112
rect 21611 22072 21676 22112
rect 21716 22072 21751 22112
rect 24451 22072 24460 22112
rect 24500 22072 24748 22112
rect 24788 22072 24797 22112
rect 25018 22072 25027 22112
rect 25067 22072 25516 22112
rect 25556 22072 25565 22112
rect 25738 22072 25747 22112
rect 25787 22072 29485 22112
rect 29548 22112 29588 22156
rect 29548 22072 29827 22112
rect 29867 22072 29876 22112
rect 29923 22072 29932 22112
rect 29972 22072 30028 22112
rect 30068 22072 30103 22112
rect 30307 22072 30316 22112
rect 30356 22072 30365 22112
rect 988 21988 2380 22028
rect 2420 21988 2429 22028
rect 4204 21988 5587 22028
rect 6403 21988 6412 22028
rect 6452 21988 7892 22028
rect 9148 22028 9188 22072
rect 10636 22028 10676 22072
rect 17836 22028 17876 22072
rect 9148 21988 10676 22028
rect 17251 21988 17260 22028
rect 17300 21988 17876 22028
rect 18124 22028 18164 22072
rect 30316 22028 30356 22072
rect 18124 21988 18892 22028
rect 18932 21988 18941 22028
rect 18988 21988 21484 22028
rect 21524 21988 21533 22028
rect 25891 21988 25900 22028
rect 25940 21988 30356 22028
rect 0 21944 400 21964
rect 0 21904 3340 21944
rect 3380 21904 3389 21944
rect 4343 21904 4352 21944
rect 4720 21904 4729 21944
rect 0 21884 400 21904
rect 1507 21820 1516 21860
rect 1556 21820 5068 21860
rect 5108 21820 5492 21860
rect 5452 21776 5492 21820
rect 5547 21776 5587 21988
rect 18988 21944 19028 21988
rect 8620 21904 9676 21944
rect 9716 21904 9725 21944
rect 12117 21904 12126 21944
rect 12494 21904 12503 21944
rect 13507 21904 13516 21944
rect 13556 21904 16396 21944
rect 16436 21904 16445 21944
rect 16963 21904 16972 21944
rect 17012 21904 19028 21944
rect 19891 21904 19900 21944
rect 20268 21904 20277 21944
rect 27665 21904 27674 21944
rect 28042 21904 28051 21944
rect 5833 21820 6412 21860
rect 6452 21820 6461 21860
rect 874 21736 883 21776
rect 923 21736 2572 21776
rect 2612 21736 2621 21776
rect 5434 21736 5443 21776
rect 5483 21736 5492 21776
rect 5539 21736 5548 21776
rect 5588 21736 5597 21776
rect 1084 21652 1844 21692
rect 1084 21608 1124 21652
rect 1804 21608 1844 21652
rect 2956 21652 3724 21692
rect 3764 21652 3773 21692
rect 4483 21652 4492 21692
rect 4532 21652 4541 21692
rect 4771 21652 4780 21692
rect 4820 21652 4894 21692
rect 2956 21608 2996 21652
rect 4492 21608 4532 21652
rect 4854 21608 4894 21652
rect 5164 21652 5176 21692
rect 5216 21652 5225 21692
rect 5609 21652 5656 21692
rect 5696 21652 5740 21692
rect 5780 21652 5789 21692
rect 5164 21608 5204 21652
rect 5833 21608 5873 21820
rect 5993 21736 6115 21776
rect 6164 21736 6173 21776
rect 6473 21736 6595 21776
rect 6644 21736 6653 21776
rect 6953 21736 6988 21776
rect 7028 21736 7084 21776
rect 7124 21736 7604 21776
rect 7651 21736 7660 21776
rect 7700 21736 7756 21776
rect 7796 21736 7831 21776
rect 7564 21692 7604 21736
rect 6019 21652 6028 21692
rect 6068 21652 6807 21692
rect 6847 21652 7220 21692
rect 7564 21652 8036 21692
rect 8218 21652 8227 21692
rect 8276 21652 8407 21692
rect 7180 21608 7220 21652
rect 7996 21608 8036 21652
rect 8620 21608 8660 21904
rect 8716 21820 9716 21860
rect 10051 21820 10060 21860
rect 10100 21820 15572 21860
rect 17443 21820 17452 21860
rect 17492 21820 26188 21860
rect 26228 21820 26237 21860
rect 8716 21776 8756 21820
rect 9676 21776 9716 21820
rect 15532 21776 15572 21820
rect 8707 21736 8716 21776
rect 8756 21736 8765 21776
rect 9449 21736 9532 21776
rect 9572 21736 9580 21776
rect 9620 21736 9629 21776
rect 9676 21736 11443 21776
rect 11483 21736 11492 21776
rect 13193 21736 13324 21776
rect 13364 21736 13373 21776
rect 13699 21736 13708 21776
rect 13748 21736 15043 21776
rect 15083 21736 15244 21776
rect 15284 21736 15293 21776
rect 15532 21736 18076 21776
rect 18116 21736 18125 21776
rect 18778 21736 18787 21776
rect 18827 21736 20140 21776
rect 20180 21736 20189 21776
rect 23980 21736 24268 21776
rect 24308 21736 24317 21776
rect 24691 21736 24700 21776
rect 24740 21736 24940 21776
rect 24980 21736 24989 21776
rect 25385 21736 25516 21776
rect 25556 21736 25565 21776
rect 27523 21736 27532 21776
rect 27572 21736 28012 21776
rect 28052 21736 28061 21776
rect 9532 21692 9572 21736
rect 8803 21652 8812 21692
rect 8852 21652 9043 21692
rect 9083 21652 9092 21692
rect 9282 21652 9572 21692
rect 9667 21652 9676 21692
rect 9716 21652 10100 21692
rect 10243 21652 10252 21692
rect 10292 21652 10963 21692
rect 11003 21652 11012 21692
rect 13411 21652 13420 21692
rect 13460 21652 15956 21692
rect 16003 21652 16012 21692
rect 16052 21652 16061 21692
rect 16195 21652 16204 21692
rect 16244 21652 16375 21692
rect 16963 21652 16972 21692
rect 17012 21652 17143 21692
rect 17314 21652 17356 21692
rect 17396 21652 17405 21692
rect 17722 21652 17731 21692
rect 17771 21652 17780 21692
rect 18761 21652 18892 21692
rect 18932 21652 20428 21692
rect 20468 21652 20477 21692
rect 20611 21652 20620 21692
rect 20660 21652 21580 21692
rect 21620 21652 21629 21692
rect 9282 21608 9322 21652
rect 10060 21608 10100 21652
rect 15916 21608 15956 21652
rect 16012 21608 16052 21652
rect 17314 21608 17354 21652
rect 17740 21608 17780 21652
rect 18892 21608 18932 21652
rect 23980 21650 24020 21736
rect 23962 21610 23971 21650
rect 24011 21610 24020 21650
rect 24412 21652 24556 21692
rect 24596 21652 24605 21692
rect 25315 21652 25324 21692
rect 25364 21652 26092 21692
rect 26132 21652 26141 21692
rect 26371 21652 26380 21692
rect 26420 21652 27764 21692
rect 24412 21608 24452 21652
rect 27724 21608 27764 21652
rect 1066 21568 1075 21608
rect 1115 21568 1124 21608
rect 1306 21568 1315 21608
rect 1355 21568 1364 21608
rect 1411 21568 1420 21608
rect 1460 21568 1469 21608
rect 1786 21568 1795 21608
rect 1835 21568 1844 21608
rect 2275 21568 2284 21608
rect 2324 21568 2572 21608
rect 2612 21568 2668 21608
rect 2708 21568 2717 21608
rect 2800 21568 2809 21608
rect 2849 21568 2858 21608
rect 2947 21568 2956 21608
rect 2996 21568 3005 21608
rect 3130 21568 3139 21608
rect 3188 21568 3319 21608
rect 3401 21568 3436 21608
rect 3476 21568 3523 21608
rect 3563 21568 3581 21608
rect 3629 21568 3638 21608
rect 3678 21568 3820 21608
rect 3860 21568 4204 21608
rect 4244 21568 4253 21608
rect 4354 21568 4363 21608
rect 4403 21568 4532 21608
rect 4579 21568 4588 21608
rect 4628 21568 4759 21608
rect 4854 21568 4865 21608
rect 4905 21568 4914 21608
rect 4963 21568 4972 21608
rect 5012 21568 5021 21608
rect 5129 21568 5164 21608
rect 5204 21568 5213 21608
rect 5338 21573 5347 21608
rect 5288 21568 5347 21573
rect 5387 21568 5396 21608
rect 5794 21568 5803 21608
rect 5843 21568 5873 21608
rect 6307 21568 6316 21608
rect 6356 21568 6499 21608
rect 6539 21568 6548 21608
rect 6691 21568 6700 21608
rect 6740 21568 7084 21608
rect 7124 21568 7133 21608
rect 7180 21568 7301 21608
rect 7341 21568 7454 21608
rect 7494 21568 7503 21608
rect 7756 21599 7796 21608
rect 0 21524 400 21544
rect 1171 21526 1180 21566
rect 1220 21526 1229 21566
rect 0 21484 1036 21524
rect 1076 21484 1085 21524
rect 0 21464 400 21484
rect 1180 21440 1220 21526
rect 1324 21440 1364 21568
rect 931 21400 940 21440
rect 980 21400 1220 21440
rect 1315 21400 1324 21440
rect 1364 21400 1373 21440
rect 1420 21356 1460 21568
rect 1507 21484 1516 21524
rect 1556 21484 1565 21524
rect 1411 21316 1420 21356
rect 1460 21316 1469 21356
rect 0 21104 400 21124
rect 0 21064 1228 21104
rect 1268 21064 1277 21104
rect 0 21044 400 21064
rect 1516 20852 1556 21484
rect 1804 21440 1844 21568
rect 2818 21524 2858 21568
rect 2083 21484 2092 21524
rect 2132 21484 2476 21524
rect 2516 21484 2525 21524
rect 2572 21484 2691 21524
rect 2731 21484 2740 21524
rect 2818 21484 2860 21524
rect 2900 21484 2909 21524
rect 3010 21484 4483 21524
rect 4523 21484 4532 21524
rect 4675 21484 4684 21524
rect 4724 21484 4855 21524
rect 2572 21440 2612 21484
rect 1804 21400 2516 21440
rect 2563 21400 2572 21440
rect 2612 21400 2621 21440
rect 2476 21356 2516 21400
rect 3010 21356 3050 21484
rect 4492 21440 4532 21484
rect 4972 21440 5012 21568
rect 5288 21533 5381 21568
rect 5288 21524 5328 21533
rect 6019 21526 6028 21566
rect 6068 21526 6116 21566
rect 6076 21524 6116 21526
rect 7996 21568 8140 21608
rect 8180 21568 8189 21608
rect 8620 21568 8728 21608
rect 8768 21568 8777 21608
rect 8899 21568 8908 21608
rect 8948 21568 9238 21608
rect 9278 21568 9322 21608
rect 9370 21599 9620 21608
rect 7756 21524 7796 21559
rect 7891 21526 7900 21566
rect 7940 21526 7949 21566
rect 9370 21559 9379 21599
rect 9419 21583 9620 21599
rect 9676 21599 9908 21608
rect 9419 21568 9580 21583
rect 9419 21559 9428 21568
rect 9370 21558 9428 21559
rect 9571 21543 9580 21568
rect 9620 21543 9629 21583
rect 9676 21568 9859 21599
rect 5059 21484 5068 21524
rect 5108 21484 5328 21524
rect 5900 21484 5909 21524
rect 5949 21484 5972 21524
rect 6076 21484 6124 21524
rect 6164 21484 6173 21524
rect 6403 21484 6412 21524
rect 6452 21484 7203 21524
rect 7243 21484 7468 21524
rect 7508 21484 7517 21524
rect 7709 21484 7756 21524
rect 7796 21484 7805 21524
rect 3331 21400 3340 21440
rect 3380 21400 3956 21440
rect 4492 21400 4972 21440
rect 5012 21400 5021 21440
rect 3916 21356 3956 21400
rect 5932 21356 5972 21484
rect 6019 21400 6028 21440
rect 6068 21400 7652 21440
rect 7612 21356 7652 21400
rect 7900 21356 7940 21526
rect 8026 21484 8035 21524
rect 8075 21484 8084 21524
rect 8227 21484 8236 21524
rect 8276 21484 8563 21524
rect 8603 21484 8612 21524
rect 8044 21440 8084 21484
rect 9676 21440 9716 21568
rect 9850 21559 9859 21568
rect 9899 21559 9908 21599
rect 10060 21599 10388 21608
rect 10060 21568 10339 21599
rect 9850 21558 9908 21559
rect 10330 21559 10339 21568
rect 10379 21559 10388 21599
rect 10531 21568 10540 21608
rect 10580 21568 11116 21608
rect 11168 21568 11287 21608
rect 11486 21568 11596 21608
rect 11648 21568 11732 21608
rect 11779 21568 11788 21608
rect 11828 21568 11959 21608
rect 12713 21568 12844 21608
rect 12884 21568 12893 21608
rect 13097 21568 13228 21608
rect 13268 21568 13277 21608
rect 13507 21568 13516 21608
rect 13556 21568 13655 21608
rect 13695 21568 13704 21608
rect 13865 21568 13900 21608
rect 13940 21568 13996 21608
rect 14036 21568 14045 21608
rect 14249 21568 14371 21608
rect 14420 21568 15331 21608
rect 15371 21568 15380 21608
rect 15593 21568 15628 21608
rect 15668 21568 15724 21608
rect 15764 21568 15773 21608
rect 15907 21568 15916 21608
rect 15956 21568 15965 21608
rect 16012 21568 16108 21608
rect 16148 21568 16157 21608
rect 16291 21568 16300 21608
rect 16340 21568 16396 21608
rect 16436 21568 16471 21608
rect 16579 21568 16588 21608
rect 16628 21568 16637 21608
rect 16684 21568 16780 21608
rect 16820 21568 16829 21608
rect 16937 21568 17068 21608
rect 17108 21568 17117 21608
rect 17296 21568 17305 21608
rect 17345 21568 17354 21608
rect 17410 21568 17419 21608
rect 17459 21568 17468 21608
rect 17514 21568 17644 21608
rect 17685 21568 17694 21608
rect 17740 21568 17810 21608
rect 10330 21558 10388 21559
rect 10003 21484 10012 21524
rect 10052 21484 10061 21524
rect 10483 21484 10492 21524
rect 10532 21484 10732 21524
rect 10772 21484 10781 21524
rect 10012 21440 10052 21484
rect 8044 21400 8812 21440
rect 8852 21400 8861 21440
rect 8995 21400 9004 21440
rect 9044 21400 9716 21440
rect 9955 21400 9964 21440
rect 10004 21400 10052 21440
rect 11692 21440 11732 21568
rect 16588 21524 16628 21568
rect 16684 21524 16724 21568
rect 17428 21524 17468 21568
rect 17770 21524 17810 21568
rect 17914 21599 17972 21608
rect 17914 21559 17923 21599
rect 17963 21559 17972 21599
rect 18883 21568 18892 21608
rect 18932 21568 18941 21608
rect 19721 21568 19852 21608
rect 19892 21568 19901 21608
rect 20227 21568 20236 21608
rect 20276 21568 20285 21608
rect 20506 21568 20515 21608
rect 20555 21568 20716 21608
rect 20756 21568 20765 21608
rect 20969 21568 21100 21608
rect 21140 21568 21149 21608
rect 21466 21568 21475 21608
rect 21515 21568 21868 21608
rect 21908 21568 22444 21608
rect 22484 21568 22493 21608
rect 22627 21568 22636 21608
rect 22676 21568 23596 21608
rect 23636 21568 23645 21608
rect 23770 21568 23779 21608
rect 23819 21568 23876 21608
rect 24067 21568 24076 21608
rect 24137 21568 24247 21608
rect 24394 21568 24403 21608
rect 24443 21568 24452 21608
rect 24538 21599 24652 21608
rect 17914 21558 17972 21559
rect 13673 21484 13795 21524
rect 13844 21484 13853 21524
rect 13987 21484 13996 21524
rect 14036 21484 14188 21524
rect 14228 21484 14237 21524
rect 14633 21484 14764 21524
rect 14804 21484 14947 21524
rect 14987 21484 14996 21524
rect 15401 21484 15523 21524
rect 15572 21484 15581 21524
rect 16099 21484 16108 21524
rect 16148 21484 16628 21524
rect 16675 21484 16684 21524
rect 16724 21484 16733 21524
rect 16867 21484 16876 21524
rect 16916 21484 17187 21524
rect 17227 21484 17236 21524
rect 17391 21484 17468 21524
rect 17530 21484 17539 21524
rect 17588 21484 17719 21524
rect 17770 21484 17836 21524
rect 17876 21484 17885 21524
rect 17391 21440 17431 21484
rect 17932 21440 17972 21558
rect 20236 21524 20276 21568
rect 23836 21524 23876 21568
rect 24538 21559 24547 21599
rect 24587 21568 24652 21599
rect 24692 21568 24727 21608
rect 25097 21568 25123 21608
rect 25163 21568 25228 21608
rect 25268 21568 25804 21608
rect 25844 21568 25853 21608
rect 27305 21568 27427 21608
rect 27476 21568 27485 21608
rect 27724 21568 27811 21608
rect 27851 21568 27860 21608
rect 28771 21568 28780 21608
rect 28820 21568 29923 21608
rect 29963 21568 29972 21608
rect 30298 21568 30307 21608
rect 30347 21568 30988 21608
rect 31028 21568 31037 21608
rect 24587 21559 24596 21568
rect 24538 21558 24596 21559
rect 18019 21484 18028 21524
rect 18068 21484 18604 21524
rect 18644 21484 18653 21524
rect 19075 21484 19084 21524
rect 19124 21484 19459 21524
rect 19499 21484 19508 21524
rect 20236 21484 20620 21524
rect 20660 21484 20669 21524
rect 22752 21484 23500 21524
rect 23540 21484 23549 21524
rect 23836 21484 23884 21524
rect 23924 21484 23933 21524
rect 24259 21484 24268 21524
rect 24308 21484 24460 21524
rect 24500 21484 24509 21524
rect 11692 21400 14668 21440
rect 14708 21400 14717 21440
rect 15907 21400 15916 21440
rect 15956 21400 17431 21440
rect 17923 21400 17932 21440
rect 17972 21400 17981 21440
rect 18508 21400 19220 21440
rect 19267 21400 19276 21440
rect 19316 21400 20716 21440
rect 20756 21400 20765 21440
rect 22819 21400 22828 21440
rect 22868 21400 23404 21440
rect 23444 21400 23453 21440
rect 24041 21400 24172 21440
rect 24212 21400 24221 21440
rect 25001 21400 25095 21440
rect 25172 21400 25181 21440
rect 2057 21316 2188 21356
rect 2228 21316 2237 21356
rect 2476 21316 3050 21356
rect 3130 21316 3139 21356
rect 3179 21316 3436 21356
rect 3476 21316 3485 21356
rect 3802 21316 3811 21356
rect 3851 21316 3860 21356
rect 3916 21316 5164 21356
rect 5204 21316 5213 21356
rect 5731 21316 5740 21356
rect 5780 21316 5972 21356
rect 6787 21316 6796 21356
rect 6836 21316 7084 21356
rect 7124 21316 7133 21356
rect 7363 21316 7372 21356
rect 7412 21316 7459 21356
rect 7499 21316 7543 21356
rect 7612 21316 11692 21356
rect 11732 21316 11741 21356
rect 11971 21316 11980 21356
rect 12020 21316 12460 21356
rect 12500 21316 12509 21356
rect 15715 21316 15724 21356
rect 15764 21316 15895 21356
rect 16579 21316 16588 21356
rect 16628 21316 16876 21356
rect 16916 21316 16925 21356
rect 17059 21316 17068 21356
rect 17108 21316 18364 21356
rect 18404 21316 18413 21356
rect 3820 21188 3860 21316
rect 18508 21272 18548 21400
rect 19075 21316 19084 21356
rect 19124 21316 19133 21356
rect 4291 21232 4300 21272
rect 4340 21232 15148 21272
rect 15188 21232 15197 21272
rect 17731 21232 17740 21272
rect 17780 21232 18548 21272
rect 19084 21188 19124 21316
rect 19180 21272 19220 21400
rect 27628 21356 27668 21504
rect 30144 21484 30796 21524
rect 30836 21484 30845 21524
rect 30307 21400 30316 21440
rect 30356 21400 30508 21440
rect 30548 21400 30557 21440
rect 30761 21400 30892 21440
rect 30932 21400 30941 21440
rect 20899 21316 20908 21356
rect 20948 21316 21388 21356
rect 21428 21316 21437 21356
rect 23657 21316 23779 21356
rect 23828 21316 23837 21356
rect 27628 21316 30604 21356
rect 30644 21316 30653 21356
rect 19180 21232 30508 21272
rect 30548 21232 30557 21272
rect 3103 21148 3112 21188
rect 3480 21148 3489 21188
rect 3715 21148 3724 21188
rect 3764 21148 3860 21188
rect 7843 21148 7852 21188
rect 7892 21148 8236 21188
rect 8276 21148 8285 21188
rect 10877 21148 10886 21188
rect 11254 21148 11263 21188
rect 18651 21148 18660 21188
rect 19028 21148 19037 21188
rect 19084 21148 23308 21188
rect 23348 21148 23357 21188
rect 26425 21148 26434 21188
rect 26802 21148 26811 21188
rect 27235 21148 27244 21188
rect 27284 21148 30316 21188
rect 30356 21148 30365 21188
rect 2947 21064 2956 21104
rect 2996 21064 6028 21104
rect 6068 21064 6077 21104
rect 6316 21064 9100 21104
rect 9140 21064 9149 21104
rect 19843 21064 19852 21104
rect 19892 21064 22924 21104
rect 22964 21064 22973 21104
rect 23020 21064 30452 21104
rect 6316 21020 6356 21064
rect 23020 21020 23060 21064
rect 1891 20980 1900 21020
rect 1940 20980 2228 21020
rect 2188 20936 2228 20980
rect 5404 20980 6124 21020
rect 6164 20980 6173 21020
rect 6307 20980 6316 21020
rect 6356 20980 6365 21020
rect 6700 20980 7372 21020
rect 7412 20980 7564 21020
rect 7604 20980 7613 21020
rect 7747 20980 7756 21020
rect 7796 20980 7939 21020
rect 7979 20980 7988 21020
rect 8995 20980 9004 21020
rect 9044 20980 9053 21020
rect 9187 20980 9196 21020
rect 9236 20980 10348 21020
rect 10388 20980 10397 21020
rect 13219 20980 13228 21020
rect 13268 20980 14764 21020
rect 14804 20980 14868 21020
rect 16771 20980 16780 21020
rect 16820 20980 16829 21020
rect 17827 20980 17836 21020
rect 17876 20980 17885 21020
rect 18115 20980 18124 21020
rect 18164 20980 23060 21020
rect 24547 20980 24556 21020
rect 24596 20980 24605 21020
rect 25097 20980 25228 21020
rect 25268 20980 25277 21020
rect 25996 20980 29740 21020
rect 29780 20980 29789 21020
rect 29945 20980 30028 21020
rect 30068 20980 30076 21020
rect 30116 20980 30125 21020
rect 1673 20896 1804 20936
rect 1844 20896 1853 20936
rect 2170 20896 2179 20936
rect 2219 20896 2228 20936
rect 3340 20896 3916 20936
rect 3956 20896 5012 20936
rect 5059 20896 5068 20936
rect 5108 20896 5164 20936
rect 5204 20896 5239 20936
rect 713 20812 748 20852
rect 788 20812 844 20852
rect 884 20812 893 20852
rect 1066 20843 1132 20852
rect 1066 20803 1075 20843
rect 1115 20812 1132 20843
rect 1172 20812 1255 20852
rect 1315 20812 1324 20852
rect 1364 20812 1556 20852
rect 1891 20812 1900 20852
rect 1940 20812 2083 20852
rect 2132 20812 2606 20852
rect 2650 20812 2659 20852
rect 2708 20812 2839 20852
rect 1115 20803 1124 20812
rect 1066 20802 1124 20803
rect 2566 20768 2606 20812
rect 3340 20768 3380 20896
rect 4972 20852 5012 20896
rect 5404 20852 5444 20980
rect 3593 20843 3724 20852
rect 3593 20812 3667 20843
rect 3658 20803 3667 20812
rect 3707 20812 3724 20843
rect 3764 20812 4148 20852
rect 4972 20812 5395 20852
rect 5435 20812 5444 20852
rect 6076 20896 6412 20936
rect 6452 20896 6461 20936
rect 3707 20803 3716 20812
rect 3658 20802 3716 20803
rect 4108 20768 4148 20812
rect 6076 20768 6116 20896
rect 6700 20852 6740 20980
rect 9004 20936 9044 20980
rect 6787 20896 6796 20936
rect 6836 20896 7013 20936
rect 7075 20896 7084 20936
rect 7124 20896 7133 20936
rect 8044 20896 9044 20936
rect 9763 20896 9772 20936
rect 9812 20896 10348 20936
rect 10388 20896 10397 20936
rect 12796 20896 13132 20936
rect 13172 20896 13181 20936
rect 13228 20896 13324 20936
rect 13364 20896 13373 20936
rect 6207 20812 6220 20852
rect 6260 20812 6281 20852
rect 6241 20768 6281 20812
rect 6604 20812 6740 20852
rect 6604 20768 6644 20812
rect 6973 20768 7013 20896
rect 7084 20768 7124 20896
rect 7267 20812 7276 20852
rect 7316 20812 7447 20852
rect 7756 20812 7948 20852
rect 7988 20812 7997 20852
rect 7756 20768 7796 20812
rect 8044 20779 8084 20896
rect 8131 20812 8140 20852
rect 8180 20812 8756 20852
rect 9257 20812 9388 20852
rect 9428 20812 9437 20852
rect 9859 20812 9868 20852
rect 9908 20812 10004 20852
rect 809 20728 940 20768
rect 980 20728 989 20768
rect 1168 20728 1177 20768
rect 1217 20728 1226 20768
rect 1481 20728 1507 20768
rect 1547 20728 1612 20768
rect 1652 20728 2188 20768
rect 2228 20728 2467 20768
rect 2507 20728 2516 20768
rect 2566 20728 2956 20768
rect 2996 20728 3005 20768
rect 3181 20728 3190 20768
rect 3230 20728 3340 20768
rect 3380 20728 3389 20768
rect 3523 20728 3532 20768
rect 3572 20728 3581 20768
rect 3760 20728 3769 20768
rect 3809 20728 3956 20768
rect 4090 20728 4099 20768
rect 4139 20728 4148 20768
rect 4195 20728 4204 20768
rect 4244 20728 5164 20768
rect 5204 20728 5213 20768
rect 5513 20728 5590 20768
rect 5630 20728 5644 20768
rect 5684 20728 5693 20768
rect 5827 20728 5836 20768
rect 5876 20728 5885 20768
rect 6010 20728 6019 20768
rect 6059 20728 6116 20768
rect 6210 20728 6219 20768
rect 6259 20728 6281 20768
rect 6403 20728 6412 20768
rect 6452 20728 6461 20768
rect 6595 20728 6604 20768
rect 6644 20728 6653 20768
rect 6778 20728 6787 20768
rect 6827 20728 6836 20768
rect 6946 20728 6955 20768
rect 6995 20728 7013 20768
rect 7066 20728 7075 20768
rect 7115 20728 7124 20768
rect 7171 20728 7180 20768
rect 7220 20728 7351 20768
rect 7481 20728 7564 20768
rect 7604 20728 7612 20768
rect 7652 20728 7661 20768
rect 7747 20728 7756 20768
rect 7796 20728 7805 20768
rect 7930 20728 7939 20768
rect 7979 20728 7988 20768
rect 8035 20739 8044 20779
rect 8084 20739 8093 20779
rect 8716 20768 8756 20812
rect 9964 20768 10004 20812
rect 11212 20812 11924 20852
rect 0 20684 400 20704
rect 0 20644 748 20684
rect 788 20644 797 20684
rect 0 20624 400 20644
rect 940 20600 980 20728
rect 1186 20684 1226 20728
rect 3532 20684 3572 20728
rect 3916 20684 3956 20728
rect 4204 20684 4244 20728
rect 1186 20644 2860 20684
rect 2900 20644 2909 20684
rect 3532 20644 3724 20684
rect 3764 20644 3773 20684
rect 3916 20644 4244 20684
rect 5836 20684 5876 20728
rect 5836 20644 6356 20684
rect 940 20560 1340 20600
rect 2371 20560 2380 20600
rect 2420 20560 2995 20600
rect 3035 20560 3044 20600
rect 3427 20560 3436 20600
rect 3476 20560 3916 20600
rect 3956 20560 3965 20600
rect 4483 20560 4492 20600
rect 4532 20560 4780 20600
rect 4820 20560 4829 20600
rect 5923 20560 5932 20600
rect 5972 20560 5981 20600
rect 259 20392 268 20432
rect 308 20392 1132 20432
rect 1172 20392 1181 20432
rect 1300 20348 1340 20560
rect 1411 20476 1420 20516
rect 1460 20476 5588 20516
rect 1699 20392 1708 20432
rect 1748 20392 2764 20432
rect 2804 20392 2813 20432
rect 3427 20392 3436 20432
rect 3476 20392 3668 20432
rect 4343 20392 4352 20432
rect 4720 20392 4729 20432
rect 931 20308 940 20348
rect 980 20308 1172 20348
rect 0 20264 400 20284
rect 1132 20264 1172 20308
rect 1300 20308 2380 20348
rect 2420 20308 2429 20348
rect 2947 20308 2956 20348
rect 2996 20308 3465 20348
rect 0 20224 1076 20264
rect 1123 20224 1132 20264
rect 1172 20224 1181 20264
rect 0 20204 400 20224
rect 1036 20180 1076 20224
rect 960 20140 1036 20180
rect 1076 20140 1085 20180
rect 1300 20096 1340 20308
rect 2179 20224 2188 20264
rect 2228 20224 2371 20264
rect 2411 20224 2420 20264
rect 3425 20180 3465 20308
rect 3628 20264 3668 20392
rect 5548 20348 5588 20476
rect 5932 20432 5972 20560
rect 6316 20432 6356 20644
rect 6412 20516 6452 20728
rect 6796 20684 6836 20728
rect 7948 20684 7988 20728
rect 6499 20644 6508 20684
rect 6548 20644 6836 20684
rect 7843 20644 7852 20684
rect 7892 20644 7988 20684
rect 8140 20728 8189 20768
rect 8229 20728 8238 20768
rect 8314 20728 8323 20768
rect 8363 20728 8372 20768
rect 8491 20728 8500 20768
rect 8540 20728 8549 20768
rect 8698 20728 8707 20768
rect 8747 20728 8756 20768
rect 9545 20728 9676 20768
rect 9716 20728 9725 20768
rect 9859 20728 9868 20768
rect 9908 20728 9917 20768
rect 9964 20728 10156 20768
rect 10196 20728 10205 20768
rect 10889 20728 11020 20768
rect 11060 20728 11069 20768
rect 8140 20600 8180 20728
rect 8332 20684 8372 20728
rect 8323 20644 8332 20684
rect 8372 20644 8419 20684
rect 6691 20560 6700 20600
rect 6740 20560 6988 20600
rect 7028 20560 7037 20600
rect 7337 20560 7459 20600
rect 7508 20560 8180 20600
rect 8509 20516 8549 20728
rect 9868 20684 9908 20728
rect 8995 20644 9004 20684
rect 9055 20644 9175 20684
rect 9868 20644 10484 20684
rect 10531 20644 10540 20684
rect 10580 20644 10964 20684
rect 8681 20560 8803 20600
rect 8852 20560 8861 20600
rect 9091 20560 9100 20600
rect 9140 20560 9148 20600
rect 9188 20560 9271 20600
rect 9763 20560 9772 20600
rect 9812 20560 10003 20600
rect 10043 20560 10052 20600
rect 10444 20516 10484 20644
rect 10924 20600 10964 20644
rect 11212 20600 11252 20812
rect 11884 20768 11924 20812
rect 12796 20810 12836 20896
rect 13228 20852 13268 20896
rect 14668 20852 14708 20980
rect 16780 20936 16820 20980
rect 14755 20896 14764 20936
rect 14804 20896 14860 20936
rect 14900 20896 14935 20936
rect 15340 20896 15532 20936
rect 15572 20896 15581 20936
rect 16780 20896 17452 20936
rect 17492 20896 17501 20936
rect 15340 20852 15380 20896
rect 13036 20812 13268 20852
rect 13388 20812 13397 20852
rect 13437 20812 13460 20852
rect 13507 20812 13516 20852
rect 13556 20812 13601 20852
rect 13699 20812 13708 20852
rect 13748 20812 13791 20852
rect 14083 20812 14092 20852
rect 14132 20812 14284 20852
rect 14324 20812 14333 20852
rect 14668 20812 14860 20852
rect 14900 20812 14909 20852
rect 15017 20812 15052 20852
rect 15092 20812 15139 20852
rect 15179 20812 15197 20852
rect 15331 20812 15340 20852
rect 15380 20812 15389 20852
rect 16270 20812 16396 20852
rect 16436 20812 16445 20852
rect 16492 20812 16780 20852
rect 16820 20812 16829 20852
rect 12787 20770 12796 20810
rect 12836 20770 12845 20810
rect 13036 20768 13076 20812
rect 11587 20728 11596 20768
rect 11636 20728 11704 20768
rect 11744 20728 11767 20768
rect 11863 20728 11872 20768
rect 11912 20728 11924 20768
rect 12028 20728 12322 20768
rect 12362 20728 12371 20768
rect 12922 20728 12931 20768
rect 12971 20728 12980 20768
rect 13027 20728 13036 20768
rect 13076 20728 13085 20768
rect 13193 20728 13291 20768
rect 13364 20728 13373 20768
rect 12028 20600 12068 20728
rect 12940 20684 12980 20728
rect 13420 20684 13460 20812
rect 13516 20768 13556 20812
rect 13751 20768 13791 20812
rect 16270 20768 16310 20812
rect 16492 20768 16532 20812
rect 16876 20768 16916 20896
rect 17836 20852 17876 20980
rect 24556 20936 24596 20980
rect 18403 20896 18412 20936
rect 18452 20896 19316 20936
rect 17059 20812 17068 20852
rect 17108 20812 17251 20852
rect 17300 20812 17309 20852
rect 17818 20812 17827 20852
rect 17867 20812 17876 20852
rect 18010 20812 18019 20852
rect 18059 20812 18115 20852
rect 18473 20812 18595 20852
rect 18644 20812 18653 20852
rect 18028 20768 18068 20812
rect 19276 20810 19316 20896
rect 19258 20801 19316 20810
rect 13505 20728 13514 20768
rect 13554 20728 13563 20768
rect 13742 20728 13751 20768
rect 13791 20728 13800 20768
rect 13882 20728 13891 20768
rect 13931 20728 13940 20768
rect 13987 20728 13996 20768
rect 14036 20728 14167 20768
rect 14371 20728 14380 20768
rect 14420 20728 14467 20768
rect 14507 20728 14551 20768
rect 14851 20728 14860 20768
rect 14900 20728 14999 20768
rect 15039 20728 15048 20768
rect 15235 20728 15244 20768
rect 15284 20728 15415 20768
rect 16003 20728 16012 20768
rect 16052 20728 16120 20768
rect 16160 20728 16183 20768
rect 16270 20728 16295 20768
rect 16335 20728 16344 20768
rect 16474 20728 16483 20768
rect 16523 20728 16532 20768
rect 16596 20728 16684 20768
rect 16724 20728 16727 20768
rect 16767 20728 16776 20768
rect 16858 20728 16867 20768
rect 16907 20728 16916 20768
rect 16963 20728 16972 20768
rect 17012 20728 17143 20768
rect 17443 20728 17452 20768
rect 17492 20728 17635 20768
rect 17675 20728 17684 20768
rect 18019 20728 18028 20768
rect 18068 20728 18077 20768
rect 18281 20728 18403 20768
rect 18452 20728 18461 20768
rect 18730 20728 18739 20768
rect 18779 20728 18788 20768
rect 19258 20761 19267 20801
rect 19307 20761 19316 20801
rect 20140 20896 20332 20936
rect 20372 20896 20381 20936
rect 20794 20896 20803 20936
rect 20843 20896 20852 20936
rect 20140 20768 20180 20896
rect 20812 20852 20852 20896
rect 20297 20812 20428 20852
rect 20468 20812 20852 20852
rect 20908 20896 24364 20936
rect 24404 20896 24413 20936
rect 24556 20896 25132 20936
rect 25172 20896 25612 20936
rect 25652 20896 25661 20936
rect 19258 20760 19316 20761
rect 20024 20728 20033 20768
rect 20073 20728 20180 20768
rect 20332 20768 20372 20812
rect 20908 20768 20948 20896
rect 21196 20812 21812 20852
rect 20489 20728 20620 20768
rect 20660 20728 20948 20768
rect 21004 20801 21128 20810
rect 21004 20770 21088 20801
rect 13900 20684 13940 20728
rect 14999 20684 15039 20728
rect 12893 20644 12940 20684
rect 12980 20644 12989 20684
rect 13097 20644 13123 20684
rect 13163 20644 13228 20684
rect 13268 20644 13277 20684
rect 13411 20644 13420 20684
rect 13460 20644 13469 20684
rect 13900 20644 14036 20684
rect 14999 20644 15916 20684
rect 15995 20644 18316 20684
rect 18356 20644 18365 20684
rect 13996 20600 14036 20644
rect 18748 20600 18788 20728
rect 20332 20719 20372 20728
rect 21004 20684 21044 20770
rect 21196 20768 21236 20812
rect 21772 20768 21812 20812
rect 22060 20812 22732 20852
rect 22772 20812 22781 20852
rect 22915 20812 22924 20852
rect 22964 20812 23203 20852
rect 23243 20812 24556 20852
rect 24596 20812 24605 20852
rect 21088 20752 21128 20761
rect 21178 20728 21187 20768
rect 21227 20728 21236 20768
rect 21283 20728 21292 20768
rect 21332 20728 21661 20768
rect 21701 20728 21716 20768
rect 21763 20728 21772 20768
rect 21812 20728 21964 20768
rect 22004 20728 22013 20768
rect 21676 20684 21716 20728
rect 22060 20684 22100 20812
rect 25996 20768 26036 20980
rect 27113 20896 27244 20936
rect 27284 20896 27293 20936
rect 29923 20896 29932 20936
rect 29972 20896 30260 20936
rect 30220 20852 30260 20896
rect 30412 20852 30452 21064
rect 30499 20980 30508 21020
rect 30548 20980 30604 21020
rect 30644 20980 30679 21020
rect 30761 20896 30892 20936
rect 30932 20896 30941 20936
rect 29376 20812 29548 20852
rect 29588 20812 29597 20852
rect 30220 20812 30316 20852
rect 30356 20812 30365 20852
rect 30412 20812 30740 20852
rect 30700 20768 30740 20812
rect 22217 20728 22348 20768
rect 22388 20728 22397 20768
rect 22458 20728 22467 20768
rect 22507 20728 22516 20768
rect 22576 20728 22585 20768
rect 22625 20728 22636 20768
rect 22676 20728 22765 20768
rect 23273 20728 23308 20768
rect 23348 20728 23404 20768
rect 23444 20728 23453 20768
rect 23587 20728 23596 20768
rect 23675 20728 23767 20768
rect 23827 20728 23836 20768
rect 23876 20728 24172 20768
rect 24212 20728 24259 20768
rect 24299 20728 24652 20768
rect 24692 20728 24931 20768
rect 24971 20728 24980 20768
rect 25233 20728 25242 20768
rect 25282 20728 26036 20768
rect 26083 20728 26092 20768
rect 26132 20728 26263 20768
rect 26371 20728 26380 20768
rect 26420 20728 26429 20768
rect 26956 20728 27532 20768
rect 27572 20728 27581 20768
rect 29033 20728 29155 20768
rect 29204 20728 29213 20768
rect 29445 20728 29740 20768
rect 29780 20728 29789 20768
rect 29923 20728 29932 20768
rect 29972 20728 30103 20768
rect 30377 20728 30508 20768
rect 30548 20728 30557 20768
rect 30691 20728 30700 20768
rect 30740 20728 30749 20768
rect 19411 20644 19420 20684
rect 19460 20644 19564 20684
rect 19604 20644 19613 20684
rect 19747 20644 19756 20684
rect 19796 20644 20276 20684
rect 21004 20644 21580 20684
rect 21620 20644 21629 20684
rect 21676 20644 22100 20684
rect 22467 20684 22507 20728
rect 26380 20684 26420 20728
rect 22467 20644 22732 20684
rect 22772 20644 22781 20684
rect 24233 20644 24364 20684
rect 24404 20644 24413 20684
rect 24561 20644 24570 20684
rect 24610 20644 25844 20684
rect 25891 20644 25900 20684
rect 25940 20644 26420 20684
rect 20236 20600 20276 20644
rect 25804 20600 25844 20644
rect 26956 20600 26996 20728
rect 29445 20684 29485 20728
rect 27043 20644 27052 20684
rect 27092 20644 28108 20684
rect 28148 20644 28157 20684
rect 28963 20644 28972 20684
rect 29012 20644 29485 20684
rect 29530 20644 29539 20684
rect 29579 20644 30220 20684
rect 30260 20644 30269 20684
rect 10906 20560 10915 20600
rect 10955 20560 10964 20600
rect 11203 20560 11212 20600
rect 11252 20560 11261 20600
rect 11465 20560 11539 20600
rect 11579 20560 11596 20600
rect 11636 20560 11645 20600
rect 11875 20560 11884 20600
rect 11924 20560 12028 20600
rect 12068 20560 12077 20600
rect 12499 20560 12508 20600
rect 12548 20560 12844 20600
rect 12884 20560 12893 20600
rect 13594 20560 13603 20600
rect 13643 20560 13900 20600
rect 13940 20560 13949 20600
rect 13996 20560 15724 20600
rect 15764 20560 15773 20600
rect 16387 20560 16396 20600
rect 16436 20560 17164 20600
rect 17204 20560 17213 20600
rect 17338 20560 17347 20600
rect 17387 20560 17932 20600
rect 17972 20560 17981 20600
rect 18106 20560 18115 20600
rect 18164 20560 18788 20600
rect 18931 20560 18940 20600
rect 18980 20560 18988 20600
rect 19028 20560 19111 20600
rect 19267 20560 19276 20600
rect 19316 20560 20131 20600
rect 20171 20560 20180 20600
rect 20227 20560 20236 20600
rect 20276 20560 20407 20600
rect 20467 20560 20476 20600
rect 20516 20560 20525 20600
rect 21185 20560 21292 20600
rect 21347 20560 21365 20600
rect 21466 20560 21475 20600
rect 21515 20560 21524 20600
rect 21667 20560 21676 20600
rect 21716 20560 22252 20600
rect 22292 20560 22636 20600
rect 22676 20560 22685 20600
rect 24905 20560 25027 20600
rect 25076 20560 25085 20600
rect 25289 20560 25420 20600
rect 25460 20560 25469 20600
rect 25804 20560 26996 20600
rect 20476 20516 20516 20560
rect 6412 20476 8140 20516
rect 8180 20476 8189 20516
rect 8509 20476 9388 20516
rect 9428 20476 9676 20516
rect 9716 20476 9725 20516
rect 10444 20476 21388 20516
rect 21428 20476 21437 20516
rect 9676 20432 9716 20476
rect 5932 20392 6220 20432
rect 6260 20392 6269 20432
rect 6316 20392 8620 20432
rect 8660 20392 8669 20432
rect 9676 20392 11884 20432
rect 11924 20392 11933 20432
rect 12117 20392 12126 20432
rect 12494 20392 12503 20432
rect 13324 20392 17068 20432
rect 17108 20392 17117 20432
rect 18979 20392 18988 20432
rect 19028 20392 19660 20432
rect 19700 20392 19709 20432
rect 19891 20392 19900 20432
rect 20268 20392 20277 20432
rect 13324 20348 13364 20392
rect 4060 20308 5068 20348
rect 5108 20308 5117 20348
rect 5405 20308 5452 20348
rect 5492 20308 5501 20348
rect 5548 20308 13364 20348
rect 13411 20308 13420 20348
rect 13460 20308 13748 20348
rect 13795 20308 13804 20348
rect 13844 20308 14132 20348
rect 15139 20308 15148 20348
rect 15188 20308 20620 20348
rect 20660 20308 20669 20348
rect 4060 20264 4100 20308
rect 5452 20264 5492 20308
rect 3619 20224 3628 20264
rect 3668 20224 3677 20264
rect 4051 20224 4060 20264
rect 4100 20224 4109 20264
rect 4588 20224 4916 20264
rect 5434 20224 5443 20264
rect 5483 20224 5492 20264
rect 5548 20224 6559 20264
rect 7651 20224 7660 20264
rect 7700 20224 8660 20264
rect 8899 20224 8908 20264
rect 8948 20224 9338 20264
rect 9449 20224 9571 20264
rect 9620 20224 9629 20264
rect 10435 20224 10444 20264
rect 10484 20224 10493 20264
rect 10627 20224 10636 20264
rect 10676 20224 11153 20264
rect 11875 20224 11884 20264
rect 11924 20224 13652 20264
rect 4588 20180 4628 20224
rect 1594 20140 1603 20180
rect 1643 20140 3244 20180
rect 3284 20140 3293 20180
rect 3416 20140 3425 20180
rect 3465 20140 3474 20180
rect 4108 20140 4628 20180
rect 4876 20180 4916 20224
rect 5548 20180 5588 20224
rect 6519 20222 6559 20224
rect 6519 20182 6616 20222
rect 6656 20182 6665 20222
rect 8620 20180 8660 20224
rect 9298 20180 9338 20224
rect 10444 20180 10484 20224
rect 4876 20140 5068 20180
rect 5108 20140 5117 20180
rect 5443 20140 5452 20180
rect 5492 20140 5588 20180
rect 6844 20140 7267 20180
rect 7307 20140 7695 20180
rect 8035 20140 8044 20180
rect 8084 20140 8564 20180
rect 8620 20140 9148 20180
rect 9188 20140 9197 20180
rect 9298 20140 9524 20180
rect 9667 20140 9676 20180
rect 9716 20140 9783 20180
rect 9823 20140 9847 20180
rect 9955 20140 9964 20180
rect 10004 20140 10484 20180
rect 10684 20140 10924 20180
rect 10964 20140 10973 20180
rect 4108 20096 4148 20140
rect 6844 20138 6884 20140
rect 5818 20098 5827 20138
rect 5867 20098 6068 20138
rect 835 20056 844 20096
rect 884 20056 893 20096
rect 1108 20093 1132 20096
rect 844 19928 884 20056
rect 977 20053 986 20093
rect 1026 20056 1132 20093
rect 1172 20056 1181 20096
rect 1282 20056 1291 20096
rect 1331 20056 1340 20096
rect 1508 20056 1517 20096
rect 1557 20056 1603 20096
rect 1673 20056 1771 20096
rect 1844 20056 1853 20096
rect 1961 20056 1996 20096
rect 2036 20056 2092 20096
rect 2132 20056 2141 20096
rect 2266 20056 2275 20096
rect 2315 20056 2324 20096
rect 2563 20056 2572 20096
rect 2623 20056 2743 20096
rect 2860 20056 3052 20096
rect 3092 20056 3101 20096
rect 3280 20056 3289 20096
rect 3329 20056 3340 20096
rect 3380 20056 3469 20096
rect 3593 20056 3724 20096
rect 3764 20056 3773 20096
rect 3907 20056 3916 20096
rect 3956 20056 4148 20096
rect 4195 20056 4204 20096
rect 4244 20056 4253 20096
rect 4378 20056 4387 20096
rect 4427 20056 4436 20096
rect 4483 20056 4492 20096
rect 4532 20056 4535 20096
rect 4575 20056 4663 20096
rect 4771 20056 4780 20096
rect 4820 20056 4829 20096
rect 4876 20056 5092 20096
rect 5132 20056 5141 20096
rect 5242 20056 5251 20096
rect 5291 20056 5300 20096
rect 1026 20053 1148 20056
rect 1300 19928 1340 20056
rect 1516 20012 1556 20056
rect 2284 20012 2324 20056
rect 1402 19972 1411 20012
rect 1451 19972 1460 20012
rect 1507 19972 1516 20012
rect 1556 19972 1565 20012
rect 1699 19972 1708 20012
rect 1748 19972 1891 20012
rect 1931 19972 1940 20012
rect 2083 19972 2092 20012
rect 2132 19972 2324 20012
rect 844 19888 1340 19928
rect 1420 19928 1460 19972
rect 2860 19928 2900 20056
rect 3724 20038 3764 20047
rect 4204 20012 4244 20056
rect 4396 20012 4436 20056
rect 2947 19972 2956 20012
rect 2996 19972 3127 20012
rect 3178 20003 3236 20012
rect 3178 19963 3187 20003
rect 3227 19963 3236 20003
rect 3811 19972 3820 20012
rect 3860 19972 4012 20012
rect 4052 19972 4244 20012
rect 4349 19972 4396 20012
rect 4436 19972 4445 20012
rect 4553 19972 4675 20012
rect 4724 19972 4733 20012
rect 3178 19962 3236 19963
rect 1420 19888 1652 19928
rect 2083 19888 2092 19928
rect 2132 19888 2900 19928
rect 0 19844 400 19864
rect 1612 19844 1652 19888
rect 3196 19844 3236 19962
rect 4204 19928 4244 19972
rect 4780 19928 4820 20056
rect 4876 20012 4916 20056
rect 5260 20012 5300 20056
rect 4867 19972 4876 20012
rect 4916 19972 4925 20012
rect 5155 19972 5164 20012
rect 5204 19972 5300 20012
rect 5356 20056 5368 20096
rect 5408 20056 5417 20096
rect 5530 20056 5539 20096
rect 5579 20056 5588 20096
rect 5652 20056 5661 20096
rect 5701 20056 5727 20096
rect 5356 19928 5396 20056
rect 5548 20012 5588 20056
rect 5687 20012 5727 20056
rect 5501 19972 5548 20012
rect 5588 19972 5597 20012
rect 5687 19972 5740 20012
rect 5780 19972 5789 20012
rect 5836 19928 5876 20098
rect 6028 20096 6068 20098
rect 6167 20098 6403 20138
rect 6443 20098 6452 20138
rect 6826 20098 6835 20138
rect 6875 20098 6884 20138
rect 6167 20096 6207 20098
rect 7655 20096 7695 20140
rect 8524 20096 8564 20140
rect 9484 20096 9524 20140
rect 10684 20096 10724 20140
rect 11113 20096 11153 20224
rect 12425 20140 12460 20180
rect 12500 20140 12556 20180
rect 12596 20140 12605 20180
rect 12970 20140 12979 20180
rect 13019 20140 13036 20180
rect 13076 20140 13159 20180
rect 13251 20140 13324 20180
rect 13364 20140 13373 20180
rect 13251 20096 13291 20140
rect 13612 20096 13652 20224
rect 13708 20096 13748 20308
rect 14092 20264 14132 20308
rect 21484 20264 21524 20560
rect 23491 20476 23500 20516
rect 23540 20476 30412 20516
rect 30452 20476 30461 20516
rect 27665 20392 27674 20432
rect 28042 20392 28051 20432
rect 21571 20308 21580 20348
rect 21620 20308 22196 20348
rect 13795 20224 13804 20264
rect 13844 20224 14022 20264
rect 14074 20224 14083 20264
rect 14123 20224 14132 20264
rect 14476 20224 14563 20264
rect 14603 20224 14612 20264
rect 15532 20224 15724 20264
rect 15764 20224 15773 20264
rect 16099 20224 16108 20264
rect 16148 20224 16483 20264
rect 16523 20224 16532 20264
rect 16588 20224 16876 20264
rect 16916 20224 17260 20264
rect 17300 20224 17309 20264
rect 17452 20224 17836 20264
rect 17876 20224 17885 20264
rect 18595 20224 18604 20264
rect 18644 20224 18691 20264
rect 18731 20224 18775 20264
rect 19555 20224 19564 20264
rect 19604 20224 19700 20264
rect 19747 20224 19756 20264
rect 19796 20224 19852 20264
rect 19892 20224 19927 20264
rect 20236 20224 21388 20264
rect 21428 20224 21437 20264
rect 21484 20224 21580 20264
rect 21620 20224 22004 20264
rect 13982 20180 14022 20224
rect 14476 20180 14516 20224
rect 15532 20180 15572 20224
rect 13982 20140 14188 20180
rect 14228 20140 14237 20180
rect 14284 20140 14516 20180
rect 14563 20140 14572 20180
rect 14612 20140 15134 20180
rect 15174 20140 15572 20180
rect 16195 20140 16204 20180
rect 16244 20140 16253 20180
rect 6028 20056 6207 20096
rect 6691 20056 6700 20096
rect 6740 20056 6749 20096
rect 6931 20056 6940 20096
rect 6980 20056 6989 20096
rect 7171 20056 7180 20096
rect 7220 20056 7351 20096
rect 7433 20056 7468 20096
rect 7508 20056 7564 20096
rect 7604 20056 7613 20096
rect 7655 20056 7683 20096
rect 7723 20056 7732 20096
rect 7792 20056 7801 20096
rect 7841 20056 7892 20096
rect 7939 20056 7948 20096
rect 7988 20056 8035 20096
rect 8131 20056 8140 20096
rect 8180 20056 8189 20096
rect 8270 20056 8279 20096
rect 8319 20056 8332 20096
rect 8372 20056 8450 20096
rect 8515 20056 8524 20096
rect 8564 20056 8573 20096
rect 8707 20056 8716 20096
rect 8756 20056 8812 20096
rect 8852 20056 8887 20096
rect 8995 20056 9004 20096
rect 9044 20056 9175 20096
rect 9283 20056 9292 20096
rect 9332 20056 9341 20096
rect 9466 20056 9475 20096
rect 9515 20056 9524 20096
rect 10147 20056 10156 20096
rect 10196 20056 10205 20096
rect 10339 20056 10348 20096
rect 10388 20056 10539 20096
rect 10579 20056 10588 20096
rect 10650 20056 10659 20096
rect 10699 20056 10724 20096
rect 10768 20056 10777 20096
rect 10817 20056 10868 20096
rect 11011 20056 11020 20096
rect 11060 20056 11070 20096
rect 11113 20056 11139 20096
rect 11179 20056 11188 20096
rect 11248 20056 11257 20096
rect 11297 20056 11596 20096
rect 11636 20056 11645 20096
rect 11849 20056 11980 20096
rect 12020 20056 12029 20096
rect 12233 20056 12355 20096
rect 12404 20056 12413 20096
rect 12657 20056 12666 20096
rect 12706 20056 12844 20096
rect 12884 20056 12893 20096
rect 13165 20056 13174 20096
rect 13214 20056 13291 20096
rect 13363 20056 13372 20096
rect 13412 20056 13421 20096
rect 13484 20056 13493 20096
rect 13533 20056 13542 20096
rect 13603 20056 13612 20096
rect 13652 20056 13661 20096
rect 13708 20056 13982 20096
rect 14022 20056 14188 20096
rect 14228 20056 14237 20096
rect 14284 20087 14324 20140
rect 14572 20096 14612 20140
rect 16204 20096 16244 20140
rect 16588 20096 16628 20224
rect 16963 20140 16972 20180
rect 17012 20140 17143 20180
rect 16786 20101 16922 20102
rect 5923 20014 5932 20054
rect 5972 20014 5981 20054
rect 6250 20014 6259 20054
rect 6299 20014 6308 20054
rect 6519 20014 6536 20054
rect 6576 20014 6585 20054
rect 4204 19888 4532 19928
rect 4780 19888 5068 19928
rect 5108 19888 5117 19928
rect 5356 19888 5836 19928
rect 5876 19888 5885 19928
rect 4492 19844 4532 19888
rect 0 19804 1420 19844
rect 1460 19804 1469 19844
rect 1612 19804 1708 19844
rect 1748 19804 1757 19844
rect 2179 19804 2188 19844
rect 2228 19804 2572 19844
rect 2612 19804 2621 19844
rect 3010 19804 3236 19844
rect 3331 19804 3340 19844
rect 3380 19804 3427 19844
rect 3467 19804 3511 19844
rect 4378 19804 4387 19844
rect 4427 19804 4436 19844
rect 4492 19804 5740 19844
rect 5780 19804 5789 19844
rect 0 19784 400 19804
rect 3010 19592 3050 19804
rect 4396 19760 4436 19804
rect 4396 19720 5356 19760
rect 5396 19720 5405 19760
rect 3103 19636 3112 19676
rect 3480 19636 3489 19676
rect 3010 19552 3668 19592
rect 3628 19508 3668 19552
rect 1036 19468 3139 19508
rect 3179 19468 3188 19508
rect 3610 19468 3619 19508
rect 3659 19468 3668 19508
rect 0 19424 400 19444
rect 0 19384 460 19424
rect 500 19384 509 19424
rect 0 19364 400 19384
rect 1036 19340 1076 19468
rect 2371 19384 2380 19424
rect 2420 19384 2804 19424
rect 1018 19300 1027 19340
rect 1067 19300 1076 19340
rect 1219 19300 1228 19340
rect 1268 19300 1420 19340
rect 1460 19300 1469 19340
rect 1987 19300 1996 19340
rect 2036 19300 2188 19340
rect 2228 19300 2572 19340
rect 2612 19300 2621 19340
rect 2764 19256 2804 19384
rect 3916 19384 5356 19424
rect 5396 19384 5405 19424
rect 2851 19300 2860 19340
rect 2900 19300 3035 19340
rect 2995 19256 3035 19300
rect 3436 19256 3476 19265
rect 3916 19256 3956 19384
rect 5932 19340 5972 20014
rect 6115 19972 6124 20012
rect 6164 19972 6207 20012
rect 6019 19888 6028 19928
rect 6068 19888 6077 19928
rect 6028 19844 6068 19888
rect 6019 19804 6028 19844
rect 6068 19804 6115 19844
rect 6167 19760 6207 19972
rect 6028 19720 6207 19760
rect 6028 19676 6068 19720
rect 6019 19636 6028 19676
rect 6068 19636 6077 19676
rect 6263 19508 6303 20014
rect 6519 20012 6559 20014
rect 6700 20012 6740 20056
rect 6940 20012 6980 20056
rect 6403 19972 6412 20012
rect 6452 19972 6559 20012
rect 6653 19972 6693 20012
rect 6733 19972 6742 20012
rect 6898 19972 6980 20012
rect 7066 19972 7075 20012
rect 7124 19972 7255 20012
rect 7337 19972 7372 20012
rect 7412 19972 7468 20012
rect 7508 19972 7517 20012
rect 6898 19928 6938 19972
rect 6595 19888 6604 19928
rect 6644 19888 6938 19928
rect 7852 19844 7892 20056
rect 7948 20012 7988 20056
rect 7939 19972 7948 20012
rect 7988 19972 7997 20012
rect 8140 19928 8180 20056
rect 9292 20012 9332 20056
rect 9783 20014 9916 20054
rect 9956 20014 9965 20054
rect 9783 20012 9823 20014
rect 8410 19972 8419 20012
rect 8459 19972 8468 20012
rect 8611 19972 8620 20012
rect 8660 19972 9332 20012
rect 9676 19972 9823 20012
rect 10042 19972 10051 20012
rect 10091 19972 10100 20012
rect 8035 19888 8044 19928
rect 8084 19888 8180 19928
rect 8428 19928 8468 19972
rect 8428 19888 8948 19928
rect 8428 19844 8468 19888
rect 7267 19804 7276 19844
rect 7316 19804 8468 19844
rect 8681 19804 8812 19844
rect 8852 19804 8861 19844
rect 8908 19760 8948 19888
rect 9676 19760 9716 19972
rect 10060 19928 10100 19972
rect 10013 19888 10060 19928
rect 10100 19888 10109 19928
rect 10156 19844 10196 20056
rect 10348 20053 10436 20056
rect 10828 20012 10868 20056
rect 11030 20012 11070 20056
rect 13372 20012 13412 20056
rect 10243 19972 10252 20012
rect 10292 19972 10303 20012
rect 10819 19972 10828 20012
rect 10868 19972 10877 20012
rect 11030 19972 11116 20012
rect 11156 19972 11165 20012
rect 12652 19972 13412 20012
rect 13493 20012 13533 20056
rect 14456 20056 14465 20096
rect 14505 20056 14612 20096
rect 14659 20056 14668 20096
rect 14708 20056 14717 20096
rect 14764 20087 14804 20096
rect 14284 20038 14324 20047
rect 14668 20012 14708 20056
rect 13493 19972 13900 20012
rect 13940 19972 13949 20012
rect 14371 19972 14380 20012
rect 14420 19972 14708 20012
rect 15209 20056 15244 20096
rect 15284 20056 15340 20096
rect 15380 20056 15389 20096
rect 15436 20087 15532 20096
rect 14764 20012 14804 20047
rect 15476 20056 15532 20087
rect 15572 20056 15607 20096
rect 15785 20056 15883 20096
rect 15956 20056 15965 20096
rect 16097 20056 16106 20096
rect 16146 20056 16155 20096
rect 16204 20056 16387 20096
rect 16427 20056 16436 20096
rect 16588 20056 16695 20096
rect 16735 20056 16744 20096
rect 16786 20062 16877 20101
rect 15436 20038 15476 20047
rect 14764 19972 15148 20012
rect 15188 19972 15197 20012
rect 15881 19972 16003 20012
rect 16052 19972 16061 20012
rect 10263 19928 10303 19972
rect 10263 19888 10444 19928
rect 10484 19888 10493 19928
rect 12652 19844 12692 19972
rect 14668 19928 14708 19972
rect 14668 19888 15244 19928
rect 15284 19888 15293 19928
rect 9763 19804 9772 19844
rect 9812 19804 10196 19844
rect 11465 19804 11587 19844
rect 11636 19804 11645 19844
rect 12643 19804 12652 19844
rect 12692 19804 12701 19844
rect 14563 19804 14572 19844
rect 14612 19804 15139 19844
rect 15179 19804 15188 19844
rect 16108 19760 16148 20056
rect 16786 20012 16826 20062
rect 16868 20061 16877 20062
rect 16917 20061 16926 20101
rect 17452 20096 17492 20224
rect 19660 20180 19700 20224
rect 20236 20180 20276 20224
rect 18144 20140 18220 20180
rect 18260 20140 18269 20180
rect 19229 20140 19276 20180
rect 19316 20140 19325 20180
rect 19546 20140 19555 20180
rect 19595 20140 19604 20180
rect 19660 20140 20276 20180
rect 20323 20140 20332 20180
rect 20372 20140 20448 20180
rect 20515 20140 20524 20180
rect 20564 20140 20852 20180
rect 18220 20096 18260 20140
rect 19276 20096 19316 20140
rect 19564 20096 19604 20140
rect 20332 20096 20372 20140
rect 20812 20096 20852 20140
rect 17129 20056 17178 20096
rect 17218 20056 17260 20096
rect 17300 20056 17309 20096
rect 17443 20056 17452 20096
rect 17492 20056 17501 20096
rect 17801 20056 17827 20096
rect 17867 20056 17932 20096
rect 17972 20056 17981 20096
rect 18106 20056 18115 20096
rect 18155 20056 18260 20096
rect 18307 20056 18316 20096
rect 18356 20056 18359 20096
rect 18399 20056 18487 20096
rect 18595 20056 18604 20096
rect 18644 20056 18653 20096
rect 18700 20056 19084 20096
rect 19124 20056 19133 20096
rect 19258 20056 19267 20096
rect 19307 20056 19316 20096
rect 19363 20056 19372 20096
rect 19412 20056 19604 20096
rect 19747 20056 19756 20096
rect 19796 20056 19805 20096
rect 19891 20056 19900 20096
rect 19940 20056 20372 20096
rect 20419 20056 20428 20096
rect 20468 20056 20599 20096
rect 20803 20056 20812 20096
rect 20852 20056 20861 20096
rect 21562 20056 21571 20096
rect 21611 20056 21620 20096
rect 21667 20056 21676 20096
rect 21716 20056 21847 20096
rect 16195 19972 16204 20012
rect 16244 19972 16253 20012
rect 16675 19972 16684 20012
rect 16724 19972 16826 20012
rect 17068 19972 17644 20012
rect 17684 19972 17693 20012
rect 18019 19972 18028 20012
rect 18068 19972 18220 20012
rect 18260 19972 18269 20012
rect 18490 19972 18499 20012
rect 18539 19972 18548 20012
rect 16204 19928 16244 19972
rect 17068 19928 17108 19972
rect 16204 19888 17108 19928
rect 17299 19888 17308 19928
rect 17348 19888 17356 19928
rect 17396 19888 17479 19928
rect 18508 19844 18548 19972
rect 16675 19804 16684 19844
rect 16724 19804 16876 19844
rect 16916 19804 16925 19844
rect 17155 19804 17164 19844
rect 17204 19804 18548 19844
rect 18604 19760 18644 20056
rect 18700 20012 18740 20056
rect 18691 19972 18700 20012
rect 18740 19972 18749 20012
rect 8908 19720 12556 19760
rect 12596 19720 12605 19760
rect 15340 19720 15820 19760
rect 15860 19720 15869 19760
rect 16108 19720 17644 19760
rect 17684 19720 17932 19760
rect 17972 19720 18644 19760
rect 18988 19760 19028 20056
rect 19756 20012 19796 20056
rect 20428 20012 20468 20056
rect 19075 19972 19084 20012
rect 19124 19972 19564 20012
rect 19604 19972 19613 20012
rect 19756 19972 20468 20012
rect 21580 20012 21620 20056
rect 21964 20012 22004 20224
rect 22156 20180 22196 20308
rect 28588 20308 30700 20348
rect 30740 20308 30749 20348
rect 28588 20264 28628 20308
rect 23971 20224 23980 20264
rect 24020 20224 24364 20264
rect 24404 20224 24413 20264
rect 24460 20224 27244 20264
rect 27284 20224 27293 20264
rect 27340 20224 28628 20264
rect 28867 20224 28876 20264
rect 28916 20224 29932 20264
rect 29972 20224 29981 20264
rect 24460 20180 24500 20224
rect 27340 20180 27380 20224
rect 22138 20140 22147 20180
rect 22187 20140 22732 20180
rect 22772 20140 22781 20180
rect 23692 20140 23884 20180
rect 23924 20140 23933 20180
rect 23980 20140 24500 20180
rect 25123 20140 25132 20180
rect 25172 20140 25420 20180
rect 25460 20140 25469 20180
rect 25603 20140 25612 20180
rect 25652 20140 27380 20180
rect 27628 20140 29164 20180
rect 29204 20140 29212 20180
rect 29252 20140 29261 20180
rect 30211 20140 30220 20180
rect 30260 20140 30268 20180
rect 30308 20140 30391 20180
rect 23692 20096 23732 20140
rect 22426 20056 22435 20096
rect 22475 20056 22772 20096
rect 23107 20056 23116 20096
rect 23156 20056 23287 20096
rect 23683 20056 23692 20096
rect 23732 20056 23741 20096
rect 23931 20056 23940 20096
rect 23980 20056 24020 20140
rect 27628 20096 27668 20140
rect 24067 20056 24076 20096
rect 24116 20056 24119 20096
rect 24159 20056 24247 20096
rect 24355 20056 24364 20096
rect 24404 20056 24535 20096
rect 24739 20056 24748 20096
rect 24788 20056 24919 20096
rect 25018 20056 25027 20096
rect 25067 20056 25076 20096
rect 26275 20056 26284 20096
rect 26324 20056 27619 20096
rect 27659 20056 27668 20096
rect 28073 20056 28204 20096
rect 28244 20056 28253 20096
rect 28300 20087 29068 20096
rect 28300 20056 29059 20087
rect 29108 20056 29117 20096
rect 29827 20056 29836 20096
rect 29876 20056 30412 20096
rect 30452 20056 30461 20096
rect 21580 19972 21716 20012
rect 21964 19972 22051 20012
rect 22091 19972 22100 20012
rect 22505 19972 22627 20012
rect 22676 19972 22685 20012
rect 19145 19888 19276 19928
rect 19316 19888 19325 19928
rect 20323 19888 20332 19928
rect 20372 19888 21004 19928
rect 21044 19888 21053 19928
rect 21676 19844 21716 19972
rect 21763 19888 21772 19928
rect 21812 19888 21868 19928
rect 21908 19888 21943 19928
rect 22732 19844 22772 20056
rect 23806 20014 23815 20054
rect 23855 20014 23871 20054
rect 23831 20012 23871 20014
rect 25036 20012 25076 20056
rect 28300 20012 28340 20056
rect 29050 20047 29059 20056
rect 29099 20047 29108 20056
rect 29050 20046 29108 20047
rect 23017 19972 23026 20012
rect 23066 19972 23732 20012
rect 23831 19972 24172 20012
rect 24212 19972 24259 20012
rect 24299 19972 24343 20012
rect 24451 19972 24460 20012
rect 24500 19972 25076 20012
rect 27331 19972 27340 20012
rect 27380 19972 27389 20012
rect 27977 19972 28003 20012
rect 28043 19972 28108 20012
rect 28148 19972 28157 20012
rect 28201 19972 28340 20012
rect 23692 19844 23732 19972
rect 25411 19888 25420 19928
rect 25460 19888 25900 19928
rect 25940 19888 25949 19928
rect 28201 19844 28241 19972
rect 29417 19888 29548 19928
rect 29588 19888 29597 19928
rect 29801 19888 29932 19928
rect 29972 19888 29981 19928
rect 19075 19804 19084 19844
rect 19124 19804 20188 19844
rect 20228 19804 20237 19844
rect 21676 19804 22772 19844
rect 22915 19804 22924 19844
rect 22964 19804 23095 19844
rect 23692 19804 25708 19844
rect 25748 19804 26092 19844
rect 26132 19804 26860 19844
rect 26900 19804 26909 19844
rect 27139 19804 27148 19844
rect 27188 19804 28241 19844
rect 22732 19760 22772 19804
rect 18988 19720 21196 19760
rect 21236 19720 21245 19760
rect 22732 19720 25652 19760
rect 15340 19676 15380 19720
rect 6499 19636 6508 19676
rect 6548 19636 8716 19676
rect 8756 19636 8765 19676
rect 10877 19636 10886 19676
rect 11254 19636 11263 19676
rect 13411 19636 13420 19676
rect 13460 19636 15380 19676
rect 15427 19636 15436 19676
rect 15476 19636 17588 19676
rect 18651 19636 18660 19676
rect 19028 19636 19037 19676
rect 23020 19636 24460 19676
rect 24500 19636 24509 19676
rect 17548 19592 17588 19636
rect 23020 19592 23060 19636
rect 7075 19552 7084 19592
rect 7124 19552 8851 19592
rect 8995 19552 9004 19592
rect 9044 19552 15340 19592
rect 15380 19552 15389 19592
rect 16003 19552 16012 19592
rect 16052 19552 17492 19592
rect 17548 19552 23060 19592
rect 23107 19552 23116 19592
rect 23156 19552 25324 19592
rect 25364 19552 25516 19592
rect 25556 19552 25565 19592
rect 8811 19508 8851 19552
rect 17452 19508 17492 19552
rect 25612 19508 25652 19720
rect 26425 19636 26434 19676
rect 26802 19636 26811 19676
rect 25699 19552 25708 19592
rect 25748 19552 28244 19592
rect 6220 19468 6303 19508
rect 7738 19468 7747 19508
rect 7787 19468 7948 19508
rect 7988 19468 8332 19508
rect 8372 19468 8381 19508
rect 8811 19468 9955 19508
rect 9995 19468 10004 19508
rect 10252 19468 10444 19508
rect 10484 19468 10493 19508
rect 11194 19468 11203 19508
rect 11243 19468 11252 19508
rect 6220 19340 6260 19468
rect 4195 19300 4204 19340
rect 4244 19300 4820 19340
rect 4780 19256 4820 19300
rect 5164 19300 5644 19340
rect 5684 19300 5693 19340
rect 5923 19300 5932 19340
rect 5972 19300 5981 19340
rect 6154 19331 6260 19340
rect 5164 19256 5204 19300
rect 6154 19291 6163 19331
rect 6203 19300 6260 19331
rect 6316 19384 6700 19424
rect 6740 19384 7276 19424
rect 7316 19384 7325 19424
rect 7747 19384 7756 19424
rect 7796 19384 7809 19424
rect 8515 19384 8524 19424
rect 8564 19384 8573 19424
rect 6203 19291 6212 19300
rect 6154 19290 6212 19291
rect 547 19216 556 19256
rect 596 19216 887 19256
rect 927 19216 936 19256
rect 1123 19216 1132 19256
rect 1172 19216 1181 19256
rect 1481 19216 1603 19256
rect 1652 19216 1661 19256
rect 2153 19216 2284 19256
rect 2324 19216 2333 19256
rect 2394 19216 2403 19256
rect 2443 19216 2452 19256
rect 2512 19216 2521 19256
rect 2561 19216 2708 19256
rect 2755 19216 2764 19256
rect 2804 19216 2813 19256
rect 2874 19216 2883 19256
rect 2923 19216 2932 19256
rect 2986 19216 2995 19256
rect 3035 19216 3044 19256
rect 3476 19216 3820 19256
rect 3860 19216 3869 19256
rect 4169 19216 4204 19256
rect 4244 19216 4300 19256
rect 4340 19216 4349 19256
rect 4396 19216 4419 19256
rect 4459 19216 4468 19256
rect 4528 19216 4537 19256
rect 4577 19216 4724 19256
rect 4771 19216 4780 19256
rect 4820 19216 4829 19256
rect 4876 19216 4899 19256
rect 4939 19216 4948 19256
rect 5008 19216 5017 19256
rect 5057 19216 5204 19256
rect 5251 19216 5260 19256
rect 5300 19216 5452 19256
rect 5492 19216 5501 19256
rect 5578 19216 5587 19256
rect 5627 19216 5740 19256
rect 5780 19216 5789 19256
rect 5897 19216 6028 19256
rect 6068 19216 6077 19256
rect 1132 18920 1172 19216
rect 2403 19172 2443 19216
rect 2668 19172 2708 19216
rect 2883 19172 2923 19216
rect 3436 19207 3476 19216
rect 3916 19207 3956 19216
rect 4396 19172 4436 19216
rect 4684 19172 4724 19216
rect 1769 19132 1900 19172
rect 1940 19132 1949 19172
rect 2403 19132 2516 19172
rect 2668 19132 2804 19172
rect 2883 19132 3137 19172
rect 3188 19132 3197 19172
rect 3523 19132 3532 19172
rect 3572 19132 3614 19172
rect 3654 19132 3703 19172
rect 4396 19132 4588 19172
rect 4628 19132 4637 19172
rect 4684 19132 4780 19172
rect 4820 19132 4829 19172
rect 2476 18920 2516 19132
rect 2572 19048 2668 19088
rect 2708 19048 2717 19088
rect 1132 18880 2092 18920
rect 2132 18880 2420 18920
rect 2467 18880 2476 18920
rect 2516 18880 2525 18920
rect 2380 18836 2420 18880
rect 2572 18836 2612 19048
rect 2764 19004 2804 19132
rect 4876 19088 4916 19216
rect 6172 19172 6212 19290
rect 6316 19256 6356 19384
rect 6499 19300 6508 19340
rect 6548 19300 6723 19340
rect 6763 19300 6772 19340
rect 6892 19300 7084 19340
rect 7124 19300 7133 19340
rect 6892 19256 6932 19300
rect 7769 19267 7809 19384
rect 8524 19340 8564 19384
rect 8811 19340 8851 19468
rect 9475 19384 9484 19424
rect 9524 19415 9764 19424
rect 9524 19384 9724 19415
rect 9724 19366 9764 19375
rect 6256 19216 6265 19256
rect 6305 19216 6356 19256
rect 6403 19216 6412 19256
rect 6452 19216 6604 19256
rect 6644 19216 6653 19256
rect 6832 19216 6841 19256
rect 6881 19216 6932 19256
rect 6981 19216 6990 19256
rect 7030 19216 7039 19256
rect 7084 19216 7097 19256
rect 7137 19216 7146 19256
rect 7203 19216 7229 19256
rect 7269 19216 7278 19256
rect 7354 19216 7363 19256
rect 7403 19216 7420 19256
rect 7530 19216 7539 19256
rect 7579 19216 7589 19256
rect 7750 19227 7759 19267
rect 7799 19227 7809 19267
rect 7900 19300 8564 19340
rect 8698 19300 8707 19340
rect 8747 19300 8851 19340
rect 8899 19300 8908 19340
rect 8948 19300 9079 19340
rect 9196 19300 9580 19340
rect 9620 19300 9629 19340
rect 7900 19256 7940 19300
rect 9196 19256 9236 19300
rect 10252 19256 10292 19468
rect 7882 19216 7891 19256
rect 7931 19216 7940 19256
rect 7988 19216 7997 19256
rect 8037 19216 8046 19256
rect 8122 19216 8131 19256
rect 8171 19216 8180 19256
rect 8299 19216 8308 19256
rect 8372 19216 8488 19256
rect 8578 19216 8587 19256
rect 8627 19216 8756 19256
rect 8803 19216 8812 19256
rect 8852 19216 9004 19256
rect 9044 19216 9053 19256
rect 9187 19216 9196 19256
rect 9236 19216 9245 19256
rect 9379 19216 9388 19256
rect 9428 19216 9559 19256
rect 9754 19216 9763 19256
rect 9812 19216 9943 19256
rect 10232 19216 10241 19256
rect 10281 19216 10292 19256
rect 10348 19384 10732 19424
rect 10772 19384 10781 19424
rect 6988 19172 7028 19216
rect 5443 19132 5452 19172
rect 5492 19132 5836 19172
rect 5876 19132 5885 19172
rect 6172 19132 6508 19172
rect 6548 19132 6557 19172
rect 6952 19132 6988 19172
rect 7028 19132 7037 19172
rect 7084 19088 7124 19216
rect 7203 19088 7243 19216
rect 7380 19172 7420 19216
rect 7549 19172 7589 19216
rect 7996 19172 8036 19216
rect 7341 19132 7372 19172
rect 7412 19132 7421 19172
rect 7549 19132 7948 19172
rect 7988 19132 8036 19172
rect 8135 19172 8175 19216
rect 8716 19172 8756 19216
rect 10348 19172 10388 19384
rect 11212 19340 11252 19468
rect 10540 19300 11252 19340
rect 11404 19468 11788 19508
rect 11828 19468 11837 19508
rect 12835 19468 12844 19508
rect 12884 19468 13036 19508
rect 13076 19468 13111 19508
rect 14266 19468 14275 19508
rect 14315 19468 15052 19508
rect 15092 19468 15101 19508
rect 15226 19468 15235 19508
rect 15275 19468 15284 19508
rect 16186 19468 16195 19508
rect 16235 19468 16244 19508
rect 16553 19468 16675 19508
rect 16724 19468 16733 19508
rect 16867 19468 16876 19508
rect 16916 19468 17300 19508
rect 17443 19468 17452 19508
rect 17492 19468 17501 19508
rect 20585 19468 20716 19508
rect 20756 19468 20765 19508
rect 22339 19468 22348 19508
rect 22388 19468 22684 19508
rect 22724 19468 22733 19508
rect 25612 19468 28108 19508
rect 28148 19468 28157 19508
rect 10540 19256 10580 19300
rect 11404 19256 11444 19468
rect 10793 19216 10828 19256
rect 10868 19216 10924 19256
rect 10964 19216 10973 19256
rect 11192 19216 11201 19256
rect 11241 19216 11444 19256
rect 11500 19384 11692 19424
rect 11732 19384 11741 19424
rect 12451 19384 12460 19424
rect 12500 19384 12748 19424
rect 12788 19384 12797 19424
rect 11500 19256 11540 19384
rect 13027 19300 13036 19340
rect 13076 19300 14036 19340
rect 13996 19256 14036 19300
rect 14725 19300 14956 19340
rect 14996 19300 15005 19340
rect 14574 19256 14614 19265
rect 14725 19256 14765 19300
rect 15244 19256 15284 19468
rect 16204 19424 16244 19468
rect 17260 19424 17300 19468
rect 16204 19384 17204 19424
rect 17260 19384 18604 19424
rect 18644 19384 18653 19424
rect 20515 19384 20524 19424
rect 20564 19384 22156 19424
rect 22196 19384 22205 19424
rect 22339 19384 22348 19424
rect 22388 19384 22397 19424
rect 23177 19384 23308 19424
rect 23348 19384 23828 19424
rect 24067 19384 24076 19424
rect 24116 19384 26804 19424
rect 26851 19384 26860 19424
rect 26900 19384 28052 19424
rect 15532 19256 15572 19265
rect 16492 19256 16532 19265
rect 16972 19256 17012 19265
rect 17164 19256 17204 19384
rect 22348 19340 22388 19384
rect 23260 19340 23300 19384
rect 23788 19340 23828 19384
rect 17251 19300 17260 19340
rect 17300 19300 17731 19340
rect 17771 19300 17780 19340
rect 17923 19300 17932 19340
rect 17972 19300 18103 19340
rect 19276 19300 22388 19340
rect 22780 19300 22924 19340
rect 22964 19300 22973 19340
rect 23242 19331 23300 19340
rect 17463 19256 17503 19300
rect 19276 19256 19316 19300
rect 22780 19256 22820 19300
rect 23242 19291 23251 19331
rect 23291 19291 23300 19331
rect 23683 19300 23692 19340
rect 23732 19300 23741 19340
rect 23788 19300 24980 19340
rect 25123 19300 25132 19340
rect 25172 19300 26217 19340
rect 26275 19300 26284 19340
rect 26324 19300 26380 19340
rect 26420 19300 26455 19340
rect 23242 19290 23300 19291
rect 23692 19256 23732 19300
rect 10540 19207 10580 19216
rect 11500 19207 11540 19216
rect 11596 19216 11635 19256
rect 11675 19216 11684 19256
rect 11779 19216 11788 19256
rect 11828 19216 11836 19256
rect 11876 19216 11959 19256
rect 12521 19216 12652 19256
rect 12692 19216 12701 19256
rect 13027 19216 13036 19256
rect 13076 19216 13172 19256
rect 13219 19216 13228 19256
rect 13268 19216 13399 19256
rect 13507 19216 13516 19256
rect 13556 19216 13804 19256
rect 13844 19216 13853 19256
rect 13987 19216 13996 19256
rect 14036 19216 14045 19256
rect 14179 19216 14188 19256
rect 14228 19216 14270 19256
rect 14310 19216 14359 19256
rect 14443 19216 14572 19256
rect 14614 19216 14621 19256
rect 14716 19216 14725 19256
rect 14765 19216 14774 19256
rect 14842 19216 14851 19256
rect 14891 19216 14900 19256
rect 14947 19216 14956 19256
rect 14996 19216 15284 19256
rect 15523 19216 15532 19256
rect 15572 19216 15703 19256
rect 16045 19216 16054 19256
rect 16094 19216 16300 19256
rect 16340 19216 16349 19256
rect 16457 19216 16492 19256
rect 16532 19216 16588 19256
rect 16628 19216 16637 19256
rect 16771 19216 16780 19256
rect 16820 19216 16972 19256
rect 17146 19216 17155 19256
rect 17195 19216 17204 19256
rect 17454 19216 17463 19256
rect 17503 19216 17512 19256
rect 17597 19216 17611 19256
rect 17651 19216 17660 19256
rect 17827 19216 17836 19256
rect 17876 19216 18007 19256
rect 18115 19216 18124 19256
rect 18164 19216 18260 19256
rect 18307 19216 18316 19256
rect 18356 19216 18365 19256
rect 18857 19216 18988 19256
rect 19028 19216 19037 19256
rect 19267 19216 19276 19256
rect 19316 19216 19325 19256
rect 20227 19216 20236 19256
rect 20276 19216 20285 19256
rect 20515 19216 20524 19256
rect 20564 19216 20573 19256
rect 20842 19216 20851 19256
rect 20891 19216 20948 19256
rect 20995 19216 21004 19256
rect 21044 19216 21196 19256
rect 21236 19216 21245 19256
rect 21754 19216 21763 19256
rect 21803 19216 21812 19256
rect 21859 19216 21868 19256
rect 21908 19216 21917 19256
rect 22147 19216 22156 19256
rect 22196 19216 22348 19256
rect 22388 19216 22397 19256
rect 22531 19216 22540 19256
rect 22580 19216 22711 19256
rect 22771 19216 22780 19256
rect 22820 19216 22829 19256
rect 22985 19216 23116 19256
rect 23156 19216 23165 19256
rect 23344 19216 23353 19256
rect 23393 19216 23444 19256
rect 23491 19216 23500 19256
rect 23540 19216 23549 19256
rect 23683 19216 23692 19256
rect 23732 19216 23779 19256
rect 23945 19216 24076 19256
rect 24116 19216 24125 19256
rect 24172 19216 24195 19256
rect 24235 19216 24244 19256
rect 24304 19216 24313 19256
rect 24353 19216 24404 19256
rect 24451 19216 24460 19256
rect 24500 19216 24631 19256
rect 11596 19172 11636 19216
rect 11836 19172 11876 19216
rect 13132 19172 13172 19216
rect 13228 19172 13268 19216
rect 14574 19207 14614 19216
rect 14860 19172 14900 19216
rect 15532 19207 15572 19216
rect 16492 19207 16532 19216
rect 16972 19172 17012 19216
rect 17620 19172 17660 19216
rect 18220 19172 18260 19216
rect 8135 19132 8620 19172
rect 8660 19132 8669 19172
rect 8716 19132 9044 19172
rect 9475 19132 9484 19172
rect 9524 19132 9676 19172
rect 9716 19132 9725 19172
rect 10330 19132 10339 19172
rect 10379 19132 10388 19172
rect 11587 19132 11596 19172
rect 11636 19132 11645 19172
rect 11836 19132 13076 19172
rect 13123 19132 13132 19172
rect 13172 19132 13181 19172
rect 13228 19132 13708 19172
rect 13748 19132 13757 19172
rect 14860 19132 14923 19172
rect 15113 19132 15233 19172
rect 15284 19132 15293 19172
rect 15715 19132 15724 19172
rect 15764 19132 16190 19172
rect 16230 19132 16239 19172
rect 16664 19132 16673 19172
rect 16724 19132 16844 19172
rect 16972 19132 17068 19172
rect 17108 19132 17117 19172
rect 17225 19132 17260 19172
rect 17300 19132 17356 19172
rect 17396 19132 17405 19172
rect 17620 19132 17644 19172
rect 17684 19132 17693 19172
rect 18211 19132 18220 19172
rect 18260 19132 18269 19172
rect 8135 19088 8175 19132
rect 3331 19048 3340 19088
rect 3380 19048 3820 19088
rect 3860 19048 3869 19088
rect 4387 19048 4396 19088
rect 4436 19048 4684 19088
rect 4724 19048 4733 19088
rect 4876 19048 6979 19088
rect 7019 19048 7028 19088
rect 7075 19048 7084 19088
rect 7124 19048 7133 19088
rect 7203 19048 7564 19088
rect 7604 19048 7613 19088
rect 7747 19048 7756 19088
rect 7796 19048 8175 19088
rect 2764 18964 4204 19004
rect 4244 18964 4253 19004
rect 4343 18880 4352 18920
rect 4720 18880 4729 18920
rect 991 18796 2324 18836
rect 2380 18796 2612 18836
rect 2851 18796 2860 18836
rect 2900 18796 3284 18836
rect 547 18628 556 18668
rect 596 18628 787 18668
rect 827 18628 836 18668
rect 796 18500 836 18628
rect 991 18584 1031 18796
rect 1324 18712 1804 18752
rect 1844 18712 1940 18752
rect 1324 18668 1364 18712
rect 1108 18628 1364 18668
rect 1411 18628 1420 18668
rect 1460 18628 1612 18668
rect 1652 18628 1661 18668
rect 1108 18584 1148 18628
rect 1900 18584 1940 18712
rect 2284 18668 2324 18796
rect 3244 18752 3284 18796
rect 3226 18712 3235 18752
rect 3275 18712 3284 18752
rect 3331 18712 3340 18752
rect 3380 18712 3511 18752
rect 3715 18712 3724 18752
rect 3764 18712 3895 18752
rect 4649 18712 4780 18752
rect 4820 18712 4829 18752
rect 2249 18628 2380 18668
rect 2420 18628 2923 18668
rect 3003 18628 3052 18668
rect 3092 18628 3134 18668
rect 3174 18628 3183 18668
rect 3820 18628 4204 18668
rect 4244 18628 4253 18668
rect 2284 18584 2324 18628
rect 2883 18584 2923 18628
rect 3820 18584 3860 18628
rect 4876 18584 4916 19048
rect 7084 19004 7124 19048
rect 6499 18964 6508 19004
rect 6548 18964 6658 19004
rect 7084 18964 8332 19004
rect 8372 18964 8524 19004
rect 8564 18964 8573 19004
rect 8631 18964 8908 19004
rect 8948 18964 8957 19004
rect 6403 18880 6412 18920
rect 6452 18880 6559 18920
rect 6519 18794 6559 18880
rect 6490 18754 6499 18794
rect 6539 18754 6559 18794
rect 5033 18712 5059 18752
rect 5099 18712 5164 18752
rect 5204 18712 5213 18752
rect 5443 18712 5452 18752
rect 5492 18712 5882 18752
rect 5356 18628 5548 18668
rect 5588 18628 5740 18668
rect 5780 18628 5789 18668
rect 5356 18584 5396 18628
rect 5842 18584 5882 18712
rect 6028 18712 6316 18752
rect 6356 18712 6365 18752
rect 6618 18740 6658 18964
rect 8631 18920 8671 18964
rect 6787 18880 6796 18920
rect 6836 18880 7660 18920
rect 7700 18880 8671 18920
rect 9004 18920 9044 19132
rect 13036 19088 13076 19132
rect 9763 19048 9772 19088
rect 9812 19048 9955 19088
rect 9995 19048 10004 19088
rect 10051 19048 10060 19088
rect 10100 19048 10444 19088
rect 10484 19048 10493 19088
rect 10601 19048 10723 19088
rect 10772 19048 10781 19088
rect 11011 19048 11020 19088
rect 11060 19048 11069 19088
rect 11273 19048 11404 19088
rect 11444 19048 11453 19088
rect 11683 19048 11692 19088
rect 11732 19048 12739 19088
rect 12779 19048 12788 19088
rect 13036 19048 13411 19088
rect 13451 19048 13516 19088
rect 13556 19048 13620 19088
rect 14467 19048 14476 19088
rect 14516 19048 14764 19088
rect 14804 19048 14813 19088
rect 11020 19004 11060 19048
rect 14883 19004 14923 19132
rect 15034 19048 15043 19088
rect 15092 19048 15223 19088
rect 15331 19048 15340 19088
rect 15380 19048 15436 19088
rect 15476 19048 15511 19088
rect 15785 19048 15859 19088
rect 15899 19048 15916 19088
rect 15956 19048 15965 19088
rect 16156 19004 16196 19132
rect 16387 19048 16396 19088
rect 16436 19048 16876 19088
rect 16916 19048 16925 19088
rect 18211 19048 18220 19088
rect 18260 19048 18269 19088
rect 9091 18964 9100 19004
rect 9140 18964 10828 19004
rect 10868 18964 10877 19004
rect 11020 18964 11308 19004
rect 11348 18964 11357 19004
rect 12931 18964 12940 19004
rect 12980 18964 14804 19004
rect 14883 18964 15532 19004
rect 15572 18964 15581 19004
rect 16156 18964 16684 19004
rect 16724 18964 16733 19004
rect 14764 18920 14804 18964
rect 18220 18920 18260 19048
rect 18316 19004 18356 19216
rect 18988 19172 19028 19207
rect 20236 19172 20276 19216
rect 18691 19132 18700 19172
rect 18740 19132 18892 19172
rect 18932 19132 18941 19172
rect 18988 19132 20428 19172
rect 20468 19132 20477 19172
rect 20524 19088 20564 19216
rect 20908 19172 20948 19216
rect 20899 19132 20908 19172
rect 20948 19132 20957 19172
rect 19555 19048 19564 19088
rect 19604 19048 19613 19088
rect 20428 19048 20564 19088
rect 20606 19048 21100 19088
rect 21140 19048 21149 19088
rect 18316 18964 19468 19004
rect 19508 18964 19517 19004
rect 19564 18920 19604 19048
rect 9004 18880 9292 18920
rect 9332 18880 10540 18920
rect 10580 18880 10589 18920
rect 10636 18880 11404 18920
rect 11444 18880 11453 18920
rect 12117 18880 12126 18920
rect 12494 18880 12503 18920
rect 14764 18880 15436 18920
rect 15476 18880 15485 18920
rect 15964 18880 17300 18920
rect 17539 18880 17548 18920
rect 17588 18880 18260 18920
rect 18316 18880 19604 18920
rect 19891 18880 19900 18920
rect 20268 18880 20277 18920
rect 10636 18836 10676 18880
rect 8035 18796 8044 18836
rect 8084 18796 10676 18836
rect 10819 18796 10828 18836
rect 10868 18796 14956 18836
rect 14996 18796 15284 18836
rect 10732 18752 10772 18761
rect 15244 18752 15284 18796
rect 6028 18584 6068 18712
rect 6616 18710 6658 18740
rect 6844 18712 7180 18752
rect 7220 18712 7948 18752
rect 7988 18712 8948 18752
rect 9667 18712 9676 18752
rect 9716 18712 10444 18752
rect 10484 18712 10493 18752
rect 10772 18712 10924 18752
rect 10964 18712 10973 18752
rect 12547 18712 12556 18752
rect 12596 18712 12691 18752
rect 12731 18712 12740 18752
rect 13507 18712 13516 18752
rect 13556 18712 14598 18752
rect 15235 18712 15244 18752
rect 15284 18712 15293 18752
rect 6607 18670 6616 18710
rect 6656 18670 6665 18710
rect 6211 18628 6220 18668
rect 6260 18628 6269 18668
rect 6220 18584 6260 18628
rect 6844 18626 6884 18712
rect 8908 18668 8948 18712
rect 10732 18703 10772 18712
rect 10924 18668 10964 18712
rect 14558 18668 14598 18712
rect 6826 18586 6835 18626
rect 6875 18586 6884 18626
rect 7084 18628 7276 18668
rect 7316 18628 7325 18668
rect 7397 18628 8203 18668
rect 973 18544 982 18584
rect 1022 18544 1031 18584
rect 1090 18544 1099 18584
rect 1139 18544 1148 18584
rect 1315 18544 1324 18584
rect 1364 18544 1708 18584
rect 1748 18544 1757 18584
rect 1891 18544 1900 18584
rect 1965 18544 2071 18584
rect 2275 18544 2284 18584
rect 2324 18544 2333 18584
rect 2380 18544 2403 18584
rect 2443 18544 2452 18584
rect 2515 18544 2524 18584
rect 2564 18544 2573 18584
rect 2753 18544 2773 18584
rect 2813 18544 2822 18584
rect 2883 18544 2981 18584
rect 3021 18544 3030 18584
rect 3139 18544 3148 18584
rect 3188 18575 3476 18584
rect 3188 18544 3436 18575
rect 1108 18500 1148 18544
rect 2380 18500 2420 18544
rect 2524 18500 2564 18544
rect 2753 18530 2804 18544
rect 796 18460 1148 18500
rect 1210 18460 1219 18500
rect 1259 18460 1268 18500
rect 1411 18460 1420 18500
rect 1460 18460 1516 18500
rect 1556 18460 1591 18500
rect 1696 18460 1804 18500
rect 1867 18460 1876 18500
rect 2083 18460 2092 18500
rect 2132 18460 2188 18500
rect 2228 18460 2263 18500
rect 2356 18460 2380 18500
rect 2420 18460 2429 18500
rect 2476 18460 2564 18500
rect 2621 18460 2668 18500
rect 2708 18460 2717 18500
rect 1228 18416 1268 18460
rect 2476 18416 2516 18460
rect 2668 18416 2708 18460
rect 1219 18376 1228 18416
rect 1268 18376 1315 18416
rect 2467 18376 2476 18416
rect 2516 18376 2525 18416
rect 2659 18376 2668 18416
rect 2708 18376 2717 18416
rect 2764 18332 2804 18530
rect 3523 18544 3532 18584
rect 3572 18544 3628 18584
rect 3668 18544 3703 18584
rect 3802 18544 3811 18584
rect 3851 18544 3860 18584
rect 4003 18544 4012 18584
rect 4052 18544 4108 18584
rect 4148 18544 4183 18584
rect 4282 18544 4291 18584
rect 4331 18544 4340 18584
rect 4876 18544 4972 18584
rect 5012 18544 5021 18584
rect 5347 18544 5356 18584
rect 5396 18544 5405 18584
rect 5513 18544 5644 18584
rect 5684 18544 5693 18584
rect 5842 18544 5861 18584
rect 5901 18544 5910 18584
rect 6019 18544 6028 18584
rect 6068 18544 6077 18584
rect 6173 18544 6219 18584
rect 6259 18544 6268 18584
rect 6473 18544 6543 18584
rect 6583 18544 6604 18584
rect 6644 18544 6653 18584
rect 7084 18575 7124 18628
rect 7397 18584 7437 18628
rect 8163 18584 8203 18628
rect 8908 18628 9964 18668
rect 10004 18628 10013 18668
rect 10060 18628 10348 18668
rect 10388 18628 10397 18668
rect 10924 18628 11828 18668
rect 13603 18628 13612 18668
rect 13652 18628 14036 18668
rect 14549 18628 14558 18668
rect 14598 18628 15807 18668
rect 8908 18584 8948 18628
rect 10060 18584 10100 18628
rect 10924 18584 10964 18628
rect 11788 18584 11828 18628
rect 13996 18584 14036 18628
rect 15148 18584 15188 18628
rect 15767 18584 15807 18628
rect 15964 18584 16004 18880
rect 16195 18796 16204 18836
rect 16244 18796 17108 18836
rect 16090 18712 16099 18752
rect 16139 18712 16972 18752
rect 17012 18712 17021 18752
rect 17068 18668 17108 18796
rect 17260 18752 17300 18880
rect 18316 18752 18356 18880
rect 20428 18836 20468 19048
rect 19555 18796 19564 18836
rect 19604 18796 20468 18836
rect 20606 18752 20646 19048
rect 21772 19004 21812 19216
rect 21868 19172 21908 19216
rect 23404 19172 23444 19216
rect 23500 19172 23540 19216
rect 24172 19172 24212 19216
rect 21868 19132 22348 19172
rect 22388 19132 22397 19172
rect 23395 19132 23404 19172
rect 23444 19132 23453 19172
rect 23500 19132 23692 19172
rect 23732 19132 23741 19172
rect 23884 19132 24212 19172
rect 24364 19172 24404 19216
rect 24940 19172 24980 19300
rect 26177 19256 26217 19300
rect 25193 19216 25324 19256
rect 25364 19216 25373 19256
rect 26168 19216 26177 19256
rect 26217 19216 26226 19256
rect 26371 19229 26380 19256
rect 26284 19216 26380 19229
rect 26420 19216 26429 19256
rect 26537 19216 26668 19256
rect 26708 19216 26717 19256
rect 26284 19189 26420 19216
rect 26284 19172 26324 19189
rect 24364 19132 24844 19172
rect 24884 19132 24893 19172
rect 24940 19132 26324 19172
rect 22025 19048 22156 19088
rect 22196 19048 22205 19088
rect 23011 19048 23020 19088
rect 23060 19048 23191 19088
rect 23369 19048 23500 19088
rect 23540 19048 23549 19088
rect 23884 19004 23924 19132
rect 26764 19088 26804 19384
rect 27427 19300 27436 19340
rect 27476 19300 27676 19340
rect 27716 19300 27725 19340
rect 28012 19261 28052 19384
rect 27139 19216 27148 19256
rect 27188 19216 27475 19256
rect 27515 19216 27524 19256
rect 28001 19221 28010 19261
rect 28050 19221 28059 19261
rect 28204 19256 28244 19552
rect 28649 19384 28684 19424
rect 28724 19384 28780 19424
rect 28820 19384 28829 19424
rect 28195 19216 28204 19256
rect 28244 19216 28253 19256
rect 28387 19216 28396 19256
rect 28436 19216 28445 19256
rect 28579 19216 28588 19256
rect 28628 19216 28637 19256
rect 28396 19172 28436 19216
rect 27331 19132 27340 19172
rect 27380 19132 28436 19172
rect 23971 19048 23980 19088
rect 24020 19048 24940 19088
rect 24980 19048 24989 19088
rect 25987 19048 25996 19088
rect 26036 19048 26708 19088
rect 26764 19048 28396 19088
rect 28436 19048 28445 19088
rect 26668 19004 26708 19048
rect 21772 18964 23788 19004
rect 23828 18964 23837 19004
rect 23884 18964 24556 19004
rect 24596 18964 26228 19004
rect 26668 18964 27532 19004
rect 27572 18964 27581 19004
rect 20707 18880 20716 18920
rect 20756 18880 23060 18920
rect 23020 18836 23060 18880
rect 26188 18836 26228 18964
rect 27665 18880 27674 18920
rect 28042 18880 28051 18920
rect 28588 18836 28628 19216
rect 29033 19048 29164 19088
rect 29204 19048 29213 19088
rect 29417 19048 29548 19088
rect 29588 19048 29597 19088
rect 23020 18796 25996 18836
rect 26036 18796 26045 18836
rect 26188 18796 28628 18836
rect 17242 18712 17251 18752
rect 17291 18712 17300 18752
rect 18298 18712 18307 18752
rect 18347 18712 18356 18752
rect 18595 18712 18604 18752
rect 18644 18712 18932 18752
rect 18979 18712 18988 18752
rect 19028 18712 20646 18752
rect 22409 18712 22540 18752
rect 22580 18712 22589 18752
rect 24451 18712 24460 18752
rect 24500 18712 25132 18752
rect 25172 18712 25181 18752
rect 27427 18712 27436 18752
rect 27476 18712 27916 18752
rect 27956 18712 27965 18752
rect 18892 18668 18932 18712
rect 16553 18628 16588 18668
rect 16628 18628 16640 18668
rect 17068 18628 17131 18668
rect 17251 18628 17260 18668
rect 17300 18628 17684 18668
rect 18010 18628 18019 18668
rect 18059 18628 18499 18668
rect 18539 18628 18548 18668
rect 18604 18628 18796 18668
rect 18836 18628 18845 18668
rect 18892 18628 19180 18668
rect 19220 18628 23252 18668
rect 24931 18628 24940 18668
rect 24980 18628 25315 18668
rect 25355 18628 25364 18668
rect 27148 18628 28684 18668
rect 28724 18628 28733 18668
rect 16600 18584 16640 18628
rect 17091 18584 17131 18628
rect 17644 18584 17684 18628
rect 18604 18584 18644 18628
rect 18892 18584 18932 18628
rect 23212 18584 23252 18628
rect 3436 18526 3476 18535
rect 2874 18460 2883 18500
rect 2923 18460 2932 18500
rect 2755 18292 2764 18332
rect 2804 18292 2813 18332
rect 2883 18080 2923 18460
rect 4108 18416 4148 18544
rect 4300 18500 4340 18544
rect 6971 18533 6980 18573
rect 7020 18533 7029 18573
rect 4300 18460 5164 18500
rect 5204 18460 5213 18500
rect 5417 18460 5548 18500
rect 5588 18460 5597 18500
rect 5770 18491 6068 18500
rect 5770 18451 5779 18491
rect 5819 18460 6068 18491
rect 6665 18460 6700 18500
rect 6740 18460 6796 18500
rect 6836 18460 6845 18500
rect 5819 18451 5828 18460
rect 5770 18450 5828 18451
rect 4108 18376 5452 18416
rect 5492 18376 5501 18416
rect 4972 18292 5212 18332
rect 5252 18292 5261 18332
rect 3103 18124 3112 18164
rect 3480 18124 3489 18164
rect 2371 18040 2380 18080
rect 2420 18040 2429 18080
rect 2883 18040 3380 18080
rect 2380 17996 2420 18040
rect 3340 17996 3380 18040
rect 617 17956 739 17996
rect 788 17956 797 17996
rect 1987 17956 1996 17996
rect 2036 17956 3242 17996
rect 3322 17956 3331 17996
rect 3371 17956 3380 17996
rect 3715 17956 3724 17996
rect 3764 17956 3811 17996
rect 3851 17956 3895 17996
rect 3202 17912 3242 17956
rect 1507 17872 1516 17912
rect 1556 17872 1565 17912
rect 1699 17872 1708 17912
rect 1748 17872 1996 17912
rect 2036 17872 2045 17912
rect 2371 17872 2380 17912
rect 2420 17872 2429 17912
rect 3202 17872 3903 17912
rect 4867 17872 4876 17912
rect 4916 17872 4925 17912
rect 1516 17828 1556 17872
rect 2380 17828 2420 17872
rect 1219 17788 1228 17828
rect 1268 17788 1556 17828
rect 1673 17788 1804 17828
rect 1844 17788 1853 17828
rect 2275 17788 2284 17828
rect 2324 17788 2333 17828
rect 2380 17788 2595 17828
rect 2635 17788 3075 17828
rect 3115 17788 3124 17828
rect 1036 17744 1076 17753
rect 2284 17744 2324 17788
rect 809 17704 940 17744
rect 980 17704 989 17744
rect 1076 17704 1132 17744
rect 1172 17704 1207 17744
rect 1402 17704 1411 17744
rect 1451 17704 1612 17744
rect 1652 17704 1661 17744
rect 1987 17704 1996 17744
rect 2036 17704 2045 17744
rect 2179 17704 2188 17744
rect 2228 17704 2237 17744
rect 2284 17704 2476 17744
rect 2516 17704 2525 17744
rect 2704 17704 2713 17744
rect 2753 17704 2804 17744
rect 2851 17704 2860 17744
rect 2900 17704 2956 17744
rect 2996 17704 3031 17744
rect 3113 17704 3193 17744
rect 3233 17704 3244 17744
rect 3284 17704 3293 17744
rect 1036 17695 1076 17704
rect 728 17620 737 17660
rect 777 17620 884 17660
rect 844 17492 884 17620
rect 809 17452 940 17492
rect 980 17452 1804 17492
rect 1844 17452 1853 17492
rect 1996 17408 2036 17704
rect 2188 17660 2228 17704
rect 2764 17660 2804 17704
rect 3340 17660 3380 17872
rect 3628 17744 3668 17753
rect 3668 17704 3724 17744
rect 3764 17704 3799 17744
rect 3628 17695 3668 17704
rect 3863 17660 3903 17872
rect 4732 17788 4780 17828
rect 4820 17788 4829 17828
rect 2188 17620 2668 17660
rect 2708 17620 2717 17660
rect 2764 17620 2956 17660
rect 2996 17620 3005 17660
rect 3139 17620 3148 17660
rect 3188 17620 3329 17660
rect 3369 17620 3380 17660
rect 3800 17620 3809 17660
rect 3849 17620 3903 17660
rect 4108 17744 4148 17753
rect 4732 17744 4772 17788
rect 4876 17744 4916 17872
rect 4972 17786 5012 18292
rect 6028 18248 6068 18460
rect 6973 18416 7013 18533
rect 7084 18526 7124 18535
rect 7258 18575 7316 18584
rect 7258 18535 7267 18575
rect 7307 18535 7316 18575
rect 7362 18544 7371 18584
rect 7411 18544 7437 18584
rect 7258 18534 7316 18535
rect 6202 18376 6211 18416
rect 6251 18376 7013 18416
rect 6970 18292 6979 18332
rect 7019 18292 7028 18332
rect 6988 18248 7028 18292
rect 6028 18208 6260 18248
rect 6403 18208 6412 18248
rect 6452 18208 7028 18248
rect 7276 18248 7316 18534
rect 7480 18533 7489 18573
rect 7529 18533 7547 18573
rect 7651 18544 7660 18584
rect 7700 18544 7708 18584
rect 7748 18544 7831 18584
rect 7913 18544 8023 18584
rect 8084 18544 8093 18584
rect 8154 18544 8163 18584
rect 8203 18544 8227 18584
rect 8419 18544 8428 18584
rect 8468 18544 8599 18584
rect 8656 18544 8665 18584
rect 8705 18544 8852 18584
rect 8899 18544 8908 18584
rect 8948 18544 8957 18584
rect 9091 18544 9100 18584
rect 9140 18544 9271 18584
rect 9475 18544 9484 18584
rect 9524 18544 9688 18584
rect 9728 18544 9737 18584
rect 9859 18544 9868 18584
rect 9908 18544 9917 18584
rect 10051 18544 10060 18584
rect 10100 18544 10109 18584
rect 10330 18544 10339 18584
rect 10379 18544 10732 18584
rect 10772 18544 10781 18584
rect 10924 18544 11107 18584
rect 11147 18544 11156 18584
rect 11491 18544 11500 18584
rect 11540 18544 11549 18584
rect 11784 18544 11793 18584
rect 11833 18544 11842 18584
rect 12023 18544 12115 18584
rect 12155 18544 12740 18584
rect 13123 18544 13132 18584
rect 13172 18544 13303 18584
rect 13498 18544 13507 18584
rect 13556 18544 13687 18584
rect 13769 18544 13804 18584
rect 13844 18544 13900 18584
rect 13940 18544 13949 18584
rect 13996 18544 14039 18584
rect 14079 18544 14088 18584
rect 14153 18544 14284 18584
rect 14324 18544 14333 18584
rect 14633 18544 14764 18584
rect 14804 18544 14813 18584
rect 14860 18575 14956 18584
rect 7507 18500 7547 18533
rect 8163 18500 8203 18544
rect 8812 18500 8852 18544
rect 9868 18500 9908 18544
rect 11500 18500 11540 18544
rect 12023 18500 12063 18544
rect 7507 18460 7700 18500
rect 7843 18460 7852 18500
rect 7892 18460 7901 18500
rect 8131 18460 8140 18500
rect 8180 18460 8203 18500
rect 8323 18460 8332 18500
rect 8372 18460 8381 18500
rect 8554 18491 8620 18500
rect 7660 18416 7700 18460
rect 7651 18376 7660 18416
rect 7700 18376 7709 18416
rect 7852 18332 7892 18460
rect 7939 18376 7948 18416
rect 7988 18376 8119 18416
rect 7555 18292 7564 18332
rect 7604 18292 7892 18332
rect 8332 18332 8372 18460
rect 8554 18451 8563 18491
rect 8603 18460 8620 18491
rect 8660 18460 8743 18500
rect 8812 18460 9388 18500
rect 9428 18460 9437 18500
rect 9514 18460 9523 18500
rect 9563 18460 9572 18500
rect 9868 18460 10156 18500
rect 10196 18460 11020 18500
rect 11060 18460 11069 18500
rect 11116 18460 12063 18500
rect 8603 18451 8612 18460
rect 8554 18450 8612 18451
rect 9532 18416 9572 18460
rect 11116 18416 11156 18460
rect 12700 18416 12740 18544
rect 12874 18502 12883 18542
rect 12923 18502 12935 18542
rect 14900 18544 14956 18575
rect 14996 18544 15031 18584
rect 15130 18575 15188 18584
rect 14860 18526 14900 18535
rect 15130 18535 15139 18575
rect 15179 18535 15188 18575
rect 15305 18544 15436 18584
rect 15476 18544 15485 18584
rect 15758 18544 15767 18584
rect 15807 18544 15816 18584
rect 15964 18544 16012 18584
rect 16052 18544 16061 18584
rect 16195 18544 16204 18584
rect 16244 18544 16324 18584
rect 16364 18544 16375 18584
rect 16474 18544 16483 18584
rect 16523 18544 16532 18584
rect 16591 18544 16600 18584
rect 16640 18544 16649 18584
rect 16695 18544 16766 18584
rect 16806 18544 16815 18584
rect 16858 18544 16867 18584
rect 16907 18544 16916 18584
rect 17083 18544 17092 18584
rect 17132 18544 17141 18584
rect 17242 18544 17251 18584
rect 17291 18544 17300 18584
rect 17359 18544 17368 18584
rect 17408 18544 17417 18584
rect 15130 18534 15188 18535
rect 12895 18500 12935 18502
rect 12895 18460 13324 18500
rect 13364 18460 13420 18500
rect 13460 18460 13469 18500
rect 14057 18460 14179 18500
rect 14228 18460 14237 18500
rect 14371 18460 14380 18500
rect 14420 18460 14551 18500
rect 15235 18460 15244 18500
rect 15284 18460 15331 18500
rect 15371 18460 15415 18500
rect 15715 18460 15724 18500
rect 15764 18460 15907 18500
rect 15947 18460 15956 18500
rect 16492 18416 16532 18544
rect 16695 18500 16735 18544
rect 16876 18500 16916 18544
rect 16675 18460 16684 18500
rect 16724 18460 16735 18500
rect 16867 18460 16876 18500
rect 16916 18460 16963 18500
rect 17260 18416 17300 18544
rect 9065 18376 9100 18416
rect 9140 18376 9196 18416
rect 9236 18376 9245 18416
rect 9292 18376 9572 18416
rect 10409 18376 10435 18416
rect 10475 18376 10540 18416
rect 10580 18376 10589 18416
rect 10723 18376 10732 18416
rect 10772 18376 11156 18416
rect 11491 18376 11500 18416
rect 11540 18376 12076 18416
rect 12116 18376 12125 18416
rect 12700 18376 17300 18416
rect 9292 18332 9332 18376
rect 17368 18332 17408 18544
rect 17526 18533 17535 18573
rect 17575 18542 17584 18573
rect 17632 18544 17641 18584
rect 17681 18544 17690 18584
rect 18211 18544 18220 18584
rect 18260 18544 18644 18584
rect 18874 18544 18883 18584
rect 18923 18544 18932 18584
rect 18979 18544 18988 18584
rect 19028 18544 20620 18584
rect 20660 18544 20669 18584
rect 20803 18544 20812 18584
rect 20852 18544 21091 18584
rect 21131 18544 21140 18584
rect 22025 18544 22102 18584
rect 22142 18544 22156 18584
rect 22196 18544 22205 18584
rect 17575 18533 17588 18542
rect 22327 18536 22336 18576
rect 22376 18536 22388 18576
rect 22531 18544 22540 18584
rect 22580 18544 22589 18584
rect 22793 18544 22828 18584
rect 22868 18544 22924 18584
rect 22964 18544 22973 18584
rect 23194 18544 23203 18584
rect 23243 18544 23252 18584
rect 25690 18544 25699 18584
rect 25739 18544 26284 18584
rect 26324 18544 26333 18584
rect 17544 18502 17588 18533
rect 17548 18500 17588 18502
rect 22348 18500 22388 18536
rect 17548 18460 17644 18500
rect 17684 18460 17693 18500
rect 20160 18460 20332 18500
rect 20372 18460 20381 18500
rect 20995 18460 21004 18500
rect 21044 18460 21907 18500
rect 21947 18460 21956 18500
rect 22348 18460 22444 18500
rect 22484 18460 22493 18500
rect 20297 18376 20428 18416
rect 20468 18376 20477 18416
rect 20681 18376 20812 18416
rect 20852 18376 20861 18416
rect 22540 18332 22580 18544
rect 27148 18500 27188 18628
rect 27523 18544 27532 18584
rect 27572 18544 27820 18584
rect 27860 18544 27869 18584
rect 27994 18544 28003 18584
rect 28043 18544 28340 18584
rect 28457 18544 28588 18584
rect 28628 18544 28637 18584
rect 28771 18544 28780 18584
rect 28820 18544 28951 18584
rect 29059 18544 29068 18584
rect 29108 18544 29260 18584
rect 29300 18544 29309 18584
rect 28300 18500 28340 18544
rect 24480 18460 24692 18500
rect 24739 18460 24748 18500
rect 24788 18460 25324 18500
rect 25364 18460 25373 18500
rect 26976 18460 27188 18500
rect 27235 18460 27244 18500
rect 27284 18460 28108 18500
rect 28148 18460 28157 18500
rect 28300 18460 28972 18500
rect 29012 18460 29021 18500
rect 8332 18292 8524 18332
rect 8564 18292 8573 18332
rect 8812 18292 9100 18332
rect 9140 18292 9149 18332
rect 9283 18292 9292 18332
rect 9332 18292 9341 18332
rect 9571 18292 9580 18332
rect 9620 18292 9964 18332
rect 10004 18292 10013 18332
rect 10627 18292 10636 18332
rect 10676 18292 11020 18332
rect 11060 18292 11069 18332
rect 11849 18292 11980 18332
rect 12020 18292 12029 18332
rect 12163 18292 12172 18332
rect 12212 18292 12988 18332
rect 13028 18292 13037 18332
rect 14441 18292 14476 18332
rect 14516 18292 14563 18332
rect 14603 18292 14621 18332
rect 16867 18292 16876 18332
rect 16916 18292 17068 18332
rect 17108 18292 17117 18332
rect 17251 18292 17260 18332
rect 17300 18292 17408 18332
rect 18691 18292 18700 18332
rect 18740 18292 20140 18332
rect 20180 18292 20189 18332
rect 20707 18292 20716 18332
rect 20756 18292 21196 18332
rect 21236 18292 21292 18332
rect 21332 18292 21341 18332
rect 22540 18292 23212 18332
rect 23252 18292 23596 18332
rect 23636 18292 23645 18332
rect 8812 18248 8852 18292
rect 24652 18248 24692 18460
rect 27331 18376 27340 18416
rect 27380 18376 28204 18416
rect 28244 18376 28253 18416
rect 28553 18376 28684 18416
rect 28724 18376 28733 18416
rect 24835 18292 24844 18332
rect 24884 18292 27572 18332
rect 27619 18292 27628 18332
rect 27668 18292 27799 18332
rect 28108 18292 28924 18332
rect 28964 18292 28973 18332
rect 27532 18248 27572 18292
rect 28108 18248 28148 18292
rect 7276 18208 8044 18248
rect 8084 18208 8852 18248
rect 8899 18208 8908 18248
rect 8948 18208 11500 18248
rect 11540 18208 11549 18248
rect 16099 18208 16108 18248
rect 16148 18208 20524 18248
rect 20564 18208 20573 18248
rect 24652 18208 26900 18248
rect 27532 18208 28148 18248
rect 5452 18040 6124 18080
rect 6164 18040 6173 18080
rect 5452 17996 5492 18040
rect 5434 17956 5443 17996
rect 5483 17956 5492 17996
rect 6220 17996 6260 18208
rect 8131 18124 8140 18164
rect 8180 18124 9196 18164
rect 9236 18124 9245 18164
rect 9580 18124 10732 18164
rect 10772 18124 10781 18164
rect 10877 18124 10886 18164
rect 11254 18124 11263 18164
rect 18651 18124 18660 18164
rect 19028 18124 19037 18164
rect 26425 18124 26434 18164
rect 26802 18124 26811 18164
rect 9580 17996 9620 18124
rect 6220 17956 6452 17996
rect 6412 17912 6452 17956
rect 7372 17956 9620 17996
rect 9676 18040 11692 18080
rect 11732 18040 11741 18080
rect 15427 18040 15436 18080
rect 15476 18040 16780 18080
rect 16820 18040 16829 18080
rect 17731 18040 17740 18080
rect 17780 18040 21004 18080
rect 21044 18040 21053 18080
rect 7372 17912 7412 17956
rect 9676 17912 9716 18040
rect 10723 17956 10732 17996
rect 10772 17956 11587 17996
rect 11627 17956 11636 17996
rect 12067 17956 12076 17996
rect 12116 17956 13612 17996
rect 13652 17956 13661 17996
rect 15523 17956 15532 17996
rect 15572 17956 15916 17996
rect 15956 17956 15965 17996
rect 17539 17956 17548 17996
rect 17588 17956 23060 17996
rect 23578 17956 23587 17996
rect 23627 17956 26092 17996
rect 26132 17956 26141 17996
rect 23020 17912 23060 17956
rect 26860 17912 26900 18208
rect 5059 17872 5068 17912
rect 5108 17872 5239 17912
rect 6403 17872 6412 17912
rect 6452 17872 6461 17912
rect 6595 17872 6604 17912
rect 6644 17903 7060 17912
rect 6644 17872 7020 17903
rect 7363 17872 7372 17912
rect 7412 17872 7421 17912
rect 7555 17872 7564 17912
rect 7604 17872 7613 17912
rect 8707 17872 8716 17912
rect 8756 17872 9676 17912
rect 9716 17872 9725 17912
rect 11692 17872 12844 17912
rect 12884 17872 12893 17912
rect 13516 17872 14188 17912
rect 14228 17872 14358 17912
rect 14755 17872 14764 17912
rect 14804 17872 14813 17912
rect 17923 17872 17932 17912
rect 17972 17872 17981 17912
rect 18508 17872 20332 17912
rect 20372 17872 20381 17912
rect 21187 17872 21196 17912
rect 21236 17872 21245 17912
rect 23020 17872 24268 17912
rect 24308 17872 24317 17912
rect 25123 17872 25132 17912
rect 25172 17872 26036 17912
rect 26851 17872 26860 17912
rect 26900 17872 26909 17912
rect 27427 17872 27436 17912
rect 27476 17872 27628 17912
rect 27668 17872 27677 17912
rect 27881 17872 28012 17912
rect 28052 17872 28061 17912
rect 7020 17854 7060 17863
rect 7564 17828 7604 17872
rect 11692 17828 11732 17872
rect 13516 17828 13556 17872
rect 5068 17788 5164 17828
rect 5204 17788 5213 17828
rect 5405 17788 5452 17828
rect 5492 17788 5501 17828
rect 5797 17788 5836 17828
rect 5876 17788 5885 17828
rect 6377 17788 6508 17828
rect 6548 17788 6557 17828
rect 6691 17788 6700 17828
rect 6740 17788 6749 17828
rect 7480 17788 7604 17828
rect 7708 17788 7756 17828
rect 7796 17788 10292 17828
rect 4963 17746 4972 17786
rect 5012 17746 5021 17786
rect 4714 17704 4723 17744
rect 4763 17704 4772 17744
rect 4836 17704 4845 17744
rect 4885 17704 4916 17744
rect 2249 17536 2380 17576
rect 2420 17536 2429 17576
rect 2851 17536 2860 17576
rect 2900 17536 3031 17576
rect 3523 17536 3532 17576
rect 3572 17536 3581 17576
rect 4003 17536 4012 17576
rect 4052 17536 4061 17576
rect 3532 17492 3572 17536
rect 2563 17452 2572 17492
rect 2612 17452 3628 17492
rect 3668 17452 3732 17492
rect 4012 17408 4052 17536
rect 4108 17492 4148 17704
rect 5068 17660 5108 17788
rect 5452 17744 5492 17788
rect 5290 17704 5299 17744
rect 5339 17704 5381 17744
rect 5434 17704 5443 17744
rect 5483 17704 5492 17744
rect 5539 17715 5548 17755
rect 5588 17715 5597 17755
rect 5836 17744 5876 17788
rect 6700 17744 6740 17788
rect 7480 17777 7520 17788
rect 7468 17744 7520 17777
rect 7708 17744 7748 17788
rect 9719 17746 9788 17788
rect 10252 17744 10292 17788
rect 10540 17788 11732 17828
rect 12160 17788 12268 17828
rect 12331 17788 12340 17828
rect 12451 17788 12460 17828
rect 12500 17788 12596 17828
rect 12643 17788 12652 17828
rect 12692 17788 13155 17828
rect 13195 17788 13204 17828
rect 13498 17788 13507 17828
rect 13547 17788 13556 17828
rect 14158 17828 14198 17872
rect 14764 17828 14804 17872
rect 17932 17828 17972 17872
rect 14158 17788 14668 17828
rect 14708 17788 14717 17828
rect 14764 17788 15044 17828
rect 10540 17744 10580 17788
rect 11884 17744 11924 17753
rect 12556 17744 12596 17788
rect 5547 17704 5588 17715
rect 5826 17704 5835 17744
rect 5875 17704 5884 17744
rect 5962 17704 5971 17744
rect 6011 17704 6020 17744
rect 6089 17704 6189 17744
rect 6260 17704 6269 17744
rect 6342 17704 6351 17744
rect 6391 17704 6548 17744
rect 6634 17704 6643 17744
rect 6683 17704 6740 17744
rect 6857 17704 6979 17744
rect 7028 17704 7037 17744
rect 7178 17704 7276 17744
rect 7340 17704 7358 17744
rect 7450 17704 7459 17744
rect 7499 17737 7520 17744
rect 7499 17704 7508 17737
rect 7567 17704 7576 17744
rect 7616 17704 7625 17744
rect 7706 17704 7715 17744
rect 7755 17704 7764 17744
rect 7834 17704 7843 17744
rect 7883 17704 7892 17744
rect 8215 17704 8224 17744
rect 8264 17704 8564 17744
rect 8611 17704 8620 17744
rect 8660 17704 9016 17744
rect 9056 17704 9065 17744
rect 9187 17704 9196 17744
rect 9236 17704 9367 17744
rect 9562 17704 9571 17744
rect 9611 17704 9620 17744
rect 5059 17620 5068 17660
rect 5108 17620 5117 17660
rect 4522 17536 4531 17576
rect 4571 17536 4780 17576
rect 4820 17536 4829 17576
rect 5341 17492 5381 17704
rect 5547 17660 5587 17704
rect 5722 17693 5780 17702
rect 5722 17660 5731 17693
rect 5443 17620 5452 17660
rect 5492 17620 5587 17660
rect 5644 17653 5731 17660
rect 5771 17653 5780 17693
rect 5644 17620 5780 17653
rect 5980 17660 6020 17704
rect 6508 17660 6548 17704
rect 7576 17660 7616 17704
rect 5980 17620 6412 17660
rect 6452 17620 6461 17660
rect 6508 17620 6796 17660
rect 6836 17620 6845 17660
rect 7529 17620 7564 17660
rect 7604 17620 7616 17660
rect 7852 17660 7892 17704
rect 8524 17660 8564 17704
rect 9580 17660 9620 17704
rect 9868 17704 9955 17744
rect 9995 17704 10004 17744
rect 10243 17704 10252 17744
rect 10292 17704 10301 17744
rect 10531 17704 10540 17744
rect 10580 17704 10589 17744
rect 10723 17704 10732 17744
rect 10772 17704 10781 17744
rect 11095 17704 11104 17744
rect 11144 17704 11308 17744
rect 11348 17704 11357 17744
rect 11657 17704 11788 17744
rect 11828 17704 11837 17744
rect 12067 17704 12076 17744
rect 12116 17704 12172 17744
rect 12212 17704 12247 17744
rect 12403 17704 12412 17744
rect 12452 17704 12461 17744
rect 12547 17704 12556 17744
rect 12596 17704 12605 17744
rect 12739 17704 12748 17744
rect 12788 17704 12980 17744
rect 13027 17704 13036 17744
rect 13076 17704 13085 17744
rect 13193 17704 13273 17744
rect 13313 17704 13324 17744
rect 13364 17704 13381 17744
rect 13421 17704 13430 17744
rect 13516 17704 13612 17744
rect 13652 17704 13783 17744
rect 13882 17704 13891 17744
rect 13931 17704 13940 17744
rect 7852 17620 8044 17660
rect 8084 17620 8093 17660
rect 8524 17620 8908 17660
rect 8948 17620 8957 17660
rect 9580 17620 9676 17660
rect 9716 17620 9725 17660
rect 5644 17576 5684 17620
rect 9868 17576 9908 17704
rect 10540 17660 10580 17704
rect 10060 17620 10580 17660
rect 10732 17660 10772 17704
rect 11884 17660 11924 17704
rect 12412 17660 12452 17704
rect 12940 17660 12980 17704
rect 13036 17660 13076 17704
rect 13516 17660 13556 17704
rect 13900 17660 13940 17704
rect 10732 17620 11212 17660
rect 11252 17620 11261 17660
rect 11395 17620 11404 17660
rect 11444 17620 11582 17660
rect 11622 17620 11631 17660
rect 11884 17620 12172 17660
rect 12212 17620 12221 17660
rect 12412 17620 12692 17660
rect 12931 17620 12940 17660
rect 12980 17620 12989 17660
rect 13036 17620 13556 17660
rect 13690 17620 13699 17660
rect 13739 17620 13940 17660
rect 13982 17715 13996 17755
rect 14036 17715 14045 17755
rect 14158 17744 14198 17788
rect 15004 17744 15044 17788
rect 15373 17788 15820 17828
rect 15860 17788 15869 17828
rect 16012 17788 17972 17828
rect 18019 17788 18028 17828
rect 18068 17788 18164 17828
rect 15373 17744 15413 17788
rect 16012 17744 16052 17788
rect 18124 17744 18164 17788
rect 18508 17744 18548 17872
rect 18761 17788 18892 17828
rect 18932 17788 18941 17828
rect 19564 17788 20372 17828
rect 20681 17788 20812 17828
rect 20852 17788 20861 17828
rect 19468 17744 19508 17753
rect 5539 17536 5548 17576
rect 5588 17536 5684 17576
rect 5731 17536 5740 17576
rect 5780 17536 7363 17576
rect 7403 17536 7412 17576
rect 8371 17536 8380 17576
rect 8420 17536 8524 17576
rect 8564 17536 8573 17576
rect 8842 17536 8851 17576
rect 8891 17536 8948 17576
rect 9859 17536 9868 17576
rect 9908 17536 9917 17576
rect 8908 17492 8948 17536
rect 10060 17492 10100 17620
rect 10147 17536 10156 17576
rect 10196 17536 10327 17576
rect 10505 17536 10540 17576
rect 10580 17536 10636 17576
rect 10676 17536 10685 17576
rect 11251 17536 11260 17576
rect 11300 17536 11500 17576
rect 11540 17536 11549 17576
rect 11945 17536 11980 17576
rect 12020 17536 12076 17576
rect 12116 17536 12125 17576
rect 12259 17536 12268 17576
rect 12308 17536 12556 17576
rect 12596 17536 12605 17576
rect 4108 17452 5276 17492
rect 5341 17452 5588 17492
rect 8899 17452 8908 17492
rect 8948 17452 8957 17492
rect 9763 17452 9772 17492
rect 9812 17452 10100 17492
rect 12652 17492 12692 17620
rect 13982 17576 14022 17715
rect 14140 17704 14149 17744
rect 14189 17704 14198 17744
rect 14261 17704 14270 17744
rect 14310 17704 14319 17744
rect 14443 17704 14452 17744
rect 14516 17704 14632 17744
rect 14764 17704 14773 17744
rect 14813 17704 14822 17744
rect 14890 17735 14948 17744
rect 14270 17660 14310 17704
rect 14766 17660 14806 17704
rect 14890 17695 14899 17735
rect 14939 17695 14948 17735
rect 14995 17704 15004 17744
rect 15044 17704 15053 17744
rect 15355 17704 15364 17744
rect 15404 17704 15413 17744
rect 15514 17704 15523 17744
rect 15563 17704 15572 17744
rect 14890 17694 14948 17695
rect 14908 17660 14948 17694
rect 15532 17660 15572 17704
rect 14270 17620 14572 17660
rect 14612 17620 14621 17660
rect 14726 17620 14764 17660
rect 14804 17620 14813 17660
rect 14908 17620 15284 17660
rect 15331 17620 15340 17660
rect 15380 17620 15572 17660
rect 15628 17704 15640 17744
rect 15680 17704 15689 17744
rect 15802 17704 15811 17744
rect 15851 17704 15860 17744
rect 15924 17704 15933 17744
rect 15973 17704 16052 17744
rect 16094 17704 16103 17744
rect 16143 17704 16153 17744
rect 16195 17704 16204 17744
rect 16244 17704 16291 17744
rect 16331 17704 16375 17744
rect 16457 17704 16588 17744
rect 16628 17704 16637 17744
rect 16762 17704 16771 17744
rect 16820 17704 16951 17744
rect 17263 17704 17272 17744
rect 17312 17704 17410 17744
rect 17450 17704 17481 17744
rect 17924 17704 17933 17744
rect 17973 17704 18019 17744
rect 18115 17704 18124 17744
rect 18164 17704 18173 17744
rect 18394 17704 18403 17744
rect 18443 17704 18452 17744
rect 18499 17704 18508 17744
rect 18548 17704 18557 17744
rect 18857 17704 18988 17744
rect 19028 17704 19037 17744
rect 19337 17704 19468 17744
rect 19508 17704 19517 17744
rect 15244 17576 15284 17620
rect 12876 17536 12940 17576
rect 12980 17536 13036 17576
rect 13076 17536 13111 17576
rect 13219 17536 13228 17576
rect 13268 17536 14022 17576
rect 14153 17536 14275 17576
rect 14324 17536 14333 17576
rect 15235 17536 15244 17576
rect 15284 17536 15293 17576
rect 12652 17452 13324 17492
rect 13364 17452 13373 17492
rect 1996 17368 3052 17408
rect 3092 17368 3820 17408
rect 3860 17368 4052 17408
rect 4343 17368 4352 17408
rect 4720 17368 4729 17408
rect 4775 17368 5060 17408
rect 1219 17284 1228 17324
rect 1268 17284 2516 17324
rect 2476 17240 2516 17284
rect 4775 17240 4815 17368
rect 4867 17284 4876 17324
rect 4916 17284 4925 17324
rect 4876 17240 4916 17284
rect 5020 17240 5060 17368
rect 5236 17324 5276 17452
rect 5548 17408 5588 17452
rect 5539 17368 5548 17408
rect 5588 17368 5597 17408
rect 8428 17368 10100 17408
rect 8428 17324 8468 17368
rect 5236 17284 8468 17324
rect 8515 17284 8524 17324
rect 8564 17284 9908 17324
rect 835 17200 844 17240
rect 884 17200 1612 17240
rect 1652 17200 1661 17240
rect 1722 17200 2380 17240
rect 2420 17200 2429 17240
rect 2476 17200 3148 17240
rect 3188 17200 3197 17240
rect 3401 17200 3436 17240
rect 3476 17200 3532 17240
rect 3572 17200 3581 17240
rect 4684 17200 4815 17240
rect 4867 17200 4876 17240
rect 4916 17200 4963 17240
rect 5020 17200 5300 17240
rect 5635 17200 5644 17240
rect 5684 17200 6307 17240
rect 6347 17200 6356 17240
rect 6403 17200 6412 17240
rect 6452 17200 9772 17240
rect 9812 17200 9821 17240
rect 1722 17156 1762 17200
rect 809 17116 929 17156
rect 980 17116 989 17156
rect 1228 17116 1420 17156
rect 1460 17116 1469 17156
rect 1562 17116 1612 17156
rect 1652 17116 1722 17156
rect 1762 17116 1771 17156
rect 1891 17116 1900 17156
rect 1940 17116 2071 17156
rect 2356 17116 2476 17156
rect 2516 17116 2525 17156
rect 3052 17116 3148 17156
rect 3188 17116 3197 17156
rect 3244 17116 4204 17156
rect 4244 17116 4253 17156
rect 1123 17032 1132 17072
rect 1172 17032 1181 17072
rect 1228 17063 1268 17116
rect 2092 17072 2155 17077
rect 2356 17072 2396 17116
rect 3052 17072 3092 17116
rect 3244 17072 3284 17116
rect 4684 17072 4724 17200
rect 5260 17198 5300 17200
rect 5260 17158 5368 17198
rect 5408 17158 5417 17198
rect 9868 17156 9908 17284
rect 10060 17240 10100 17368
rect 11308 17368 11884 17408
rect 11924 17368 11933 17408
rect 12117 17368 12126 17408
rect 12494 17368 12503 17408
rect 10060 17200 10924 17240
rect 10964 17200 10973 17240
rect 11308 17156 11348 17368
rect 11692 17284 12556 17324
rect 12596 17284 12605 17324
rect 15139 17284 15148 17324
rect 15188 17284 15476 17324
rect 11692 17240 11732 17284
rect 15436 17240 15476 17284
rect 11674 17200 11683 17240
rect 11723 17200 11732 17240
rect 11779 17200 11788 17240
rect 11828 17200 11971 17240
rect 12011 17200 12020 17240
rect 12076 17200 12835 17240
rect 12875 17200 13228 17240
rect 13268 17200 13277 17240
rect 13961 17200 14083 17240
rect 14132 17200 14804 17240
rect 15418 17200 15427 17240
rect 15467 17200 15476 17240
rect 4771 17116 4780 17156
rect 4820 17116 4862 17156
rect 5059 17116 5068 17156
rect 5108 17116 5117 17156
rect 5827 17116 5836 17156
rect 5876 17116 6220 17156
rect 6260 17116 6347 17156
rect 7324 17116 7372 17156
rect 7412 17116 7421 17156
rect 8035 17116 8044 17156
rect 8084 17116 8332 17156
rect 8372 17116 8381 17156
rect 8716 17116 9292 17156
rect 9332 17116 9341 17156
rect 9868 17116 10732 17156
rect 10772 17116 10781 17156
rect 11266 17116 11348 17156
rect 11395 17116 11404 17156
rect 11444 17116 11467 17156
rect 11933 17116 11980 17156
rect 12020 17116 12029 17156
rect 4780 17072 4820 17116
rect 5068 17072 5108 17116
rect 6147 17072 6187 17116
rect 7324 17072 7364 17116
rect 8716 17072 8756 17116
rect 8860 17072 8903 17073
rect 8980 17072 9020 17116
rect 9868 17072 9908 17116
rect 11266 17072 11306 17116
rect 11404 17072 11444 17116
rect 11980 17072 12020 17116
rect 1132 16904 1172 17032
rect 1373 17032 1411 17072
rect 1451 17032 1460 17072
rect 1507 17032 1516 17072
rect 1556 17032 1687 17072
rect 1987 17048 1996 17072
rect 1228 17014 1268 17023
rect 1420 16988 1460 17032
rect 1411 16948 1420 16988
rect 1460 16948 1469 16988
rect 1516 16904 1556 17032
rect 1889 17008 1996 17048
rect 2036 17008 2045 17072
rect 2092 17063 2180 17072
rect 2092 17023 2131 17063
rect 2171 17023 2180 17063
rect 2227 17032 2236 17072
rect 2276 17032 2285 17072
rect 2338 17032 2347 17072
rect 2387 17032 2396 17072
rect 2563 17032 2572 17072
rect 2612 17032 2743 17072
rect 3043 17032 3052 17072
rect 3092 17032 3101 17072
rect 3226 17032 3235 17072
rect 3275 17032 3284 17072
rect 3427 17032 3436 17072
rect 3476 17032 3485 17072
rect 3532 17032 3628 17072
rect 3668 17032 3677 17072
rect 3907 17032 3916 17072
rect 3956 17032 3965 17072
rect 4012 17032 4103 17072
rect 4143 17032 4152 17072
rect 4282 17032 4291 17072
rect 4331 17032 4724 17072
rect 4766 17032 4775 17072
rect 4815 17032 4824 17072
rect 4954 17032 4963 17072
rect 5003 17032 5012 17072
rect 5068 17032 5116 17072
rect 5156 17032 5165 17072
rect 5415 17032 5452 17072
rect 5492 17032 5501 17072
rect 5698 17032 5707 17072
rect 5780 17032 5887 17072
rect 6138 17032 6147 17072
rect 6187 17032 6196 17072
rect 6307 17032 6316 17072
rect 6356 17032 6460 17072
rect 6500 17032 6509 17072
rect 6569 17032 6604 17072
rect 6644 17032 6700 17072
rect 6740 17032 6749 17072
rect 6796 17032 7180 17072
rect 7220 17032 7229 17072
rect 7306 17063 7364 17072
rect 2092 17022 2180 17023
rect 2092 17007 2155 17022
rect 2115 16946 2155 17007
rect 2236 16988 2276 17032
rect 3436 16988 3476 17032
rect 3532 16988 3572 17032
rect 2236 16948 2324 16988
rect 2083 16906 2092 16946
rect 2132 16906 2155 16946
rect 1132 16864 1708 16904
rect 1748 16864 1757 16904
rect 2284 16820 2324 16948
rect 2435 16948 2453 16988
rect 2493 16948 2502 16988
rect 2659 16948 2668 16988
rect 2708 16948 2839 16988
rect 2956 16948 3476 16988
rect 3523 16948 3532 16988
rect 3572 16948 3581 16988
rect 2435 16904 2475 16948
rect 2956 16904 2996 16948
rect 2435 16864 2476 16904
rect 2516 16864 2525 16904
rect 2947 16864 2956 16904
rect 2996 16864 3005 16904
rect 809 16780 931 16820
rect 980 16780 989 16820
rect 2284 16780 2380 16820
rect 2420 16780 2429 16820
rect 2956 16780 3772 16820
rect 3812 16780 3821 16820
rect 796 16444 1996 16484
rect 2036 16444 2045 16484
rect 2554 16444 2563 16484
rect 2603 16444 2764 16484
rect 2804 16444 2813 16484
rect 796 16274 836 16444
rect 1132 16360 1420 16400
rect 1460 16360 1469 16400
rect 1900 16360 2668 16400
rect 2708 16360 2717 16400
rect 1132 16316 1172 16360
rect 1900 16316 1940 16360
rect 1123 16276 1132 16316
rect 1172 16276 1181 16316
rect 1306 16276 1315 16316
rect 1355 16276 1612 16316
rect 1652 16276 1661 16316
rect 1882 16276 1891 16316
rect 1931 16276 1940 16316
rect 2081 16276 2092 16316
rect 2132 16276 2601 16316
rect 787 16234 796 16274
rect 836 16234 845 16274
rect 2081 16232 2121 16276
rect 922 16192 931 16232
rect 971 16192 980 16232
rect 1027 16192 1036 16232
rect 1076 16192 1228 16232
rect 1268 16192 1277 16232
rect 1577 16192 1699 16232
rect 1748 16192 1757 16232
rect 2072 16192 2081 16232
rect 2121 16192 2130 16232
rect 2256 16192 2378 16232
rect 2420 16192 2436 16232
rect 940 16148 980 16192
rect 2561 16148 2601 16276
rect 2860 16232 2900 16241
rect 2956 16232 2996 16780
rect 3103 16612 3112 16652
rect 3480 16612 3489 16652
rect 3628 16360 3820 16400
rect 3860 16360 3869 16400
rect 3628 16316 3668 16360
rect 3916 16316 3956 17032
rect 4012 16988 4052 17032
rect 4972 16988 5012 17032
rect 5279 16990 5288 17030
rect 5328 16990 5348 17030
rect 5308 16988 5348 16990
rect 5452 16988 5492 17032
rect 5578 16990 5587 17030
rect 5627 16990 5636 17030
rect 6010 16990 6019 17030
rect 6059 16990 6068 17030
rect 4003 16948 4012 16988
rect 4052 16948 4061 16988
rect 4972 16948 5068 16988
rect 5108 16948 5117 16988
rect 5308 16948 5396 16988
rect 5452 16948 5462 16988
rect 5502 16948 5511 16988
rect 5356 16946 5396 16948
rect 5356 16906 5408 16946
rect 5368 16736 5408 16906
rect 5583 16904 5623 16990
rect 6028 16988 6068 16990
rect 5705 16948 5836 16988
rect 5876 16948 5885 16988
rect 6028 16948 6124 16988
rect 6164 16948 6173 16988
rect 5583 16864 5873 16904
rect 5368 16696 5740 16736
rect 5780 16696 5789 16736
rect 5833 16652 5873 16864
rect 5923 16822 5932 16862
rect 5972 16822 5981 16862
rect 5932 16736 5972 16822
rect 5923 16696 5932 16736
rect 5972 16696 5981 16736
rect 5833 16612 5972 16652
rect 5932 16568 5972 16612
rect 5923 16528 5932 16568
rect 5972 16528 5981 16568
rect 4867 16444 4876 16484
rect 4916 16444 5012 16484
rect 4387 16360 4396 16400
rect 4436 16360 4874 16400
rect 3427 16276 3436 16316
rect 3476 16276 3524 16316
rect 3610 16276 3619 16316
rect 3659 16276 3668 16316
rect 3811 16276 3820 16316
rect 3860 16276 3956 16316
rect 4099 16276 4108 16316
rect 4148 16276 4244 16316
rect 4576 16276 4684 16316
rect 4747 16276 4756 16316
rect 3484 16232 3524 16276
rect 4204 16232 4244 16276
rect 4834 16232 4874 16360
rect 4972 16316 5012 16444
rect 6796 16400 6836 17032
rect 7306 17023 7315 17063
rect 7355 17023 7364 17063
rect 7721 17032 7852 17072
rect 7892 17032 7901 17072
rect 8105 17032 8179 17072
rect 8219 17032 8236 17072
rect 8276 17032 8285 17072
rect 8332 17032 8380 17072
rect 8420 17032 8429 17072
rect 8686 17032 8695 17072
rect 8735 17032 8756 17072
rect 8836 17032 8845 17072
rect 8885 17032 8903 17072
rect 8962 17032 8971 17072
rect 9011 17032 9020 17072
rect 9091 17032 9100 17072
rect 9140 17032 9257 17072
rect 9297 17032 9306 17072
rect 9418 17032 9427 17072
rect 9467 17032 9484 17072
rect 9524 17032 9607 17072
rect 9663 17032 9672 17072
rect 9712 17032 9721 17072
rect 9859 17032 9868 17072
rect 9908 17032 9917 17072
rect 10147 17032 10156 17072
rect 10196 17032 10648 17072
rect 10688 17032 10828 17072
rect 10868 17032 10877 17072
rect 11011 17032 11020 17072
rect 11060 17032 11069 17072
rect 11248 17032 11257 17072
rect 11297 17032 11306 17072
rect 11362 17032 11371 17072
rect 11411 17032 11444 17072
rect 11587 17032 11596 17072
rect 11636 17032 11767 17072
rect 11962 17032 11971 17072
rect 12011 17032 12020 17072
rect 12076 17063 12116 17200
rect 12250 17147 12460 17156
rect 12250 17107 12259 17147
rect 12299 17116 12460 17147
rect 12500 17116 12509 17156
rect 12643 17116 12652 17156
rect 12692 17116 12788 17156
rect 13027 17116 13036 17156
rect 13087 17116 13207 17156
rect 13694 17116 13996 17156
rect 14036 17116 14045 17156
rect 14371 17116 14380 17156
rect 14420 17116 14516 17156
rect 12299 17107 12308 17116
rect 12250 17106 12308 17107
rect 12748 17072 12788 17116
rect 13694 17114 13734 17116
rect 13650 17105 13734 17114
rect 7306 17022 7364 17023
rect 7411 16990 7420 17030
rect 7460 16990 7484 17030
rect 7444 16988 7484 16990
rect 6953 16948 7084 16988
rect 7124 16948 7133 16988
rect 7444 16948 7948 16988
rect 7988 16948 7997 16988
rect 8332 16904 8372 17032
rect 8863 16988 8903 17032
rect 9672 16988 9712 17032
rect 8515 16948 8524 16988
rect 8564 16948 8695 16988
rect 8803 16948 8812 16988
rect 8852 16948 9100 16988
rect 9140 16948 9149 16988
rect 9667 16948 9676 16988
rect 9716 16948 9759 16988
rect 9955 16948 9964 16988
rect 10004 16948 10348 16988
rect 10388 16948 10483 16988
rect 10523 16948 10548 16988
rect 7267 16864 7276 16904
rect 7316 16864 8372 16904
rect 8419 16864 8428 16904
rect 8468 16864 8620 16904
rect 8660 16864 8669 16904
rect 8995 16864 9004 16904
rect 9044 16864 9196 16904
rect 9236 16864 9245 16904
rect 9859 16864 9868 16904
rect 9908 16864 9917 16904
rect 8332 16820 8372 16864
rect 9868 16820 9908 16864
rect 8332 16780 9868 16820
rect 9908 16780 9917 16820
rect 11020 16736 11060 17032
rect 12346 17032 12355 17072
rect 12395 17032 12404 17072
rect 12076 17014 12116 17023
rect 12364 16988 12404 17032
rect 12523 17021 12532 17061
rect 12572 17021 12581 17061
rect 12730 17032 12739 17072
rect 12779 17032 12980 17072
rect 13193 17032 13324 17072
rect 13364 17032 13373 17072
rect 13650 17065 13651 17105
rect 13691 17074 13734 17105
rect 13691 17065 13700 17074
rect 14476 17072 14516 17116
rect 14764 17114 14804 17200
rect 15628 17156 15668 17704
rect 15820 17660 15860 17704
rect 15820 17620 16012 17660
rect 16052 17620 16061 17660
rect 16113 17492 16153 17704
rect 17281 17660 17321 17704
rect 17933 17660 17973 17704
rect 16675 17620 16684 17660
rect 16724 17620 17321 17660
rect 17513 17620 17596 17660
rect 17636 17620 17644 17660
rect 17684 17620 17693 17660
rect 17923 17620 17932 17660
rect 17972 17620 17981 17660
rect 16195 17536 16204 17576
rect 16244 17536 16396 17576
rect 16436 17536 16445 17576
rect 16675 17536 16684 17576
rect 16724 17536 17107 17576
rect 17147 17536 17156 17576
rect 16113 17452 16204 17492
rect 16244 17452 16253 17492
rect 18412 17324 18452 17704
rect 19468 17695 19508 17704
rect 19564 17576 19604 17788
rect 20332 17744 20372 17788
rect 21196 17744 21236 17872
rect 25996 17828 26036 17872
rect 19978 17704 19987 17744
rect 20027 17704 20084 17744
rect 20201 17704 20332 17744
rect 20372 17704 20381 17744
rect 20515 17704 20524 17744
rect 20564 17704 21236 17744
rect 21340 17788 22243 17828
rect 22283 17788 22292 17828
rect 22348 17788 23500 17828
rect 23540 17788 23549 17828
rect 23779 17788 23788 17828
rect 23828 17788 24172 17828
rect 24212 17788 24221 17828
rect 24355 17788 24364 17828
rect 24404 17788 25900 17828
rect 25940 17788 25949 17828
rect 25996 17788 27532 17828
rect 27572 17788 27581 17828
rect 19171 17536 19180 17576
rect 19220 17536 19604 17576
rect 20044 17492 20084 17704
rect 21340 17660 21380 17788
rect 21449 17704 21580 17744
rect 21620 17704 21629 17744
rect 21737 17704 21868 17744
rect 21908 17704 21917 17744
rect 21580 17686 21620 17695
rect 21964 17660 22004 17788
rect 22348 17744 22388 17788
rect 22051 17704 22060 17744
rect 22100 17704 22103 17744
rect 22143 17704 22231 17744
rect 22339 17704 22348 17744
rect 22388 17704 22397 17744
rect 23107 17704 23116 17744
rect 23156 17704 23224 17744
rect 23264 17704 23287 17744
rect 23390 17704 23399 17744
rect 23439 17704 23448 17744
rect 23578 17704 23587 17744
rect 23627 17704 23788 17744
rect 23828 17704 23837 17744
rect 23962 17704 23971 17744
rect 24011 17704 24020 17744
rect 24451 17704 24460 17744
rect 24500 17704 24739 17744
rect 24779 17704 24788 17744
rect 25699 17704 25708 17744
rect 25760 17704 25879 17744
rect 25987 17704 25996 17744
rect 26036 17704 26045 17744
rect 26659 17704 26668 17744
rect 26708 17704 27244 17744
rect 27284 17704 27293 17744
rect 27427 17704 27436 17744
rect 27476 17704 27485 17744
rect 23399 17660 23439 17704
rect 20467 17620 20476 17660
rect 20516 17620 21380 17660
rect 21475 17620 21484 17660
rect 21524 17620 21533 17660
rect 21964 17620 22636 17660
rect 22676 17620 22685 17660
rect 23299 17620 23308 17660
rect 23348 17620 23439 17660
rect 21484 17576 21524 17620
rect 23980 17576 24020 17704
rect 25996 17660 26036 17704
rect 27436 17660 27476 17704
rect 24931 17620 24940 17660
rect 24980 17620 26036 17660
rect 27043 17620 27052 17660
rect 27092 17620 27476 17660
rect 20131 17536 20140 17576
rect 20180 17536 20311 17576
rect 20441 17536 20524 17576
rect 20564 17536 20572 17576
rect 20612 17536 20621 17576
rect 21484 17536 22156 17576
rect 22196 17536 22205 17576
rect 22313 17536 22435 17576
rect 22484 17536 22493 17576
rect 23050 17536 23059 17576
rect 23099 17536 23212 17576
rect 23252 17536 23261 17576
rect 23491 17536 23500 17576
rect 23540 17536 24940 17576
rect 24980 17536 24989 17576
rect 25546 17536 25555 17576
rect 25595 17536 25604 17576
rect 27209 17536 27340 17576
rect 27380 17536 27389 17576
rect 25564 17492 25604 17536
rect 18691 17452 18700 17492
rect 18740 17452 20620 17492
rect 20660 17452 20669 17492
rect 23587 17452 23596 17492
rect 23636 17452 25604 17492
rect 19891 17368 19900 17408
rect 20268 17368 20277 17408
rect 27665 17368 27674 17408
rect 28042 17368 28051 17408
rect 18412 17284 21868 17324
rect 21908 17284 21917 17324
rect 16867 17200 16876 17240
rect 16916 17200 17068 17240
rect 17108 17200 17117 17240
rect 17162 17200 18316 17240
rect 18356 17200 18365 17240
rect 19555 17200 19564 17240
rect 19604 17200 19852 17240
rect 19892 17200 19901 17240
rect 17162 17156 17202 17200
rect 14746 17074 14755 17114
rect 14795 17074 14804 17114
rect 15052 17116 15148 17156
rect 15188 17116 15197 17156
rect 15256 17116 15668 17156
rect 13650 17056 13700 17065
rect 13987 17032 13996 17072
rect 14036 17032 14045 17072
rect 14153 17032 14284 17072
rect 14324 17032 14333 17072
rect 14458 17032 14467 17072
rect 14507 17032 14516 17072
rect 14860 17032 14881 17072
rect 14921 17032 14930 17072
rect 11146 16979 11348 16988
rect 11146 16939 11155 16979
rect 11195 16948 11348 16979
rect 11482 16948 11491 16988
rect 11531 16948 11692 16988
rect 11732 16948 11741 16988
rect 12355 16948 12364 16988
rect 12404 16948 12451 16988
rect 11195 16939 11204 16948
rect 11146 16938 11204 16939
rect 11308 16904 11348 16948
rect 12541 16904 12581 17021
rect 12940 16988 12980 17032
rect 12940 16948 13420 16988
rect 13460 16948 13469 16988
rect 11308 16864 11500 16904
rect 11540 16864 11549 16904
rect 12541 16864 12556 16904
rect 12596 16864 12605 16904
rect 13027 16780 13036 16820
rect 13076 16780 13085 16820
rect 13673 16780 13804 16820
rect 13844 16780 13853 16820
rect 13036 16736 13076 16780
rect 13996 16736 14036 17032
rect 14860 16988 14900 17032
rect 15052 16988 15092 17116
rect 15256 17072 15296 17116
rect 15628 17072 15668 17116
rect 15820 17116 16012 17156
rect 16052 17116 16061 17156
rect 16483 17116 16492 17156
rect 16532 17116 16541 17156
rect 16771 17116 16780 17156
rect 16820 17116 17202 17156
rect 17482 17116 17491 17156
rect 17531 17116 17836 17156
rect 17876 17116 17885 17156
rect 17932 17116 18220 17156
rect 18260 17116 18269 17156
rect 15820 17072 15860 17116
rect 16492 17072 16532 17116
rect 17932 17072 17972 17116
rect 20236 17072 20276 17284
rect 20323 17200 20332 17240
rect 20372 17200 23871 17240
rect 20419 17116 20428 17156
rect 20468 17116 21004 17156
rect 21044 17116 21053 17156
rect 21955 17116 21964 17156
rect 22004 17116 22444 17156
rect 22484 17116 23156 17156
rect 23116 17114 23156 17116
rect 23116 17105 23179 17114
rect 23116 17074 23130 17105
rect 15178 17032 15187 17072
rect 15227 17032 15296 17072
rect 15341 17021 15356 17061
rect 15396 17021 15405 17061
rect 15528 17032 15537 17072
rect 15577 17032 15586 17072
rect 15628 17032 15667 17072
rect 15707 17032 15752 17072
rect 15802 17032 15811 17072
rect 15851 17032 15860 17072
rect 15341 16988 15381 17021
rect 15534 16988 15574 17032
rect 15712 16988 15752 17032
rect 15907 17021 15916 17061
rect 15956 17021 15965 17061
rect 16429 17032 16438 17072
rect 16478 17032 16532 17072
rect 16579 17032 16588 17072
rect 16628 17032 16637 17072
rect 16771 17032 16780 17072
rect 16820 17032 16829 17072
rect 16964 17032 16973 17072
rect 17013 17032 17059 17072
rect 17148 17032 17157 17072
rect 17197 17032 17206 17072
rect 17609 17032 17686 17072
rect 17726 17032 17740 17072
rect 17780 17032 17789 17072
rect 17923 17032 17932 17072
rect 17972 17032 17981 17072
rect 18115 17032 18124 17072
rect 18164 17032 18173 17072
rect 18490 17032 18499 17072
rect 18539 17032 18700 17072
rect 18740 17032 18749 17072
rect 18988 17063 19180 17072
rect 14371 16948 14380 16988
rect 14420 16948 14900 16988
rect 15043 16948 15052 16988
rect 15092 16948 15101 16988
rect 15235 16948 15244 16988
rect 15284 16948 15381 16988
rect 15490 16948 15532 16988
rect 15572 16948 15581 16988
rect 15712 16948 15764 16988
rect 14755 16864 14764 16904
rect 14804 16864 14956 16904
rect 14996 16864 15005 16904
rect 15724 16820 15764 16948
rect 15916 16904 15956 17021
rect 16588 16988 16628 17032
rect 16169 16948 16243 16988
rect 16283 16948 16300 16988
rect 16340 16948 16349 16988
rect 16483 16948 16492 16988
rect 16532 16948 16628 16988
rect 16780 16904 16820 17032
rect 16972 16988 17012 17032
rect 17164 16988 17204 17032
rect 16963 16948 16972 16988
rect 17012 16948 17021 16988
rect 17155 16948 17164 16988
rect 17204 16948 17244 16988
rect 18124 16904 18164 17032
rect 19028 17032 19180 17063
rect 19220 17032 19229 17072
rect 19337 17032 19468 17072
rect 19508 17032 19517 17072
rect 19817 17032 19948 17072
rect 19988 17032 19997 17072
rect 20057 17032 20066 17072
rect 20106 17032 20276 17072
rect 20489 17032 20620 17072
rect 20660 17032 20669 17072
rect 20777 17032 20899 17072
rect 20948 17032 20957 17072
rect 22084 17032 22093 17072
rect 22133 17032 22156 17072
rect 22196 17032 22273 17072
rect 22339 17032 22348 17072
rect 22388 17032 22397 17072
rect 22889 17032 23020 17072
rect 23060 17032 23069 17072
rect 23129 17065 23130 17074
rect 23170 17065 23179 17105
rect 23129 17056 23179 17065
rect 23369 17032 23404 17072
rect 23444 17032 23500 17072
rect 23540 17032 23549 17072
rect 18988 17014 19028 17023
rect 22348 16988 22388 17032
rect 23404 16988 23444 17032
rect 19433 16948 19564 16988
rect 19604 16948 19613 16988
rect 21100 16948 21716 16988
rect 21859 16948 21868 16988
rect 21908 16948 23444 16988
rect 23831 16988 23871 17200
rect 23980 17200 25708 17240
rect 25748 17200 25757 17240
rect 25891 17200 25900 17240
rect 25940 17200 28492 17240
rect 28532 17200 28541 17240
rect 23980 17072 24020 17200
rect 24451 17116 24460 17156
rect 24500 17116 25556 17156
rect 27331 17116 27340 17156
rect 27380 17116 28099 17156
rect 28139 17116 28148 17156
rect 25516 17072 25556 17116
rect 23962 17032 23971 17072
rect 24011 17032 24020 17072
rect 24460 17063 24500 17072
rect 24547 17032 24556 17072
rect 24596 17032 24940 17072
rect 24980 17032 25132 17072
rect 25172 17032 25181 17072
rect 25289 17032 25324 17072
rect 25364 17032 25420 17072
rect 25460 17032 25469 17072
rect 25512 17032 25521 17072
rect 25561 17032 25570 17072
rect 27523 17032 27532 17072
rect 27572 17032 27715 17072
rect 27755 17032 27764 17072
rect 24460 16988 24500 17023
rect 23831 16948 24364 16988
rect 24404 16948 24413 16988
rect 24460 16948 24844 16988
rect 24884 16948 24893 16988
rect 25027 16948 25036 16988
rect 25076 16948 26284 16988
rect 26324 16948 26333 16988
rect 27427 16948 27436 16988
rect 27476 16948 27485 16988
rect 21100 16904 21140 16948
rect 21676 16904 21716 16948
rect 15916 16864 16588 16904
rect 16628 16864 16637 16904
rect 16780 16864 17740 16904
rect 17780 16864 17789 16904
rect 18124 16864 19756 16904
rect 19796 16864 19805 16904
rect 19852 16864 21140 16904
rect 21283 16864 21292 16904
rect 21332 16864 21580 16904
rect 21620 16864 21629 16904
rect 21676 16864 22732 16904
rect 22772 16864 22781 16904
rect 22828 16864 26324 16904
rect 14458 16780 14467 16820
rect 14507 16780 15628 16820
rect 15668 16780 15677 16820
rect 15724 16780 16012 16820
rect 16052 16780 16061 16820
rect 17801 16780 17932 16820
rect 17972 16780 17981 16820
rect 19852 16736 19892 16864
rect 22828 16820 22868 16864
rect 26284 16820 26324 16864
rect 20131 16780 20140 16820
rect 20180 16780 21676 16820
rect 21716 16780 21725 16820
rect 21859 16780 21868 16820
rect 21908 16780 22868 16820
rect 23020 16780 23740 16820
rect 23780 16780 23789 16820
rect 24739 16780 24748 16820
rect 24788 16780 25804 16820
rect 25844 16780 25853 16820
rect 26057 16780 26188 16820
rect 26228 16780 26237 16820
rect 26284 16780 28108 16820
rect 28148 16780 28157 16820
rect 23020 16736 23060 16780
rect 10787 16696 11060 16736
rect 13027 16696 13036 16736
rect 13076 16696 13123 16736
rect 13411 16696 13420 16736
rect 13460 16696 19892 16736
rect 19939 16696 19948 16736
rect 19988 16696 23060 16736
rect 8323 16612 8332 16652
rect 8372 16612 10444 16652
rect 10484 16612 10493 16652
rect 6892 16528 7589 16568
rect 8515 16528 8524 16568
rect 8564 16528 10156 16568
rect 10196 16528 10205 16568
rect 5155 16360 5164 16400
rect 5204 16360 5644 16400
rect 5684 16360 5693 16400
rect 6787 16360 6796 16400
rect 6836 16360 6845 16400
rect 6892 16316 6932 16528
rect 7363 16444 7372 16484
rect 7412 16444 7421 16484
rect 7023 16360 7276 16400
rect 7316 16360 7325 16400
rect 4963 16276 4972 16316
rect 5012 16276 5021 16316
rect 5178 16276 5187 16316
rect 5227 16276 5548 16316
rect 5588 16276 5597 16316
rect 5705 16276 5740 16316
rect 5780 16276 5836 16316
rect 5876 16276 5885 16316
rect 6124 16276 6316 16316
rect 6379 16276 6487 16316
rect 6691 16276 6700 16316
rect 6740 16276 6892 16316
rect 6932 16276 6941 16316
rect 6124 16232 6164 16276
rect 7023 16274 7063 16360
rect 7372 16316 7412 16444
rect 7549 16400 7589 16528
rect 10787 16484 10827 16696
rect 10877 16612 10886 16652
rect 11254 16612 11263 16652
rect 12940 16612 16108 16652
rect 16148 16612 16157 16652
rect 18651 16612 18660 16652
rect 19028 16612 19037 16652
rect 21283 16612 21292 16652
rect 21332 16612 25324 16652
rect 25364 16612 25373 16652
rect 26425 16612 26434 16652
rect 26802 16612 26811 16652
rect 11212 16528 11596 16568
rect 11636 16528 11645 16568
rect 10787 16444 10819 16484
rect 10859 16444 10868 16484
rect 11212 16400 11252 16528
rect 12940 16484 12980 16612
rect 11308 16444 12980 16484
rect 7549 16360 7604 16400
rect 7651 16360 7660 16400
rect 7700 16360 8135 16400
rect 8175 16360 8184 16400
rect 8227 16360 8236 16400
rect 8276 16360 8660 16400
rect 8794 16360 8803 16400
rect 8843 16360 9044 16400
rect 10435 16360 10444 16400
rect 10484 16360 10493 16400
rect 10604 16391 10636 16400
rect 10676 16360 10775 16400
rect 11203 16360 11212 16400
rect 11252 16360 11261 16400
rect 7564 16316 7604 16360
rect 7171 16276 7180 16316
rect 7220 16276 7229 16316
rect 7372 16276 7520 16316
rect 7564 16276 7616 16316
rect 8227 16276 8236 16316
rect 8276 16276 8524 16316
rect 8564 16276 8573 16316
rect 7018 16234 7027 16274
rect 7067 16234 7076 16274
rect 7180 16232 7220 16276
rect 7480 16232 7520 16276
rect 7576 16241 7616 16276
rect 7576 16232 7652 16241
rect 8620 16232 8660 16360
rect 9004 16316 9044 16360
rect 10444 16316 10484 16360
rect 10604 16342 10644 16351
rect 11308 16316 11348 16444
rect 11452 16360 11692 16400
rect 11732 16360 11741 16400
rect 8995 16276 9004 16316
rect 9044 16276 9140 16316
rect 9100 16232 9140 16276
rect 10282 16307 10484 16316
rect 10282 16267 10291 16307
rect 10331 16276 10484 16307
rect 11011 16276 11020 16316
rect 11060 16276 11308 16316
rect 11348 16276 11357 16316
rect 10331 16267 10340 16276
rect 11452 16274 11492 16360
rect 12940 16316 12980 16444
rect 13036 16528 13324 16568
rect 13364 16528 13373 16568
rect 15436 16528 16012 16568
rect 16052 16528 16061 16568
rect 19747 16528 19756 16568
rect 19796 16528 22628 16568
rect 23011 16528 23020 16568
rect 23060 16528 23924 16568
rect 25411 16528 25420 16568
rect 25460 16528 28724 16568
rect 13036 16400 13076 16528
rect 15436 16484 15476 16528
rect 22588 16484 22628 16528
rect 23884 16484 23924 16528
rect 15427 16444 15436 16484
rect 15476 16444 15485 16484
rect 15610 16444 15619 16484
rect 15668 16444 15799 16484
rect 17443 16444 17452 16484
rect 17492 16444 17972 16484
rect 19363 16444 19372 16484
rect 19412 16444 19421 16484
rect 21571 16444 21580 16484
rect 21620 16444 22156 16484
rect 22196 16444 22205 16484
rect 22339 16444 22348 16484
rect 22388 16444 22444 16484
rect 22484 16444 22519 16484
rect 22588 16444 23500 16484
rect 23540 16444 23549 16484
rect 23875 16444 23884 16484
rect 23924 16444 28300 16484
rect 28340 16444 28349 16484
rect 13027 16360 13036 16400
rect 13076 16360 13085 16400
rect 13155 16360 13420 16400
rect 13460 16360 13469 16400
rect 13795 16360 13804 16400
rect 13844 16360 13853 16400
rect 14179 16360 14188 16400
rect 14228 16360 15092 16400
rect 13155 16316 13195 16360
rect 11753 16276 11884 16316
rect 11924 16276 12263 16316
rect 10282 16266 10340 16267
rect 11434 16234 11443 16274
rect 11483 16234 11492 16274
rect 2900 16192 2996 16232
rect 3343 16192 3352 16232
rect 3392 16192 3401 16232
rect 3475 16192 3484 16232
rect 3524 16192 3533 16232
rect 3715 16192 3724 16232
rect 3764 16192 3840 16232
rect 4099 16192 4108 16232
rect 4148 16192 4157 16232
rect 4204 16192 4227 16232
rect 4267 16192 4276 16232
rect 4336 16192 4345 16232
rect 4385 16192 4396 16232
rect 4436 16192 4525 16232
rect 4579 16192 4588 16232
rect 4628 16192 4637 16232
rect 4816 16192 4825 16232
rect 4865 16192 4894 16232
rect 5068 16192 5077 16232
rect 5117 16192 5126 16232
rect 5290 16192 5299 16232
rect 5339 16192 5348 16232
rect 5574 16192 5583 16232
rect 5623 16192 5782 16232
rect 5866 16192 5875 16232
rect 5915 16192 6164 16232
rect 6211 16192 6220 16232
rect 6260 16192 6269 16232
rect 6448 16192 6457 16232
rect 6497 16192 6604 16232
rect 6644 16192 6653 16232
rect 6726 16192 6735 16232
rect 6775 16192 6938 16232
rect 7180 16192 7204 16232
rect 7244 16192 7267 16232
rect 7354 16192 7363 16232
rect 7403 16192 7412 16232
rect 7471 16192 7480 16232
rect 7520 16192 7529 16232
rect 7576 16192 7612 16232
rect 7745 16192 7754 16232
rect 7794 16192 7803 16232
rect 7901 16192 7917 16232
rect 7957 16192 7966 16232
rect 8070 16192 8079 16232
rect 8119 16192 8236 16232
rect 8276 16192 8285 16232
rect 8362 16192 8371 16232
rect 8411 16192 8420 16232
rect 8611 16192 8620 16232
rect 8660 16192 8669 16232
rect 8794 16192 8803 16232
rect 8852 16192 8983 16232
rect 9100 16192 9331 16232
rect 9371 16192 9380 16232
rect 10147 16192 10156 16232
rect 10196 16192 10205 16232
rect 10384 16192 10393 16232
rect 10433 16192 10444 16232
rect 10484 16192 10573 16232
rect 10618 16192 10627 16232
rect 10667 16192 10676 16232
rect 10723 16192 10732 16232
rect 10772 16192 10972 16232
rect 11012 16192 11021 16232
rect 11142 16192 11151 16232
rect 11191 16192 11212 16232
rect 11252 16192 11322 16232
rect 11539 16192 11548 16232
rect 11588 16192 11597 16232
rect 11718 16192 11727 16232
rect 11767 16192 11788 16232
rect 11828 16192 11898 16232
rect 11971 16192 11980 16232
rect 12045 16192 12151 16232
rect 2860 16183 2900 16192
rect 3361 16148 3401 16192
rect 3724 16148 3764 16192
rect 4108 16148 4148 16192
rect 940 16108 1556 16148
rect 2552 16108 2561 16148
rect 2612 16108 2732 16148
rect 3361 16108 3628 16148
rect 3668 16108 4148 16148
rect 4361 16108 4492 16148
rect 4532 16108 4541 16148
rect 1516 16064 1556 16108
rect 1289 16024 1411 16064
rect 1460 16024 1469 16064
rect 1516 16024 2179 16064
rect 2219 16024 2228 16064
rect 2275 16024 2284 16064
rect 2324 16024 2333 16064
rect 2633 16024 2764 16064
rect 2804 16024 2813 16064
rect 2956 16024 3187 16064
rect 3227 16024 3236 16064
rect 3331 16024 3340 16064
rect 3380 16024 4012 16064
rect 4052 16024 4061 16064
rect 2284 15980 2324 16024
rect 2956 15980 2996 16024
rect 4588 15980 4628 16192
rect 4854 16148 4894 16192
rect 5077 16148 5117 16192
rect 4854 16108 4916 16148
rect 5030 16108 5068 16148
rect 5108 16108 5117 16148
rect 5303 16148 5343 16192
rect 5742 16148 5782 16192
rect 6220 16148 6260 16192
rect 5303 16108 5684 16148
rect 5742 16108 6124 16148
rect 6164 16108 6173 16148
rect 6220 16108 6316 16148
rect 6356 16108 6365 16148
rect 4876 15980 4916 16108
rect 5644 16064 5684 16108
rect 6466 16064 6506 16192
rect 6898 16148 6938 16192
rect 6898 16108 6988 16148
rect 7028 16108 7037 16148
rect 5644 16024 6124 16064
rect 6164 16024 6506 16064
rect 6787 16024 6796 16064
rect 6836 16024 7267 16064
rect 7307 16024 7316 16064
rect 5530 15982 5539 16022
rect 5579 15982 5588 16022
rect 6682 15982 6691 16022
rect 6731 15982 6740 16022
rect 5548 15980 5588 15982
rect 2284 15940 2956 15980
rect 2996 15940 3005 15980
rect 4588 15940 4820 15980
rect 4876 15940 5164 15980
rect 5204 15940 5213 15980
rect 5548 15940 6220 15980
rect 6260 15940 6269 15980
rect 2467 15856 2476 15896
rect 2516 15856 2525 15896
rect 4343 15856 4352 15896
rect 4720 15856 4729 15896
rect 2476 15812 2516 15856
rect 1996 15772 2516 15812
rect 2563 15772 2572 15812
rect 2612 15772 2996 15812
rect 1996 15728 2036 15772
rect 2572 15728 2612 15772
rect 2956 15728 2996 15772
rect 3436 15772 4394 15812
rect 3436 15728 3476 15772
rect 1027 15688 1036 15728
rect 1076 15688 1507 15728
rect 1547 15688 1556 15728
rect 1603 15688 1612 15728
rect 1652 15688 1708 15728
rect 1748 15688 1783 15728
rect 1978 15688 1987 15728
rect 2027 15688 2036 15728
rect 2092 15688 2612 15728
rect 2947 15688 2956 15728
rect 2996 15688 3005 15728
rect 3305 15688 3436 15728
rect 3476 15688 3485 15728
rect 3881 15688 4003 15728
rect 4052 15688 4061 15728
rect 0 15644 400 15664
rect 0 15604 1420 15644
rect 1460 15604 1469 15644
rect 0 15584 400 15604
rect 2092 15560 2132 15688
rect 2275 15604 2284 15644
rect 2324 15604 2367 15644
rect 2327 15560 2367 15604
rect 2476 15604 2668 15644
rect 2708 15604 2717 15644
rect 2851 15604 2860 15644
rect 2900 15604 3092 15644
rect 3209 15604 3233 15644
rect 3273 15604 3340 15644
rect 3380 15604 3389 15644
rect 3706 15604 3715 15644
rect 3755 15604 4052 15644
rect 2476 15560 2516 15604
rect 3052 15560 3092 15604
rect 4012 15560 4052 15604
rect 4354 15560 4394 15772
rect 4780 15728 4820 15940
rect 6700 15896 6740 15982
rect 7372 15980 7412 16192
rect 7612 16183 7652 16192
rect 7756 16148 7796 16192
rect 7926 16148 7966 16192
rect 8380 16148 8420 16192
rect 7716 16108 7756 16148
rect 7796 16108 7805 16148
rect 7926 16108 7948 16148
rect 7988 16108 7997 16148
rect 8380 16108 9100 16148
rect 9140 16108 9532 16148
rect 9572 16108 9676 16148
rect 9716 16108 9964 16148
rect 10004 16108 10013 16148
rect 8380 16064 8420 16108
rect 10156 16064 10196 16192
rect 10636 16148 10676 16192
rect 10243 16108 10252 16148
rect 10292 16108 10676 16148
rect 10972 16148 11012 16192
rect 11548 16148 11588 16192
rect 10972 16108 11588 16148
rect 12223 16148 12263 16276
rect 12586 16307 12652 16316
rect 12586 16267 12595 16307
rect 12635 16276 12652 16307
rect 12692 16276 12775 16316
rect 12931 16276 12940 16316
rect 12980 16276 12989 16316
rect 13153 16276 13195 16316
rect 13276 16276 13556 16316
rect 12635 16267 12644 16276
rect 13153 16274 13193 16276
rect 12586 16266 12644 16267
rect 13114 16234 13123 16274
rect 13163 16234 13193 16274
rect 13276 16232 13316 16276
rect 12329 16192 12460 16232
rect 12500 16192 12509 16232
rect 12691 16192 12700 16232
rect 12740 16192 12749 16232
rect 12802 16192 12811 16232
rect 12851 16192 12940 16232
rect 12980 16192 12991 16232
rect 13260 16192 13269 16232
rect 13309 16192 13318 16232
rect 12223 16108 12500 16148
rect 11713 16066 11800 16106
rect 11840 16066 11849 16106
rect 11713 16064 11753 16066
rect 7555 16024 7564 16064
rect 7604 16024 8420 16064
rect 9235 16024 9244 16064
rect 9284 16024 9428 16064
rect 9475 16024 9484 16064
rect 9524 16024 10060 16064
rect 10100 16024 10109 16064
rect 10156 16024 11753 16064
rect 12355 16024 12364 16064
rect 12404 16024 12413 16064
rect 6979 15940 6988 15980
rect 7028 15940 7412 15980
rect 9388 15980 9428 16024
rect 12364 15980 12404 16024
rect 9388 15940 11308 15980
rect 11348 15940 11357 15980
rect 11587 15940 11596 15980
rect 11636 15940 12404 15980
rect 12460 15980 12500 16108
rect 12700 16064 12740 16192
rect 13381 16165 13411 16205
rect 13451 16165 13460 16205
rect 13381 16148 13421 16165
rect 13516 16148 13556 16276
rect 13694 16276 13708 16316
rect 13748 16276 13757 16316
rect 13694 16232 13734 16276
rect 13804 16232 13844 16360
rect 14083 16276 14092 16316
rect 14132 16276 14228 16316
rect 13606 16192 13615 16232
rect 13655 16192 13734 16232
rect 13786 16192 13795 16232
rect 13835 16192 13844 16232
rect 13891 16203 13900 16243
rect 13940 16203 13949 16243
rect 14188 16232 14228 16276
rect 15052 16232 15092 16360
rect 15295 16360 15820 16400
rect 15860 16360 16820 16400
rect 17347 16360 17356 16400
rect 17396 16360 17405 16400
rect 17500 16360 17876 16400
rect 15295 16243 15335 16360
rect 15523 16276 15532 16316
rect 15572 16276 16052 16316
rect 16099 16276 16108 16316
rect 16148 16276 16532 16316
rect 13900 16148 13940 16203
rect 13315 16108 13324 16148
rect 13364 16108 13421 16148
rect 13507 16108 13516 16148
rect 13556 16108 13940 16148
rect 13996 16192 14045 16232
rect 14085 16192 14094 16232
rect 14170 16192 14179 16232
rect 14219 16192 14228 16232
rect 14345 16192 14356 16232
rect 14396 16192 14476 16232
rect 14516 16192 14525 16232
rect 14659 16192 14668 16232
rect 14708 16192 14884 16232
rect 14924 16192 14933 16232
rect 15034 16192 15043 16232
rect 15083 16192 15092 16232
rect 15151 16192 15160 16232
rect 15200 16192 15209 16232
rect 15283 16203 15292 16243
rect 15332 16203 15341 16243
rect 16012 16232 16052 16276
rect 16492 16232 16532 16276
rect 16670 16276 16684 16316
rect 16724 16276 16733 16316
rect 16670 16232 16710 16276
rect 16780 16232 16820 16360
rect 17356 16316 17396 16360
rect 17500 16316 17540 16360
rect 17836 16316 17876 16360
rect 17129 16276 17260 16316
rect 17300 16276 17309 16316
rect 17356 16276 17540 16316
rect 17596 16276 17644 16316
rect 17684 16276 17693 16316
rect 17818 16276 17827 16316
rect 17867 16276 17876 16316
rect 17932 16316 17972 16444
rect 19372 16400 19412 16444
rect 19084 16360 19412 16400
rect 20297 16360 20428 16400
rect 20468 16360 20477 16400
rect 20524 16360 21484 16400
rect 21524 16360 21533 16400
rect 21754 16360 21763 16400
rect 21803 16360 22252 16400
rect 22292 16360 22301 16400
rect 24259 16360 24268 16400
rect 24308 16360 25420 16400
rect 25460 16360 25469 16400
rect 26179 16360 26188 16400
rect 26228 16360 27188 16400
rect 17932 16276 18028 16316
rect 18068 16276 18077 16316
rect 17596 16232 17636 16276
rect 19084 16274 19124 16360
rect 19241 16276 19372 16316
rect 19412 16276 19421 16316
rect 19564 16276 20236 16316
rect 20276 16276 20285 16316
rect 19018 16234 19027 16274
rect 19067 16234 19124 16274
rect 19564 16232 19604 16276
rect 20524 16232 20564 16360
rect 21868 16276 22348 16316
rect 22388 16276 22772 16316
rect 22819 16276 22828 16316
rect 22868 16276 23596 16316
rect 23636 16276 23645 16316
rect 23884 16276 24596 16316
rect 25699 16276 25708 16316
rect 25748 16276 26420 16316
rect 26729 16276 26860 16316
rect 26900 16276 26909 16316
rect 21868 16232 21908 16276
rect 22732 16232 22772 16276
rect 23212 16232 23252 16276
rect 15418 16192 15427 16232
rect 15467 16192 15476 16232
rect 15622 16192 15631 16232
rect 15671 16192 15680 16232
rect 15728 16192 15737 16232
rect 15777 16192 15786 16232
rect 15894 16192 15903 16232
rect 15943 16192 15956 16232
rect 16002 16192 16011 16232
rect 16051 16192 16060 16232
rect 16108 16192 16137 16232
rect 16177 16192 16186 16232
rect 16378 16192 16387 16232
rect 16427 16192 16436 16232
rect 16492 16192 16505 16232
rect 16545 16192 16554 16232
rect 16600 16192 16665 16232
rect 16705 16192 16714 16232
rect 16762 16192 16771 16232
rect 16811 16192 16820 16232
rect 16867 16192 16876 16232
rect 16945 16192 17047 16232
rect 17107 16192 17116 16232
rect 17156 16192 17165 16232
rect 17321 16192 17431 16232
rect 17492 16192 17501 16232
rect 17578 16192 17587 16232
rect 17627 16192 17636 16232
rect 17683 16192 17692 16232
rect 17732 16192 17741 16232
rect 17827 16192 17836 16232
rect 17876 16192 17932 16232
rect 17972 16192 18007 16232
rect 18499 16192 18508 16232
rect 18560 16192 18679 16232
rect 19555 16192 19564 16232
rect 19604 16192 19613 16232
rect 19721 16223 19852 16232
rect 19721 16192 19843 16223
rect 19892 16192 19901 16232
rect 20131 16192 20140 16232
rect 20180 16192 20564 16232
rect 20777 16192 20908 16232
rect 20948 16192 20957 16232
rect 21065 16192 21187 16232
rect 21236 16192 21245 16232
rect 21868 16192 21964 16232
rect 22004 16192 22013 16232
rect 22060 16192 22085 16232
rect 22125 16192 22134 16232
rect 22478 16192 22487 16232
rect 22527 16192 22536 16232
rect 22588 16223 22676 16232
rect 13996 16148 14036 16192
rect 15160 16148 15200 16192
rect 15436 16148 15476 16192
rect 15640 16148 15680 16192
rect 13996 16108 14380 16148
rect 14420 16108 15200 16148
rect 15341 16108 15476 16148
rect 15593 16108 15628 16148
rect 15668 16108 15680 16148
rect 13996 16064 14036 16108
rect 12700 16024 13076 16064
rect 13481 16024 13603 16064
rect 13652 16024 13661 16064
rect 13708 16024 14036 16064
rect 14266 16024 14275 16064
rect 14315 16024 14324 16064
rect 13036 15980 13076 16024
rect 13708 15980 13748 16024
rect 14284 15980 14324 16024
rect 12460 15940 12940 15980
rect 12980 15940 12989 15980
rect 13036 15940 13324 15980
rect 13364 15940 13373 15980
rect 13699 15940 13708 15980
rect 13748 15940 13757 15980
rect 14284 15940 14668 15980
rect 14708 15940 14717 15980
rect 6700 15856 7852 15896
rect 7892 15856 8812 15896
rect 8852 15856 8861 15896
rect 12117 15856 12126 15896
rect 12494 15856 12503 15896
rect 12988 15856 14284 15896
rect 14324 15856 14333 15896
rect 4867 15772 4876 15812
rect 4916 15772 6356 15812
rect 6316 15728 6356 15772
rect 4474 15688 4483 15728
rect 4523 15688 4820 15728
rect 4867 15688 4876 15728
rect 4916 15688 5356 15728
rect 5396 15688 5405 15728
rect 5609 15688 5740 15728
rect 5780 15688 5789 15728
rect 6298 15688 6307 15728
rect 6347 15688 6356 15728
rect 7276 15772 7660 15812
rect 7700 15772 7709 15812
rect 7948 15772 8524 15812
rect 8564 15772 11060 15812
rect 5155 15604 5164 15644
rect 5204 15604 5243 15644
rect 5443 15604 5452 15644
rect 5492 15604 5876 15644
rect 5203 15560 5243 15604
rect 5836 15560 5876 15604
rect 6067 15604 6124 15644
rect 6164 15604 6173 15644
rect 6403 15604 6412 15644
rect 6452 15604 7180 15644
rect 7220 15604 7229 15644
rect 6067 15560 6107 15604
rect 7276 15560 7316 15772
rect 7625 15688 7756 15728
rect 7796 15688 7805 15728
rect 7363 15604 7372 15644
rect 7412 15604 7421 15644
rect 7651 15604 7660 15644
rect 7700 15604 7709 15644
rect 7372 15560 7412 15604
rect 7660 15560 7700 15604
rect 7948 15560 7988 15772
rect 11020 15728 11060 15772
rect 8035 15688 8044 15728
rect 8084 15688 8140 15728
rect 8180 15688 8215 15728
rect 8279 15688 8428 15728
rect 8468 15688 8477 15728
rect 8611 15688 8620 15728
rect 8660 15688 10444 15728
rect 10484 15688 10493 15728
rect 10627 15688 10636 15728
rect 10676 15688 10732 15728
rect 10772 15688 10807 15728
rect 11020 15688 12028 15728
rect 12068 15688 12077 15728
rect 8279 15644 8319 15688
rect 12988 15644 13028 15856
rect 15341 15812 15381 16108
rect 15746 16064 15786 16192
rect 15916 16148 15956 16192
rect 16108 16148 16148 16192
rect 16396 16148 16436 16192
rect 15916 16108 15982 16148
rect 16099 16108 16108 16148
rect 16148 16108 16157 16148
rect 16396 16108 16492 16148
rect 16532 16108 16541 16148
rect 15427 16024 15436 16064
rect 15476 16024 15786 16064
rect 15942 16064 15982 16108
rect 16600 16064 16640 16192
rect 17116 16148 17156 16192
rect 17692 16148 17732 16192
rect 19834 16183 19843 16192
rect 19883 16183 19892 16192
rect 19834 16182 19892 16183
rect 22060 16148 22100 16192
rect 15942 16024 16640 16064
rect 16695 16108 17156 16148
rect 17539 16108 17548 16148
rect 17588 16108 17732 16148
rect 18124 16108 19132 16148
rect 19172 16108 19181 16148
rect 19939 16108 19948 16148
rect 19988 16108 20332 16148
rect 20372 16108 20381 16148
rect 20524 16108 21292 16148
rect 21332 16108 21341 16148
rect 21955 16108 21964 16148
rect 22004 16108 22100 16148
rect 16695 15980 16735 16108
rect 18124 16064 18164 16108
rect 16858 16024 16867 16064
rect 16907 16024 16972 16064
rect 17012 16024 17047 16064
rect 17164 16024 18164 16064
rect 18346 16024 18355 16064
rect 18395 16024 18404 16064
rect 18595 16024 18604 16064
rect 18644 16024 18835 16064
rect 18875 16024 18884 16064
rect 19699 16024 19708 16064
rect 19748 16024 19756 16064
rect 19796 16024 19879 16064
rect 17164 15980 17204 16024
rect 18364 15980 18404 16024
rect 20524 15980 20564 16108
rect 22487 16064 22527 16192
rect 21929 16024 22060 16064
rect 22100 16024 22527 16064
rect 22588 16183 22627 16223
rect 22667 16183 22676 16223
rect 22723 16192 22732 16232
rect 22772 16192 22781 16232
rect 23203 16192 23212 16232
rect 23252 16192 23261 16232
rect 23369 16192 23491 16232
rect 23540 16192 23549 16232
rect 22588 16182 22676 16183
rect 22588 15980 22628 16182
rect 23884 16148 23924 16276
rect 24556 16232 24596 16276
rect 26380 16232 26420 16276
rect 27148 16232 27188 16360
rect 27619 16276 27628 16316
rect 27668 16276 28532 16316
rect 27436 16232 27476 16241
rect 27964 16232 28004 16276
rect 28492 16232 28532 16276
rect 28684 16274 28724 16528
rect 28771 16360 28780 16400
rect 28820 16360 29068 16400
rect 29108 16360 29117 16400
rect 28675 16234 28684 16274
rect 28724 16234 28733 16274
rect 24110 16192 24119 16232
rect 24159 16192 24168 16232
rect 24250 16223 24308 16232
rect 23587 16108 23596 16148
rect 23636 16108 23692 16148
rect 23732 16108 23924 16148
rect 24119 16064 24159 16192
rect 24250 16183 24259 16223
rect 24299 16183 24308 16223
rect 24355 16192 24364 16232
rect 24404 16192 24413 16232
rect 24547 16192 24556 16232
rect 24596 16192 25228 16232
rect 25268 16192 25277 16232
rect 25891 16192 25900 16232
rect 25940 16192 26092 16232
rect 26132 16192 26141 16232
rect 26362 16192 26371 16232
rect 26411 16192 26420 16232
rect 26467 16192 26476 16232
rect 26516 16192 26647 16232
rect 26755 16192 26764 16232
rect 26804 16192 26956 16232
rect 26996 16192 27005 16232
rect 27148 16192 27436 16232
rect 27946 16192 27955 16232
rect 27995 16192 28004 16232
rect 28169 16192 28300 16232
rect 28340 16192 28349 16232
rect 28483 16192 28492 16232
rect 28532 16192 28541 16232
rect 28867 16192 28876 16232
rect 28916 16192 28925 16232
rect 24250 16182 24308 16183
rect 24266 16064 24306 16182
rect 24364 16148 24404 16192
rect 27436 16183 27476 16192
rect 28876 16148 28916 16192
rect 24364 16108 24556 16148
rect 24596 16108 24605 16148
rect 25219 16108 25228 16148
rect 25268 16108 27380 16148
rect 27340 16064 27380 16108
rect 28012 16108 28916 16148
rect 28012 16064 28052 16108
rect 23491 16024 23500 16064
rect 23540 16024 24159 16064
rect 24259 16024 24268 16064
rect 24308 16024 24317 16064
rect 25411 16024 25420 16064
rect 25460 16024 25708 16064
rect 25748 16024 25757 16064
rect 27340 16024 28052 16064
rect 28099 16024 28108 16064
rect 28148 16024 28279 16064
rect 28361 16024 28396 16064
rect 28436 16024 28492 16064
rect 28532 16024 28541 16064
rect 28771 16024 28780 16064
rect 28820 16024 28829 16064
rect 28780 15980 28820 16024
rect 16003 15940 16012 15980
rect 16052 15940 16492 15980
rect 16532 15940 16735 15980
rect 16867 15940 16876 15980
rect 16916 15940 17204 15980
rect 18019 15940 18028 15980
rect 18068 15940 18404 15980
rect 19555 15940 19564 15980
rect 19604 15940 20564 15980
rect 21955 15940 21964 15980
rect 22004 15940 22628 15980
rect 25996 15940 28820 15980
rect 16073 15856 16204 15896
rect 16244 15856 17972 15896
rect 19891 15856 19900 15896
rect 20268 15856 20277 15896
rect 23779 15856 23788 15896
rect 23828 15856 25268 15896
rect 13123 15772 13132 15812
rect 13172 15772 13700 15812
rect 15341 15772 16052 15812
rect 13660 15728 13700 15772
rect 16012 15728 16052 15772
rect 8044 15604 8319 15644
rect 8428 15604 8524 15644
rect 8564 15604 8573 15644
rect 8707 15604 8716 15644
rect 8756 15604 8765 15644
rect 8986 15604 8995 15644
rect 9035 15604 9044 15644
rect 9379 15604 9388 15644
rect 9428 15604 9772 15644
rect 9812 15604 9821 15644
rect 9955 15604 9964 15644
rect 10004 15635 10868 15644
rect 10004 15604 10819 15635
rect 8044 15560 8084 15604
rect 8428 15560 8468 15604
rect 8716 15560 8756 15604
rect 643 15520 652 15560
rect 692 15520 931 15560
rect 971 15520 980 15560
rect 1097 15520 1228 15560
rect 1268 15520 1277 15560
rect 1400 15520 1409 15560
rect 1449 15520 1612 15560
rect 1652 15520 1661 15560
rect 1708 15551 1748 15560
rect 1891 15520 1900 15560
rect 1940 15520 2132 15560
rect 2179 15520 2188 15560
rect 2228 15520 2237 15560
rect 2318 15520 2327 15560
rect 2367 15520 2376 15560
rect 2458 15520 2467 15560
rect 2507 15520 2516 15560
rect 2563 15520 2572 15560
rect 2612 15520 2621 15560
rect 2851 15520 2860 15560
rect 2900 15520 2909 15560
rect 3043 15520 3052 15560
rect 3092 15520 3101 15560
rect 3532 15551 3572 15560
rect 1219 15352 1228 15392
rect 1268 15352 1516 15392
rect 1556 15352 1565 15392
rect 1708 15308 1748 15511
rect 2188 15392 2228 15520
rect 2572 15476 2612 15520
rect 2860 15476 2900 15520
rect 3785 15520 3820 15560
rect 3860 15520 3916 15560
rect 3956 15520 3965 15560
rect 4012 15520 4151 15560
rect 4191 15520 4200 15560
rect 4354 15520 4396 15560
rect 4436 15520 4567 15560
rect 4963 15520 4972 15560
rect 5012 15520 5021 15560
rect 5194 15520 5203 15560
rect 5243 15520 5252 15560
rect 5347 15520 5356 15560
rect 5396 15520 5405 15560
rect 5539 15520 5548 15560
rect 5588 15520 5719 15560
rect 5827 15520 5836 15560
rect 5876 15520 5885 15560
rect 6058 15520 6067 15560
rect 6107 15520 6116 15560
rect 6202 15520 6211 15560
rect 6260 15520 6391 15560
rect 6510 15520 6519 15560
rect 6559 15520 6568 15560
rect 6665 15520 6796 15560
rect 6836 15520 6845 15560
rect 6970 15520 6979 15560
rect 7019 15520 7084 15560
rect 7124 15520 7159 15560
rect 7267 15520 7276 15560
rect 7316 15520 7325 15560
rect 7372 15520 7493 15560
rect 7533 15520 7542 15560
rect 7651 15520 7660 15560
rect 7700 15520 7747 15560
rect 7834 15520 7843 15560
rect 7883 15520 7988 15560
rect 8035 15520 8044 15560
rect 8084 15520 8093 15560
rect 8419 15520 8428 15560
rect 8468 15520 8477 15560
rect 8669 15520 8683 15560
rect 8723 15520 8756 15560
rect 8899 15520 8908 15560
rect 8948 15520 8957 15560
rect 2371 15436 2380 15476
rect 2420 15436 2612 15476
rect 2659 15436 2668 15476
rect 2708 15436 2717 15476
rect 2860 15436 2956 15476
rect 2996 15436 3127 15476
rect 2188 15352 2572 15392
rect 2612 15352 2621 15392
rect 2668 15308 2708 15436
rect 1708 15268 2708 15308
rect 0 15224 400 15244
rect 3052 15224 3092 15436
rect 3532 15392 3572 15511
rect 4169 15436 4291 15476
rect 4340 15436 4349 15476
rect 3532 15352 3956 15392
rect 3226 15268 3235 15308
rect 3275 15268 3820 15308
rect 3860 15268 3869 15308
rect 3916 15224 3956 15352
rect 0 15184 2476 15224
rect 2516 15184 2525 15224
rect 3052 15184 3572 15224
rect 3916 15184 4780 15224
rect 4820 15184 4829 15224
rect 0 15164 400 15184
rect 3532 15140 3572 15184
rect 3103 15100 3112 15140
rect 3480 15100 3489 15140
rect 3532 15100 4012 15140
rect 4052 15100 4061 15140
rect 4972 14972 5012 15520
rect 5356 15476 5396 15520
rect 5082 15436 5091 15476
rect 5131 15436 5396 15476
rect 5824 15436 5932 15476
rect 5995 15436 6004 15476
rect 6124 15436 6412 15476
rect 6452 15436 6461 15476
rect 5356 15392 5396 15436
rect 6124 15392 6164 15436
rect 6519 15392 6559 15520
rect 8044 15476 8084 15520
rect 8227 15478 8236 15518
rect 8276 15478 8285 15518
rect 7386 15436 7395 15476
rect 7435 15436 8084 15476
rect 8236 15392 8276 15478
rect 8419 15436 8428 15476
rect 8468 15436 8803 15476
rect 8843 15436 8852 15476
rect 5356 15352 6164 15392
rect 6307 15352 6316 15392
rect 6356 15352 6559 15392
rect 7843 15352 7852 15392
rect 7892 15352 8276 15392
rect 5443 15268 5452 15308
rect 5492 15268 5548 15308
rect 5588 15268 5623 15308
rect 5731 15268 5740 15308
rect 5780 15268 6508 15308
rect 6548 15268 6557 15308
rect 6691 15268 6700 15308
rect 6740 15268 6979 15308
rect 7019 15268 7028 15308
rect 8563 15268 8572 15308
rect 8612 15268 8812 15308
rect 8852 15268 8861 15308
rect 8908 15224 8948 15520
rect 9004 15476 9044 15604
rect 9580 15560 9620 15604
rect 10810 15595 10819 15604
rect 10859 15595 10868 15635
rect 10915 15604 10924 15644
rect 10964 15604 11007 15644
rect 11299 15604 11308 15644
rect 11348 15604 11636 15644
rect 12344 15604 12353 15644
rect 12393 15604 13028 15644
rect 13180 15688 13228 15728
rect 13268 15688 13516 15728
rect 13556 15688 13565 15728
rect 13660 15688 13804 15728
rect 13844 15688 13853 15728
rect 13982 15688 14860 15728
rect 14900 15688 14909 15728
rect 15427 15688 15436 15728
rect 15476 15688 15956 15728
rect 16003 15688 16012 15728
rect 16052 15688 16061 15728
rect 10810 15594 10868 15595
rect 10920 15560 10960 15604
rect 9091 15520 9100 15560
rect 9140 15520 9283 15560
rect 9323 15520 9332 15560
rect 9562 15520 9571 15560
rect 9611 15520 9620 15560
rect 10051 15520 10060 15560
rect 10100 15520 10109 15560
rect 10243 15520 10252 15560
rect 10317 15520 10423 15560
rect 10492 15520 10523 15560
rect 10563 15520 10572 15560
rect 10678 15520 10687 15560
rect 10727 15520 10736 15560
rect 10902 15520 10911 15560
rect 10951 15520 10960 15560
rect 11083 15520 11092 15560
rect 11156 15520 11272 15560
rect 11380 15520 11452 15560
rect 11492 15520 11501 15560
rect 9004 15436 9187 15476
rect 9227 15436 9236 15476
rect 9667 15436 9676 15476
rect 9716 15436 9724 15476
rect 9764 15436 9847 15476
rect 9955 15436 9964 15476
rect 10004 15436 10013 15476
rect 9964 15392 10004 15436
rect 8515 15184 8524 15224
rect 8564 15184 8948 15224
rect 9004 15352 10004 15392
rect 9004 15056 9044 15352
rect 10060 15308 10100 15520
rect 10492 15476 10532 15520
rect 10684 15476 10724 15520
rect 10170 15436 10179 15476
rect 10219 15436 10348 15476
rect 10388 15436 10397 15476
rect 10492 15436 10540 15476
rect 10580 15436 10589 15476
rect 10684 15436 10732 15476
rect 10772 15436 10781 15476
rect 11380 15392 11420 15520
rect 11596 15476 11636 15604
rect 13180 15602 13220 15688
rect 13180 15562 13219 15602
rect 13259 15562 13268 15602
rect 13982 15560 14022 15688
rect 14158 15604 14284 15644
rect 14324 15604 14333 15644
rect 15139 15604 15148 15644
rect 15188 15604 15380 15644
rect 15497 15604 15628 15644
rect 15668 15604 15677 15644
rect 14158 15560 14198 15604
rect 15340 15560 15380 15604
rect 15916 15560 15956 15688
rect 16108 15560 16148 15856
rect 16876 15772 17836 15812
rect 17876 15772 17885 15812
rect 16876 15728 16916 15772
rect 17932 15728 17972 15856
rect 18403 15772 18412 15812
rect 18452 15772 21676 15812
rect 21716 15772 21725 15812
rect 22924 15772 24268 15812
rect 24308 15772 24317 15812
rect 16858 15688 16867 15728
rect 16907 15688 16916 15728
rect 17251 15688 17260 15728
rect 17300 15688 17827 15728
rect 17867 15688 17876 15728
rect 17923 15688 17932 15728
rect 17972 15688 18316 15728
rect 18356 15688 18365 15728
rect 20419 15688 20428 15728
rect 20468 15688 21154 15728
rect 21763 15688 21772 15728
rect 21812 15688 21964 15728
rect 22004 15688 22013 15728
rect 22217 15688 22339 15728
rect 22388 15688 22397 15728
rect 21114 15644 21154 15688
rect 22924 15644 22964 15772
rect 25228 15728 25268 15856
rect 23011 15688 23020 15728
rect 23060 15688 23252 15728
rect 23299 15688 23308 15728
rect 23348 15688 23357 15728
rect 23500 15688 23788 15728
rect 23828 15688 23837 15728
rect 24809 15688 24940 15728
rect 24980 15688 24989 15728
rect 25210 15688 25219 15728
rect 25259 15688 25268 15728
rect 25769 15688 25900 15728
rect 25940 15688 25949 15728
rect 23212 15644 23252 15688
rect 17240 15604 17249 15644
rect 17289 15604 17726 15644
rect 17766 15604 17775 15644
rect 17923 15604 17932 15644
rect 17972 15604 17981 15644
rect 18176 15604 18220 15644
rect 18260 15604 18269 15644
rect 18508 15604 19180 15644
rect 19220 15604 19229 15644
rect 19363 15604 19372 15644
rect 19412 15604 19421 15644
rect 19468 15604 19852 15644
rect 19892 15604 19901 15644
rect 20044 15604 21004 15644
rect 21044 15604 21053 15644
rect 21105 15604 21114 15644
rect 21154 15604 22156 15644
rect 22196 15604 22205 15644
rect 22540 15604 22636 15644
rect 22676 15604 22685 15644
rect 22793 15604 22842 15644
rect 22882 15604 22924 15644
rect 22964 15604 22973 15644
rect 23194 15604 23203 15644
rect 23243 15604 23252 15644
rect 17260 15560 17300 15604
rect 17932 15560 17972 15604
rect 18223 15560 18263 15604
rect 18508 15560 18548 15604
rect 19372 15560 19412 15604
rect 19468 15560 19508 15604
rect 11875 15520 11884 15560
rect 11947 15520 12055 15560
rect 12163 15520 12172 15560
rect 12212 15520 12343 15560
rect 12547 15520 12556 15560
rect 12596 15520 12605 15560
rect 12652 15551 12692 15560
rect 11770 15478 11779 15518
rect 11819 15478 11828 15518
rect 11587 15436 11596 15476
rect 11636 15436 11645 15476
rect 10540 15352 11420 15392
rect 11491 15352 11500 15392
rect 11540 15352 11692 15392
rect 11732 15352 11741 15392
rect 10540 15308 10580 15352
rect 10060 15268 10348 15308
rect 10388 15268 10397 15308
rect 10522 15268 10531 15308
rect 10571 15268 10580 15308
rect 9475 15184 9484 15224
rect 9524 15184 10540 15224
rect 10580 15184 10589 15224
rect 9379 15100 9388 15140
rect 9428 15100 10444 15140
rect 10484 15100 10493 15140
rect 10877 15100 10886 15140
rect 11254 15100 11263 15140
rect 5742 15016 9044 15056
rect 9475 15016 9484 15056
rect 9524 15016 11596 15056
rect 11636 15016 11645 15056
rect 929 14932 1804 14972
rect 1844 14932 1853 14972
rect 4666 14932 4675 14972
rect 4715 14932 4876 14972
rect 4916 14932 4925 14972
rect 4972 14932 5068 14972
rect 5108 14932 5117 14972
rect 0 14804 400 14824
rect 929 14804 969 14932
rect 3139 14848 3148 14888
rect 3188 14848 3197 14888
rect 3994 14848 4003 14888
rect 4043 14848 5381 14888
rect 3148 14804 3188 14848
rect 0 14764 969 14804
rect 1018 14764 1027 14804
rect 1076 14764 1207 14804
rect 2083 14764 2092 14804
rect 2132 14764 2141 14804
rect 2938 14764 2947 14804
rect 2987 14764 3188 14804
rect 4387 14764 4396 14804
rect 4436 14764 5012 14804
rect 0 14744 400 14764
rect 4972 14720 5012 14764
rect 5341 14720 5381 14848
rect 5742 14804 5782 15016
rect 6691 14932 6700 14972
rect 6740 14932 7028 14972
rect 7075 14932 7084 14972
rect 7124 14932 9964 14972
rect 10004 14932 10013 14972
rect 5980 14848 6932 14888
rect 5980 14804 6020 14848
rect 5452 14764 5782 14804
rect 5827 14764 5836 14804
rect 5876 14764 5885 14804
rect 5971 14764 5980 14804
rect 6020 14764 6029 14804
rect 6281 14764 6403 14804
rect 6452 14764 6461 14804
rect 6595 14764 6604 14804
rect 6644 14764 6796 14804
rect 6836 14764 6845 14804
rect 5452 14720 5492 14764
rect 5836 14720 5876 14764
rect 2537 14680 2563 14720
rect 2603 14680 2668 14720
rect 2708 14680 2717 14720
rect 3017 14680 3148 14720
rect 3188 14680 3197 14720
rect 3264 14680 3273 14720
rect 3313 14680 3380 14720
rect 3427 14680 3436 14720
rect 3476 14680 3628 14720
rect 3668 14680 3677 14720
rect 3811 14680 3820 14720
rect 3860 14680 3869 14720
rect 3994 14680 4003 14720
rect 4043 14680 4204 14720
rect 4244 14680 4253 14720
rect 4300 14680 4481 14720
rect 4521 14680 4530 14720
rect 4579 14680 4588 14720
rect 4628 14680 4759 14720
rect 4963 14680 4972 14720
rect 5012 14680 5021 14720
rect 5155 14680 5164 14720
rect 5204 14680 5213 14720
rect 5294 14680 5303 14720
rect 5343 14680 5381 14720
rect 5434 14680 5443 14720
rect 5483 14680 5492 14720
rect 5539 14680 5548 14720
rect 5588 14680 5719 14720
rect 5789 14680 5824 14720
rect 5864 14680 5876 14720
rect 5923 14680 5932 14720
rect 5972 14680 6263 14720
rect 6303 14680 6312 14720
rect 3340 14636 3380 14680
rect 3820 14636 3860 14680
rect 3340 14596 3724 14636
rect 3764 14596 3773 14636
rect 3820 14596 4108 14636
rect 4148 14596 4157 14636
rect 521 14512 652 14552
rect 692 14512 701 14552
rect 2659 14512 2668 14552
rect 2708 14512 3628 14552
rect 3668 14512 3677 14552
rect 4300 14468 4340 14680
rect 5164 14636 5204 14680
rect 5164 14596 5635 14636
rect 5675 14596 5684 14636
rect 6389 14552 6429 14764
rect 6892 14720 6932 14848
rect 6988 14804 7028 14932
rect 7171 14848 7180 14888
rect 7220 14848 7892 14888
rect 8515 14848 8524 14888
rect 8564 14848 8947 14888
rect 8987 14848 8996 14888
rect 9187 14848 9196 14888
rect 9236 14848 10916 14888
rect 11011 14848 11020 14888
rect 11060 14848 11191 14888
rect 7852 14804 7892 14848
rect 10876 14804 10916 14848
rect 11788 14804 11828 15478
rect 12233 15268 12355 15308
rect 12404 15268 12413 15308
rect 12556 14972 12596 15520
rect 12931 15520 12940 15560
rect 12980 15520 12989 15560
rect 13411 15520 13420 15560
rect 13460 15520 13469 15560
rect 13603 15520 13612 15560
rect 13652 15520 13844 15560
rect 13891 15520 13900 15560
rect 13940 15520 14022 15560
rect 14128 15520 14137 15560
rect 14177 15520 14198 15560
rect 14244 15520 14253 15560
rect 14293 15520 14324 15560
rect 14371 15520 14380 15560
rect 14441 15520 14551 15560
rect 14659 15520 14668 15560
rect 14733 15520 14839 15560
rect 15034 15520 15043 15560
rect 15083 15520 15244 15560
rect 15284 15520 15293 15560
rect 15340 15520 15532 15560
rect 15572 15520 15581 15560
rect 15715 15520 15724 15560
rect 15764 15520 15773 15560
rect 15907 15520 15916 15560
rect 15956 15520 15965 15560
rect 16099 15520 16108 15560
rect 16148 15520 16157 15560
rect 16666 15520 16675 15560
rect 16715 15520 16724 15560
rect 17251 15520 17260 15560
rect 17300 15520 17376 15560
rect 17443 15520 17452 15560
rect 17492 15520 17501 15560
rect 17548 15551 17588 15560
rect 12652 15308 12692 15511
rect 12787 15478 12796 15518
rect 12836 15478 12845 15518
rect 12796 15392 12836 15478
rect 12940 15476 12980 15520
rect 13114 15478 13123 15518
rect 13163 15478 13178 15518
rect 12893 15436 12938 15476
rect 12978 15436 12987 15476
rect 13138 15392 13178 15478
rect 13420 15476 13460 15520
rect 13804 15476 13844 15520
rect 14284 15476 14324 15520
rect 14693 15476 14733 15520
rect 15724 15476 15764 15520
rect 16108 15476 16148 15520
rect 16684 15476 16724 15520
rect 13420 15436 13708 15476
rect 13748 15436 13757 15476
rect 13804 15436 13877 15476
rect 14010 15436 14019 15476
rect 14059 15436 14198 15476
rect 14275 15436 14284 15476
rect 14324 15436 14349 15476
rect 14563 15436 14572 15476
rect 14612 15436 14621 15476
rect 14693 15448 15140 15476
rect 14693 15436 15091 15448
rect 12796 15352 12844 15392
rect 12884 15352 12893 15392
rect 13027 15352 13036 15392
rect 13076 15352 13085 15392
rect 13138 15352 13460 15392
rect 13507 15352 13516 15392
rect 13556 15352 13610 15392
rect 12652 15268 12940 15308
rect 12980 15268 12989 15308
rect 12556 14932 12844 14972
rect 12884 14932 12893 14972
rect 13036 14804 13076 15352
rect 13420 15308 13460 15352
rect 13411 15268 13420 15308
rect 13460 15268 13469 15308
rect 13570 15224 13610 15352
rect 13837 15308 13877 15436
rect 14158 15392 14198 15436
rect 14158 15352 14476 15392
rect 14516 15352 14525 15392
rect 13837 15268 14188 15308
rect 14228 15268 14237 15308
rect 13570 15184 13996 15224
rect 14036 15184 14045 15224
rect 14572 15056 14612 15436
rect 15082 15408 15091 15436
rect 15131 15408 15140 15448
rect 15724 15436 16148 15476
rect 16396 15436 16724 15476
rect 16396 15392 16436 15436
rect 17452 15392 17492 15520
rect 17932 15551 18068 15560
rect 17932 15520 18028 15551
rect 17548 15476 17588 15511
rect 18214 15520 18223 15560
rect 18263 15520 18272 15560
rect 18336 15520 18345 15560
rect 18385 15520 18452 15560
rect 18499 15520 18508 15560
rect 18548 15520 18557 15560
rect 18691 15520 18700 15560
rect 18740 15520 18743 15560
rect 18783 15520 18871 15560
rect 18979 15520 18988 15560
rect 19028 15520 19084 15560
rect 19124 15520 19159 15560
rect 19234 15520 19243 15560
rect 19283 15520 19412 15560
rect 19459 15520 19468 15560
rect 19508 15520 19517 15560
rect 19660 15520 19708 15560
rect 19748 15520 19757 15560
rect 19817 15520 19887 15560
rect 19927 15520 19948 15560
rect 19988 15520 19997 15560
rect 18028 15502 18068 15511
rect 18412 15476 18452 15520
rect 19660 15476 19700 15520
rect 20044 15476 20084 15604
rect 22156 15560 22196 15604
rect 22540 15560 22580 15604
rect 23310 15571 23350 15688
rect 20419 15520 20428 15560
rect 20468 15520 20599 15560
rect 20659 15520 20668 15560
rect 20708 15520 20717 15560
rect 20794 15520 20803 15560
rect 20843 15520 20852 15560
rect 20899 15520 20908 15560
rect 20948 15520 21079 15560
rect 21283 15520 21292 15560
rect 21332 15520 21484 15560
rect 21524 15520 21533 15560
rect 21737 15520 21823 15560
rect 21863 15520 21868 15560
rect 21908 15520 21917 15560
rect 22018 15520 22027 15560
rect 22067 15520 22196 15560
rect 22243 15520 22252 15560
rect 22292 15520 22423 15560
rect 22522 15520 22531 15560
rect 22571 15520 22580 15560
rect 22627 15520 22636 15560
rect 22676 15520 22685 15560
rect 23292 15531 23301 15571
rect 23341 15531 23350 15571
rect 23500 15560 23540 15688
rect 25996 15644 26036 15940
rect 27665 15856 27674 15896
rect 28042 15856 28051 15896
rect 28291 15772 28300 15812
rect 28340 15772 28780 15812
rect 28820 15772 28829 15812
rect 26947 15688 26956 15728
rect 26996 15688 28972 15728
rect 29012 15688 29021 15728
rect 23683 15604 23692 15644
rect 23732 15604 24116 15644
rect 24076 15560 24116 15604
rect 24556 15604 26036 15644
rect 27523 15604 27532 15644
rect 27572 15604 29300 15644
rect 24556 15560 24596 15604
rect 27820 15560 27860 15604
rect 29260 15560 29300 15604
rect 23491 15520 23500 15560
rect 23540 15520 23549 15560
rect 23700 15520 23788 15560
rect 23828 15520 23831 15560
rect 23871 15520 23880 15560
rect 23949 15551 24020 15560
rect 20170 15478 20179 15518
rect 20219 15478 20276 15518
rect 20236 15476 20276 15478
rect 20668 15476 20708 15520
rect 20812 15476 20852 15520
rect 22636 15476 22676 15520
rect 23949 15511 23971 15551
rect 24011 15511 24020 15551
rect 24067 15520 24076 15560
rect 24116 15520 24125 15560
rect 24538 15520 24547 15560
rect 24587 15520 24596 15560
rect 24643 15520 24652 15560
rect 24692 15520 24748 15560
rect 24788 15520 24823 15560
rect 25289 15520 25420 15560
rect 25460 15520 25469 15560
rect 25577 15520 25708 15560
rect 25748 15520 25757 15560
rect 26284 15520 26764 15560
rect 26804 15520 26813 15560
rect 27689 15520 27811 15560
rect 27860 15520 27869 15560
rect 28099 15520 28108 15560
rect 28148 15520 28195 15560
rect 28235 15520 28279 15560
rect 28378 15551 28396 15560
rect 23949 15510 24020 15511
rect 23949 15476 23989 15510
rect 17548 15436 17932 15476
rect 17972 15436 17981 15476
rect 18403 15436 18412 15476
rect 18452 15436 18604 15476
rect 18644 15436 18653 15476
rect 18761 15436 18883 15476
rect 18932 15436 18941 15476
rect 19075 15436 19084 15476
rect 19124 15436 19363 15476
rect 19403 15436 19412 15476
rect 19555 15436 19564 15476
rect 19604 15436 19613 15476
rect 19660 15436 19756 15476
rect 19796 15436 19805 15476
rect 20035 15436 20044 15476
rect 20084 15436 20093 15476
rect 20236 15436 20332 15476
rect 20372 15436 20381 15476
rect 20428 15436 20547 15476
rect 20587 15436 20596 15476
rect 20668 15436 20756 15476
rect 20803 15436 20812 15476
rect 20852 15436 20899 15476
rect 21475 15436 21484 15476
rect 21524 15436 21706 15476
rect 21746 15436 21755 15476
rect 21955 15436 21964 15476
rect 22004 15436 22147 15476
rect 22187 15436 22196 15476
rect 22476 15436 22540 15476
rect 22580 15436 23500 15476
rect 23540 15436 23989 15476
rect 15235 15352 15244 15392
rect 15284 15352 16436 15392
rect 16483 15352 16492 15392
rect 16532 15352 16647 15392
rect 16687 15352 16696 15392
rect 17452 15352 18028 15392
rect 18068 15352 18077 15392
rect 18892 15308 18932 15436
rect 19564 15392 19604 15436
rect 20428 15392 20468 15436
rect 20716 15392 20756 15436
rect 24652 15392 24692 15520
rect 26284 15476 26324 15520
rect 28378 15511 28387 15551
rect 28436 15520 28567 15560
rect 28745 15520 28780 15560
rect 28820 15520 28876 15560
rect 28916 15520 28925 15560
rect 29059 15520 29068 15560
rect 29108 15520 29117 15560
rect 29251 15520 29260 15560
rect 29300 15520 29309 15560
rect 28427 15511 28436 15520
rect 28378 15510 28436 15511
rect 25219 15436 25228 15476
rect 25268 15436 26275 15476
rect 26315 15436 26324 15476
rect 28032 15436 28300 15476
rect 28340 15436 28349 15476
rect 28483 15436 28492 15476
rect 28532 15436 28540 15476
rect 28580 15436 28663 15476
rect 19171 15352 19180 15392
rect 19220 15352 19604 15392
rect 19939 15352 19948 15392
rect 19988 15352 20044 15392
rect 20084 15352 20119 15392
rect 20419 15352 20428 15392
rect 20468 15352 20477 15392
rect 20707 15352 20716 15392
rect 20756 15352 20765 15392
rect 21571 15352 21580 15392
rect 21620 15352 22444 15392
rect 22484 15352 22493 15392
rect 23875 15352 23884 15392
rect 23924 15352 24364 15392
rect 24404 15352 24692 15392
rect 16387 15268 16396 15308
rect 16436 15268 17251 15308
rect 17291 15268 17300 15308
rect 18211 15268 18220 15308
rect 18260 15268 18269 15308
rect 18892 15268 19276 15308
rect 19316 15268 19325 15308
rect 19555 15268 19564 15308
rect 19604 15268 19756 15308
rect 19796 15268 19805 15308
rect 20515 15268 20524 15308
rect 20564 15268 22828 15308
rect 22868 15268 22877 15308
rect 23849 15268 23980 15308
rect 24020 15268 28972 15308
rect 29012 15268 29021 15308
rect 18220 15224 18260 15268
rect 17443 15184 17452 15224
rect 17492 15184 18260 15224
rect 18508 15184 26284 15224
rect 26324 15184 26333 15224
rect 18508 15140 18548 15184
rect 15139 15100 15148 15140
rect 15188 15100 18548 15140
rect 18651 15100 18660 15140
rect 19028 15100 19037 15140
rect 20035 15100 20044 15140
rect 20084 15100 22252 15140
rect 22292 15100 22301 15140
rect 23212 15100 24116 15140
rect 26425 15100 26434 15140
rect 26802 15100 26811 15140
rect 23212 15056 23252 15100
rect 24076 15056 24116 15100
rect 14572 15016 16004 15056
rect 16291 15016 16300 15056
rect 16340 15016 19564 15056
rect 19604 15016 23252 15056
rect 23299 15016 23308 15056
rect 23348 15016 23788 15056
rect 23828 15016 24020 15056
rect 24076 15016 27148 15056
rect 27188 15016 27197 15056
rect 15964 14972 16004 15016
rect 13315 14932 13324 14972
rect 13364 14932 13612 14972
rect 13652 14932 13661 14972
rect 14825 14932 14956 14972
rect 14996 14932 15005 14972
rect 15964 14932 17443 14972
rect 17483 14932 17492 14972
rect 17801 14932 17932 14972
rect 17972 14932 17981 14972
rect 18115 14932 18124 14972
rect 18164 14932 18604 14972
rect 18644 14932 18653 14972
rect 18953 14932 19084 14972
rect 19124 14932 19133 14972
rect 19180 14932 19756 14972
rect 19796 14932 19805 14972
rect 20515 14932 20524 14972
rect 20564 14932 20812 14972
rect 20852 14932 20861 14972
rect 21833 14932 21964 14972
rect 22004 14932 22013 14972
rect 22371 14932 23500 14972
rect 23540 14932 23549 14972
rect 19180 14888 19220 14932
rect 14851 14848 14860 14888
rect 14900 14848 15427 14888
rect 15467 14848 15476 14888
rect 15619 14848 15628 14888
rect 15668 14848 16628 14888
rect 6988 14764 7315 14804
rect 7529 14764 7651 14804
rect 7700 14764 7709 14804
rect 7843 14764 7852 14804
rect 7892 14764 7901 14804
rect 8995 14764 9004 14804
rect 9044 14764 9149 14804
rect 7275 14720 7315 14764
rect 9109 14762 9149 14764
rect 9244 14764 9292 14804
rect 9332 14764 9341 14804
rect 9449 14764 9484 14804
rect 9524 14764 9571 14804
rect 9611 14764 9629 14804
rect 9763 14764 9772 14804
rect 9812 14764 10060 14804
rect 10100 14764 10109 14804
rect 10531 14764 10540 14804
rect 10603 14764 10711 14804
rect 10876 14764 10964 14804
rect 11107 14764 11116 14804
rect 11156 14764 11287 14804
rect 11779 14764 11788 14804
rect 11828 14764 11837 14804
rect 11971 14764 11980 14804
rect 12020 14764 12029 14804
rect 12617 14764 12652 14804
rect 12692 14764 12748 14804
rect 12788 14764 12797 14804
rect 13036 14764 13172 14804
rect 9109 14753 9188 14762
rect 9109 14722 9148 14753
rect 6499 14680 6508 14720
rect 6548 14680 6557 14720
rect 6691 14680 6700 14720
rect 6740 14680 6973 14720
rect 7013 14680 7028 14720
rect 7075 14680 7084 14720
rect 7124 14680 7133 14720
rect 7275 14680 7511 14720
rect 7551 14680 7560 14720
rect 7747 14680 7756 14720
rect 7796 14680 7805 14720
rect 8023 14680 8032 14720
rect 8072 14680 8620 14720
rect 8660 14680 8669 14720
rect 8777 14680 8854 14720
rect 8894 14680 8908 14720
rect 8948 14680 9065 14720
rect 9244 14720 9284 14764
rect 10924 14762 10964 14764
rect 10924 14722 10952 14762
rect 10992 14722 11001 14762
rect 11980 14720 12020 14764
rect 13132 14720 13172 14764
rect 13900 14764 13996 14804
rect 14036 14764 14045 14804
rect 14554 14764 14563 14804
rect 14603 14764 14764 14804
rect 14804 14764 14813 14804
rect 15043 14764 15052 14804
rect 15092 14764 15572 14804
rect 13900 14720 13940 14764
rect 15532 14762 15572 14764
rect 15532 14753 15752 14762
rect 15532 14722 15712 14753
rect 9148 14704 9188 14713
rect 9235 14680 9244 14720
rect 9284 14680 9293 14720
rect 9439 14680 9448 14720
rect 9488 14680 9497 14720
rect 9667 14680 9676 14720
rect 9716 14680 9847 14720
rect 9955 14680 9964 14720
rect 10004 14680 10013 14720
rect 10147 14680 10156 14720
rect 10196 14680 10327 14720
rect 10435 14680 10444 14720
rect 10484 14680 10493 14720
rect 10652 14680 10661 14720
rect 10701 14680 10723 14720
rect 10788 14680 10797 14720
rect 10837 14680 10868 14720
rect 11443 14680 11452 14720
rect 11492 14680 11501 14720
rect 11578 14680 11587 14720
rect 11627 14680 11636 14720
rect 11683 14680 11692 14720
rect 11732 14680 11863 14720
rect 11971 14680 11980 14720
rect 12020 14680 12067 14720
rect 12163 14680 12172 14720
rect 12212 14680 12343 14720
rect 12756 14680 12844 14720
rect 12884 14680 12887 14720
rect 12927 14680 12936 14720
rect 13018 14711 13076 14720
rect 6508 14636 6548 14680
rect 6988 14636 7028 14680
rect 7084 14636 7124 14680
rect 7756 14636 7796 14680
rect 9025 14636 9065 14680
rect 9453 14636 9493 14680
rect 9964 14636 10004 14680
rect 6508 14596 6604 14636
rect 6644 14596 6653 14636
rect 6979 14596 6988 14636
rect 7028 14596 7037 14636
rect 7084 14596 7564 14636
rect 7604 14596 7613 14636
rect 7756 14596 8852 14636
rect 9025 14596 9580 14636
rect 9620 14596 9629 14636
rect 9763 14596 9772 14636
rect 9812 14596 10004 14636
rect 6389 14512 6787 14552
rect 6827 14512 6836 14552
rect 8179 14512 8188 14552
rect 8228 14512 8236 14552
rect 8276 14512 8359 14552
rect 8537 14512 8620 14552
rect 8699 14512 8717 14552
rect 8812 14468 8852 14596
rect 10444 14552 10484 14680
rect 10657 14636 10697 14680
rect 10627 14596 10636 14636
rect 10676 14596 10697 14636
rect 10828 14636 10868 14680
rect 11242 14638 11251 14678
rect 11291 14638 11306 14678
rect 10828 14596 11116 14636
rect 11156 14596 11165 14636
rect 9091 14512 9100 14552
rect 9140 14512 10348 14552
rect 10388 14512 10397 14552
rect 10444 14512 11020 14552
rect 11060 14512 11069 14552
rect 11266 14468 11306 14638
rect 11452 14636 11492 14680
rect 11596 14636 11636 14680
rect 13018 14671 13027 14711
rect 13067 14671 13076 14711
rect 13123 14680 13132 14720
rect 13172 14680 13315 14720
rect 13355 14680 13364 14720
rect 13411 14680 13420 14720
rect 13460 14680 13612 14720
rect 13652 14680 13661 14720
rect 13891 14680 13900 14720
rect 13940 14680 13949 14720
rect 14001 14680 14019 14720
rect 14059 14680 14068 14720
rect 14128 14680 14137 14720
rect 14177 14680 14188 14720
rect 14228 14680 14317 14720
rect 14362 14711 14420 14720
rect 13018 14670 13076 14671
rect 13036 14636 13076 14670
rect 13420 14636 13460 14680
rect 14001 14636 14041 14680
rect 14362 14671 14371 14711
rect 14411 14671 14420 14711
rect 14563 14680 14572 14720
rect 14612 14680 14668 14720
rect 14708 14680 14743 14720
rect 14947 14680 14956 14720
rect 14996 14680 15005 14720
rect 15139 14680 15148 14720
rect 15188 14680 15319 14720
rect 16396 14720 16436 14729
rect 16588 14720 16628 14848
rect 18124 14848 19220 14888
rect 19337 14848 19468 14888
rect 19508 14848 19517 14888
rect 19939 14848 19948 14888
rect 19988 14848 20812 14888
rect 20852 14848 20861 14888
rect 20995 14848 21004 14888
rect 21044 14848 21974 14888
rect 16675 14764 16684 14804
rect 16724 14764 16733 14804
rect 16684 14720 16724 14764
rect 18124 14720 18164 14848
rect 18307 14764 18316 14804
rect 18356 14764 18812 14804
rect 19747 14764 19756 14804
rect 19796 14764 19805 14804
rect 20236 14764 21044 14804
rect 21091 14764 21100 14804
rect 21140 14764 21332 14804
rect 18772 14762 18812 14764
rect 18772 14753 18836 14762
rect 18772 14722 18787 14753
rect 15712 14704 15752 14713
rect 15802 14680 15811 14720
rect 15851 14680 15860 14720
rect 15977 14680 16097 14720
rect 16148 14680 16157 14720
rect 16265 14680 16396 14720
rect 16436 14680 16445 14720
rect 16579 14680 16588 14720
rect 16628 14680 16637 14720
rect 16684 14680 16780 14720
rect 16820 14680 16829 14720
rect 17129 14680 17260 14720
rect 17300 14680 17309 14720
rect 17434 14680 17443 14720
rect 17492 14680 17623 14720
rect 17923 14680 17932 14720
rect 17972 14680 17981 14720
rect 18115 14680 18124 14720
rect 18164 14680 18173 14720
rect 18403 14680 18412 14720
rect 18452 14680 18461 14720
rect 18516 14680 18604 14720
rect 18644 14680 18647 14720
rect 18687 14680 18696 14720
rect 18778 14713 18787 14722
rect 18827 14713 18836 14753
rect 19756 14720 19796 14764
rect 20236 14720 20276 14764
rect 21004 14720 21044 14764
rect 21292 14762 21332 14764
rect 21433 14764 21580 14804
rect 21620 14764 21629 14804
rect 21292 14753 21380 14762
rect 21292 14722 21340 14753
rect 18778 14712 18836 14713
rect 18878 14680 18887 14720
rect 18927 14680 19028 14720
rect 19075 14680 19084 14720
rect 19124 14680 19220 14720
rect 19267 14680 19276 14720
rect 19316 14680 19796 14720
rect 20218 14680 20227 14720
rect 20267 14680 20276 14720
rect 20404 14680 20524 14720
rect 20575 14680 20584 14720
rect 20707 14680 20716 14720
rect 20756 14680 20765 14720
rect 20842 14680 20851 14720
rect 20891 14680 20900 14720
rect 20956 14680 20965 14720
rect 21005 14680 21174 14720
rect 21433 14720 21473 14764
rect 21934 14720 21974 14848
rect 22371 14804 22411 14932
rect 23980 14888 24020 15016
rect 29068 14972 29108 15520
rect 24067 14932 24076 14972
rect 24116 14932 25900 14972
rect 25940 14932 25949 14972
rect 26476 14932 27092 14972
rect 28003 14932 28012 14972
rect 28052 14932 28396 14972
rect 28436 14932 28445 14972
rect 28963 14932 28972 14972
rect 29012 14932 29108 14972
rect 23020 14848 23583 14888
rect 23971 14848 23980 14888
rect 24020 14848 24029 14888
rect 23020 14804 23060 14848
rect 22362 14764 22371 14804
rect 22411 14764 22420 14804
rect 22531 14764 22540 14804
rect 22580 14764 22724 14804
rect 22444 14720 22509 14723
rect 22684 14720 22724 14764
rect 21340 14704 21380 14713
rect 21427 14680 21436 14720
rect 21476 14680 21485 14720
rect 21545 14680 21676 14720
rect 21716 14680 21725 14720
rect 21807 14680 21816 14720
rect 21856 14680 21872 14720
rect 21916 14680 21925 14720
rect 21965 14680 21974 14720
rect 22121 14680 22252 14720
rect 22292 14680 22301 14720
rect 22433 14680 22444 14720
rect 22509 14680 22609 14720
rect 22666 14680 22675 14720
rect 22715 14680 22724 14720
rect 22780 14764 23020 14804
rect 23060 14764 23069 14804
rect 23145 14764 23154 14804
rect 23194 14764 23203 14804
rect 23260 14764 23308 14804
rect 23348 14764 23357 14804
rect 14362 14670 14420 14671
rect 14380 14636 14420 14670
rect 14956 14636 14996 14680
rect 15820 14636 15860 14680
rect 16396 14671 16436 14680
rect 17932 14636 17972 14680
rect 18412 14636 18452 14680
rect 18988 14636 19028 14680
rect 19180 14636 19220 14680
rect 11452 14596 11500 14636
rect 11540 14596 11549 14636
rect 11596 14596 12076 14636
rect 12116 14596 12125 14636
rect 12451 14596 12460 14636
rect 12500 14596 12980 14636
rect 13036 14596 13460 14636
rect 13516 14596 13623 14636
rect 13663 14596 13942 14636
rect 14001 14596 14284 14636
rect 14324 14596 14333 14636
rect 14380 14596 14764 14636
rect 14804 14596 14996 14636
rect 15427 14596 15436 14636
rect 15476 14596 15860 14636
rect 17260 14596 18220 14636
rect 18260 14596 18269 14636
rect 18412 14596 18892 14636
rect 18932 14596 18941 14636
rect 18988 14596 19084 14636
rect 19124 14596 19133 14636
rect 19180 14596 19468 14636
rect 19508 14596 19517 14636
rect 19843 14596 19852 14636
rect 19892 14596 20332 14636
rect 20372 14596 20381 14636
rect 12940 14552 12980 14596
rect 13516 14552 13556 14596
rect 13902 14552 13942 14596
rect 17260 14552 17300 14596
rect 20716 14552 20756 14680
rect 20860 14636 20900 14680
rect 21004 14636 21044 14680
rect 21676 14636 21716 14680
rect 20860 14596 20908 14636
rect 20948 14596 20957 14636
rect 21004 14596 21332 14636
rect 21571 14596 21580 14636
rect 21620 14596 21716 14636
rect 21292 14552 21332 14596
rect 11587 14512 11596 14552
rect 11636 14512 12412 14552
rect 12452 14512 12748 14552
rect 12788 14512 12797 14552
rect 12940 14512 13556 14552
rect 13673 14512 13804 14552
rect 13844 14512 13853 14552
rect 13902 14512 15244 14552
rect 15284 14512 15293 14552
rect 15946 14512 15955 14552
rect 15995 14512 16195 14552
rect 16235 14512 16244 14552
rect 16291 14512 16300 14552
rect 16340 14512 16471 14552
rect 16553 14512 16684 14552
rect 16724 14512 16733 14552
rect 17251 14512 17260 14552
rect 17300 14512 17309 14552
rect 17635 14512 17644 14552
rect 17684 14512 18268 14552
rect 18308 14512 18644 14552
rect 18787 14512 18796 14552
rect 18836 14512 19852 14552
rect 19892 14512 19901 14552
rect 20131 14512 20140 14552
rect 20180 14512 20189 14552
rect 20707 14512 20716 14552
rect 20756 14512 20765 14552
rect 21065 14512 21187 14552
rect 21236 14512 21245 14552
rect 21292 14512 21676 14552
rect 21716 14512 21725 14552
rect 748 14428 1420 14468
rect 1460 14428 4340 14468
rect 4771 14428 4780 14468
rect 4820 14428 6517 14468
rect 0 14384 400 14404
rect 0 14344 596 14384
rect 0 14324 400 14344
rect 556 14132 596 14344
rect 748 14216 788 14428
rect 6477 14384 6517 14428
rect 7084 14428 8756 14468
rect 8812 14428 10495 14468
rect 11266 14428 14860 14468
rect 14900 14428 14909 14468
rect 7084 14384 7124 14428
rect 4343 14344 4352 14384
rect 4720 14344 4729 14384
rect 6477 14344 7124 14384
rect 8716 14384 8756 14428
rect 8716 14344 9100 14384
rect 9140 14344 9149 14384
rect 3235 14260 3244 14300
rect 3284 14260 3916 14300
rect 3956 14260 3965 14300
rect 4195 14260 4204 14300
rect 4244 14260 4253 14300
rect 4867 14260 4876 14300
rect 4916 14260 5492 14300
rect 4204 14216 4244 14260
rect 730 14176 739 14216
rect 779 14176 788 14216
rect 1097 14176 1228 14216
rect 1268 14176 1277 14216
rect 3043 14176 3052 14216
rect 3092 14176 3101 14216
rect 3715 14176 3724 14216
rect 3764 14176 3773 14216
rect 4186 14176 4195 14216
rect 4235 14176 4291 14216
rect 4841 14176 4972 14216
rect 5012 14176 5021 14216
rect 3052 14132 3092 14176
rect 3724 14132 3764 14176
rect 556 14092 1612 14132
rect 1652 14092 1661 14132
rect 3052 14092 3572 14132
rect 3724 14092 4052 14132
rect 3532 14048 3572 14092
rect 547 14008 556 14048
rect 596 14008 844 14048
rect 884 14008 893 14048
rect 1027 14008 1036 14048
rect 1076 14008 1900 14048
rect 1940 14008 1949 14048
rect 2563 14008 2572 14048
rect 2612 14008 2753 14048
rect 2793 14008 2802 14048
rect 2851 14008 2860 14048
rect 2900 14008 2956 14048
rect 2996 14008 3031 14048
rect 3113 14008 3244 14048
rect 3284 14008 3293 14048
rect 3523 14008 3532 14048
rect 3572 14008 3581 14048
rect 4012 14037 4052 14092
rect 4354 14123 5108 14132
rect 4354 14092 5059 14123
rect 4354 14048 4394 14092
rect 5020 14083 5059 14092
rect 5099 14083 5108 14123
rect 5020 14082 5108 14083
rect 5164 14092 5356 14132
rect 5396 14092 5405 14132
rect 0 13964 400 13984
rect 0 13924 940 13964
rect 980 13924 989 13964
rect 0 13904 400 13924
rect 1027 13840 1036 13880
rect 1076 13840 2036 13880
rect 2083 13840 2092 13880
rect 2132 13840 2263 13880
rect 1996 13796 2036 13840
rect 1996 13756 3148 13796
rect 3188 13756 3436 13796
rect 3476 13756 3485 13796
rect 3103 13588 3112 13628
rect 3480 13588 3489 13628
rect 0 13544 400 13564
rect 0 13504 844 13544
rect 884 13504 893 13544
rect 0 13484 400 13504
rect 2441 13420 2563 13460
rect 2612 13420 2621 13460
rect 2572 13292 2612 13420
rect 2572 13252 3284 13292
rect 3244 13208 3284 13252
rect 3532 13208 3572 14008
rect 4012 13997 4028 14037
rect 4068 13997 4077 14037
rect 4218 14008 4227 14048
rect 4267 14008 4276 14048
rect 4330 14008 4339 14048
rect 4379 14008 4394 14048
rect 4474 14008 4483 14048
rect 4523 14008 4532 14048
rect 4596 14008 4605 14048
rect 4645 14008 4684 14048
rect 4724 14008 4771 14048
rect 4811 14008 4820 14048
rect 4876 14039 4916 14048
rect 4227 13964 4267 14008
rect 4227 13924 4300 13964
rect 4340 13924 4349 13964
rect 4492 13880 4532 14008
rect 4876 13964 4916 13999
rect 5020 13964 5060 14082
rect 5164 14048 5204 14092
rect 5452 14048 5492 14260
rect 5836 14260 6356 14300
rect 5836 14216 5876 14260
rect 6316 14216 6356 14260
rect 7180 14260 7468 14300
rect 7508 14260 7517 14300
rect 7878 14260 10348 14300
rect 10388 14260 10397 14300
rect 7180 14216 7220 14260
rect 5818 14176 5827 14216
rect 5867 14176 5876 14216
rect 6115 14176 6124 14216
rect 6164 14176 6260 14216
rect 6316 14176 6508 14216
rect 6548 14176 6557 14216
rect 7171 14176 7180 14216
rect 7220 14176 7229 14216
rect 7275 14176 7372 14216
rect 7412 14176 7421 14216
rect 6220 14132 6260 14176
rect 7275 14132 7315 14176
rect 7878 14132 7918 14260
rect 10455 14216 10495 14428
rect 12117 14344 12126 14384
rect 12494 14344 12503 14384
rect 18604 14300 18644 14512
rect 20140 14468 20180 14512
rect 21832 14468 21872 14680
rect 21934 14636 21974 14680
rect 21934 14596 21964 14636
rect 22004 14596 22021 14636
rect 22780 14552 22820 14764
rect 22915 14680 22924 14720
rect 22964 14680 23095 14720
rect 23154 14636 23194 14764
rect 23260 14720 23300 14764
rect 23543 14753 23583 14848
rect 23645 14764 23692 14804
rect 23732 14764 23741 14804
rect 23254 14680 23263 14720
rect 23303 14680 23312 14720
rect 23692 14720 23732 14764
rect 24141 14720 24181 14729
rect 24652 14720 24692 14932
rect 26476 14804 26516 14932
rect 27052 14888 27092 14932
rect 26947 14848 26956 14888
rect 26996 14848 27005 14888
rect 27052 14848 28876 14888
rect 28916 14848 28925 14888
rect 29705 14848 29836 14888
rect 29876 14848 29885 14888
rect 26304 14764 26516 14804
rect 26563 14764 26572 14804
rect 26612 14764 26621 14804
rect 26572 14720 26612 14764
rect 23543 14704 23583 14713
rect 23644 14711 23732 14720
rect 23644 14671 23683 14711
rect 23723 14671 23732 14711
rect 23779 14680 23788 14720
rect 23828 14680 23884 14720
rect 23924 14680 24141 14720
rect 24248 14680 24257 14720
rect 24297 14680 24306 14720
rect 24360 14680 24369 14720
rect 24409 14680 24692 14720
rect 25018 14680 25027 14720
rect 25067 14680 25076 14720
rect 25123 14680 25132 14720
rect 25172 14680 26612 14720
rect 26956 14720 26996 14848
rect 27139 14764 27148 14804
rect 27188 14764 28196 14804
rect 28156 14720 28196 14764
rect 26956 14680 27340 14720
rect 27380 14680 27389 14720
rect 28138 14680 28147 14720
rect 28187 14680 28684 14720
rect 28724 14680 28733 14720
rect 29513 14680 29644 14720
rect 29684 14680 29693 14720
rect 24141 14671 24181 14680
rect 23644 14670 23732 14671
rect 23644 14636 23684 14670
rect 23154 14596 23684 14636
rect 24266 14552 24306 14680
rect 25036 14636 25076 14680
rect 24521 14596 24643 14636
rect 24692 14596 24701 14636
rect 25036 14596 27820 14636
rect 27860 14596 28348 14636
rect 28388 14596 28397 14636
rect 22025 14512 22060 14552
rect 22100 14512 22156 14552
rect 22196 14512 22205 14552
rect 22339 14512 22348 14552
rect 22388 14512 22780 14552
rect 22820 14512 22829 14552
rect 23011 14512 23020 14552
rect 23060 14512 23116 14552
rect 23156 14512 23191 14552
rect 24266 14512 25516 14552
rect 25556 14512 25565 14552
rect 24266 14468 24306 14512
rect 20140 14428 21388 14468
rect 21428 14428 21437 14468
rect 21832 14428 22540 14468
rect 22580 14428 22589 14468
rect 23299 14428 23308 14468
rect 23348 14428 24306 14468
rect 19891 14344 19900 14384
rect 20268 14344 20277 14384
rect 23587 14344 23596 14384
rect 23636 14344 24884 14384
rect 27665 14344 27674 14384
rect 28042 14344 28051 14384
rect 10627 14260 10636 14300
rect 10676 14260 10685 14300
rect 12695 14260 12748 14300
rect 12788 14260 15942 14300
rect 18604 14260 20180 14300
rect 10636 14216 10676 14260
rect 8026 14176 8035 14216
rect 8075 14176 9236 14216
rect 9322 14176 9331 14216
rect 9371 14176 9388 14216
rect 9428 14176 9511 14216
rect 9667 14176 9676 14216
rect 9716 14176 9763 14216
rect 9803 14176 9847 14216
rect 10455 14176 10540 14216
rect 10580 14176 10589 14216
rect 10636 14176 10868 14216
rect 5635 14092 5644 14132
rect 5684 14092 6068 14132
rect 6115 14092 6124 14132
rect 6164 14092 6173 14132
rect 6220 14092 6548 14132
rect 6028 14048 6068 14092
rect 6124 14048 6164 14092
rect 6508 14048 6548 14092
rect 6892 14092 7315 14132
rect 7397 14092 7918 14132
rect 6892 14048 6932 14092
rect 7397 14048 7437 14092
rect 9196 14048 9236 14176
rect 9571 14092 9580 14132
rect 9620 14092 10004 14132
rect 10147 14092 10156 14132
rect 10196 14092 10263 14132
rect 10303 14092 10327 14132
rect 10627 14092 10636 14132
rect 10676 14092 10685 14132
rect 9964 14048 10004 14092
rect 10636 14048 10676 14092
rect 10828 14048 10868 14176
rect 12556 14176 12595 14216
rect 12635 14176 12644 14216
rect 12556 14132 12596 14176
rect 11299 14092 11308 14132
rect 11348 14092 11540 14132
rect 12499 14092 12508 14132
rect 12548 14092 12596 14132
rect 11500 14048 11540 14092
rect 12855 14048 12895 14260
rect 13978 14176 13987 14216
rect 14027 14176 14380 14216
rect 14420 14176 14429 14216
rect 14659 14176 14668 14216
rect 14708 14176 15235 14216
rect 15275 14176 15284 14216
rect 15902 14132 15942 14260
rect 20140 14216 20180 14260
rect 20236 14260 22004 14300
rect 15994 14176 16003 14216
rect 16043 14176 16300 14216
rect 16340 14176 16349 14216
rect 16570 14176 16579 14216
rect 16619 14176 16628 14216
rect 18883 14176 18892 14216
rect 18932 14176 19124 14216
rect 19171 14176 19180 14216
rect 19220 14176 19372 14216
rect 19412 14176 19421 14216
rect 20131 14176 20140 14216
rect 20180 14176 20189 14216
rect 13324 14092 13516 14132
rect 13556 14092 13565 14132
rect 13660 14092 13708 14132
rect 13748 14092 13757 14132
rect 14188 14092 14764 14132
rect 14804 14092 14813 14132
rect 15235 14092 15244 14132
rect 15284 14092 15572 14132
rect 15893 14092 15902 14132
rect 15942 14092 15951 14132
rect 16003 14092 16012 14132
rect 16052 14092 16061 14132
rect 13324 14048 13364 14092
rect 5146 14008 5155 14048
rect 5195 14008 5204 14048
rect 5323 14008 5332 14048
rect 5372 14008 5396 14048
rect 5452 14008 5495 14048
rect 5535 14008 5544 14048
rect 5731 14008 5740 14048
rect 5780 14008 5911 14048
rect 6019 14008 6028 14048
rect 6068 14008 6077 14048
rect 6124 14008 6220 14048
rect 6260 14008 6269 14048
rect 6370 14008 6379 14048
rect 6419 14008 6430 14048
rect 6490 14008 6499 14048
rect 6539 14008 6548 14048
rect 6595 14008 6604 14048
rect 6644 14008 6775 14048
rect 6883 14008 6892 14048
rect 6932 14008 6941 14048
rect 7132 14008 7141 14048
rect 7181 14008 7437 14048
rect 7507 14039 7573 14048
rect 5356 13964 5396 14008
rect 4867 13924 4876 13964
rect 4916 13924 4963 13964
rect 5020 13924 5117 13964
rect 5356 13924 5635 13964
rect 5675 13924 5836 13964
rect 5876 13924 5885 13964
rect 4195 13840 4204 13880
rect 4244 13840 4532 13880
rect 5077 13880 5117 13924
rect 6390 13880 6430 14008
rect 7507 14006 7533 14039
rect 6988 13966 7014 14006
rect 7054 13966 7063 14006
rect 7489 13999 7533 14006
rect 7489 13990 7573 13999
rect 7642 14039 7700 14048
rect 7642 13999 7651 14039
rect 7691 13999 7700 14039
rect 7747 14008 7756 14048
rect 7800 14008 7927 14048
rect 8035 14008 8044 14048
rect 8084 14008 8188 14048
rect 8228 14008 8237 14048
rect 8323 14008 8332 14048
rect 8372 14008 8503 14048
rect 9088 14039 9128 14048
rect 7642 13998 7700 13999
rect 9178 14008 9187 14048
rect 9227 14008 9236 14048
rect 9283 14008 9292 14048
rect 9332 14008 9431 14048
rect 9471 14008 9480 14048
rect 9667 14008 9676 14048
rect 9716 14008 9725 14048
rect 9946 14008 9955 14048
rect 9995 14008 10004 14048
rect 10051 14008 10060 14048
rect 10100 14008 10231 14048
rect 10435 14008 10444 14048
rect 10484 14008 10493 14048
rect 10589 14008 10634 14048
rect 10674 14008 10683 14048
rect 10810 14039 10868 14048
rect 7489 13966 7547 13990
rect 6988 13964 7028 13966
rect 7489 13964 7529 13966
rect 6691 13924 6700 13964
rect 6740 13924 7028 13964
rect 7171 13924 7180 13964
rect 7220 13924 7529 13964
rect 7656 13880 7696 13998
rect 9088 13880 9128 13999
rect 9676 13964 9716 14008
rect 9449 13924 9571 13964
rect 9620 13924 9629 13964
rect 9676 13924 10252 13964
rect 10292 13924 10301 13964
rect 10444 13880 10484 14008
rect 10810 13999 10819 14039
rect 10859 13999 10868 14039
rect 10963 14008 10972 14048
rect 11012 14008 11404 14048
rect 11444 14008 11453 14048
rect 11500 14008 11519 14048
rect 11559 14008 11568 14048
rect 11683 14008 11692 14048
rect 11732 14008 11741 14048
rect 11875 14008 11884 14048
rect 11924 14008 12055 14048
rect 12137 14008 12268 14048
rect 12308 14008 12317 14048
rect 12617 14008 12739 14048
rect 12788 14008 12797 14048
rect 12844 14039 12895 14048
rect 10810 13998 10868 13999
rect 11692 13964 11732 14008
rect 12884 14008 12895 14039
rect 13315 14008 13324 14048
rect 13364 14008 13373 14048
rect 13498 14008 13507 14048
rect 13547 14008 13556 14048
rect 12844 13990 12884 13999
rect 13516 13964 13556 14008
rect 13660 14006 13700 14092
rect 14188 14048 14228 14092
rect 15532 14048 15572 14092
rect 16012 14048 16052 14092
rect 16588 14048 16628 14176
rect 19084 14132 19124 14176
rect 20236 14132 20276 14260
rect 21964 14216 22004 14260
rect 23020 14260 23212 14300
rect 23252 14260 24788 14300
rect 23020 14216 23060 14260
rect 24748 14216 24788 14260
rect 20611 14176 20620 14216
rect 20660 14176 21716 14216
rect 21946 14176 21955 14216
rect 21995 14176 22004 14216
rect 22243 14176 22252 14216
rect 22292 14176 23060 14216
rect 23875 14176 23884 14216
rect 23924 14176 23933 14216
rect 24041 14176 24163 14216
rect 24212 14176 24221 14216
rect 24739 14176 24748 14216
rect 24788 14176 24797 14216
rect 16876 14092 18700 14132
rect 18740 14092 18749 14132
rect 19084 14092 19627 14132
rect 16876 14048 16916 14092
rect 13884 14008 13893 14048
rect 13933 14008 13996 14048
rect 14036 14008 14073 14048
rect 14170 14039 14228 14048
rect 13651 13966 13660 14006
rect 13700 13966 13709 14006
rect 14170 13999 14179 14039
rect 14219 13999 14228 14039
rect 14345 14008 14476 14048
rect 14516 14008 14525 14048
rect 14572 14008 14903 14048
rect 14943 14008 14952 14048
rect 15139 14008 15148 14048
rect 15188 14008 15476 14048
rect 15523 14008 15532 14048
rect 15572 14008 15581 14048
rect 15760 14008 15769 14048
rect 15809 14008 16052 14048
rect 16099 14008 16108 14048
rect 16148 14008 16157 14048
rect 16204 14039 16396 14048
rect 14170 13998 14228 13999
rect 11692 13924 12460 13964
rect 12500 13924 12509 13964
rect 13315 13924 13324 13964
rect 13364 13924 13556 13964
rect 13786 13924 13795 13964
rect 13835 13924 13844 13964
rect 13804 13880 13844 13924
rect 14188 13880 14228 13998
rect 14572 13964 14612 14008
rect 15436 13964 15476 14008
rect 14563 13924 14572 13964
rect 14612 13924 14621 13964
rect 14921 13924 15043 13964
rect 15092 13924 15101 13964
rect 15427 13924 15436 13964
rect 15476 13924 15485 13964
rect 15619 13924 15628 13964
rect 15691 13924 15828 13964
rect 15651 13880 15691 13924
rect 16113 13880 16153 14008
rect 16244 14008 16396 14039
rect 16436 14008 16628 14048
rect 16867 14008 16876 14048
rect 16916 14008 16925 14048
rect 17513 14008 17644 14048
rect 17684 14008 17693 14048
rect 18137 14008 18220 14048
rect 18260 14008 18268 14048
rect 18308 14008 18317 14048
rect 18403 14008 18412 14048
rect 18452 14008 18569 14048
rect 18609 14008 18618 14048
rect 18665 14008 18739 14048
rect 18779 14008 18796 14048
rect 18836 14008 18845 14048
rect 18891 14008 18988 14048
rect 19028 14008 19037 14048
rect 19216 14008 19225 14048
rect 19265 14008 19292 14048
rect 16204 13990 16244 13999
rect 18891 13964 18931 14008
rect 16771 13924 16780 13964
rect 16826 13924 16951 13964
rect 17545 13924 17554 13964
rect 17594 13924 17740 13964
rect 17780 13924 17789 13964
rect 18403 13924 18412 13964
rect 18452 13924 18461 13964
rect 18508 13924 18931 13964
rect 19098 13924 19107 13964
rect 19147 13924 19156 13964
rect 5077 13840 6508 13880
rect 6548 13840 6557 13880
rect 7459 13840 7468 13880
rect 7508 13840 8948 13880
rect 9088 13840 10156 13880
rect 10196 13840 10205 13880
rect 10444 13840 11404 13880
rect 11444 13840 11453 13880
rect 12931 13840 12940 13880
rect 12980 13840 13132 13880
rect 13172 13840 13181 13880
rect 13498 13840 13507 13880
rect 13547 13840 13844 13880
rect 13900 13840 14228 13880
rect 14275 13840 14284 13880
rect 14324 13840 14420 13880
rect 14467 13840 14476 13880
rect 14516 13840 15691 13880
rect 15953 13840 16012 13880
rect 16052 13840 17644 13880
rect 17684 13840 17693 13880
rect 8908 13796 8948 13840
rect 13900 13796 13940 13840
rect 14380 13796 14420 13840
rect 5827 13756 5836 13796
rect 5876 13756 6220 13796
rect 6260 13756 8140 13796
rect 8180 13756 8189 13796
rect 8515 13756 8524 13796
rect 8564 13756 8803 13796
rect 8843 13756 8852 13796
rect 8908 13756 9772 13796
rect 9812 13756 9821 13796
rect 10121 13756 10252 13796
rect 10292 13756 10540 13796
rect 10580 13756 10589 13796
rect 10819 13756 10828 13796
rect 10868 13756 10877 13796
rect 12355 13756 12364 13796
rect 12404 13756 12508 13796
rect 12548 13756 12557 13796
rect 13507 13756 13516 13796
rect 13556 13756 13940 13796
rect 14266 13756 14275 13796
rect 14315 13756 14324 13796
rect 14380 13756 17452 13796
rect 17492 13756 17501 13796
rect 10828 13712 10868 13756
rect 14284 13712 14324 13756
rect 18412 13712 18452 13924
rect 18508 13880 18548 13924
rect 18499 13840 18508 13880
rect 18548 13840 18557 13880
rect 19107 13796 19147 13924
rect 19252 13880 19292 14008
rect 19337 13966 19468 14006
rect 19508 13966 19517 14006
rect 19587 13964 19627 14092
rect 19756 14092 19948 14132
rect 19988 14092 19997 14132
rect 20140 14092 20276 14132
rect 20332 14092 20524 14132
rect 20564 14092 20573 14132
rect 21196 14092 21379 14132
rect 21419 14092 21428 14132
rect 21548 14092 21580 14132
rect 21620 14092 21629 14132
rect 19756 14048 19796 14092
rect 20140 14048 20180 14092
rect 20332 14048 20372 14092
rect 21196 14048 21236 14092
rect 21548 14048 21588 14092
rect 21676 14048 21716 14176
rect 23884 14132 23924 14176
rect 24844 14132 24884 14344
rect 25987 14176 25996 14216
rect 26036 14176 26804 14216
rect 29443 14176 29452 14216
rect 29492 14176 29644 14216
rect 29684 14176 29693 14216
rect 21859 14092 21868 14132
rect 21908 14092 22540 14132
rect 22580 14092 22589 14132
rect 23154 14092 23596 14132
rect 23636 14092 23645 14132
rect 23884 14092 24116 14132
rect 24634 14092 24643 14132
rect 24683 14092 24884 14132
rect 25315 14092 25324 14132
rect 25364 14092 25900 14132
rect 25940 14092 26612 14132
rect 19696 14008 19705 14048
rect 19745 14008 19796 14048
rect 19843 14008 19852 14048
rect 19892 14008 19901 14048
rect 19980 14008 20044 14048
rect 20084 14008 20140 14048
rect 20180 14008 20189 14048
rect 20323 14008 20332 14048
rect 20372 14008 20381 14048
rect 20506 14008 20515 14048
rect 20555 14008 20564 14048
rect 20611 14008 20620 14048
rect 20660 14008 20669 14048
rect 20803 14008 20812 14048
rect 20852 14008 20983 14048
rect 21142 14008 21151 14048
rect 21191 14008 21236 14048
rect 21302 14008 21388 14048
rect 21428 14039 21473 14048
rect 21428 14008 21433 14039
rect 19578 13924 19587 13964
rect 19627 13924 19636 13964
rect 19252 13840 19756 13880
rect 19796 13840 19805 13880
rect 18787 13756 18796 13796
rect 18836 13756 18845 13796
rect 18979 13756 18988 13796
rect 19028 13756 19147 13796
rect 18796 13712 18836 13756
rect 19852 13712 19892 14008
rect 20524 13964 20564 14008
rect 20227 13924 20236 13964
rect 20276 13924 20564 13964
rect 20620 13964 20660 14008
rect 21522 14008 21531 14048
rect 21571 14008 21588 14048
rect 21658 14039 21716 14048
rect 21433 13990 21473 13999
rect 21658 13999 21667 14039
rect 21707 13999 21716 14039
rect 21763 14008 21772 14048
rect 21812 14008 22060 14048
rect 22100 14008 22109 14048
rect 22313 14008 22444 14048
rect 22484 14008 22493 14048
rect 22627 14008 22636 14048
rect 22676 14008 22685 14048
rect 22788 14008 22797 14048
rect 22837 14008 22868 14048
rect 21658 13998 21716 13999
rect 22636 13964 22676 14008
rect 20620 13955 21196 13964
rect 20620 13924 21043 13955
rect 21034 13915 21043 13924
rect 21083 13924 21196 13955
rect 21236 13924 21245 13964
rect 22147 13924 22156 13964
rect 22196 13924 22732 13964
rect 22772 13924 22781 13964
rect 21083 13915 21092 13924
rect 21034 13914 21092 13915
rect 22828 13880 22868 14008
rect 22915 13966 22924 14006
rect 22964 13966 22973 14006
rect 21187 13840 21196 13880
rect 21236 13840 21908 13880
rect 22819 13840 22828 13880
rect 22868 13840 22877 13880
rect 20611 13756 20620 13796
rect 20660 13756 20852 13796
rect 20899 13756 20908 13796
rect 20948 13756 21196 13796
rect 21236 13756 21245 13796
rect 7459 13672 7468 13712
rect 7508 13672 9868 13712
rect 9908 13672 10156 13712
rect 10196 13672 10205 13712
rect 10252 13672 11444 13712
rect 11875 13672 11884 13712
rect 11924 13672 12884 13712
rect 13315 13672 13324 13712
rect 13364 13672 14324 13712
rect 18403 13672 18412 13712
rect 18452 13672 18461 13712
rect 18796 13672 19124 13712
rect 19171 13672 19180 13712
rect 19220 13672 19892 13712
rect 10252 13628 10292 13672
rect 11404 13628 11444 13672
rect 12844 13628 12884 13672
rect 6051 13588 6412 13628
rect 6452 13588 10292 13628
rect 10877 13588 10886 13628
rect 11254 13588 11263 13628
rect 11404 13588 12788 13628
rect 12844 13588 18452 13628
rect 18651 13588 18660 13628
rect 19028 13588 19037 13628
rect 3811 13420 3820 13460
rect 3860 13420 3869 13460
rect 5702 13420 5932 13460
rect 5972 13420 5981 13460
rect 3820 13292 3860 13420
rect 4762 13336 4771 13376
rect 4811 13336 4820 13376
rect 5059 13336 5068 13376
rect 5108 13336 5588 13376
rect 4780 13292 4820 13336
rect 5548 13292 5588 13336
rect 3820 13252 4628 13292
rect 4780 13252 5347 13292
rect 5387 13252 5396 13292
rect 5539 13252 5548 13292
rect 5588 13252 5597 13292
rect 4588 13208 4628 13252
rect 5702 13250 5742 13420
rect 5818 13252 5827 13292
rect 5876 13252 6007 13292
rect 5683 13210 5692 13250
rect 5732 13210 5742 13250
rect 643 13168 652 13208
rect 692 13168 940 13208
rect 980 13168 989 13208
rect 1795 13168 1804 13208
rect 1844 13168 2275 13208
rect 2315 13168 2324 13208
rect 2371 13168 2380 13208
rect 2420 13168 2551 13208
rect 2938 13168 2947 13208
rect 2996 13168 3127 13208
rect 3235 13168 3244 13208
rect 3284 13168 3293 13208
rect 3514 13168 3523 13208
rect 3563 13168 3572 13208
rect 3619 13168 3628 13208
rect 3668 13168 3916 13208
rect 3956 13168 3965 13208
rect 4474 13168 4483 13208
rect 4523 13168 4532 13208
rect 4579 13168 4588 13208
rect 4628 13168 4972 13208
rect 5012 13168 5021 13208
rect 5218 13168 5227 13208
rect 5267 13168 5276 13208
rect 5321 13168 5452 13208
rect 5492 13168 5501 13208
rect 0 13124 400 13144
rect 4492 13124 4532 13168
rect 5236 13124 5276 13168
rect 5702 13124 5742 13210
rect 6051 13208 6091 13588
rect 12748 13544 12788 13588
rect 6307 13504 6316 13544
rect 6356 13504 6452 13544
rect 8611 13504 8620 13544
rect 8660 13504 12706 13544
rect 12748 13504 14476 13544
rect 14516 13504 14525 13544
rect 6412 13460 6452 13504
rect 8620 13460 8660 13504
rect 11308 13460 11348 13504
rect 12666 13460 12706 13504
rect 18412 13460 18452 13588
rect 19084 13460 19124 13672
rect 20812 13628 20852 13756
rect 21868 13712 21908 13840
rect 21868 13672 22636 13712
rect 22676 13672 22685 13712
rect 19459 13588 19468 13628
rect 19508 13588 20716 13628
rect 20756 13588 20765 13628
rect 20812 13588 20908 13628
rect 20948 13588 22484 13628
rect 20323 13504 20332 13544
rect 20372 13504 20524 13544
rect 20564 13504 20573 13544
rect 6412 13420 8660 13460
rect 9130 13420 9139 13460
rect 9179 13420 11060 13460
rect 11299 13420 11308 13460
rect 11348 13420 11357 13460
rect 12346 13420 12355 13460
rect 12395 13420 12556 13460
rect 12596 13420 12605 13460
rect 12666 13420 13612 13460
rect 13652 13420 14188 13460
rect 14228 13420 14572 13460
rect 14612 13420 14621 13460
rect 15593 13420 15724 13460
rect 15764 13420 15773 13460
rect 18394 13420 18403 13460
rect 18443 13420 18452 13460
rect 19075 13420 19084 13460
rect 19124 13420 19133 13460
rect 19459 13420 19468 13460
rect 19508 13420 19639 13460
rect 19939 13420 19948 13460
rect 19988 13420 20236 13460
rect 20276 13420 20620 13460
rect 20660 13420 20669 13460
rect 20777 13420 20812 13460
rect 20852 13420 20899 13460
rect 20939 13420 20957 13460
rect 21667 13420 21676 13460
rect 21716 13420 21763 13460
rect 21803 13420 21847 13460
rect 6185 13252 6220 13292
rect 6260 13252 6307 13292
rect 6347 13252 6365 13292
rect 6412 13208 6452 13420
rect 11020 13376 11060 13420
rect 22444 13376 22484 13588
rect 22924 13460 22964 13966
rect 23154 13964 23194 14092
rect 24076 14048 24116 14092
rect 26572 14048 26612 14092
rect 26764 14048 26804 14176
rect 23395 14008 23404 14048
rect 23444 14008 23575 14048
rect 23657 14008 23743 14048
rect 23783 14008 23788 14048
rect 23828 14008 23837 14048
rect 24067 14008 24076 14048
rect 24116 14008 24125 14048
rect 24233 14008 24364 14048
rect 24404 14008 24413 14048
rect 24536 14008 24545 14048
rect 24585 14008 24748 14048
rect 24788 14008 24797 14048
rect 24844 14039 24884 14048
rect 23242 13966 23251 14006
rect 23291 13966 23348 14006
rect 23110 13924 23119 13964
rect 23159 13924 23194 13964
rect 23011 13840 23020 13880
rect 23060 13840 23069 13880
rect 23020 13628 23060 13840
rect 23308 13712 23348 13966
rect 25577 14008 25708 14048
rect 25748 14008 25757 14048
rect 26563 14008 26572 14048
rect 26612 14008 26621 14048
rect 26755 14008 26764 14048
rect 26804 14008 26813 14048
rect 26921 14008 26956 14048
rect 26996 14008 27052 14048
rect 27092 14008 27101 14048
rect 27514 14008 27523 14048
rect 27572 14008 27703 14048
rect 24844 13964 24884 13999
rect 23561 13955 23692 13964
rect 23561 13924 23635 13955
rect 23626 13915 23635 13924
rect 23675 13924 23692 13955
rect 23732 13924 23741 13964
rect 23788 13924 24884 13964
rect 26851 13924 26860 13964
rect 26900 13924 27148 13964
rect 27188 13924 27197 13964
rect 28800 13924 29836 13964
rect 29876 13924 29885 13964
rect 23675 13915 23684 13924
rect 23626 13914 23684 13915
rect 23788 13880 23828 13924
rect 23779 13840 23788 13880
rect 23828 13840 23837 13880
rect 23884 13840 26764 13880
rect 26804 13840 26813 13880
rect 28867 13840 28876 13880
rect 28916 13840 29644 13880
rect 29684 13840 29693 13880
rect 23491 13756 23500 13796
rect 23540 13756 23671 13796
rect 23884 13712 23924 13840
rect 24739 13756 24748 13796
rect 24788 13756 25036 13796
rect 25076 13756 25085 13796
rect 25315 13756 25324 13796
rect 25364 13756 25900 13796
rect 25940 13756 25949 13796
rect 28937 13756 29068 13796
rect 29108 13756 29117 13796
rect 23308 13672 23924 13712
rect 23020 13588 24172 13628
rect 24212 13588 24221 13628
rect 26425 13588 26434 13628
rect 26802 13588 26811 13628
rect 22697 13420 22828 13460
rect 22868 13420 22877 13460
rect 22924 13420 23308 13460
rect 23348 13420 23404 13460
rect 23444 13420 23453 13460
rect 23683 13420 23692 13460
rect 23732 13420 24028 13460
rect 24068 13420 24077 13460
rect 24521 13420 24652 13460
rect 24692 13420 24701 13460
rect 25708 13420 28780 13460
rect 28820 13420 28829 13460
rect 25708 13376 25748 13420
rect 7267 13336 7276 13376
rect 7316 13336 9379 13376
rect 9419 13336 9428 13376
rect 9484 13336 10964 13376
rect 11020 13336 17780 13376
rect 18115 13336 18124 13376
rect 18164 13336 18316 13376
rect 18356 13336 18365 13376
rect 18691 13336 18700 13376
rect 18740 13336 19316 13376
rect 19843 13336 19852 13376
rect 19892 13336 20044 13376
rect 20084 13336 20948 13376
rect 21065 13336 21196 13376
rect 21236 13336 21245 13376
rect 22217 13336 22348 13376
rect 22388 13336 22397 13376
rect 22444 13336 22772 13376
rect 9484 13292 9524 13336
rect 10924 13292 10964 13336
rect 6499 13252 6508 13292
rect 6548 13252 6679 13292
rect 7363 13252 7372 13292
rect 7412 13252 7852 13292
rect 7892 13252 7948 13292
rect 7988 13252 7997 13292
rect 8515 13252 8524 13292
rect 8564 13252 9524 13292
rect 9664 13252 10060 13292
rect 10100 13252 10109 13292
rect 10243 13252 10252 13292
rect 10298 13252 10423 13292
rect 10906 13252 10915 13292
rect 10955 13252 10964 13292
rect 11020 13252 11788 13292
rect 11828 13252 11837 13292
rect 12355 13252 12364 13292
rect 12404 13252 12692 13292
rect 13075 13252 13084 13292
rect 13124 13252 13228 13292
rect 13268 13252 13277 13292
rect 13324 13252 13516 13292
rect 13556 13252 13565 13292
rect 13626 13252 13635 13292
rect 13675 13252 13804 13292
rect 13844 13252 13853 13292
rect 14755 13252 14764 13292
rect 14804 13252 14996 13292
rect 15139 13252 15148 13292
rect 15188 13252 16204 13292
rect 16244 13252 16436 13292
rect 16867 13252 16876 13292
rect 16916 13252 17187 13292
rect 17227 13252 17236 13292
rect 9664 13241 9704 13252
rect 8428 13208 8468 13217
rect 5921 13168 5930 13208
rect 5970 13168 5979 13208
rect 6051 13168 6167 13208
rect 6207 13168 6216 13208
rect 6403 13168 6412 13208
rect 6452 13168 6461 13208
rect 6508 13168 6691 13208
rect 6731 13168 6740 13208
rect 6787 13168 6796 13208
rect 6836 13168 6967 13208
rect 7211 13168 7276 13208
rect 7316 13168 7342 13208
rect 7382 13168 7391 13208
rect 5932 13124 5972 13168
rect 6508 13124 6548 13168
rect 7450 13140 7459 13180
rect 7499 13140 7508 13180
rect 0 13084 1132 13124
rect 1172 13084 1181 13124
rect 3139 13084 3148 13124
rect 3188 13084 3831 13124
rect 3871 13084 3880 13124
rect 4492 13084 4780 13124
rect 4820 13084 4829 13124
rect 5236 13084 5742 13124
rect 5923 13084 5932 13124
rect 5972 13084 6017 13124
rect 6211 13084 6220 13124
rect 6260 13084 6548 13124
rect 6953 13084 7002 13124
rect 7042 13084 7084 13124
rect 7124 13084 7133 13124
rect 0 13064 400 13084
rect 7468 13040 7508 13140
rect 7564 13168 7852 13208
rect 7892 13168 7948 13208
rect 7988 13168 7997 13208
rect 8899 13168 8908 13208
rect 8956 13168 9079 13208
rect 11020 13208 11060 13252
rect 12652 13208 12692 13252
rect 13324 13208 13364 13252
rect 14956 13208 14996 13252
rect 16396 13208 16436 13252
rect 17740 13208 17780 13336
rect 17980 13252 19220 13292
rect 17980 13250 18020 13252
rect 9664 13192 9704 13201
rect 9754 13168 9763 13208
rect 9812 13168 9943 13208
rect 10342 13168 10351 13208
rect 10391 13168 10484 13208
rect 10531 13168 10540 13208
rect 10580 13168 10775 13208
rect 10815 13168 10824 13208
rect 11011 13168 11020 13208
rect 11060 13168 11069 13208
rect 11587 13168 11596 13208
rect 11636 13168 11704 13208
rect 11744 13168 11767 13208
rect 12205 13168 12214 13208
rect 12254 13168 12460 13208
rect 12500 13168 12509 13208
rect 12919 13168 12928 13208
rect 12968 13168 13364 13208
rect 13507 13168 13516 13208
rect 13556 13168 13652 13208
rect 13744 13168 13753 13208
rect 13793 13168 13844 13208
rect 14057 13168 14188 13208
rect 14228 13168 14237 13208
rect 14284 13168 14307 13208
rect 14347 13168 14371 13208
rect 14416 13168 14425 13208
rect 14465 13168 14476 13208
rect 14516 13168 14711 13208
rect 14751 13168 14760 13208
rect 14842 13168 14851 13208
rect 14891 13168 14900 13208
rect 14947 13168 14956 13208
rect 14996 13168 15005 13208
rect 15226 13168 15235 13208
rect 15275 13168 15340 13208
rect 15380 13168 15415 13208
rect 15537 13168 15546 13208
rect 15586 13168 15724 13208
rect 15764 13168 15773 13208
rect 16108 13199 16148 13208
rect 1219 13000 1228 13040
rect 1268 13000 1612 13040
rect 1652 13000 1661 13040
rect 5897 13000 6019 13040
rect 6068 13000 6077 13040
rect 6307 13000 6316 13040
rect 6356 13000 6892 13040
rect 6932 13000 6941 13040
rect 7459 13000 7468 13040
rect 7508 13000 7517 13040
rect 7564 12956 7604 13168
rect 8428 13124 8468 13168
rect 8035 13084 8044 13124
rect 8084 13084 8468 13124
rect 10444 13124 10484 13168
rect 12652 13159 12692 13168
rect 10444 13084 10828 13124
rect 10868 13084 10877 13124
rect 11098 13084 11107 13124
rect 11147 13084 11212 13124
rect 11252 13084 11287 13124
rect 11388 13084 11404 13124
rect 11444 13084 11539 13124
rect 11579 13084 12353 13124
rect 12393 13084 12556 13124
rect 12596 13084 12605 13124
rect 13315 13084 13324 13124
rect 13364 13084 13420 13124
rect 13460 13084 13495 13124
rect 13612 13040 13652 13168
rect 13804 13124 13844 13168
rect 14284 13124 14324 13168
rect 13795 13084 13804 13124
rect 13844 13084 13853 13124
rect 14275 13084 14284 13124
rect 14324 13084 14333 13124
rect 14860 13040 14900 13168
rect 16387 13168 16396 13208
rect 16436 13168 16445 13208
rect 16937 13168 17068 13208
rect 17108 13168 17117 13208
rect 17296 13168 17305 13208
rect 17345 13168 17548 13208
rect 17588 13168 17597 13208
rect 17740 13159 17780 13168
rect 17851 13241 17891 13250
rect 17945 13210 17954 13250
rect 17994 13210 18020 13250
rect 15034 13084 15043 13124
rect 15083 13084 15244 13124
rect 15284 13084 15293 13124
rect 15340 13084 15628 13124
rect 15668 13084 15677 13124
rect 15881 13084 16012 13124
rect 16052 13084 16061 13124
rect 15340 13040 15380 13084
rect 16108 13040 16148 13159
rect 17851 13124 17891 13201
rect 18787 13168 18796 13208
rect 18836 13168 18967 13208
rect 19075 13168 19084 13208
rect 19124 13168 19133 13208
rect 16963 13084 16972 13124
rect 17012 13084 17356 13124
rect 17396 13084 17405 13124
rect 17827 13084 17836 13124
rect 17876 13084 17891 13124
rect 19084 13040 19124 13168
rect 19180 13124 19220 13252
rect 19276 13208 19316 13336
rect 20908 13292 20948 13336
rect 19660 13252 19852 13292
rect 19892 13252 19901 13292
rect 20323 13252 20332 13292
rect 20372 13252 20381 13292
rect 20716 13252 20812 13292
rect 20852 13252 20861 13292
rect 20908 13252 21044 13292
rect 22531 13252 22540 13292
rect 22580 13252 22597 13292
rect 19660 13208 19700 13252
rect 20332 13208 20372 13252
rect 20716 13208 20756 13252
rect 21004 13250 21044 13252
rect 21004 13241 21130 13250
rect 21004 13210 21090 13241
rect 19267 13168 19276 13208
rect 19316 13168 19325 13208
rect 19459 13168 19468 13208
rect 19508 13168 19517 13208
rect 19651 13168 19660 13208
rect 19700 13168 19709 13208
rect 19843 13168 19852 13208
rect 19892 13168 19901 13208
rect 20035 13168 20044 13208
rect 20084 13168 20236 13208
rect 20276 13168 20372 13208
rect 20515 13168 20524 13208
rect 20564 13168 20573 13208
rect 20707 13168 20716 13208
rect 20756 13168 20765 13208
rect 20898 13168 20907 13208
rect 20947 13168 20956 13208
rect 22540 13208 22580 13252
rect 22732 13208 22772 13336
rect 22929 13336 25748 13376
rect 28609 13336 28684 13376
rect 28724 13336 28733 13376
rect 22929 13292 22969 13336
rect 22924 13252 22969 13292
rect 23299 13252 23308 13292
rect 23348 13252 23775 13292
rect 24509 13252 24556 13292
rect 24596 13252 24940 13292
rect 24980 13252 24989 13292
rect 25891 13252 25900 13292
rect 25940 13252 25987 13292
rect 26027 13252 26071 13292
rect 27744 13252 28396 13292
rect 28436 13252 28445 13292
rect 21090 13192 21130 13201
rect 21244 13181 21272 13208
rect 21196 13168 21272 13181
rect 21312 13168 21321 13208
rect 21374 13168 21388 13208
rect 21428 13168 21437 13208
rect 21548 13168 21575 13208
rect 21615 13168 21624 13208
rect 21762 13168 21771 13208
rect 21811 13168 21868 13208
rect 21908 13168 21942 13208
rect 21994 13168 22003 13208
rect 22043 13168 22076 13208
rect 22121 13168 22156 13208
rect 22196 13168 22252 13208
rect 22292 13168 22301 13208
rect 22378 13168 22387 13208
rect 22427 13168 22436 13208
rect 22492 13168 22501 13208
rect 22541 13168 22580 13208
rect 22723 13168 22732 13208
rect 22772 13168 22781 13208
rect 22924 13205 22964 13252
rect 23735 13250 23775 13252
rect 23735 13241 23780 13250
rect 23735 13210 23740 13241
rect 19468 13124 19508 13168
rect 19852 13124 19892 13168
rect 20524 13124 20564 13168
rect 19180 13084 19756 13124
rect 19796 13084 19805 13124
rect 19852 13084 20236 13124
rect 20276 13084 20716 13124
rect 20756 13084 20765 13124
rect 19852 13040 19892 13084
rect 10042 13000 10051 13040
rect 10091 13000 10444 13040
rect 10484 13000 10493 13040
rect 11779 13000 11788 13040
rect 11828 13000 12019 13040
rect 12059 13000 12068 13040
rect 12163 13000 12172 13040
rect 12212 13000 12556 13040
rect 12596 13000 12605 13040
rect 12931 13000 12940 13040
rect 12980 13000 13652 13040
rect 13699 13000 13708 13040
rect 13748 13000 14092 13040
rect 14132 13000 14188 13040
rect 14228 13000 14292 13040
rect 14860 13000 15148 13040
rect 15188 13000 15197 13040
rect 15322 13000 15331 13040
rect 15371 13000 15380 13040
rect 15427 13000 15436 13040
rect 15476 13000 16148 13040
rect 18700 13000 19892 13040
rect 9868 12958 9907 12998
rect 9947 12958 9956 12998
rect 9868 12956 9908 12958
rect 18700 12956 18740 13000
rect 20908 12956 20948 13168
rect 21196 13141 21284 13168
rect 21196 13124 21236 13141
rect 20995 13084 21004 13124
rect 21044 13084 21236 13124
rect 21374 13040 21414 13168
rect 21548 13124 21588 13168
rect 22036 13124 22076 13168
rect 22396 13124 22436 13168
rect 22908 13165 22917 13205
rect 22957 13165 22966 13205
rect 23098 13168 23107 13208
rect 23156 13168 23287 13208
rect 23465 13168 23596 13208
rect 23636 13168 23645 13208
rect 24556 13208 24596 13252
rect 28609 13250 28649 13336
rect 28733 13252 28780 13292
rect 28820 13252 28829 13292
rect 28609 13210 28627 13250
rect 28667 13210 28676 13250
rect 28780 13208 28820 13252
rect 23740 13192 23780 13201
rect 24163 13168 24172 13208
rect 24212 13168 24221 13208
rect 24355 13168 24364 13208
rect 24404 13168 24413 13208
rect 24538 13168 24547 13208
rect 24587 13168 24596 13208
rect 24643 13168 24652 13208
rect 24692 13168 24748 13208
rect 24788 13168 24823 13208
rect 25018 13168 25027 13208
rect 25067 13168 25076 13208
rect 25123 13168 25132 13208
rect 25172 13168 25324 13208
rect 25364 13168 25373 13208
rect 27139 13168 27148 13208
rect 27188 13168 27523 13208
rect 27572 13168 27581 13208
rect 28771 13168 28780 13208
rect 28820 13168 28829 13208
rect 28963 13168 28972 13208
rect 29012 13168 29143 13208
rect 24172 13124 24212 13168
rect 24364 13124 24404 13168
rect 25036 13124 25076 13168
rect 21548 13084 21580 13124
rect 21620 13084 21629 13124
rect 22036 13084 22060 13124
rect 22100 13084 22109 13124
rect 22236 13084 22252 13124
rect 22292 13084 22732 13124
rect 22772 13084 22781 13124
rect 23081 13084 23212 13124
rect 23252 13084 23261 13124
rect 23409 13084 23418 13124
rect 23458 13084 23788 13124
rect 23828 13084 23837 13124
rect 23923 13084 23932 13124
rect 23972 13084 23980 13124
rect 24020 13084 24103 13124
rect 24172 13084 24268 13124
rect 24308 13084 24317 13124
rect 24364 13084 24652 13124
rect 24692 13084 24701 13124
rect 24989 13084 25036 13124
rect 25076 13084 25085 13124
rect 25411 13084 25420 13124
rect 25460 13084 25603 13124
rect 25643 13084 25652 13124
rect 27532 13040 27572 13168
rect 27898 13084 27907 13124
rect 27947 13084 28204 13124
rect 28244 13084 28253 13124
rect 21091 13000 21100 13040
rect 21140 13000 21414 13040
rect 22099 13000 22108 13040
rect 22148 13000 23350 13040
rect 23395 13000 23404 13040
rect 23444 13000 24500 13040
rect 25411 13000 25420 13040
rect 25460 13000 25556 13040
rect 27264 13000 27340 13040
rect 27380 13000 27389 13040
rect 27532 13000 28435 13040
rect 28475 13000 28484 13040
rect 3907 12916 3916 12956
rect 3956 12916 7180 12956
rect 7220 12916 7604 12956
rect 9772 12916 9908 12956
rect 11203 12916 11212 12956
rect 11252 12916 18740 12956
rect 19459 12916 19468 12956
rect 19508 12916 19756 12956
rect 19796 12916 22732 12956
rect 22772 12916 22781 12956
rect 4343 12832 4352 12872
rect 4720 12832 4729 12872
rect 643 12748 652 12788
rect 692 12748 884 12788
rect 0 12704 400 12724
rect 844 12704 884 12748
rect 3580 12748 5108 12788
rect 5923 12748 5932 12788
rect 5972 12748 6356 12788
rect 3580 12704 3620 12748
rect 0 12664 460 12704
rect 500 12664 509 12704
rect 826 12664 835 12704
rect 875 12664 884 12704
rect 1673 12664 1804 12704
rect 1844 12664 2035 12704
rect 2075 12664 2084 12704
rect 2947 12664 2956 12704
rect 2996 12664 3043 12704
rect 3083 12664 3127 12704
rect 3532 12664 3571 12704
rect 3611 12664 3620 12704
rect 4579 12664 4588 12704
rect 4628 12664 4780 12704
rect 4820 12664 4829 12704
rect 0 12644 400 12664
rect 844 12620 884 12664
rect 3532 12620 3572 12664
rect 844 12580 1364 12620
rect 1324 12536 1364 12580
rect 2188 12580 2380 12620
rect 2420 12580 2429 12620
rect 2740 12580 3572 12620
rect 3628 12580 4492 12620
rect 4532 12580 4541 12620
rect 4876 12580 4972 12620
rect 5012 12580 5021 12620
rect 2188 12536 2228 12580
rect 2740 12536 2780 12580
rect 3628 12536 3668 12580
rect 4204 12536 4244 12580
rect 4876 12536 4916 12580
rect 5068 12536 5108 12748
rect 6316 12704 6356 12748
rect 6412 12748 6796 12788
rect 6836 12748 6845 12788
rect 7555 12748 7564 12788
rect 7604 12748 9676 12788
rect 9716 12748 9725 12788
rect 6412 12704 6452 12748
rect 5827 12664 5836 12704
rect 5876 12664 6028 12704
rect 6068 12664 6077 12704
rect 6298 12664 6307 12704
rect 6347 12664 6356 12704
rect 6403 12664 6412 12704
rect 6452 12664 6461 12704
rect 6508 12664 7084 12704
rect 7124 12664 7133 12704
rect 6508 12620 6548 12664
rect 5539 12580 5548 12620
rect 5588 12580 5780 12620
rect 5740 12536 5780 12580
rect 6209 12580 6548 12620
rect 6680 12580 6689 12620
rect 6729 12580 6796 12620
rect 6836 12580 6860 12620
rect 6979 12580 6988 12620
rect 7028 12580 7075 12620
rect 7171 12580 7180 12620
rect 7220 12580 7267 12620
rect 6209 12536 6249 12580
rect 809 12496 940 12536
rect 980 12496 989 12536
rect 1315 12496 1324 12536
rect 1364 12496 1373 12536
rect 1577 12496 1708 12536
rect 1748 12496 1757 12536
rect 2170 12496 2179 12536
rect 2219 12496 2228 12536
rect 2284 12527 2324 12536
rect 2722 12496 2731 12536
rect 2771 12496 2780 12536
rect 2947 12496 2956 12536
rect 2996 12496 3127 12536
rect 3436 12496 3668 12536
rect 3757 12496 3766 12536
rect 3806 12496 3916 12536
rect 3956 12496 3965 12536
rect 4186 12496 4195 12536
rect 4235 12496 4244 12536
rect 4291 12496 4300 12536
rect 4340 12496 4471 12536
rect 4738 12496 4747 12536
rect 4787 12496 4916 12536
rect 4963 12496 4972 12536
rect 5012 12496 5021 12536
rect 5068 12496 5164 12536
rect 5204 12496 5635 12536
rect 5675 12496 5684 12536
rect 5731 12496 5740 12536
rect 5780 12496 5789 12536
rect 6200 12496 6209 12536
rect 6249 12496 6258 12536
rect 6377 12496 6508 12536
rect 6548 12496 6557 12536
rect 6883 12496 6892 12536
rect 6932 12496 6941 12536
rect 6988 12527 7028 12580
rect 7180 12536 7220 12580
rect 7948 12536 7988 12748
rect 9772 12704 9812 12916
rect 23310 12872 23350 13000
rect 24460 12956 24500 13000
rect 25516 12956 25556 13000
rect 27340 12956 27380 13000
rect 24460 12916 25172 12956
rect 25516 12916 27380 12956
rect 27436 12916 28492 12956
rect 28532 12916 28541 12956
rect 25132 12872 25172 12916
rect 27436 12872 27476 12916
rect 12117 12832 12126 12872
rect 12494 12832 12503 12872
rect 12940 12832 13804 12872
rect 13844 12832 13853 12872
rect 16579 12832 16588 12872
rect 16628 12832 18356 12872
rect 19891 12832 19900 12872
rect 20268 12832 20277 12872
rect 23310 12832 25076 12872
rect 25132 12832 27476 12872
rect 27665 12832 27674 12872
rect 28042 12832 28051 12872
rect 12940 12788 12980 12832
rect 18316 12788 18356 12832
rect 12172 12748 12980 12788
rect 13036 12748 16108 12788
rect 16148 12748 16157 12788
rect 17059 12748 17068 12788
rect 17108 12748 18260 12788
rect 18316 12748 19988 12788
rect 21187 12748 21196 12788
rect 21236 12748 21524 12788
rect 8428 12664 9100 12704
rect 9140 12664 9149 12704
rect 9274 12664 9283 12704
rect 9323 12664 9332 12704
rect 9754 12664 9763 12704
rect 9803 12664 9812 12704
rect 9859 12664 9868 12704
rect 9908 12664 10867 12704
rect 10907 12664 10916 12704
rect 11395 12664 11404 12704
rect 11444 12664 11500 12704
rect 11540 12664 11575 12704
rect 8035 12580 8044 12620
rect 8084 12580 8129 12620
rect 8201 12580 8332 12620
rect 8372 12580 8381 12620
rect 8044 12536 8084 12580
rect 8428 12536 8468 12664
rect 9292 12620 9332 12664
rect 8585 12580 8716 12620
rect 8756 12580 8765 12620
rect 8908 12580 9004 12620
rect 9044 12580 9053 12620
rect 9292 12580 9956 12620
rect 11192 12580 11201 12620
rect 11241 12580 11404 12620
rect 11444 12580 11453 12620
rect 11945 12580 11971 12620
rect 12011 12580 12076 12620
rect 12116 12580 12125 12620
rect 8908 12536 8948 12580
rect 9916 12536 9956 12580
rect 12172 12536 12212 12748
rect 13036 12704 13076 12748
rect 12547 12664 12556 12704
rect 12596 12664 13076 12704
rect 13289 12664 13420 12704
rect 13460 12664 13469 12704
rect 13699 12664 13708 12704
rect 13748 12664 13757 12704
rect 13708 12620 13748 12664
rect 13516 12580 13748 12620
rect 13795 12580 13804 12620
rect 13844 12580 13853 12620
rect 13516 12536 13556 12580
rect 13796 12536 13836 12580
rect 13900 12536 13940 12748
rect 18220 12704 18260 12748
rect 19948 12704 19988 12748
rect 14947 12664 14956 12704
rect 14996 12664 15091 12704
rect 15131 12664 15140 12704
rect 15881 12664 16012 12704
rect 16052 12664 16061 12704
rect 16169 12664 16291 12704
rect 16340 12664 16349 12704
rect 16745 12664 16876 12704
rect 16916 12664 16925 12704
rect 17513 12664 17644 12704
rect 17684 12664 17693 12704
rect 18202 12664 18211 12704
rect 18251 12664 18260 12704
rect 19066 12664 19075 12704
rect 19115 12664 19124 12704
rect 19939 12664 19948 12704
rect 19988 12664 19997 12704
rect 20515 12664 20524 12704
rect 20564 12664 20611 12704
rect 20651 12664 20695 12704
rect 21091 12664 21100 12704
rect 21140 12664 21388 12704
rect 21428 12664 21437 12704
rect 19084 12620 19124 12664
rect 20620 12620 20660 12664
rect 21484 12620 21524 12748
rect 23779 12664 23788 12704
rect 23828 12664 24692 12704
rect 24809 12664 24940 12704
rect 24980 12664 24989 12704
rect 14170 12611 14188 12620
rect 14170 12571 14179 12611
rect 14228 12580 14359 12620
rect 15340 12580 15532 12620
rect 15572 12580 15581 12620
rect 15715 12580 15724 12620
rect 15764 12580 16190 12620
rect 16230 12580 16239 12620
rect 16387 12580 16396 12620
rect 16436 12580 17438 12620
rect 17492 12580 17638 12620
rect 17740 12580 19124 12620
rect 19564 12580 19660 12620
rect 19700 12580 19709 12620
rect 20620 12580 21140 12620
rect 21466 12580 21475 12620
rect 21515 12580 21524 12620
rect 21580 12580 22540 12620
rect 22580 12580 22589 12620
rect 14219 12571 14228 12580
rect 14170 12570 14228 12571
rect 15340 12536 15380 12580
rect 2284 12452 2324 12487
rect 1132 12412 2324 12452
rect 2842 12412 2851 12452
rect 2891 12412 3052 12452
rect 3092 12412 3101 12452
rect 1132 12368 1172 12412
rect 3436 12368 3476 12496
rect 4745 12412 4780 12452
rect 4820 12412 4867 12452
rect 4907 12412 4925 12452
rect 1123 12328 1132 12368
rect 1172 12328 1181 12368
rect 2563 12328 2572 12368
rect 2612 12328 3476 12368
rect 4972 12368 5012 12496
rect 6508 12478 6548 12487
rect 6892 12452 6932 12496
rect 7171 12496 7180 12536
rect 7220 12496 7229 12536
rect 7366 12496 7375 12536
rect 7415 12496 7468 12536
rect 7508 12496 7555 12536
rect 7843 12496 7852 12536
rect 7892 12496 7988 12536
rect 8033 12496 8042 12536
rect 8082 12496 8091 12536
rect 8140 12496 8236 12536
rect 8276 12496 8285 12536
rect 8419 12496 8428 12536
rect 8468 12496 8477 12536
rect 8600 12496 8609 12536
rect 8649 12496 8660 12536
rect 8803 12496 8812 12536
rect 8852 12496 8948 12536
rect 8995 12496 9004 12536
rect 9044 12496 9100 12536
rect 9140 12496 9175 12536
rect 9435 12496 9444 12536
rect 6988 12478 7028 12487
rect 8140 12452 8180 12496
rect 8620 12452 8660 12496
rect 9484 12452 9524 12536
rect 9571 12496 9580 12536
rect 9620 12496 9751 12536
rect 9907 12496 9916 12536
rect 9956 12496 9965 12536
rect 10051 12496 10060 12536
rect 10100 12496 10292 12536
rect 11053 12496 11062 12536
rect 11102 12496 11212 12536
rect 11252 12496 11261 12536
rect 11500 12527 11884 12536
rect 5059 12412 5068 12452
rect 5108 12412 6412 12452
rect 6452 12412 6461 12452
rect 6595 12412 6604 12452
rect 6644 12412 6932 12452
rect 7075 12412 7084 12452
rect 7124 12412 8084 12452
rect 8131 12412 8140 12452
rect 8180 12412 8189 12452
rect 8611 12412 8620 12452
rect 8660 12412 8696 12452
rect 9484 12412 10156 12452
rect 10196 12412 10205 12452
rect 8044 12368 8084 12412
rect 10252 12368 10292 12496
rect 11540 12496 11884 12527
rect 11924 12496 11933 12536
rect 11980 12496 12172 12536
rect 12212 12496 12221 12536
rect 12730 12496 12739 12536
rect 12779 12496 12788 12536
rect 12837 12496 12846 12536
rect 12886 12496 12940 12536
rect 12980 12496 13026 12536
rect 13507 12496 13516 12536
rect 13556 12496 13565 12536
rect 13744 12496 13753 12536
rect 13793 12496 13836 12536
rect 13882 12496 13891 12536
rect 13931 12496 13940 12536
rect 13996 12527 14036 12536
rect 11500 12478 11540 12487
rect 11980 12368 12020 12496
rect 12748 12452 12788 12496
rect 14266 12496 14275 12536
rect 14315 12496 14324 12536
rect 12739 12412 12748 12452
rect 12788 12412 12835 12452
rect 13642 12443 13700 12452
rect 13642 12403 13651 12443
rect 13691 12403 13700 12443
rect 13642 12402 13700 12403
rect 4972 12328 7276 12368
rect 7316 12328 7325 12368
rect 8044 12328 10348 12368
rect 10388 12328 10452 12368
rect 11020 12328 12020 12368
rect 13660 12368 13700 12402
rect 13660 12328 13804 12368
rect 13844 12328 13853 12368
rect 6682 12244 6691 12284
rect 6731 12244 6740 12284
rect 7721 12244 7852 12284
rect 7892 12244 7901 12284
rect 8035 12244 8044 12284
rect 8084 12244 9148 12284
rect 9188 12244 9196 12284
rect 9236 12244 9245 12284
rect 9667 12244 9676 12284
rect 9716 12244 10732 12284
rect 10772 12244 10781 12284
rect 6700 12116 6740 12244
rect 11020 12200 11060 12328
rect 11194 12244 11203 12284
rect 11243 12244 11252 12284
rect 13018 12244 13027 12284
rect 13067 12244 13076 12284
rect 13769 12244 13891 12284
rect 13940 12244 13949 12284
rect 3103 12076 3112 12116
rect 3480 12076 3489 12116
rect 6307 12076 6316 12116
rect 6356 12076 6740 12116
rect 9388 12160 11060 12200
rect 11212 12200 11252 12244
rect 11212 12160 12652 12200
rect 12692 12160 12701 12200
rect 2956 11992 5548 12032
rect 5588 11992 5597 12032
rect 1411 11908 1420 11948
rect 1460 11908 1469 11948
rect 1420 11864 1460 11908
rect 2956 11864 2996 11992
rect 3331 11908 3340 11948
rect 3380 11908 3764 11948
rect 6857 11908 6883 11948
rect 6923 11908 6988 11948
rect 7028 11908 7037 11948
rect 7459 11908 7468 11948
rect 7508 11908 8332 11948
rect 8372 11908 8381 11948
rect 988 11824 1132 11864
rect 1172 11824 1460 11864
rect 2908 11824 2996 11864
rect 3043 11824 3052 11864
rect 3092 11824 3668 11864
rect 988 11780 1028 11824
rect 2908 11780 2948 11824
rect 3628 11780 3668 11824
rect 970 11740 979 11780
rect 1019 11740 1028 11780
rect 1411 11740 1420 11780
rect 1460 11740 2324 11780
rect 2371 11740 2380 11780
rect 2420 11740 2551 11780
rect 2908 11740 3148 11780
rect 3188 11740 3197 11780
rect 3610 11740 3619 11780
rect 3659 11740 3668 11780
rect 2284 11696 2324 11740
rect 2908 11738 2948 11740
rect 2890 11698 2899 11738
rect 2939 11698 2948 11738
rect 3724 11696 3764 11908
rect 6892 11864 6932 11908
rect 3820 11824 4204 11864
rect 4244 11824 4253 11864
rect 6700 11824 6932 11864
rect 3820 11780 3860 11824
rect 6700 11780 6740 11824
rect 3811 11740 3820 11780
rect 3860 11740 3869 11780
rect 6089 11740 6220 11780
rect 6260 11740 6269 11780
rect 6442 11771 6740 11780
rect 6442 11731 6451 11771
rect 6491 11740 6740 11771
rect 6787 11740 6796 11780
rect 6836 11740 6898 11780
rect 6938 11740 7468 11780
rect 7508 11740 7517 11780
rect 8419 11740 8428 11780
rect 8468 11740 8564 11780
rect 6491 11731 6500 11740
rect 6442 11730 6500 11731
rect 8524 11696 8564 11740
rect 9388 11696 9428 12160
rect 10877 12076 10886 12116
rect 11254 12076 11263 12116
rect 10444 11992 12940 12032
rect 12980 11992 12989 12032
rect 10444 11948 10484 11992
rect 9571 11908 9580 11948
rect 9620 11908 10388 11948
rect 10435 11908 10444 11948
rect 10484 11908 10493 11948
rect 10636 11908 12460 11948
rect 12500 11908 12509 11948
rect 12617 11908 12748 11948
rect 12788 11908 12797 11948
rect 10051 11824 10060 11864
rect 10100 11824 10109 11864
rect 10060 11780 10100 11824
rect 9964 11740 10100 11780
rect 10147 11740 10156 11780
rect 10196 11740 10205 11780
rect 9964 11696 10004 11740
rect 10156 11696 10196 11740
rect 10348 11696 10388 11908
rect 10636 11696 10676 11908
rect 10828 11824 12980 11864
rect 10828 11696 10868 11824
rect 11209 11740 11218 11780
rect 11258 11740 11731 11780
rect 11771 11740 11780 11780
rect 12451 11740 12460 11780
rect 12500 11740 12509 11780
rect 12460 11696 12500 11740
rect 12940 11696 12980 11824
rect 13036 11780 13076 12244
rect 13996 12116 14036 12487
rect 13315 12076 13324 12116
rect 13364 12076 14036 12116
rect 14284 11948 14324 12496
rect 14443 12485 14452 12525
rect 14492 12485 14516 12525
rect 15209 12496 15286 12536
rect 15326 12496 15340 12536
rect 15380 12496 15389 12536
rect 15610 12496 15619 12536
rect 15659 12496 15668 12536
rect 15715 12496 15724 12536
rect 15764 12496 15773 12536
rect 16492 12527 16588 12536
rect 13987 11908 13996 11948
rect 14036 11908 14324 11948
rect 14476 11948 14516 12485
rect 15628 11948 15668 12496
rect 15724 12032 15764 12496
rect 16532 12496 16588 12527
rect 16628 12496 16663 12536
rect 16841 12496 16972 12536
rect 17012 12496 17021 12536
rect 17129 12496 17209 12536
rect 17249 12496 17260 12536
rect 17300 12496 17309 12536
rect 17740 12527 17780 12580
rect 18508 12536 18644 12538
rect 19564 12536 19604 12580
rect 21100 12536 21140 12580
rect 21580 12536 21620 12580
rect 24652 12536 24692 12664
rect 25036 12620 25076 12832
rect 25385 12664 25507 12704
rect 25556 12664 25565 12704
rect 25036 12580 25460 12620
rect 25420 12536 25460 12580
rect 16492 12478 16532 12487
rect 18499 12496 18508 12536
rect 18548 12498 18700 12536
rect 18548 12496 18557 12498
rect 18604 12496 18700 12498
rect 18740 12496 18749 12536
rect 18883 12496 18892 12536
rect 18932 12496 19276 12536
rect 19316 12496 19372 12536
rect 19412 12496 19421 12536
rect 19555 12496 19564 12536
rect 19604 12496 19613 12536
rect 19747 12496 19756 12536
rect 19796 12496 19927 12536
rect 20131 12496 20140 12536
rect 20180 12496 20276 12536
rect 20323 12496 20332 12536
rect 20372 12496 20524 12536
rect 20564 12496 20573 12536
rect 20707 12496 20716 12536
rect 20756 12496 20887 12536
rect 21091 12496 21100 12536
rect 21140 12496 21149 12536
rect 21283 12496 21292 12536
rect 21332 12496 21620 12536
rect 21850 12496 21859 12536
rect 21908 12496 22039 12536
rect 24643 12496 24652 12536
rect 24692 12496 24701 12536
rect 24931 12496 24940 12536
rect 24980 12496 25076 12536
rect 25121 12496 25130 12536
rect 25170 12533 25179 12536
rect 25170 12496 25268 12533
rect 25402 12496 25411 12536
rect 25451 12496 25460 12536
rect 25708 12536 25748 12832
rect 25891 12664 25900 12704
rect 25940 12664 26036 12704
rect 26729 12664 26860 12704
rect 26900 12664 26909 12704
rect 27331 12664 27340 12704
rect 27380 12664 27764 12704
rect 28073 12664 28204 12704
rect 28244 12664 28253 12704
rect 25996 12620 26036 12664
rect 27724 12620 27764 12664
rect 25795 12580 25804 12620
rect 25844 12580 25940 12620
rect 25996 12580 26708 12620
rect 26836 12580 26956 12620
rect 27007 12580 27016 12620
rect 27235 12580 27244 12620
rect 27284 12580 27380 12620
rect 27427 12580 27436 12620
rect 27476 12580 27614 12620
rect 27654 12580 27663 12620
rect 27724 12580 28148 12620
rect 25900 12536 25940 12580
rect 26668 12536 26708 12580
rect 27340 12536 27380 12580
rect 28108 12536 28148 12580
rect 25708 12496 25719 12536
rect 25759 12496 25768 12536
rect 25882 12527 25940 12536
rect 17740 12478 17780 12487
rect 17059 12412 17068 12452
rect 17131 12412 17239 12452
rect 18409 12412 18418 12452
rect 18458 12412 19084 12452
rect 19124 12412 19133 12452
rect 19756 12368 19796 12496
rect 18115 12328 18124 12368
rect 18164 12328 19796 12368
rect 20236 12368 20276 12496
rect 20716 12452 20756 12496
rect 21292 12452 21332 12496
rect 25036 12452 25076 12496
rect 25132 12493 25268 12496
rect 25228 12452 25268 12493
rect 25882 12487 25891 12527
rect 25931 12487 25940 12527
rect 26035 12496 26044 12536
rect 26084 12496 26188 12536
rect 26228 12496 26237 12536
rect 26650 12496 26659 12536
rect 26699 12496 26708 12536
rect 26755 12496 26764 12536
rect 26804 12496 26935 12536
rect 27043 12496 27052 12536
rect 27092 12496 27095 12536
rect 27135 12496 27223 12536
rect 27331 12496 27340 12536
rect 27380 12496 27389 12536
rect 27689 12496 27820 12536
rect 27860 12496 27869 12536
rect 27916 12527 28003 12536
rect 25882 12486 25940 12487
rect 27956 12496 28003 12527
rect 28099 12496 28108 12536
rect 28148 12496 28157 12536
rect 28204 12496 28281 12536
rect 28321 12496 28330 12536
rect 27916 12452 27956 12487
rect 28204 12452 28244 12496
rect 20716 12412 21332 12452
rect 23116 12443 23156 12452
rect 23273 12412 23404 12452
rect 23444 12412 23453 12452
rect 24905 12412 25036 12452
rect 25076 12412 25085 12452
rect 25228 12412 25804 12452
rect 25844 12412 25853 12452
rect 27212 12412 27221 12452
rect 27261 12412 27270 12452
rect 27427 12412 27436 12452
rect 27476 12412 27607 12452
rect 27907 12412 27916 12452
rect 27956 12412 27965 12452
rect 28099 12412 28108 12452
rect 28148 12412 28244 12452
rect 23116 12394 23156 12403
rect 20236 12328 21196 12368
rect 21236 12328 21245 12368
rect 17434 12244 17443 12284
rect 17483 12244 17492 12284
rect 19747 12244 19756 12284
rect 19796 12244 19852 12284
rect 19892 12244 19927 12284
rect 20131 12244 20140 12284
rect 20180 12244 20189 12284
rect 20899 12244 20908 12284
rect 20948 12244 21100 12284
rect 21140 12244 21772 12284
rect 21812 12244 21821 12284
rect 23587 12244 23596 12284
rect 23636 12244 23980 12284
rect 24020 12244 24029 12284
rect 15811 12160 15820 12200
rect 15860 12160 17068 12200
rect 17108 12160 17117 12200
rect 17452 12032 17492 12244
rect 20140 12200 20180 12244
rect 25036 12200 25076 12412
rect 27221 12368 27261 12412
rect 27221 12328 27244 12368
rect 27284 12328 27308 12368
rect 28387 12328 28396 12368
rect 28436 12328 28492 12368
rect 28532 12328 28567 12368
rect 28745 12328 28876 12368
rect 28916 12328 28925 12368
rect 25411 12244 25420 12284
rect 25460 12244 25708 12284
rect 25748 12244 25757 12284
rect 27497 12244 27532 12284
rect 27572 12244 27619 12284
rect 27659 12244 27677 12284
rect 20140 12160 20236 12200
rect 20276 12160 20285 12200
rect 25036 12160 27724 12200
rect 27764 12160 27773 12200
rect 18651 12076 18660 12116
rect 19028 12076 19037 12116
rect 19651 12076 19660 12116
rect 19700 12076 22828 12116
rect 22868 12076 22877 12116
rect 15724 11992 15860 12032
rect 14476 11908 14764 11948
rect 14804 11908 14813 11948
rect 15628 11908 15724 11948
rect 15764 11908 15773 11948
rect 15820 11864 15860 11992
rect 17314 11992 17492 12032
rect 15052 11824 15860 11864
rect 16460 11855 16684 11864
rect 15052 11780 15092 11824
rect 16500 11824 16684 11855
rect 16724 11824 16733 11864
rect 16460 11806 16500 11815
rect 17314 11780 17354 11992
rect 25036 11948 25076 12160
rect 26425 12076 26434 12116
rect 26802 12076 26811 12116
rect 25516 11992 26284 12032
rect 26324 11992 27916 12032
rect 27956 11992 27965 12032
rect 25516 11948 25556 11992
rect 17417 11908 17443 11948
rect 17483 11908 17548 11948
rect 17588 11908 17597 11948
rect 19267 11908 19276 11948
rect 19316 11908 19372 11948
rect 19412 11908 19447 11948
rect 21283 11908 21292 11948
rect 21332 11908 22732 11948
rect 22772 11908 22781 11948
rect 24067 11908 24076 11948
rect 24116 11908 25076 11948
rect 25507 11908 25516 11948
rect 25556 11908 25565 11948
rect 27244 11908 28876 11948
rect 28916 11908 28925 11948
rect 17443 11824 17452 11864
rect 17492 11824 19028 11864
rect 22723 11824 22732 11864
rect 22772 11824 23924 11864
rect 13036 11740 13635 11780
rect 13675 11740 13684 11780
rect 14092 11740 14420 11780
rect 14092 11696 14132 11740
rect 14380 11696 14420 11740
rect 14476 11740 15092 11780
rect 15139 11740 15148 11780
rect 15188 11740 15236 11780
rect 15305 11740 15436 11780
rect 15476 11740 15485 11780
rect 15811 11740 15820 11780
rect 15866 11740 15991 11780
rect 16963 11740 16972 11780
rect 17012 11740 17164 11780
rect 17204 11740 17213 11780
rect 17314 11740 17492 11780
rect 1165 11656 1174 11696
rect 1214 11656 1228 11696
rect 1268 11656 1354 11696
rect 1498 11656 1507 11696
rect 1547 11656 1556 11696
rect 1603 11656 1612 11696
rect 1652 11656 1708 11696
rect 1748 11656 2039 11696
rect 2079 11656 2088 11696
rect 2170 11656 2179 11696
rect 2219 11656 2228 11696
rect 2275 11656 2284 11696
rect 2324 11656 2333 11696
rect 3032 11656 3041 11696
rect 3081 11656 3092 11696
rect 3220 11656 3340 11696
rect 3391 11656 3400 11696
rect 3475 11656 3484 11696
rect 3524 11656 3533 11696
rect 3715 11656 3724 11696
rect 3764 11656 3773 11696
rect 4140 11656 4204 11696
rect 4244 11656 4300 11696
rect 4340 11656 4396 11696
rect 4436 11656 4445 11696
rect 4841 11656 4972 11696
rect 5012 11656 5021 11696
rect 5098 11656 5107 11696
rect 5147 11656 5164 11696
rect 5204 11656 5287 11696
rect 5364 11656 5452 11696
rect 5492 11656 5495 11696
rect 5535 11656 5544 11696
rect 5626 11656 5635 11696
rect 5675 11656 5684 11696
rect 5731 11656 5740 11696
rect 5780 11656 5911 11696
rect 6185 11656 6316 11696
rect 6356 11656 6365 11696
rect 6544 11656 6553 11696
rect 6593 11656 6604 11696
rect 6644 11656 6733 11696
rect 6979 11656 6988 11696
rect 7028 11656 7037 11696
rect 7625 11656 7756 11696
rect 7796 11656 7805 11696
rect 7913 11656 8044 11696
rect 8084 11656 8093 11696
rect 8404 11656 8413 11696
rect 8453 11656 8468 11696
rect 8515 11656 8524 11696
rect 8564 11656 8573 11696
rect 8873 11656 9004 11696
rect 9044 11656 9053 11696
rect 9379 11656 9388 11696
rect 9428 11656 9437 11696
rect 9763 11656 9772 11696
rect 9812 11656 9821 11696
rect 9946 11656 9955 11696
rect 9995 11656 10004 11696
rect 10141 11656 10150 11696
rect 10190 11656 10243 11696
rect 10348 11656 10455 11696
rect 10495 11656 10504 11696
rect 10627 11656 10636 11696
rect 10676 11656 10685 11696
rect 10819 11656 10828 11696
rect 10868 11656 10877 11696
rect 11299 11656 11308 11696
rect 11348 11656 11500 11696
rect 11540 11656 11549 11696
rect 11849 11656 11980 11696
rect 12020 11656 12029 11696
rect 12163 11656 12172 11696
rect 12212 11656 12364 11696
rect 12404 11656 12413 11696
rect 12460 11656 12796 11696
rect 12836 11656 12845 11696
rect 12931 11656 12940 11696
rect 12980 11656 13228 11696
rect 13268 11656 13277 11696
rect 13507 11656 13516 11696
rect 13556 11656 13565 11696
rect 13708 11656 13733 11696
rect 13773 11656 13782 11696
rect 13891 11656 13900 11696
rect 13940 11656 13949 11696
rect 14083 11656 14092 11696
rect 14132 11656 14141 11696
rect 14188 11656 14275 11696
rect 14315 11656 14324 11696
rect 14371 11656 14380 11696
rect 14420 11656 14429 11696
rect 1516 11612 1556 11656
rect 2188 11612 2228 11656
rect 3052 11612 3092 11656
rect 1516 11572 1612 11612
rect 1652 11572 2228 11612
rect 2284 11572 2900 11612
rect 3043 11572 3052 11612
rect 3092 11572 3137 11612
rect 2284 11528 2324 11572
rect 2860 11528 2900 11572
rect 3484 11528 3524 11656
rect 5644 11612 5684 11656
rect 6988 11612 7028 11656
rect 8428 11612 8468 11656
rect 5059 11572 5068 11612
rect 5108 11572 5684 11612
rect 5818 11572 5827 11612
rect 5867 11572 6124 11612
rect 6164 11572 6173 11612
rect 6988 11572 7604 11612
rect 8428 11572 9044 11612
rect 7564 11528 7604 11572
rect 9004 11528 9044 11572
rect 1891 11488 1900 11528
rect 1940 11488 2324 11528
rect 2380 11488 2707 11528
rect 2747 11488 2756 11528
rect 2860 11488 3139 11528
rect 3179 11488 3524 11528
rect 4099 11488 4108 11528
rect 4148 11488 4195 11528
rect 4235 11488 4279 11528
rect 4483 11488 4492 11528
rect 4532 11488 4541 11528
rect 5129 11488 5260 11528
rect 5300 11488 5309 11528
rect 7546 11488 7555 11528
rect 7595 11488 7604 11528
rect 8995 11488 9004 11528
rect 9044 11488 9484 11528
rect 9524 11488 9533 11528
rect 2380 11444 2420 11488
rect 1795 11404 1804 11444
rect 1844 11404 2420 11444
rect 4492 11444 4532 11488
rect 4492 11404 5164 11444
rect 5204 11404 5213 11444
rect 748 11320 3724 11360
rect 3764 11320 3773 11360
rect 4343 11320 4352 11360
rect 4720 11320 4729 11360
rect 748 11192 788 11320
rect 2881 11236 4108 11276
rect 4148 11236 4157 11276
rect 4204 11236 6836 11276
rect 2881 11192 2921 11236
rect 4204 11192 4244 11236
rect 739 11152 748 11192
rect 788 11152 797 11192
rect 1481 11152 1612 11192
rect 1652 11152 1661 11192
rect 2249 11152 2380 11192
rect 2420 11152 2429 11192
rect 2633 11152 2764 11192
rect 2804 11152 2813 11192
rect 2860 11152 2921 11192
rect 3043 11152 3052 11192
rect 3092 11152 3235 11192
rect 3275 11152 3284 11192
rect 4186 11152 4195 11192
rect 4235 11152 4244 11192
rect 4474 11152 4483 11192
rect 4523 11152 5452 11192
rect 5492 11152 5501 11192
rect 6490 11152 6499 11192
rect 6539 11152 6604 11192
rect 6644 11152 6679 11192
rect 2860 11108 2900 11152
rect 739 11068 748 11108
rect 788 11068 797 11108
rect 931 11068 940 11108
rect 980 11068 2900 11108
rect 748 11024 788 11068
rect 2860 11024 2900 11068
rect 2956 11068 3148 11108
rect 3188 11068 3197 11108
rect 3436 11068 4148 11108
rect 4457 11068 4588 11108
rect 4628 11068 4637 11108
rect 5068 11068 5260 11108
rect 5300 11068 5309 11108
rect 5452 11068 5828 11108
rect 2956 11024 2996 11068
rect 643 10984 652 11024
rect 692 10984 701 11024
rect 748 10984 835 11024
rect 875 10984 884 11024
rect 1123 10984 1132 11024
rect 1172 10984 1324 11024
rect 1364 10984 1373 11024
rect 1450 10984 1459 11024
rect 1499 10984 1612 11024
rect 1652 10984 1804 11024
rect 1844 10984 1853 11024
rect 1978 10984 1987 11024
rect 2027 10984 2036 11024
rect 2083 10984 2092 11024
rect 2132 10984 2263 11024
rect 2755 10984 2764 11024
rect 2804 10984 2900 11024
rect 2947 10984 2956 11024
rect 2996 10984 3005 11024
rect 3209 10984 3340 11024
rect 3380 10984 3389 11024
rect 652 10940 692 10984
rect 1132 10940 1172 10984
rect 652 10900 1172 10940
rect 1996 10856 2036 10984
rect 3436 10940 3476 11068
rect 4108 11024 4148 11068
rect 5068 11024 5108 11068
rect 5452 11024 5492 11068
rect 5788 11024 5828 11068
rect 6796 11024 6836 11236
rect 7564 11192 7604 11488
rect 9772 11360 9812 11656
rect 13516 11612 13556 11656
rect 9859 11572 9868 11612
rect 9908 11572 10100 11612
rect 10217 11572 10252 11612
rect 10292 11572 10348 11612
rect 10388 11572 10397 11612
rect 10723 11572 10732 11612
rect 10772 11572 12844 11612
rect 12884 11572 12893 11612
rect 12940 11572 13556 11612
rect 10060 11444 10100 11572
rect 12940 11528 12980 11572
rect 11002 11488 11011 11528
rect 11060 11488 11191 11528
rect 12643 11488 12652 11528
rect 12692 11488 12980 11528
rect 13027 11488 13036 11528
rect 13076 11488 13420 11528
rect 13460 11488 13469 11528
rect 10060 11404 11980 11444
rect 12020 11404 12029 11444
rect 13708 11360 13748 11656
rect 13900 11612 13940 11656
rect 14188 11612 14228 11656
rect 14476 11612 14516 11740
rect 15196 11696 15236 11740
rect 17452 11696 17492 11740
rect 14633 11656 14764 11696
rect 14804 11656 14813 11696
rect 14860 11656 14956 11696
rect 14996 11656 15005 11696
rect 15086 11656 15095 11696
rect 15135 11656 15144 11696
rect 15196 11656 15235 11696
rect 15275 11656 15284 11696
rect 15332 11656 15341 11696
rect 15381 11656 15390 11696
rect 15907 11656 15916 11696
rect 15956 11656 16300 11696
rect 16340 11656 16349 11696
rect 16474 11656 16483 11696
rect 16523 11656 16532 11696
rect 16675 11656 16684 11696
rect 16724 11656 17068 11696
rect 17108 11656 17117 11696
rect 17178 11656 17187 11696
rect 17227 11656 17236 11696
rect 17296 11656 17305 11696
rect 17345 11656 17354 11696
rect 17432 11656 17441 11696
rect 17481 11656 17492 11696
rect 13900 11572 14188 11612
rect 14228 11572 14237 11612
rect 14467 11572 14476 11612
rect 14516 11572 14525 11612
rect 14572 11572 14583 11612
rect 14623 11572 14632 11612
rect 14249 11488 14371 11528
rect 14420 11488 14429 11528
rect 14572 11444 14612 11572
rect 13795 11404 13804 11444
rect 13844 11404 14612 11444
rect 14860 11444 14900 11656
rect 15095 11612 15135 11656
rect 15340 11612 15380 11656
rect 16492 11612 16532 11656
rect 14947 11572 14956 11612
rect 14996 11572 15135 11612
rect 15235 11572 15244 11612
rect 15284 11572 16532 11612
rect 17187 11528 17227 11656
rect 17314 11612 17354 11656
rect 17620 11612 17660 11824
rect 18761 11740 18883 11780
rect 18932 11740 18941 11780
rect 17740 11696 17780 11705
rect 18988 11696 19028 11824
rect 23884 11780 23924 11824
rect 20044 11740 20236 11780
rect 20276 11740 20285 11780
rect 21955 11740 21964 11780
rect 22004 11740 22013 11780
rect 22531 11740 22540 11780
rect 22580 11740 23443 11780
rect 23483 11740 23492 11780
rect 23570 11740 23596 11780
rect 23636 11740 23657 11780
rect 23872 11740 23884 11780
rect 23924 11740 23959 11780
rect 27244 11760 27284 11908
rect 27497 11824 27628 11864
rect 27668 11824 27677 11864
rect 27907 11824 27916 11864
rect 27956 11824 27965 11864
rect 28099 11824 28108 11864
rect 28148 11824 28204 11864
rect 28244 11824 28279 11864
rect 20044 11696 20084 11740
rect 23617 11696 23657 11740
rect 23919 11696 23959 11740
rect 27341 11740 27427 11780
rect 27467 11740 27476 11780
rect 27715 11740 27724 11780
rect 27764 11740 27773 11780
rect 17731 11656 17740 11696
rect 17780 11656 17911 11696
rect 18377 11656 18508 11696
rect 18548 11656 18557 11696
rect 18612 11656 18700 11696
rect 18740 11656 18743 11696
rect 18783 11656 18792 11696
rect 18979 11656 18988 11696
rect 19028 11656 19037 11696
rect 19337 11656 19468 11696
rect 19508 11656 19517 11696
rect 20026 11656 20035 11696
rect 20075 11656 20084 11696
rect 20131 11656 20140 11696
rect 20180 11656 20812 11696
rect 20852 11656 20861 11696
rect 21178 11656 21187 11696
rect 21227 11656 21868 11696
rect 21908 11656 21917 11696
rect 23599 11656 23608 11696
rect 23648 11656 23657 11696
rect 23779 11656 23788 11696
rect 23828 11656 23837 11696
rect 23901 11656 23910 11696
rect 23950 11656 23959 11696
rect 24028 11731 24086 11738
rect 24028 11729 24116 11731
rect 24028 11689 24037 11729
rect 24077 11689 24116 11729
rect 24028 11688 24116 11689
rect 17740 11647 17780 11656
rect 23788 11612 23828 11656
rect 17314 11572 17452 11612
rect 17492 11572 17501 11612
rect 17620 11572 17644 11612
rect 17684 11572 17693 11612
rect 17923 11572 17932 11612
rect 17972 11572 18115 11612
rect 18155 11572 18164 11612
rect 20794 11572 20803 11612
rect 20843 11572 21580 11612
rect 21620 11572 21629 11612
rect 21763 11572 21772 11612
rect 21812 11572 23828 11612
rect 24076 11612 24116 11688
rect 24163 11656 24172 11696
rect 24212 11656 24268 11696
rect 24308 11656 25172 11696
rect 26947 11656 26956 11696
rect 26996 11656 27043 11696
rect 27083 11656 27148 11696
rect 27188 11656 27197 11696
rect 25132 11612 25172 11656
rect 24076 11572 24364 11612
rect 24404 11572 24413 11612
rect 25114 11572 25123 11612
rect 25163 11572 25172 11612
rect 27341 11528 27381 11740
rect 27529 11729 27668 11738
rect 27529 11698 27628 11729
rect 27529 11696 27569 11698
rect 27427 11656 27436 11696
rect 27476 11656 27569 11696
rect 27724 11696 27764 11740
rect 27916 11729 27956 11824
rect 27628 11680 27668 11689
rect 27717 11656 27726 11696
rect 27766 11656 27811 11696
rect 27916 11680 27956 11689
rect 17187 11488 19075 11528
rect 19115 11488 19124 11528
rect 20419 11488 20428 11528
rect 20468 11488 20908 11528
rect 20948 11488 20957 11528
rect 23107 11488 23116 11528
rect 23156 11488 23732 11528
rect 24809 11488 24940 11528
rect 24980 11488 24989 11528
rect 27341 11488 27532 11528
rect 27572 11488 27581 11528
rect 23692 11444 23732 11488
rect 14860 11404 17260 11444
rect 17300 11404 17309 11444
rect 19363 11404 19372 11444
rect 19412 11404 23308 11444
rect 23348 11404 23357 11444
rect 23692 11404 24460 11444
rect 24500 11404 24509 11444
rect 14860 11360 14900 11404
rect 9772 11320 10060 11360
rect 10100 11320 10109 11360
rect 10243 11320 10252 11360
rect 10292 11320 10732 11360
rect 10772 11320 11153 11360
rect 12117 11320 12126 11360
rect 12494 11320 12503 11360
rect 13708 11320 14900 11360
rect 19891 11320 19900 11360
rect 20268 11320 20277 11360
rect 21283 11320 21292 11360
rect 21332 11320 24020 11360
rect 27665 11320 27674 11360
rect 28042 11320 28051 11360
rect 8419 11236 8428 11276
rect 8468 11236 8852 11276
rect 9763 11236 9772 11276
rect 9812 11236 10636 11276
rect 10676 11236 10685 11276
rect 7241 11152 7324 11192
rect 7364 11152 7372 11192
rect 7412 11152 7421 11192
rect 7546 11152 7555 11192
rect 7595 11152 7604 11192
rect 8393 11152 8524 11192
rect 8564 11152 8573 11192
rect 7721 11068 7770 11108
rect 7810 11068 7852 11108
rect 7892 11068 7901 11108
rect 8419 11068 8428 11108
rect 8468 11068 8716 11108
rect 8756 11068 8765 11108
rect 8812 11024 8852 11236
rect 9091 11152 9100 11192
rect 9140 11152 9428 11192
rect 9571 11152 9580 11192
rect 9620 11152 9868 11192
rect 9908 11152 9917 11192
rect 10138 11152 10147 11192
rect 10187 11152 10580 11192
rect 9187 11068 9196 11108
rect 9236 11068 9245 11108
rect 9196 11024 9236 11068
rect 9388 11024 9428 11152
rect 9562 11068 9571 11108
rect 9611 11068 10100 11108
rect 10147 11068 10156 11108
rect 10196 11068 10348 11108
rect 10388 11068 10397 11108
rect 10060 11024 10100 11068
rect 10540 11024 10580 11152
rect 11113 11024 11153 11320
rect 11404 11236 12836 11276
rect 11404 11108 11444 11236
rect 11491 11152 11500 11192
rect 11540 11152 12068 11192
rect 12346 11152 12355 11192
rect 12395 11152 12556 11192
rect 12596 11152 12605 11192
rect 11404 11068 11732 11108
rect 11692 11024 11732 11068
rect 2179 10900 2188 10940
rect 2228 10900 3476 10940
rect 3614 10984 3724 11024
rect 3764 10984 3863 11024
rect 3903 10984 3924 11024
rect 4099 10984 4108 11024
rect 4148 10984 4157 11024
rect 4265 10984 4387 11024
rect 4436 10984 4445 11024
rect 4675 10984 4684 11024
rect 4735 10984 4855 11024
rect 5050 10984 5059 11024
rect 5099 10984 5108 11024
rect 5155 10984 5164 11024
rect 5204 10984 5492 11024
rect 5539 10984 5548 11024
rect 5588 10984 5596 11024
rect 5636 10984 5719 11024
rect 5788 10984 5897 11024
rect 5937 10984 5946 11024
rect 6019 10984 6028 11024
rect 6091 10984 6199 11024
rect 6595 10984 6604 11024
rect 6644 10984 6653 11024
rect 6796 10984 6988 11024
rect 7028 10984 7037 11024
rect 7171 10984 7180 11024
rect 7220 10984 7229 11024
rect 7337 10984 7459 11024
rect 7508 10984 7517 11024
rect 7660 10984 7948 11024
rect 7988 10984 7997 11024
rect 8131 10984 8140 11024
rect 8180 10984 8189 11024
rect 8314 10984 8323 11024
rect 8363 10984 8372 11024
rect 8500 10984 8620 11024
rect 8671 10984 8680 11024
rect 8803 10984 8812 11024
rect 8852 10984 8861 11024
rect 8945 10984 8954 11024
rect 8994 10984 9004 11024
rect 9044 10984 9134 11024
rect 9196 10984 9239 11024
rect 9279 10984 9288 11024
rect 9388 10984 9484 11024
rect 9524 10984 9533 11024
rect 10051 10984 10060 11024
rect 10100 10984 10109 11024
rect 10522 10984 10531 11024
rect 10571 10984 11020 11024
rect 11060 10984 11069 11024
rect 11113 10984 11128 11024
rect 11168 10984 11177 11024
rect 11683 10984 11692 11024
rect 11732 10984 11741 11024
rect 11788 10984 11875 11024
rect 11915 10984 11924 11024
rect 1987 10816 1996 10856
rect 2036 10816 2045 10856
rect 3103 10564 3112 10604
rect 3480 10564 3489 10604
rect 3614 10520 3654 10984
rect 5068 10940 5108 10984
rect 3811 10900 3820 10940
rect 3860 10900 4003 10940
rect 4043 10900 4052 10940
rect 5068 10900 5740 10940
rect 5780 10900 5789 10940
rect 5705 10816 5836 10856
rect 5876 10816 5885 10856
rect 3148 10480 3654 10520
rect 3148 10436 3188 10480
rect 6604 10436 6644 10984
rect 7180 10940 7220 10984
rect 6691 10900 6700 10940
rect 6740 10900 7220 10940
rect 7660 10604 7700 10984
rect 8140 10856 8180 10984
rect 8332 10940 8372 10984
rect 10060 10940 10100 10984
rect 11788 10940 11828 10984
rect 12028 10982 12068 11152
rect 12796 11108 12836 11236
rect 12940 11236 14380 11276
rect 14420 11236 14429 11276
rect 17731 11236 17740 11276
rect 17780 11236 23060 11276
rect 12940 11192 12980 11236
rect 12922 11152 12931 11192
rect 12971 11152 12980 11192
rect 13097 11152 13219 11192
rect 13268 11152 13277 11192
rect 13978 11152 13987 11192
rect 14027 11152 14188 11192
rect 14228 11152 14237 11192
rect 14746 11152 14755 11192
rect 14795 11152 14804 11192
rect 15043 11152 15052 11192
rect 15092 11152 16483 11192
rect 16523 11152 16532 11192
rect 16771 11152 16780 11192
rect 16820 11152 16829 11192
rect 17443 11152 17452 11192
rect 17492 11152 17740 11192
rect 17780 11152 17789 11192
rect 18010 11152 18019 11192
rect 18059 11152 18499 11192
rect 18539 11152 18700 11192
rect 18740 11152 18749 11192
rect 18892 11152 20035 11192
rect 20075 11152 20084 11192
rect 20515 11152 20524 11192
rect 20564 11152 21772 11192
rect 21812 11152 21821 11192
rect 14764 11108 14804 11152
rect 16780 11108 16820 11152
rect 12604 11068 12652 11108
rect 12692 11068 12701 11108
rect 12796 11068 14804 11108
rect 15244 11068 16204 11108
rect 16244 11068 17588 11108
rect 12604 11024 12644 11068
rect 14476 11024 14516 11068
rect 15244 11024 15284 11068
rect 17548 11024 17588 11068
rect 17932 11068 18796 11108
rect 18836 11068 18845 11108
rect 17932 11024 17972 11068
rect 18892 11024 18932 11152
rect 23020 11108 23060 11236
rect 23980 11192 24020 11320
rect 25795 11236 25804 11276
rect 25844 11236 27436 11276
rect 27476 11236 27764 11276
rect 27724 11192 27764 11236
rect 23347 11152 23356 11192
rect 23396 11152 23788 11192
rect 23828 11152 23837 11192
rect 23971 11152 23980 11192
rect 24020 11152 24029 11192
rect 24355 11152 24364 11192
rect 24404 11152 24604 11192
rect 24644 11152 24653 11192
rect 25315 11152 25324 11192
rect 25364 11152 26188 11192
rect 26228 11152 27284 11192
rect 27706 11152 27715 11192
rect 27755 11152 27764 11192
rect 19699 11068 19708 11108
rect 19748 11068 21868 11108
rect 21908 11068 21917 11108
rect 22435 11068 22444 11108
rect 22484 11068 22964 11108
rect 23020 11068 23540 11108
rect 22924 11024 22964 11068
rect 12259 10984 12268 11024
rect 12309 10984 12439 11024
rect 12595 10984 12604 11024
rect 12644 10984 12653 11024
rect 12713 10984 12844 11024
rect 12884 10984 12893 11024
rect 13411 10984 13420 11024
rect 13460 10984 13469 11024
rect 13577 10984 13708 11024
rect 13748 10984 13757 11024
rect 14056 10984 14092 11024
rect 14132 10984 14141 11024
rect 14467 10984 14476 11024
rect 14516 10984 14525 11024
rect 14947 10984 14956 11024
rect 14996 10984 15005 11024
rect 15235 10984 15244 11024
rect 15284 10984 15293 11024
rect 16003 11000 16012 11024
rect 15942 10984 16012 11000
rect 16052 10984 16061 11024
rect 16138 10984 16147 11024
rect 16187 10984 16396 11024
rect 16436 10984 16445 11024
rect 16649 10984 16780 11024
rect 16820 10984 16829 11024
rect 16963 10984 16972 11024
rect 17012 10984 17251 11024
rect 17291 10984 17300 11024
rect 17417 10984 17548 11024
rect 17588 10984 17597 11024
rect 17923 10984 17932 11024
rect 17972 10984 17981 11024
rect 18115 10984 18124 11024
rect 18164 10984 18167 11024
rect 18207 10984 18295 11024
rect 18403 10984 18412 11024
rect 18452 10984 18461 11024
rect 18508 10984 18932 11024
rect 19021 10984 19030 11024
rect 19070 10984 19180 11024
rect 19220 10984 19229 11024
rect 19433 11015 19564 11024
rect 19433 10984 19555 11015
rect 19604 10984 19613 11024
rect 20201 10984 20332 11024
rect 20372 10984 20381 11024
rect 20777 10984 20908 11024
rect 20948 10984 20957 11024
rect 21475 10984 21484 11024
rect 21524 10984 22444 11024
rect 22484 10984 22493 11024
rect 22723 10984 22732 11024
rect 22772 10984 22781 11024
rect 22915 10984 22924 11024
rect 22964 10984 22973 11024
rect 23020 11015 23252 11024
rect 23020 10984 23203 11015
rect 12019 10942 12028 10982
rect 12068 10942 12077 10982
rect 13420 10940 13460 10984
rect 8332 10900 9196 10940
rect 9236 10900 9245 10940
rect 9370 10900 9379 10940
rect 9419 10900 9772 10940
rect 9812 10900 9821 10940
rect 10060 10900 10580 10940
rect 10540 10898 10580 10900
rect 10732 10900 10963 10940
rect 11003 10900 11012 10940
rect 11177 10900 11308 10940
rect 11348 10900 11357 10940
rect 11740 10900 11828 10940
rect 12154 10900 12163 10940
rect 12212 10900 12343 10940
rect 12617 10900 12739 10940
rect 12788 10900 12797 10940
rect 13420 10900 13900 10940
rect 13940 10900 13949 10940
rect 10540 10858 10572 10898
rect 10612 10858 10621 10898
rect 8140 10816 10156 10856
rect 10196 10816 10205 10856
rect 10732 10772 10772 10900
rect 11740 10772 11780 10900
rect 11866 10816 11875 10856
rect 11915 10816 13804 10856
rect 13844 10816 13853 10856
rect 14056 10772 14096 10984
rect 14956 10940 14996 10984
rect 15942 10960 16052 10984
rect 14956 10900 15244 10940
rect 15284 10900 15293 10940
rect 15942 10856 15982 10960
rect 16204 10900 16690 10940
rect 16730 10900 16739 10940
rect 17548 10900 18307 10940
rect 18347 10900 18356 10940
rect 16204 10856 16244 10900
rect 17548 10856 17588 10900
rect 15043 10816 15052 10856
rect 15092 10816 15982 10856
rect 16186 10816 16195 10856
rect 16235 10816 16244 10856
rect 17539 10816 17548 10856
rect 17588 10816 17597 10856
rect 7747 10732 7756 10772
rect 7796 10732 7805 10772
rect 8035 10732 8044 10772
rect 8084 10732 9964 10772
rect 10004 10732 10013 10772
rect 10627 10732 10636 10772
rect 10676 10732 10772 10772
rect 11539 10732 11548 10772
rect 11588 10732 11597 10772
rect 11740 10732 14096 10772
rect 15942 10772 15982 10816
rect 15942 10732 18124 10772
rect 18164 10732 18173 10772
rect 7756 10688 7796 10732
rect 7756 10648 9100 10688
rect 9140 10648 9149 10688
rect 11548 10604 11588 10732
rect 7660 10564 9580 10604
rect 9620 10564 10252 10604
rect 10292 10564 10301 10604
rect 10877 10564 10886 10604
rect 11254 10564 11263 10604
rect 11548 10564 13228 10604
rect 13268 10564 13277 10604
rect 11548 10520 11588 10564
rect 7939 10480 7948 10520
rect 7988 10480 10444 10520
rect 10484 10480 10493 10520
rect 11548 10480 11828 10520
rect 11875 10480 11884 10520
rect 11924 10480 12788 10520
rect 1747 10396 1756 10436
rect 1796 10396 1996 10436
rect 2036 10396 2045 10436
rect 2092 10396 2956 10436
rect 2996 10396 3005 10436
rect 3130 10396 3139 10436
rect 3179 10396 3188 10436
rect 3401 10396 3532 10436
rect 3572 10396 3581 10436
rect 4474 10396 4483 10436
rect 4523 10396 4780 10436
rect 4820 10396 4829 10436
rect 6586 10396 6595 10436
rect 6635 10396 7316 10436
rect 8585 10396 8716 10436
rect 8756 10396 8765 10436
rect 9065 10396 9196 10436
rect 9236 10396 9245 10436
rect 10060 10396 11444 10436
rect 2092 10352 2132 10396
rect 922 10312 931 10352
rect 971 10312 2132 10352
rect 2515 10312 2524 10352
rect 2564 10312 3340 10352
rect 3380 10312 3389 10352
rect 3619 10312 3628 10352
rect 3668 10312 4012 10352
rect 4052 10312 4061 10352
rect 4780 10312 5068 10352
rect 5108 10312 5117 10352
rect 5347 10312 5356 10352
rect 5396 10312 5740 10352
rect 5780 10312 5789 10352
rect 4780 10268 4820 10312
rect 7276 10268 7316 10396
rect 8026 10312 8035 10352
rect 8075 10312 8084 10352
rect 8044 10268 8084 10312
rect 10060 10268 10100 10396
rect 748 10228 940 10268
rect 980 10228 989 10268
rect 1036 10228 1612 10268
rect 1652 10228 1661 10268
rect 1865 10228 1987 10268
rect 2036 10228 2045 10268
rect 2179 10228 2188 10268
rect 2228 10228 2764 10268
rect 2804 10228 2813 10268
rect 3628 10228 4204 10268
rect 4244 10228 4253 10268
rect 4396 10228 4492 10268
rect 4532 10228 4541 10268
rect 4762 10228 4771 10268
rect 4811 10228 4820 10268
rect 4867 10228 4876 10268
rect 4916 10228 4972 10268
rect 5012 10228 5047 10268
rect 5251 10228 5260 10268
rect 5300 10228 5431 10268
rect 5539 10228 5548 10268
rect 5588 10228 5780 10268
rect 748 10184 788 10228
rect 1036 10184 1076 10228
rect 1612 10184 1652 10228
rect 3628 10184 3668 10228
rect 4204 10184 4244 10228
rect 4396 10184 4436 10228
rect 5740 10184 5780 10228
rect 6316 10228 6700 10268
rect 6740 10228 6749 10268
rect 6979 10228 6988 10268
rect 7028 10228 7124 10268
rect 7267 10228 7276 10268
rect 7316 10228 7325 10268
rect 7756 10228 7852 10268
rect 7892 10228 7901 10268
rect 8044 10228 8564 10268
rect 6316 10184 6356 10228
rect 7084 10184 7124 10228
rect 7756 10184 7796 10228
rect 8524 10184 8564 10228
rect 8620 10228 10100 10268
rect 11116 10228 11308 10268
rect 11348 10228 11357 10268
rect 8620 10184 8660 10228
rect 11116 10226 11156 10228
rect 11098 10217 11156 10226
rect 739 10144 748 10184
rect 788 10144 797 10184
rect 922 10144 931 10184
rect 971 10144 1076 10184
rect 1123 10144 1132 10184
rect 1172 10144 1181 10184
rect 1507 10144 1516 10184
rect 1556 10144 1652 10184
rect 1795 10144 1804 10184
rect 1844 10144 1847 10184
rect 1887 10144 1975 10184
rect 2083 10144 2092 10184
rect 2132 10144 2141 10184
rect 2371 10144 2380 10184
rect 2420 10144 2516 10184
rect 2563 10144 2572 10184
rect 2612 10144 2851 10184
rect 2891 10144 2900 10184
rect 2947 10144 2956 10184
rect 2996 10144 3127 10184
rect 3305 10144 3436 10184
rect 3476 10144 3485 10184
rect 3619 10144 3628 10184
rect 3668 10144 3677 10184
rect 3907 10144 3916 10184
rect 3956 10144 4052 10184
rect 4099 10144 4108 10184
rect 4148 10144 4244 10184
rect 4291 10144 4300 10184
rect 4340 10144 4436 10184
rect 4482 10144 4491 10184
rect 4531 10144 4540 10184
rect 4588 10144 4631 10184
rect 4671 10144 4680 10184
rect 4867 10144 4876 10184
rect 4916 10144 4972 10184
rect 5012 10144 5047 10184
rect 5122 10144 5131 10184
rect 5204 10144 5311 10184
rect 5356 10144 5417 10184
rect 5457 10144 5466 10184
rect 5578 10144 5587 10184
rect 5627 10144 5684 10184
rect 5731 10144 5740 10184
rect 5780 10144 5789 10184
rect 5923 10144 5932 10184
rect 5977 10144 6103 10184
rect 6156 10144 6220 10184
rect 6260 10144 6307 10184
rect 6347 10144 6356 10184
rect 6403 10144 6412 10184
rect 6452 10144 6461 10184
rect 6948 10144 6957 10184
rect 6997 10144 7028 10184
rect 7084 10144 7105 10184
rect 7145 10144 7154 10184
rect 7363 10144 7372 10184
rect 7437 10144 7543 10184
rect 7738 10144 7747 10184
rect 7787 10144 7796 10184
rect 7843 10144 7852 10184
rect 7892 10144 7948 10184
rect 7988 10144 8023 10184
rect 8506 10144 8515 10184
rect 8555 10144 8564 10184
rect 8611 10144 8620 10184
rect 8660 10144 8669 10184
rect 9091 10144 9100 10184
rect 9140 10144 9244 10184
rect 9284 10144 9332 10184
rect 9379 10144 9388 10184
rect 9428 10144 9908 10184
rect 10013 10144 10045 10184
rect 10085 10144 10100 10184
rect 10147 10144 10156 10184
rect 10196 10144 10327 10184
rect 10627 10144 10636 10184
rect 10676 10144 10685 10184
rect 10732 10144 10775 10184
rect 10815 10144 10824 10184
rect 11098 10177 11107 10217
rect 11147 10177 11156 10217
rect 11098 10176 11156 10177
rect 11404 10184 11444 10396
rect 11788 10268 11828 10480
rect 12748 10436 12788 10480
rect 13708 10436 13748 10732
rect 16204 10480 16396 10520
rect 16436 10480 16445 10520
rect 16204 10436 16244 10480
rect 12058 10396 12067 10436
rect 12107 10396 12116 10436
rect 12748 10396 12884 10436
rect 13690 10396 13699 10436
rect 13739 10396 13748 10436
rect 14179 10396 14188 10436
rect 14228 10396 14764 10436
rect 14804 10396 14813 10436
rect 15436 10396 15668 10436
rect 16186 10396 16195 10436
rect 16235 10396 16244 10436
rect 16291 10396 16300 10436
rect 16340 10396 16588 10436
rect 16628 10396 16637 10436
rect 17932 10396 18316 10436
rect 18356 10396 18365 10436
rect 12076 10352 12116 10396
rect 12076 10312 12788 10352
rect 11561 10228 11683 10268
rect 11732 10228 11741 10268
rect 11788 10228 12068 10268
rect 12028 10184 12068 10228
rect 12364 10228 12643 10268
rect 12692 10228 12701 10268
rect 12364 10184 12404 10228
rect 12748 10184 12788 10312
rect 12844 10268 12884 10396
rect 13228 10312 13324 10352
rect 13364 10312 13373 10352
rect 13762 10312 13996 10352
rect 14036 10312 14045 10352
rect 14179 10312 14188 10352
rect 14228 10312 14237 10352
rect 14371 10312 14380 10352
rect 14420 10312 14429 10352
rect 13228 10268 13268 10312
rect 13762 10268 13802 10312
rect 12835 10228 12844 10268
rect 12884 10228 12893 10268
rect 13219 10228 13228 10268
rect 13268 10228 13277 10268
rect 13450 10259 13802 10268
rect 13450 10219 13459 10259
rect 13499 10228 13802 10259
rect 13499 10219 13508 10228
rect 14188 10226 14228 10312
rect 14380 10226 14420 10312
rect 15436 10226 15476 10396
rect 15628 10352 15668 10396
rect 15523 10312 15532 10352
rect 15572 10312 15581 10352
rect 15628 10312 17740 10352
rect 17780 10312 17789 10352
rect 15532 10268 15572 10312
rect 15532 10228 16690 10268
rect 16730 10228 16739 10268
rect 13450 10218 13508 10219
rect 13996 10184 14036 10193
rect 14179 10186 14188 10226
rect 14228 10186 14237 10226
rect 14371 10186 14380 10226
rect 14420 10186 14429 10226
rect 15256 10217 15476 10226
rect 11404 10144 11543 10184
rect 11583 10144 11592 10184
rect 11779 10144 11788 10184
rect 11828 10144 11837 10184
rect 12028 10144 12062 10184
rect 12102 10144 12111 10184
rect 12514 10144 12523 10184
rect 12563 10144 12596 10184
rect 12739 10144 12748 10184
rect 12788 10144 12797 10184
rect 13193 10144 13324 10184
rect 13364 10144 13373 10184
rect 13552 10144 13561 10184
rect 13601 10144 13900 10184
rect 13940 10144 13949 10184
rect 1132 10016 1172 10144
rect 2092 10100 2132 10144
rect 2476 10100 2516 10144
rect 4012 10100 4052 10144
rect 4492 10100 4532 10144
rect 1603 10060 1612 10100
rect 1652 10060 2132 10100
rect 2467 10060 2476 10100
rect 2516 10060 2525 10100
rect 4012 10060 4148 10100
rect 4387 10060 4396 10100
rect 4436 10060 4532 10100
rect 4588 10100 4628 10144
rect 4588 10060 4780 10100
rect 4820 10060 4829 10100
rect 4108 10016 4148 10060
rect 5356 10016 5396 10144
rect 5644 10100 5684 10144
rect 6412 10100 6452 10144
rect 5644 10060 6452 10100
rect 6988 10100 7028 10144
rect 6988 10060 7124 10100
rect 5644 10016 5684 10060
rect 1132 9976 1844 10016
rect 3811 9976 3820 10016
rect 3860 9976 4148 10016
rect 4195 9976 4204 10016
rect 4244 9976 5396 10016
rect 5443 9976 5452 10016
rect 5492 9976 5684 10016
rect 5731 9976 5740 10016
rect 5780 9976 5789 10016
rect 1804 9848 1844 9976
rect 5740 9932 5780 9976
rect 3427 9892 3436 9932
rect 3476 9892 5780 9932
rect 7084 9932 7124 10060
rect 7185 10018 7194 10058
rect 7234 10018 7564 10058
rect 7604 10018 7613 10058
rect 8620 10016 8660 10144
rect 9292 10100 9332 10144
rect 9292 10060 9676 10100
rect 9716 10060 9725 10100
rect 9868 10016 9908 10144
rect 10060 10100 10100 10144
rect 10060 10060 10252 10100
rect 10292 10060 10301 10100
rect 7747 9976 7756 10016
rect 7796 9976 8468 10016
rect 8515 9976 8524 10016
rect 8564 9976 8660 10016
rect 9708 9976 9772 10016
rect 9812 9976 9859 10016
rect 9899 9976 9908 10016
rect 8428 9932 8468 9976
rect 10636 9932 10676 10144
rect 10732 10100 10772 10144
rect 11788 10100 11828 10144
rect 12364 10135 12404 10144
rect 10723 10060 10732 10100
rect 10772 10060 10781 10100
rect 10963 10060 10972 10100
rect 11012 10060 11828 10100
rect 12556 10016 12596 10144
rect 13996 10100 14036 10144
rect 13027 10060 13036 10100
rect 13076 10060 13694 10100
rect 13734 10060 13743 10100
rect 13795 10060 13804 10100
rect 13844 10060 14036 10100
rect 14572 10144 14611 10184
rect 14651 10144 14660 10184
rect 14704 10144 14713 10184
rect 14753 10144 14764 10184
rect 14804 10144 14893 10184
rect 15017 10144 15139 10184
rect 15188 10144 15197 10184
rect 15296 10186 15476 10217
rect 17932 10184 17972 10396
rect 18412 10352 18452 10984
rect 18028 10312 18452 10352
rect 15256 10168 15296 10177
rect 15715 10144 15724 10184
rect 15764 10144 16012 10184
rect 16052 10144 16061 10184
rect 16138 10144 16147 10184
rect 16187 10144 16204 10184
rect 16244 10144 16327 10184
rect 16483 10144 16492 10184
rect 16532 10144 16780 10184
rect 16820 10144 16829 10184
rect 16963 10144 16972 10184
rect 17012 10144 17260 10184
rect 17300 10144 17309 10184
rect 17393 10144 17402 10184
rect 17442 10144 17548 10184
rect 17588 10144 17597 10184
rect 17923 10144 17932 10184
rect 17972 10144 17981 10184
rect 14572 10100 14612 10144
rect 18028 10100 18068 10312
rect 18508 10184 18548 10984
rect 19546 10975 19555 10984
rect 19595 10975 19604 10984
rect 19546 10974 19604 10975
rect 22732 10940 22772 10984
rect 18826 10900 18835 10940
rect 18875 10900 19124 10940
rect 20233 10900 20242 10940
rect 20282 10900 21100 10940
rect 21140 10900 21149 10940
rect 21667 10900 21676 10940
rect 21716 10900 22348 10940
rect 22388 10900 22772 10940
rect 18651 10564 18660 10604
rect 19028 10564 19037 10604
rect 19084 10436 19124 10900
rect 19363 10816 19372 10856
rect 19412 10816 19796 10856
rect 22601 10816 22723 10856
rect 22772 10816 22781 10856
rect 18979 10396 18988 10436
rect 19028 10396 19124 10436
rect 18211 10144 18220 10184
rect 18260 10144 18269 10184
rect 18394 10144 18403 10184
rect 18443 10144 18548 10184
rect 18796 10312 19604 10352
rect 14572 10060 14668 10100
rect 14708 10060 14717 10100
rect 14899 10060 14908 10100
rect 14948 10060 16012 10100
rect 16052 10060 16061 10100
rect 17587 10060 17596 10100
rect 17636 10060 18068 10100
rect 11011 9976 11020 10016
rect 11060 9976 11260 10016
rect 11300 9976 11309 10016
rect 11849 9976 11875 10016
rect 11915 9976 11980 10016
rect 12020 9976 12029 10016
rect 12259 9976 12268 10016
rect 12308 9976 12556 10016
rect 12596 9976 12605 10016
rect 13411 9976 13420 10016
rect 13460 9976 13708 10016
rect 13748 9976 13900 10016
rect 13940 9976 14900 10016
rect 7084 9892 8332 9932
rect 8372 9892 8381 9932
rect 8428 9892 10060 9932
rect 10100 9892 10109 9932
rect 10435 9892 10444 9932
rect 10484 9892 13516 9932
rect 13556 9892 13565 9932
rect 14860 9848 14900 9976
rect 15034 10007 15244 10016
rect 15034 9967 15043 10007
rect 15083 9976 15244 10007
rect 15284 9976 15293 10016
rect 16291 9976 16300 10016
rect 16340 9976 18019 10016
rect 18059 9976 18068 10016
rect 15083 9967 15092 9976
rect 15034 9966 15092 9967
rect 18220 9932 18260 10144
rect 18796 10100 18836 10312
rect 19564 10268 19604 10312
rect 18883 10228 18892 10268
rect 18932 10228 18978 10268
rect 19555 10228 19564 10268
rect 19604 10228 19613 10268
rect 19756 10248 19796 10816
rect 21571 10732 21580 10772
rect 21620 10732 21772 10772
rect 21812 10732 21821 10772
rect 20131 10480 20140 10520
rect 20180 10480 21292 10520
rect 21332 10480 21341 10520
rect 21353 10396 21484 10436
rect 21524 10396 21533 10436
rect 23020 10352 23060 10984
rect 23194 10975 23203 10984
rect 23243 10975 23252 11015
rect 23194 10974 23252 10975
rect 23500 10436 23540 11068
rect 27244 11024 27284 11152
rect 24041 10984 24172 11024
rect 24212 10984 24221 11024
rect 24329 11015 24460 11024
rect 24329 10984 24451 11015
rect 24500 10984 24509 11024
rect 26825 10984 26947 11024
rect 26996 10984 27005 11024
rect 27244 10984 27532 11024
rect 27572 10984 27581 11024
rect 27715 10984 27724 11024
rect 27764 10984 28492 11024
rect 28532 10984 28541 11024
rect 24442 10975 24451 10984
rect 24491 10975 24500 10984
rect 24442 10974 24500 10975
rect 25402 10900 25411 10940
rect 25451 10900 25612 10940
rect 25652 10900 25661 10940
rect 27139 10900 27148 10940
rect 27188 10900 27197 10940
rect 27322 10900 27331 10940
rect 27380 10900 27511 10940
rect 25027 10732 25036 10772
rect 25076 10732 25228 10772
rect 25268 10732 25277 10772
rect 26425 10564 26434 10604
rect 26802 10564 26811 10604
rect 23500 10396 24076 10436
rect 24116 10396 24125 10436
rect 21859 10312 21868 10352
rect 21908 10312 23060 10352
rect 23674 10312 23683 10352
rect 23723 10312 23732 10352
rect 27017 10312 27148 10352
rect 27188 10312 27197 10352
rect 18892 10184 18932 10228
rect 23020 10184 23060 10312
rect 23692 10184 23732 10312
rect 24163 10228 24172 10268
rect 24218 10228 24343 10268
rect 24874 10228 24883 10268
rect 24923 10228 27052 10268
rect 27092 10228 27101 10268
rect 18882 10144 18891 10184
rect 18931 10144 18940 10184
rect 19018 10144 19027 10184
rect 19067 10144 19084 10184
rect 19124 10144 19700 10184
rect 19930 10144 19939 10184
rect 19979 10144 21868 10184
rect 21908 10144 22060 10184
rect 22100 10144 22109 10184
rect 23011 10144 23020 10184
rect 23060 10144 23069 10184
rect 23273 10144 23308 10184
rect 23348 10144 23395 10184
rect 23435 10144 23444 10184
rect 23491 10144 23500 10184
rect 23540 10144 23636 10184
rect 23692 10144 24268 10184
rect 24308 10144 24317 10184
rect 24931 10144 24940 10184
rect 24980 10144 25048 10184
rect 25088 10144 25111 10184
rect 25219 10144 25228 10184
rect 25268 10144 25420 10184
rect 25460 10144 25469 10184
rect 25987 10144 25996 10184
rect 26036 10144 26956 10184
rect 26996 10144 27005 10184
rect 19660 10100 19700 10144
rect 18307 10060 18316 10100
rect 18356 10060 18836 10100
rect 18883 10060 18892 10100
rect 18932 10060 18941 10100
rect 19660 10060 22732 10100
rect 22772 10060 22781 10100
rect 18892 10016 18932 10060
rect 23596 10016 23636 10144
rect 18892 9976 19180 10016
rect 19220 9976 19229 10016
rect 19459 9976 19468 10016
rect 19508 9976 20332 10016
rect 20372 9976 21484 10016
rect 21524 9976 21533 10016
rect 22339 9976 22348 10016
rect 22388 9976 22540 10016
rect 22580 9976 22589 10016
rect 23596 9976 23884 10016
rect 23924 9976 23933 10016
rect 25961 9976 26092 10016
rect 26132 9976 26141 10016
rect 26275 9976 26284 10016
rect 26324 9976 26455 10016
rect 18220 9892 20524 9932
rect 20564 9892 21868 9932
rect 21908 9892 21917 9932
rect 1804 9808 2284 9848
rect 2324 9808 2956 9848
rect 2996 9808 3005 9848
rect 4343 9808 4352 9848
rect 4720 9808 4729 9848
rect 6307 9808 6316 9848
rect 6356 9808 8812 9848
rect 8852 9808 8861 9848
rect 8908 9808 10348 9848
rect 10388 9808 10397 9848
rect 12117 9808 12126 9848
rect 12494 9808 12503 9848
rect 12547 9808 12556 9848
rect 12596 9808 12605 9848
rect 14860 9808 15284 9848
rect 16099 9808 16108 9848
rect 16148 9808 19604 9848
rect 19891 9808 19900 9848
rect 20268 9808 20277 9848
rect 27665 9808 27674 9848
rect 28042 9808 28051 9848
rect 1132 9724 1708 9764
rect 1748 9724 1757 9764
rect 1132 9680 1172 9724
rect 1804 9680 1844 9808
rect 8908 9764 8948 9808
rect 12556 9764 12596 9808
rect 5827 9724 5836 9764
rect 5876 9724 6604 9764
rect 6644 9724 6932 9764
rect 8515 9724 8524 9764
rect 8564 9724 8948 9764
rect 9379 9724 9388 9764
rect 9428 9724 11788 9764
rect 11828 9724 11837 9764
rect 12364 9724 12596 9764
rect 1114 9640 1123 9680
rect 1163 9640 1172 9680
rect 1498 9640 1507 9680
rect 1547 9640 1844 9680
rect 1996 9640 2668 9680
rect 2708 9640 2956 9680
rect 2996 9640 3005 9680
rect 4649 9640 4780 9680
rect 4820 9640 4829 9680
rect 4954 9640 4963 9680
rect 5003 9640 5260 9680
rect 5300 9640 5309 9680
rect 6307 9640 6316 9680
rect 6356 9640 6836 9680
rect 1996 9596 2036 9640
rect 4972 9596 5012 9640
rect 931 9556 940 9596
rect 980 9556 1172 9596
rect 1713 9556 1722 9596
rect 1762 9556 2036 9596
rect 2170 9556 2179 9596
rect 2219 9556 3092 9596
rect 1132 9512 1172 9556
rect 3052 9512 3092 9556
rect 4396 9556 5012 9596
rect 4396 9512 4436 9556
rect 6796 9512 6836 9640
rect 6892 9512 6932 9724
rect 12364 9680 12404 9724
rect 7171 9640 7180 9680
rect 7220 9640 7229 9680
rect 7529 9640 7564 9680
rect 7604 9640 7660 9680
rect 7700 9640 7709 9680
rect 8201 9640 8323 9680
rect 8372 9640 8381 9680
rect 8611 9640 8620 9680
rect 8660 9640 9475 9680
rect 9515 9640 9524 9680
rect 11491 9640 11500 9680
rect 11540 9640 12020 9680
rect 12355 9640 12364 9680
rect 12404 9640 12413 9680
rect 12547 9640 12556 9680
rect 12596 9640 13123 9680
rect 13163 9640 13172 9680
rect 13315 9640 13324 9680
rect 13364 9640 13795 9680
rect 13835 9640 13844 9680
rect 13891 9640 13900 9680
rect 13940 9640 14275 9680
rect 14315 9640 14324 9680
rect 15034 9640 15043 9680
rect 15083 9640 15092 9680
rect 7180 9596 7220 9640
rect 7180 9556 7468 9596
rect 7508 9556 7517 9596
rect 8803 9556 8812 9596
rect 8852 9556 8861 9596
rect 8995 9556 9004 9596
rect 9044 9556 9163 9596
rect 10051 9556 10060 9596
rect 10100 9556 10580 9596
rect 10627 9556 10636 9596
rect 10676 9556 11692 9596
rect 11732 9556 11741 9596
rect 8812 9512 8852 9556
rect 9123 9512 9163 9556
rect 10540 9512 10580 9556
rect 11980 9512 12020 9640
rect 15052 9596 15092 9640
rect 12067 9556 12076 9596
rect 12116 9556 12740 9596
rect 12931 9556 12940 9596
rect 12980 9556 13003 9596
rect 12076 9512 12116 9556
rect 643 9472 652 9512
rect 692 9472 701 9512
rect 835 9472 844 9512
rect 884 9472 940 9512
rect 980 9472 1015 9512
rect 1123 9472 1132 9512
rect 1172 9472 1181 9512
rect 1402 9472 1411 9512
rect 1451 9472 1460 9512
rect 1507 9472 1516 9512
rect 1556 9472 1847 9512
rect 1887 9472 1896 9512
rect 2083 9472 2092 9512
rect 2132 9472 2141 9512
rect 3043 9472 3052 9512
rect 3092 9472 3101 9512
rect 3305 9472 3436 9512
rect 3476 9472 3485 9512
rect 3593 9472 3724 9512
rect 3764 9472 3773 9512
rect 4378 9472 4387 9512
rect 4427 9472 4436 9512
rect 4483 9472 4492 9512
rect 4532 9472 4541 9512
rect 5251 9472 5260 9512
rect 5300 9472 5684 9512
rect 5827 9472 5836 9512
rect 5876 9472 6007 9512
rect 6089 9472 6220 9512
rect 6260 9472 6269 9512
rect 6778 9472 6787 9512
rect 6827 9472 6836 9512
rect 6883 9472 6892 9512
rect 6932 9472 6941 9512
rect 7354 9472 7363 9512
rect 7403 9472 7412 9512
rect 7540 9472 7564 9512
rect 7604 9472 7671 9512
rect 7711 9472 7720 9512
rect 7843 9472 7852 9512
rect 7892 9472 8236 9512
rect 8276 9472 8428 9512
rect 8468 9472 8477 9512
rect 8698 9472 8707 9512
rect 8747 9472 8756 9512
rect 8812 9472 8948 9512
rect 9006 9472 9015 9512
rect 9055 9472 9064 9512
rect 9123 9472 9143 9512
rect 9183 9472 9192 9512
rect 9257 9472 9388 9512
rect 9428 9472 9437 9512
rect 9641 9472 9739 9512
rect 9812 9472 9821 9512
rect 9955 9472 9964 9512
rect 10004 9472 10135 9512
rect 10313 9472 10435 9512
rect 10484 9472 10493 9512
rect 10540 9472 10636 9512
rect 10676 9472 10732 9512
rect 10772 9472 10807 9512
rect 11011 9472 11020 9512
rect 11060 9472 11212 9512
rect 11252 9472 11261 9512
rect 11369 9472 11404 9512
rect 11444 9472 11500 9512
rect 11540 9472 11549 9512
rect 11962 9472 11971 9512
rect 12011 9472 12020 9512
rect 12067 9472 12076 9512
rect 12116 9472 12125 9512
rect 12451 9472 12460 9512
rect 12500 9472 12508 9512
rect 12548 9472 12631 9512
rect 12700 9511 12740 9556
rect 12963 9512 13003 9556
rect 14476 9556 14764 9596
rect 14804 9556 15092 9596
rect 14476 9512 14516 9556
rect 15244 9512 15284 9808
rect 19564 9680 19604 9808
rect 19747 9724 19756 9764
rect 19796 9724 20372 9764
rect 20419 9724 20428 9764
rect 20468 9724 24268 9764
rect 24308 9724 24317 9764
rect 15619 9640 15628 9680
rect 15668 9640 16291 9680
rect 16331 9640 16340 9680
rect 17164 9640 17932 9680
rect 17972 9640 17981 9680
rect 18281 9640 18412 9680
rect 18452 9640 18461 9680
rect 18778 9640 18787 9680
rect 18827 9640 19276 9680
rect 19316 9640 19325 9680
rect 19546 9640 19555 9680
rect 19595 9640 19604 9680
rect 20332 9680 20372 9724
rect 20332 9640 21091 9680
rect 21131 9640 21140 9680
rect 22697 9640 22819 9680
rect 22868 9640 22877 9680
rect 17164 9596 17204 9640
rect 16195 9556 16204 9596
rect 16244 9556 17204 9596
rect 17251 9556 17260 9596
rect 17300 9556 17396 9596
rect 17164 9512 17204 9556
rect 17356 9512 17396 9556
rect 17740 9556 18356 9596
rect 17740 9512 17780 9556
rect 18316 9512 18356 9556
rect 18988 9556 19988 9596
rect 21475 9556 21484 9596
rect 21524 9556 22147 9596
rect 22187 9556 22196 9596
rect 18988 9512 19028 9556
rect 12700 9488 12788 9511
rect 652 9428 692 9472
rect 1420 9428 1460 9472
rect 652 9388 980 9428
rect 1420 9388 1516 9428
rect 1556 9388 1987 9428
rect 2027 9388 2036 9428
rect 787 9220 796 9260
rect 836 9220 884 9260
rect 0 8924 400 8944
rect 0 8884 460 8924
rect 500 8884 509 8924
rect 0 8864 400 8884
rect 844 8756 884 9220
rect 940 9176 980 9388
rect 2092 9344 2132 9472
rect 4492 9428 4532 9472
rect 5644 9428 5684 9472
rect 6796 9428 6836 9472
rect 3331 9388 3340 9428
rect 3380 9388 4204 9428
rect 4244 9388 4532 9428
rect 4867 9388 4876 9428
rect 4916 9388 5164 9428
rect 5210 9388 5219 9428
rect 5644 9388 6124 9428
rect 6164 9388 6173 9428
rect 6749 9388 6796 9428
rect 6836 9388 6845 9428
rect 7372 9344 7412 9472
rect 8716 9428 8756 9472
rect 8716 9388 8812 9428
rect 8852 9388 8861 9428
rect 1708 9304 2132 9344
rect 4666 9304 4675 9344
rect 4715 9304 5356 9344
rect 5396 9304 5405 9344
rect 5539 9304 5548 9344
rect 5588 9304 7276 9344
rect 7316 9304 7412 9344
rect 1708 9260 1748 9304
rect 1699 9220 1708 9260
rect 1748 9220 1757 9260
rect 2371 9220 2380 9260
rect 2420 9220 2429 9260
rect 4051 9220 4060 9260
rect 4100 9220 5068 9260
rect 5108 9220 5117 9260
rect 6953 9220 7075 9260
rect 7124 9220 7133 9260
rect 7913 9220 8044 9260
rect 8084 9220 8093 9260
rect 2380 9176 2420 9220
rect 940 9136 2420 9176
rect 8908 9176 8948 9472
rect 9015 9344 9055 9472
rect 11980 9428 12020 9472
rect 12700 9471 12856 9488
rect 12954 9472 12963 9512
rect 13003 9472 13027 9512
rect 13123 9472 13132 9512
rect 13172 9472 13276 9512
rect 13316 9472 13325 9512
rect 13385 9472 13420 9512
rect 13460 9472 13516 9512
rect 13556 9472 13565 9512
rect 13635 9472 13694 9512
rect 13734 9472 13743 9512
rect 13865 9472 13996 9512
rect 14036 9472 14045 9512
rect 14467 9472 14476 9512
rect 14516 9472 14525 9512
rect 14604 9472 14668 9512
rect 14708 9472 14764 9512
rect 14804 9472 14813 9512
rect 15235 9472 15244 9512
rect 15284 9472 15293 9512
rect 15523 9472 15532 9512
rect 15572 9472 15724 9512
rect 15764 9472 15767 9512
rect 15807 9472 15924 9512
rect 16003 9472 16012 9512
rect 16052 9472 16183 9512
rect 16313 9472 16396 9512
rect 16436 9472 16444 9512
rect 16484 9472 16493 9512
rect 16579 9472 16588 9512
rect 16628 9472 16637 9512
rect 17164 9472 17212 9512
rect 17252 9472 17261 9512
rect 17347 9472 17356 9512
rect 17396 9472 17405 9512
rect 17539 9472 17548 9512
rect 17588 9472 17597 9512
rect 17722 9472 17731 9512
rect 17771 9472 17780 9512
rect 17827 9472 17836 9512
rect 17876 9472 17932 9512
rect 17972 9472 18007 9512
rect 18307 9472 18316 9512
rect 18356 9472 18836 9512
rect 18964 9472 18973 9512
rect 19013 9472 19028 9512
rect 19075 9472 19084 9512
rect 19124 9472 19133 9512
rect 19577 9472 19660 9512
rect 19700 9472 19708 9512
rect 19748 9472 19757 9512
rect 19843 9472 19852 9512
rect 19892 9472 19901 9512
rect 13132 9471 13220 9472
rect 12748 9470 12856 9471
rect 12748 9448 12816 9470
rect 12807 9430 12816 9448
rect 12856 9430 12865 9470
rect 13635 9428 13675 9472
rect 13996 9454 14036 9463
rect 9187 9388 9196 9428
rect 9236 9388 9283 9428
rect 9323 9388 9367 9428
rect 9667 9388 9676 9428
rect 9716 9388 9859 9428
rect 9899 9388 9908 9428
rect 10051 9388 10060 9428
rect 10100 9388 11884 9428
rect 11924 9388 11933 9428
rect 11980 9388 12652 9428
rect 12692 9388 12701 9428
rect 13219 9388 13228 9428
rect 13268 9388 13675 9428
rect 13635 9344 13675 9388
rect 9015 9304 9100 9344
rect 9140 9304 9149 9344
rect 12739 9304 12748 9344
rect 12788 9304 12797 9344
rect 13635 9304 14668 9344
rect 14708 9304 14717 9344
rect 12748 9260 12788 9304
rect 14764 9260 14804 9472
rect 15244 9428 15284 9472
rect 16588 9428 16628 9472
rect 17548 9428 17588 9472
rect 15244 9388 15907 9428
rect 15947 9388 15956 9428
rect 16099 9388 16108 9428
rect 16148 9388 16628 9428
rect 16684 9388 17204 9428
rect 17347 9388 17356 9428
rect 17396 9388 17644 9428
rect 17684 9388 17693 9428
rect 15916 9344 15956 9388
rect 16684 9344 16724 9388
rect 17164 9344 17204 9388
rect 17740 9344 17780 9472
rect 17932 9428 17972 9472
rect 18796 9428 18836 9472
rect 17932 9388 18700 9428
rect 18740 9388 18749 9428
rect 18796 9388 18988 9428
rect 19028 9388 19037 9428
rect 19084 9344 19124 9472
rect 15916 9304 16724 9344
rect 17002 9304 17011 9344
rect 17051 9304 17108 9344
rect 17164 9304 17548 9344
rect 17588 9304 17780 9344
rect 18883 9304 18892 9344
rect 18932 9304 19124 9344
rect 8995 9220 9004 9260
rect 9044 9220 9868 9260
rect 9908 9220 9917 9260
rect 12748 9220 14804 9260
rect 17068 9260 17108 9304
rect 17068 9220 17260 9260
rect 17300 9220 17309 9260
rect 17722 9220 17731 9260
rect 17771 9220 18508 9260
rect 18548 9220 18557 9260
rect 8908 9136 9292 9176
rect 9332 9136 9341 9176
rect 3103 9052 3112 9092
rect 3480 9052 3489 9092
rect 3532 9052 6316 9092
rect 6356 9052 6365 9092
rect 10877 9052 10886 9092
rect 11254 9052 11263 9092
rect 13132 9052 14572 9092
rect 14612 9052 17684 9092
rect 18651 9052 18660 9092
rect 19028 9052 19037 9092
rect 3532 9008 3572 9052
rect 2860 8968 3572 9008
rect 7363 8968 7372 9008
rect 7412 8968 8852 9008
rect 9667 8968 9676 9008
rect 9716 8968 11348 9008
rect 2860 8924 2900 8968
rect 2851 8884 2860 8924
rect 2900 8884 2909 8924
rect 3593 8884 3619 8924
rect 3659 8884 3724 8924
rect 3764 8884 3773 8924
rect 4963 8884 4972 8924
rect 5012 8884 5548 8924
rect 5588 8884 5597 8924
rect 6019 8884 6028 8924
rect 6068 8884 7892 8924
rect 7939 8884 7948 8924
rect 7988 8884 8140 8924
rect 8180 8884 8189 8924
rect 7852 8840 7892 8884
rect 8812 8840 8852 8968
rect 9763 8884 9772 8924
rect 9812 8884 10828 8924
rect 10868 8884 11252 8924
rect 5033 8800 5116 8840
rect 5156 8800 5164 8840
rect 5204 8800 5876 8840
rect 6211 8800 6220 8840
rect 6260 8831 6391 8840
rect 6260 8800 6268 8831
rect 844 8716 940 8756
rect 980 8716 989 8756
rect 2467 8716 2476 8756
rect 2516 8716 2525 8756
rect 4492 8716 4780 8756
rect 4820 8716 4829 8756
rect 4492 8672 4532 8716
rect 163 8632 172 8672
rect 212 8632 500 8672
rect 1306 8632 1315 8672
rect 1355 8632 2956 8672
rect 2996 8632 3005 8672
rect 3052 8632 3580 8672
rect 3620 8632 3629 8672
rect 3715 8632 3724 8672
rect 3764 8632 4204 8672
rect 4244 8632 4253 8672
rect 4483 8632 4492 8672
rect 4532 8632 4541 8672
rect 4675 8632 4684 8672
rect 4724 8632 4780 8672
rect 4820 8632 4855 8672
rect 5059 8632 5068 8672
rect 5108 8632 5251 8672
rect 5291 8632 5300 8672
rect 5347 8632 5356 8672
rect 5396 8632 5527 8672
rect 5609 8632 5644 8672
rect 5684 8632 5731 8672
rect 5771 8632 5789 8672
rect 0 8504 400 8524
rect 460 8504 500 8632
rect 3052 8588 3092 8632
rect 2083 8548 2092 8588
rect 2132 8548 3092 8588
rect 3148 8548 4876 8588
rect 4916 8548 4925 8588
rect 5553 8548 5562 8588
rect 5602 8548 5727 8588
rect 0 8464 500 8504
rect 0 8444 400 8464
rect 3148 8420 3188 8548
rect 3235 8464 3244 8504
rect 3284 8464 3293 8504
rect 748 8380 2572 8420
rect 2612 8380 3188 8420
rect 3244 8420 3284 8464
rect 3244 8380 3724 8420
rect 3764 8380 3773 8420
rect 0 8084 400 8104
rect 0 8044 460 8084
rect 500 8044 509 8084
rect 0 8024 400 8044
rect 748 8000 788 8380
rect 5687 8336 5727 8548
rect 5836 8504 5876 8800
rect 6308 8800 6391 8831
rect 6490 8800 6499 8840
rect 6539 8800 6548 8840
rect 7852 8800 8716 8840
rect 8756 8800 8765 8840
rect 8812 8800 9388 8840
rect 9428 8800 9437 8840
rect 9850 8800 9859 8840
rect 9899 8800 10196 8840
rect 10243 8800 10252 8840
rect 10292 8800 11156 8840
rect 6268 8782 6308 8791
rect 6508 8756 6548 8800
rect 6508 8716 6932 8756
rect 7258 8716 7267 8756
rect 7316 8716 7447 8756
rect 8297 8716 8338 8756
rect 8378 8716 8428 8756
rect 8468 8716 8852 8756
rect 6892 8672 6932 8716
rect 8812 8672 8852 8716
rect 9004 8672 9044 8800
rect 10156 8756 10196 8800
rect 9091 8716 9100 8756
rect 9140 8747 9772 8756
rect 9179 8716 9772 8747
rect 9812 8716 9821 8756
rect 10147 8716 10156 8756
rect 10196 8716 10205 8756
rect 10601 8716 10732 8756
rect 10772 8716 10781 8756
rect 9130 8707 9139 8716
rect 9179 8707 9188 8716
rect 9130 8706 9188 8707
rect 11116 8672 11156 8800
rect 11212 8672 11252 8884
rect 11308 8840 11348 8968
rect 12643 8884 12652 8924
rect 12692 8884 13036 8924
rect 13076 8884 13085 8924
rect 13132 8840 13172 9052
rect 15436 8968 17588 9008
rect 11308 8800 12844 8840
rect 12884 8800 13172 8840
rect 13306 8800 13315 8840
rect 13355 8800 13652 8840
rect 14083 8800 14092 8840
rect 14132 8800 15052 8840
rect 15092 8800 15101 8840
rect 13612 8756 13652 8800
rect 15436 8756 15476 8968
rect 17548 8924 17588 8968
rect 16282 8884 16291 8924
rect 16331 8884 17012 8924
rect 17530 8884 17539 8924
rect 17579 8884 17588 8924
rect 16300 8756 16340 8884
rect 16972 8756 17012 8884
rect 17644 8840 17684 9052
rect 19852 8924 19892 9472
rect 19948 9344 19988 9556
rect 20323 9472 20332 9512
rect 20372 9472 20620 9512
rect 20660 9472 20669 9512
rect 21379 9472 21388 9512
rect 21428 9472 21524 9512
rect 22409 9472 22540 9512
rect 22580 9472 22589 9512
rect 23110 9472 23119 9512
rect 23159 9472 23308 9512
rect 23348 9472 23357 9512
rect 20131 9388 20140 9428
rect 20180 9388 20530 9428
rect 20570 9388 20579 9428
rect 21187 9388 21196 9428
rect 21236 9388 21298 9428
rect 21338 9388 21367 9428
rect 19948 9304 20468 9344
rect 20428 9260 20468 9304
rect 20419 9220 20428 9260
rect 20468 9220 20477 9260
rect 21484 8924 21524 9472
rect 23017 9388 23026 9428
rect 23066 9388 23252 9428
rect 23212 8924 23252 9388
rect 23596 9260 23636 9724
rect 24041 9640 24172 9680
rect 24212 9640 24221 9680
rect 25027 9640 25036 9680
rect 25076 9640 25996 9680
rect 26036 9640 26045 9680
rect 26179 9640 26188 9680
rect 26228 9640 27340 9680
rect 27380 9640 27389 9680
rect 24652 9556 25900 9596
rect 25940 9556 25949 9596
rect 24652 9512 24692 9556
rect 23770 9472 23779 9512
rect 23819 9472 23828 9512
rect 23875 9472 23884 9512
rect 23924 9472 23933 9512
rect 24634 9472 24643 9512
rect 24683 9472 24692 9512
rect 24739 9472 24748 9512
rect 24788 9472 25172 9512
rect 25219 9472 25228 9512
rect 25268 9472 25411 9512
rect 25451 9472 25460 9512
rect 25987 9472 25996 9512
rect 26036 9472 26092 9512
rect 26132 9472 26167 9512
rect 26266 9472 26275 9512
rect 26324 9472 26455 9512
rect 23788 9344 23828 9472
rect 23884 9428 23924 9472
rect 23884 9388 24844 9428
rect 24884 9388 24893 9428
rect 25132 9344 25172 9472
rect 26083 9388 26092 9428
rect 26132 9388 26476 9428
rect 26516 9388 26525 9428
rect 23788 9304 24460 9344
rect 24500 9304 24509 9344
rect 25132 9304 25708 9344
rect 25748 9304 26716 9344
rect 26756 9304 26996 9344
rect 23596 9220 25612 9260
rect 25652 9220 25661 9260
rect 26425 9052 26434 9092
rect 26802 9052 26811 9092
rect 18586 8884 18595 8924
rect 18635 8884 19892 8924
rect 20009 8884 20131 8924
rect 20180 8884 20189 8924
rect 21235 8884 21244 8924
rect 21284 8884 21524 8924
rect 21571 8884 21580 8924
rect 21620 8884 21868 8924
rect 21908 8884 21917 8924
rect 23212 8884 23404 8924
rect 23444 8884 23453 8924
rect 24067 8884 24076 8924
rect 24116 8884 25708 8924
rect 25748 8884 25757 8924
rect 17356 8800 17684 8840
rect 18403 8800 18412 8840
rect 18452 8800 19508 8840
rect 19555 8800 19564 8840
rect 19604 8800 22291 8840
rect 24538 8800 24547 8840
rect 24587 8800 24596 8840
rect 26851 8800 26860 8840
rect 26900 8800 26909 8840
rect 12931 8716 12940 8756
rect 12980 8716 13228 8756
rect 13268 8716 13277 8756
rect 13603 8716 13612 8756
rect 13652 8716 14036 8756
rect 14179 8716 14188 8756
rect 14228 8716 15476 8756
rect 15529 8716 15538 8756
rect 15578 8716 16340 8756
rect 16396 8716 16492 8756
rect 16532 8716 16541 8756
rect 16954 8716 16963 8756
rect 17003 8716 17012 8756
rect 17068 8716 17260 8756
rect 17300 8716 17309 8756
rect 13132 8672 13172 8716
rect 13996 8672 14036 8716
rect 16396 8672 16436 8716
rect 17068 8672 17108 8716
rect 17356 8672 17396 8800
rect 17539 8716 17548 8756
rect 17588 8716 17597 8756
rect 17548 8672 17588 8716
rect 18412 8705 18452 8714
rect 6185 8632 6307 8672
rect 6356 8632 6365 8672
rect 6516 8632 6604 8672
rect 6644 8632 6647 8672
rect 6687 8632 6696 8672
rect 6778 8632 6787 8672
rect 6827 8632 6836 8672
rect 6883 8632 6892 8672
rect 6932 8632 6941 8672
rect 7075 8632 7084 8672
rect 7124 8632 7127 8672
rect 7167 8632 7255 8672
rect 7363 8632 7372 8672
rect 7412 8632 7543 8672
rect 7642 8632 7651 8672
rect 7691 8632 7700 8672
rect 7913 8632 7962 8672
rect 8002 8632 8044 8672
rect 8084 8632 8093 8672
rect 8393 8632 8428 8672
rect 8468 8632 8524 8672
rect 8564 8632 8573 8672
rect 8812 8632 8948 8672
rect 8995 8632 9004 8672
rect 9044 8632 9053 8672
rect 9232 8632 9241 8672
rect 9281 8632 9292 8672
rect 9332 8632 9421 8672
rect 9562 8632 9571 8672
rect 9611 8632 9620 8672
rect 9667 8632 9676 8672
rect 9716 8632 9847 8672
rect 9916 8632 10060 8672
rect 10100 8632 10109 8672
rect 10243 8632 10252 8672
rect 10292 8632 10339 8672
rect 10379 8632 10423 8672
rect 10531 8632 10540 8672
rect 10580 8632 10924 8672
rect 10964 8632 10973 8672
rect 11107 8632 11116 8672
rect 11156 8632 11165 8672
rect 11212 8632 11308 8672
rect 11348 8632 11357 8672
rect 11465 8632 11500 8672
rect 11540 8632 11596 8672
rect 11636 8632 11645 8672
rect 12451 8632 12460 8672
rect 12500 8632 12509 8672
rect 13129 8632 13138 8672
rect 13178 8632 13187 8672
rect 13258 8632 13267 8672
rect 13307 8632 13420 8672
rect 13460 8632 13469 8672
rect 13603 8632 13612 8672
rect 13652 8632 13795 8672
rect 13835 8632 13940 8672
rect 13996 8632 14524 8672
rect 14564 8632 14573 8672
rect 14659 8632 14668 8672
rect 14708 8632 14717 8672
rect 15619 8632 15628 8672
rect 15668 8632 15677 8672
rect 16121 8632 16204 8672
rect 16244 8632 16252 8672
rect 16292 8632 16301 8672
rect 16387 8632 16396 8672
rect 16436 8632 16445 8672
rect 16492 8632 16823 8672
rect 16863 8632 16872 8672
rect 17052 8632 17061 8672
rect 17101 8632 17110 8672
rect 17347 8632 17356 8672
rect 17396 8632 17405 8672
rect 17530 8632 17539 8672
rect 17579 8632 17635 8672
rect 17923 8632 17932 8672
rect 17972 8632 18028 8672
rect 18068 8632 18103 8672
rect 18508 8672 18548 8800
rect 19468 8756 19508 8800
rect 18595 8716 18604 8756
rect 18644 8716 18883 8756
rect 18923 8716 18932 8756
rect 19450 8716 19459 8756
rect 19499 8716 19508 8756
rect 19948 8716 20812 8756
rect 20852 8716 20861 8756
rect 21091 8716 21100 8756
rect 21140 8716 21292 8756
rect 21332 8716 21716 8756
rect 21859 8716 21868 8756
rect 21908 8716 22076 8756
rect 19948 8672 19988 8716
rect 21676 8681 21716 8716
rect 21676 8672 21718 8681
rect 22036 8672 22076 8716
rect 22251 8714 22291 8800
rect 24556 8756 24596 8800
rect 26860 8756 26900 8800
rect 23465 8716 23506 8756
rect 23546 8716 23596 8756
rect 23636 8716 23645 8756
rect 23875 8716 23884 8756
rect 23924 8716 24364 8756
rect 24404 8716 24413 8756
rect 24556 8716 25042 8756
rect 25082 8716 25091 8756
rect 26464 8716 26572 8756
rect 26635 8716 26644 8756
rect 26764 8716 26900 8756
rect 26956 8756 26996 9304
rect 26956 8716 27476 8756
rect 22234 8705 22292 8714
rect 6796 8588 6836 8632
rect 7660 8588 7700 8632
rect 8908 8588 8948 8632
rect 9580 8588 9620 8632
rect 9916 8588 9956 8632
rect 12460 8588 12500 8632
rect 13900 8588 13940 8632
rect 14668 8588 14708 8632
rect 5923 8548 5932 8588
rect 5972 8548 6039 8588
rect 6079 8548 6103 8588
rect 6787 8548 6796 8588
rect 6836 8548 6883 8588
rect 7433 8548 7459 8588
rect 7499 8548 7564 8588
rect 7604 8548 7613 8588
rect 7660 8548 8180 8588
rect 8908 8548 9956 8588
rect 10627 8548 10636 8588
rect 10676 8548 10685 8588
rect 11683 8548 11692 8588
rect 11732 8548 12404 8588
rect 12460 8548 13324 8588
rect 13364 8548 13373 8588
rect 13900 8548 14708 8588
rect 15628 8588 15668 8632
rect 16492 8588 16532 8632
rect 18412 8588 18452 8665
rect 18499 8632 18508 8672
rect 18548 8632 18557 8672
rect 18748 8632 19267 8672
rect 19307 8632 19316 8672
rect 19939 8632 19948 8672
rect 19988 8632 19997 8672
rect 20074 8632 20083 8672
rect 20123 8632 20428 8672
rect 20468 8632 20477 8672
rect 20611 8632 20620 8672
rect 20660 8632 20669 8672
rect 20995 8632 21004 8672
rect 21044 8632 21388 8672
rect 21428 8632 21437 8672
rect 21484 8632 21580 8672
rect 21620 8632 21629 8672
rect 21676 8632 21678 8672
rect 21763 8632 21772 8672
rect 21812 8632 21868 8672
rect 21908 8632 21943 8672
rect 22032 8632 22041 8672
rect 22081 8632 22090 8672
rect 22234 8665 22243 8705
rect 22283 8665 22292 8705
rect 24370 8672 24410 8716
rect 26764 8714 26804 8716
rect 26707 8674 26716 8714
rect 26756 8674 26804 8714
rect 26956 8672 26996 8716
rect 27436 8672 27476 8716
rect 22234 8664 22292 8665
rect 22636 8632 22684 8672
rect 22724 8632 22733 8672
rect 22865 8632 22874 8672
rect 22914 8632 23116 8672
rect 23156 8632 23165 8672
rect 23587 8632 23596 8672
rect 23636 8632 23980 8672
rect 24020 8632 24029 8672
rect 24361 8632 24370 8672
rect 24410 8632 24419 8672
rect 24490 8632 24499 8672
rect 24539 8632 24556 8672
rect 24596 8632 24679 8672
rect 24835 8632 24844 8672
rect 24884 8632 24893 8672
rect 25123 8632 25132 8672
rect 25172 8632 25181 8672
rect 25625 8632 25708 8672
rect 25748 8632 25756 8672
rect 25796 8632 25805 8672
rect 25891 8632 25900 8672
rect 25940 8632 26071 8672
rect 26467 8632 26476 8672
rect 26516 8632 26647 8672
rect 26851 8632 26860 8672
rect 26900 8632 26996 8672
rect 27043 8632 27052 8672
rect 27092 8632 27244 8672
rect 27284 8632 27293 8672
rect 27427 8632 27436 8672
rect 27476 8632 27485 8672
rect 18748 8588 18788 8632
rect 20620 8588 20660 8632
rect 21484 8588 21524 8632
rect 21678 8623 21718 8632
rect 15628 8548 16532 8588
rect 17146 8548 17155 8588
rect 17195 8548 18788 8588
rect 18970 8548 18979 8588
rect 19019 8548 20660 8588
rect 20899 8548 20908 8588
rect 20948 8548 21374 8588
rect 21414 8548 21423 8588
rect 21466 8548 21475 8588
rect 21515 8548 21524 8588
rect 22636 8588 22676 8632
rect 22636 8548 24076 8588
rect 24116 8548 24125 8588
rect 8140 8504 8180 8548
rect 5818 8464 5827 8504
rect 5867 8464 5876 8504
rect 6970 8464 6979 8504
rect 7019 8464 7747 8504
rect 7787 8464 7796 8504
rect 8009 8464 8131 8504
rect 8180 8464 8189 8504
rect 8899 8464 8908 8504
rect 8948 8464 9196 8504
rect 9236 8464 9245 8504
rect 9833 8464 9964 8504
rect 10004 8464 10013 8504
rect 7756 8420 7796 8464
rect 10636 8420 10676 8548
rect 12364 8504 12404 8548
rect 11098 8464 11107 8504
rect 11147 8464 11404 8504
rect 11444 8464 11453 8504
rect 11657 8464 11788 8504
rect 11828 8464 11837 8504
rect 12346 8464 12355 8504
rect 12395 8464 12748 8504
rect 12788 8464 12797 8504
rect 14362 8464 14371 8504
rect 14411 8464 14476 8504
rect 14516 8464 14551 8504
rect 15322 8464 15331 8504
rect 15371 8464 15532 8504
rect 15572 8464 15581 8504
rect 15628 8420 15668 8548
rect 17779 8464 17788 8504
rect 17828 8464 18124 8504
rect 18164 8464 18173 8504
rect 7756 8380 8428 8420
rect 8468 8380 8477 8420
rect 10636 8380 15668 8420
rect 20620 8420 20660 8548
rect 20803 8464 20812 8504
rect 20852 8464 21580 8504
rect 21620 8464 21629 8504
rect 22387 8464 22396 8504
rect 22436 8464 22732 8504
rect 22772 8464 22781 8504
rect 22929 8420 22969 8548
rect 24844 8504 24884 8632
rect 25132 8588 25172 8632
rect 25132 8548 26380 8588
rect 26420 8548 26429 8588
rect 23011 8464 23020 8504
rect 23060 8464 23404 8504
rect 23444 8464 23453 8504
rect 24826 8464 24835 8504
rect 24875 8464 24884 8504
rect 26467 8464 26476 8504
rect 26516 8464 27244 8504
rect 27284 8464 27293 8504
rect 20620 8380 22969 8420
rect 4343 8296 4352 8336
rect 4720 8296 4729 8336
rect 5059 8296 5068 8336
rect 5108 8296 10484 8336
rect 10444 8252 10484 8296
rect 11212 8296 11788 8336
rect 11828 8296 11837 8336
rect 12117 8296 12126 8336
rect 12494 8296 12503 8336
rect 19891 8296 19900 8336
rect 20268 8296 20277 8336
rect 27665 8296 27674 8336
rect 28042 8296 28051 8336
rect 3532 8212 5548 8252
rect 5588 8212 5597 8252
rect 6883 8212 6892 8252
rect 6932 8212 7796 8252
rect 3532 8168 3572 8212
rect 7756 8168 7796 8212
rect 10444 8212 10636 8252
rect 10676 8212 10685 8252
rect 1210 8128 1219 8168
rect 1259 8128 1420 8168
rect 1460 8128 1469 8168
rect 2083 8128 2092 8168
rect 2132 8128 2141 8168
rect 3523 8128 3532 8168
rect 3572 8128 3581 8168
rect 3811 8128 3820 8168
rect 3860 8128 3868 8168
rect 3908 8128 3991 8168
rect 4195 8128 4204 8168
rect 4244 8128 4396 8168
rect 4436 8128 5204 8168
rect 5251 8128 5260 8168
rect 5300 8128 5635 8168
rect 5675 8128 5740 8168
rect 5780 8128 5789 8168
rect 6787 8128 6796 8168
rect 6836 8128 7564 8168
rect 7604 8128 7613 8168
rect 7747 8128 7756 8168
rect 7796 8128 7805 8168
rect 8707 8128 8716 8168
rect 8756 8128 9140 8168
rect 9353 8128 9484 8168
rect 9524 8128 9533 8168
rect 9641 8128 9763 8168
rect 9812 8128 9821 8168
rect 2092 8084 2132 8128
rect 3868 8084 3908 8128
rect 5164 8084 5204 8128
rect 6796 8084 6836 8128
rect 844 8044 940 8084
rect 980 8044 989 8084
rect 1036 8044 1516 8084
rect 1556 8044 2132 8084
rect 2860 8044 3764 8084
rect 3868 8044 4532 8084
rect 4937 8044 5057 8084
rect 5108 8044 5117 8084
rect 5164 8044 5452 8084
rect 5492 8044 5501 8084
rect 5836 8044 6836 8084
rect 844 8000 884 8044
rect 1036 8000 1076 8044
rect 1324 8000 1364 8044
rect 2860 8000 2900 8044
rect 3724 8000 3764 8044
rect 4492 8000 4532 8044
rect 5836 8000 5876 8044
rect 9100 8000 9140 8128
rect 10444 8084 10484 8212
rect 11212 8168 11252 8296
rect 11692 8212 11980 8252
rect 12020 8212 12029 8252
rect 14947 8212 14956 8252
rect 14996 8212 17684 8252
rect 18019 8212 18028 8252
rect 18068 8212 21332 8252
rect 22435 8212 22444 8252
rect 22484 8212 23212 8252
rect 23252 8212 26655 8252
rect 10627 8128 10636 8168
rect 10676 8128 11252 8168
rect 11369 8128 11395 8168
rect 11435 8128 11500 8168
rect 11540 8128 11549 8168
rect 11692 8084 11732 8212
rect 11875 8128 11884 8168
rect 11924 8128 12115 8168
rect 12155 8128 12268 8168
rect 12308 8128 12324 8168
rect 13603 8128 13612 8168
rect 13652 8128 13804 8168
rect 13844 8128 13853 8168
rect 14083 8128 14092 8168
rect 14132 8128 14188 8168
rect 14228 8128 14263 8168
rect 14851 8128 14860 8168
rect 14900 8128 15436 8168
rect 15476 8128 15485 8168
rect 15538 8084 15578 8212
rect 17644 8168 17684 8212
rect 16265 8128 16396 8168
rect 16436 8128 16445 8168
rect 16666 8128 16675 8168
rect 16715 8128 16724 8168
rect 17626 8128 17635 8168
rect 17675 8128 17684 8168
rect 18883 8128 18892 8168
rect 18932 8128 19660 8168
rect 19700 8128 19709 8168
rect 21065 8128 21196 8168
rect 21236 8128 21245 8168
rect 10424 8044 10433 8084
rect 10473 8044 10484 8084
rect 11581 8044 11732 8084
rect 12067 8044 12076 8084
rect 12116 8044 12556 8084
rect 12596 8044 12605 8084
rect 14467 8044 14476 8084
rect 14516 8044 14525 8084
rect 14851 8044 14860 8084
rect 14900 8044 15148 8084
rect 15188 8044 15197 8084
rect 15388 8044 15578 8084
rect 11581 8000 11621 8044
rect 14476 8000 14516 8044
rect 15388 8000 15428 8044
rect 16684 8000 16724 8128
rect 16876 8044 18028 8084
rect 18068 8044 18077 8084
rect 19171 8044 19180 8084
rect 19220 8044 19316 8084
rect 16876 8000 16916 8044
rect 19276 8000 19316 8044
rect 20332 8044 20620 8084
rect 20660 8044 21100 8084
rect 21140 8044 21149 8084
rect 20332 8000 20372 8044
rect 21292 8000 21332 8212
rect 21379 8128 21388 8168
rect 21428 8128 21571 8168
rect 21611 8128 21620 8168
rect 23177 8128 23299 8168
rect 23348 8128 23357 8168
rect 23587 8128 23596 8168
rect 23636 8128 25795 8168
rect 25835 8128 25844 8168
rect 25891 8128 25900 8168
rect 25940 8128 26071 8168
rect 26266 8128 26275 8168
rect 26324 8128 26455 8168
rect 22435 8044 22444 8084
rect 22484 8044 22493 8084
rect 23192 8044 23201 8084
rect 23241 8044 23692 8084
rect 23732 8044 23741 8084
rect 25949 8044 25996 8084
rect 26036 8044 26045 8084
rect 26371 8044 26380 8084
rect 26420 8044 26551 8084
rect 22444 8000 22484 8044
rect 643 7960 652 8000
rect 692 7960 788 8000
rect 835 7960 844 8000
rect 884 7960 893 8000
rect 1027 7960 1036 8000
rect 1076 7960 1085 8000
rect 1181 7960 1227 8000
rect 1267 7960 1276 8000
rect 1324 7960 1403 8000
rect 1443 7960 1452 8000
rect 1603 7960 1612 8000
rect 1652 7960 1804 8000
rect 1844 7960 1853 8000
rect 1961 7960 2092 8000
rect 2132 7960 2141 8000
rect 2275 7960 2284 8000
rect 2324 7960 2611 8000
rect 2651 7960 2660 8000
rect 2797 7960 2806 8000
rect 2846 7960 2900 8000
rect 3130 7960 3139 8000
rect 3179 7960 3188 8000
rect 3235 7960 3244 8000
rect 3284 7960 3293 8000
rect 3593 7991 3724 8000
rect 3593 7960 3715 7991
rect 3764 7960 3773 8000
rect 4483 7960 4492 8000
rect 4532 7960 4541 8000
rect 4603 7960 4612 8000
rect 4652 7960 4684 8000
rect 4724 7960 4792 8000
rect 5225 7960 5356 8000
rect 5396 7960 5405 8000
rect 5827 7960 5836 8000
rect 5876 7960 5885 8000
rect 6019 7960 6028 8000
rect 6068 7960 6124 8000
rect 6164 7960 6199 8000
rect 6307 7960 6316 8000
rect 6356 7960 6487 8000
rect 6595 7960 6604 8000
rect 6644 7960 6653 8000
rect 7354 7960 7363 8000
rect 7403 7960 7948 8000
rect 7988 7960 7997 8000
rect 8131 7960 8140 8000
rect 8180 7960 8323 8000
rect 8363 7960 8372 8000
rect 8419 7960 8428 8000
rect 8468 7960 8599 8000
rect 9082 7960 9091 8000
rect 9131 7960 9140 8000
rect 9187 7960 9196 8000
rect 9236 7960 9245 8000
rect 9833 7960 9964 8000
rect 10004 7960 10013 8000
rect 10121 7960 10252 8000
rect 10292 7960 10301 8000
rect 10601 7960 10636 8000
rect 10676 7991 10772 8000
rect 10676 7960 10732 7991
rect 1228 7916 1268 7960
rect 3148 7916 3188 7960
rect 739 7876 748 7916
rect 788 7876 1172 7916
rect 1219 7876 1228 7916
rect 1268 7876 1277 7916
rect 2179 7876 2188 7916
rect 2228 7876 2237 7916
rect 2755 7876 2764 7916
rect 2804 7876 3188 7916
rect 1132 7832 1172 7876
rect 2188 7832 2228 7876
rect 3244 7832 3284 7960
rect 3706 7951 3715 7960
rect 3755 7951 3764 7960
rect 3706 7950 3764 7951
rect 4282 7918 4291 7958
rect 4331 7918 4341 7958
rect 5356 7942 5396 7951
rect 1132 7792 2228 7832
rect 2563 7792 2572 7832
rect 2612 7792 3284 7832
rect 4301 7832 4341 7918
rect 6604 7916 6644 7960
rect 9196 7916 9236 7960
rect 10819 7960 10828 8000
rect 10868 7960 10871 8000
rect 10911 7960 10999 8000
rect 11107 7960 11116 8000
rect 11156 7960 11444 8000
rect 11572 7960 11581 8000
rect 11621 7960 11630 8000
rect 11683 7960 11692 8000
rect 11732 7960 11863 8000
rect 11971 7960 11980 8000
rect 12020 7960 12259 8000
rect 12299 7960 12308 8000
rect 12355 7960 12364 8000
rect 12404 7960 12535 8000
rect 12739 7960 12748 8000
rect 12788 7960 13132 8000
rect 13172 7960 13181 8000
rect 13315 7960 13324 8000
rect 13364 7960 13420 8000
rect 13460 7960 13495 8000
rect 14249 7960 14284 8000
rect 14324 7960 14380 8000
rect 14420 7960 14429 8000
rect 14476 7960 14515 8000
rect 14555 7960 14564 8000
rect 14648 7960 14657 8000
rect 14708 7960 14828 8000
rect 14947 7960 14956 8000
rect 14996 7960 15127 8000
rect 15370 7991 15428 8000
rect 10732 7942 10772 7951
rect 11404 7916 11444 7960
rect 12364 7942 12404 7951
rect 14956 7942 14996 7951
rect 15235 7918 15244 7958
rect 15284 7918 15293 7958
rect 15370 7951 15379 7991
rect 15419 7951 15428 7991
rect 15472 7960 15481 8000
rect 15521 7960 15532 8000
rect 15572 7960 15661 8000
rect 15994 7960 16003 8000
rect 16043 7960 16052 8000
rect 16099 7960 16108 8000
rect 16148 7960 16724 8000
rect 16867 7960 16876 8000
rect 16916 7960 16925 8000
rect 17155 7960 17164 8000
rect 17204 7960 17356 8000
rect 17396 7960 17405 8000
rect 17609 7960 17740 8000
rect 17780 7960 17789 8000
rect 17993 7960 18124 8000
rect 18164 7960 18173 8000
rect 18490 7960 18499 8000
rect 18539 7960 18548 8000
rect 18595 7960 18604 8000
rect 18644 7960 18775 8000
rect 19075 7960 19084 8000
rect 19124 7960 19133 8000
rect 19258 7960 19267 8000
rect 19307 7960 19768 8000
rect 19808 7960 19817 8000
rect 20314 7960 20323 8000
rect 20363 7960 20372 8000
rect 20419 7960 20428 8000
rect 20468 7960 20477 8000
rect 20777 7960 20908 8000
rect 20948 7960 20957 8000
rect 15370 7950 15428 7951
rect 6211 7876 6220 7916
rect 6260 7888 7316 7916
rect 6260 7876 7315 7888
rect 7276 7848 7315 7876
rect 7355 7848 7364 7888
rect 8803 7876 8812 7916
rect 8852 7876 9236 7916
rect 11002 7876 11011 7916
rect 11051 7876 11156 7916
rect 11203 7876 11212 7916
rect 11252 7876 11261 7916
rect 11404 7876 12076 7916
rect 12116 7876 12125 7916
rect 14410 7907 14764 7916
rect 4301 7792 4780 7832
rect 4820 7792 4829 7832
rect 11116 7748 11156 7876
rect 11212 7832 11252 7876
rect 14410 7867 14419 7907
rect 14459 7876 14764 7907
rect 14804 7876 14813 7916
rect 14459 7867 14468 7876
rect 14410 7866 14468 7867
rect 15244 7832 15284 7918
rect 11212 7792 13612 7832
rect 13652 7792 13661 7832
rect 14668 7792 15284 7832
rect 14668 7748 14708 7792
rect 1507 7708 1516 7748
rect 1556 7708 1565 7748
rect 2057 7708 2188 7748
rect 2228 7708 2237 7748
rect 4771 7708 4780 7748
rect 4820 7708 4829 7748
rect 5050 7708 5059 7748
rect 5099 7708 6220 7748
rect 6260 7708 6269 7748
rect 7546 7708 7555 7748
rect 7595 7708 7660 7748
rect 7700 7708 7735 7748
rect 10426 7708 10435 7748
rect 10475 7708 10484 7748
rect 11116 7708 11500 7748
rect 11540 7708 11549 7748
rect 12643 7708 12652 7748
rect 12692 7708 13900 7748
rect 13940 7708 13949 7748
rect 14650 7708 14659 7748
rect 14699 7708 14708 7748
rect 0 7664 400 7684
rect 1516 7664 1556 7708
rect 4780 7664 4820 7708
rect 10444 7664 10484 7708
rect 0 7624 652 7664
rect 692 7624 701 7664
rect 1516 7624 3724 7664
rect 3764 7624 3773 7664
rect 4780 7624 8908 7664
rect 8948 7624 8957 7664
rect 10444 7624 11692 7664
rect 11732 7624 11741 7664
rect 0 7604 400 7624
rect 3103 7540 3112 7580
rect 3480 7540 3489 7580
rect 10877 7540 10886 7580
rect 11254 7540 11263 7580
rect 652 7456 2380 7496
rect 2420 7456 2429 7496
rect 3244 7456 7180 7496
rect 7220 7456 7229 7496
rect 7756 7456 10252 7496
rect 10292 7456 10301 7496
rect 0 7244 400 7264
rect 652 7244 692 7456
rect 3244 7412 3284 7456
rect 739 7372 748 7412
rect 788 7372 1708 7412
rect 1748 7372 1757 7412
rect 1804 7372 2284 7412
rect 2324 7372 2333 7412
rect 3235 7372 3244 7412
rect 3284 7372 3293 7412
rect 5225 7372 5347 7412
rect 5396 7372 6164 7412
rect 905 7288 1036 7328
rect 1076 7288 1085 7328
rect 0 7204 692 7244
rect 802 7204 844 7244
rect 884 7204 893 7244
rect 940 7204 1228 7244
rect 1268 7204 1277 7244
rect 1507 7204 1516 7244
rect 1556 7204 1565 7244
rect 0 7184 400 7204
rect 844 7160 884 7204
rect 643 7120 652 7160
rect 692 7120 701 7160
rect 840 7120 849 7160
rect 889 7120 898 7160
rect 652 7076 692 7120
rect 940 7076 980 7204
rect 1516 7160 1556 7204
rect 1804 7160 1844 7372
rect 2179 7288 2188 7328
rect 2228 7288 3340 7328
rect 3380 7288 4300 7328
rect 4340 7288 4349 7328
rect 4483 7288 4492 7328
rect 4532 7288 5260 7328
rect 5300 7288 5309 7328
rect 5635 7288 5644 7328
rect 5684 7288 5693 7328
rect 5644 7244 5684 7288
rect 2284 7204 2996 7244
rect 3043 7204 3052 7244
rect 3092 7204 4876 7244
rect 4916 7204 4925 7244
rect 5068 7204 5684 7244
rect 5731 7204 5740 7244
rect 5780 7204 5972 7244
rect 2284 7160 2324 7204
rect 2956 7202 2996 7204
rect 2956 7193 3000 7202
rect 2956 7162 2960 7193
rect 1027 7120 1036 7160
rect 1076 7120 1085 7160
rect 1217 7120 1226 7160
rect 1266 7120 1275 7160
rect 1411 7120 1420 7160
rect 1460 7120 1556 7160
rect 1603 7120 1612 7160
rect 1652 7120 1844 7160
rect 1891 7120 1900 7160
rect 1940 7120 2071 7160
rect 2275 7120 2284 7160
rect 2324 7120 2333 7160
rect 2417 7120 2426 7160
rect 2466 7149 2708 7160
rect 2842 7149 2851 7160
rect 2466 7120 2851 7149
rect 2891 7120 2904 7160
rect 4108 7160 4148 7204
rect 5068 7160 5108 7204
rect 5932 7202 5972 7204
rect 5932 7162 5980 7202
rect 6020 7162 6029 7202
rect 6124 7160 6164 7372
rect 7756 7244 7796 7456
rect 16012 7412 16052 7960
rect 18508 7412 18548 7960
rect 19084 7916 19124 7960
rect 20428 7916 20468 7960
rect 21004 7936 21036 7976
rect 21076 7936 21085 7976
rect 21292 7960 21724 8000
rect 21764 7960 21812 8000
rect 21859 7960 21868 8000
rect 21908 7960 21917 8000
rect 22217 7960 22348 8000
rect 22388 7960 22397 8000
rect 22444 7960 22492 8000
rect 22532 7960 22541 8000
rect 22627 7960 22636 8000
rect 22676 7960 22807 8000
rect 23273 7960 23404 8000
rect 23444 7960 23453 8000
rect 23500 7991 23596 8000
rect 19084 7876 19180 7916
rect 19220 7876 19229 7916
rect 19363 7876 19372 7916
rect 19412 7876 19603 7916
rect 19643 7876 19652 7916
rect 20428 7876 20812 7916
rect 20852 7876 20861 7916
rect 19258 7708 19267 7748
rect 19307 7708 20236 7748
rect 20276 7708 20285 7748
rect 20393 7708 20524 7748
rect 20564 7708 20573 7748
rect 18651 7540 18660 7580
rect 19028 7540 19037 7580
rect 8681 7372 8764 7412
rect 8804 7372 8812 7412
rect 8852 7372 8861 7412
rect 9283 7372 9292 7412
rect 9332 7372 9580 7412
rect 9620 7372 9629 7412
rect 12569 7372 12652 7412
rect 12692 7372 12700 7412
rect 12740 7372 12749 7412
rect 13865 7372 13987 7412
rect 14036 7372 14045 7412
rect 14371 7372 14380 7412
rect 14420 7372 14563 7412
rect 14603 7372 14612 7412
rect 16012 7372 16588 7412
rect 16628 7372 16637 7412
rect 17971 7372 17980 7412
rect 18020 7372 18124 7412
rect 18164 7372 18173 7412
rect 18508 7372 18748 7412
rect 18788 7372 18797 7412
rect 18883 7372 18892 7412
rect 18932 7372 19124 7412
rect 20515 7372 20524 7412
rect 20564 7372 20908 7412
rect 20948 7372 20957 7412
rect 19084 7328 19124 7372
rect 9004 7288 15052 7328
rect 15092 7288 15101 7328
rect 15235 7288 15244 7328
rect 15284 7288 16348 7328
rect 16388 7288 16397 7328
rect 19084 7288 19220 7328
rect 19555 7288 19564 7328
rect 19604 7288 19613 7328
rect 20227 7288 20236 7328
rect 20276 7288 20716 7328
rect 20756 7288 20765 7328
rect 9004 7244 9044 7288
rect 6307 7204 6316 7244
rect 6356 7204 6508 7244
rect 6548 7204 6557 7244
rect 7433 7204 7555 7244
rect 7604 7204 7613 7244
rect 7747 7204 7756 7244
rect 7796 7204 7805 7244
rect 8044 7204 8276 7244
rect 8995 7204 9004 7244
rect 9044 7204 9053 7244
rect 9196 7204 9620 7244
rect 11465 7204 11596 7244
rect 11636 7204 11645 7244
rect 11779 7204 11788 7244
rect 11828 7204 12020 7244
rect 8044 7160 8084 7204
rect 8236 7160 8276 7204
rect 9196 7160 9236 7204
rect 9580 7160 9620 7204
rect 11980 7160 12020 7204
rect 13228 7204 13324 7244
rect 13364 7204 13373 7244
rect 15139 7204 15148 7244
rect 15188 7204 18548 7244
rect 13228 7160 13268 7204
rect 14862 7160 14902 7169
rect 15532 7160 15572 7204
rect 18508 7160 18548 7204
rect 19180 7160 19220 7288
rect 19564 7244 19604 7288
rect 21004 7244 21044 7936
rect 21772 7832 21812 7960
rect 21868 7916 21908 7960
rect 23540 7960 23596 7991
rect 23636 7960 23671 8000
rect 23779 7960 23788 8000
rect 23828 7960 23959 8000
rect 24016 7960 24025 8000
rect 24065 7960 24076 8000
rect 24116 7960 24133 8000
rect 24173 7960 24276 8000
rect 24355 7960 24364 8000
rect 24404 7960 24556 8000
rect 24596 7960 24605 8000
rect 24713 7960 24844 8000
rect 24884 7960 24893 8000
rect 25603 7960 25612 8000
rect 25652 7960 25694 8000
rect 25734 7960 25783 8000
rect 25996 7991 26036 8044
rect 26177 8000 26228 8002
rect 26615 8000 26655 8212
rect 23500 7942 23540 7951
rect 26168 7960 26177 8000
rect 26217 7960 26228 8000
rect 25996 7942 26036 7951
rect 26188 7916 26228 7960
rect 26380 7991 26518 8000
rect 26380 7960 26478 7991
rect 21868 7876 22828 7916
rect 22868 7876 22877 7916
rect 23884 7876 23907 7916
rect 23947 7876 24259 7916
rect 24299 7876 24308 7916
rect 24451 7876 24460 7916
rect 24500 7876 24631 7916
rect 26179 7876 26188 7916
rect 26228 7876 26260 7916
rect 23884 7832 23924 7876
rect 26380 7832 26420 7960
rect 26606 7960 26615 8000
rect 26655 7960 26664 8000
rect 26729 7960 26860 8000
rect 26900 7960 26909 8000
rect 26478 7942 26518 7951
rect 26633 7876 26755 7916
rect 26804 7876 26813 7916
rect 26947 7876 26956 7916
rect 26996 7876 27005 7916
rect 26956 7832 26996 7876
rect 21772 7792 22540 7832
rect 22580 7792 22589 7832
rect 22636 7792 23116 7832
rect 23156 7792 23165 7832
rect 23299 7792 23308 7832
rect 23348 7792 23924 7832
rect 23980 7792 25900 7832
rect 25940 7792 25949 7832
rect 26380 7792 26996 7832
rect 27139 7792 27148 7832
rect 27188 7792 27197 7832
rect 22636 7748 22676 7792
rect 23980 7748 24020 7792
rect 21754 7708 21763 7748
rect 21803 7708 22676 7748
rect 22819 7708 22828 7748
rect 22868 7708 23020 7748
rect 23060 7708 24020 7748
rect 25123 7708 25132 7748
rect 25172 7708 25516 7748
rect 25556 7708 25565 7748
rect 26380 7664 26420 7792
rect 23491 7624 23500 7664
rect 23540 7624 25996 7664
rect 26036 7624 26420 7664
rect 26425 7540 26434 7580
rect 26802 7540 26811 7580
rect 22828 7456 25612 7496
rect 25652 7456 25661 7496
rect 22828 7412 22868 7456
rect 22819 7372 22828 7412
rect 22868 7372 22877 7412
rect 23020 7372 23788 7412
rect 23828 7372 23837 7412
rect 24355 7372 24364 7412
rect 24404 7372 26092 7412
rect 26132 7372 26141 7412
rect 23020 7328 23060 7372
rect 21298 7288 21428 7328
rect 21475 7288 21484 7328
rect 21524 7288 23060 7328
rect 23107 7288 23116 7328
rect 23156 7288 23318 7328
rect 19564 7204 19733 7244
rect 19773 7204 19782 7244
rect 20035 7204 20044 7244
rect 20084 7204 20332 7244
rect 20372 7204 20381 7244
rect 20428 7204 20524 7244
rect 20564 7204 20948 7244
rect 20995 7204 21004 7244
rect 21044 7204 21053 7244
rect 20428 7160 20468 7204
rect 20908 7160 20948 7204
rect 21298 7160 21338 7288
rect 21388 7244 21428 7288
rect 21388 7204 23020 7244
rect 23060 7204 23168 7244
rect 23128 7202 23168 7204
rect 23278 7202 23318 7288
rect 27148 7244 27188 7792
rect 25440 7204 27188 7244
rect 23128 7162 23142 7202
rect 23182 7162 23191 7202
rect 2960 7144 3000 7153
rect 3348 7120 3436 7160
rect 3476 7120 3479 7160
rect 3519 7120 3528 7160
rect 3610 7120 3619 7160
rect 3659 7120 3668 7160
rect 3715 7120 3724 7160
rect 3764 7120 3895 7160
rect 4099 7120 4108 7160
rect 4148 7120 4157 7160
rect 4204 7120 5059 7160
rect 5099 7120 5108 7160
rect 5155 7120 5164 7160
rect 5204 7120 5335 7160
rect 5635 7120 5644 7160
rect 5684 7120 5693 7160
rect 5827 7120 5836 7160
rect 5876 7120 5885 7160
rect 6106 7120 6115 7160
rect 6155 7120 6164 7160
rect 6211 7120 6220 7160
rect 6260 7120 6391 7160
rect 6473 7120 6604 7160
rect 6644 7120 6653 7160
rect 6700 7120 7415 7160
rect 7455 7120 7464 7160
rect 7651 7120 7660 7160
rect 7700 7120 7831 7160
rect 7948 7120 8084 7160
rect 8131 7120 8140 7160
rect 8180 7120 8189 7160
rect 8236 7120 8428 7160
rect 8468 7120 8477 7160
rect 8969 7120 9100 7160
rect 9140 7120 9149 7160
rect 9196 7120 9219 7160
rect 9259 7120 9268 7160
rect 9328 7120 9337 7160
rect 9377 7120 9524 7160
rect 9580 7120 9628 7160
rect 9668 7120 9677 7160
rect 9763 7120 9772 7160
rect 9812 7120 9943 7160
rect 10409 7120 10444 7160
rect 10484 7120 10540 7160
rect 10580 7120 11011 7160
rect 11051 7120 11060 7160
rect 11107 7120 11116 7160
rect 11156 7120 11308 7160
rect 11348 7120 11357 7160
rect 11561 7120 11692 7160
rect 11732 7120 11741 7160
rect 11788 7120 11811 7160
rect 11851 7120 11860 7160
rect 11920 7120 11929 7160
rect 11969 7120 12020 7160
rect 12067 7120 12076 7160
rect 12116 7120 12125 7160
rect 12259 7120 12268 7160
rect 12308 7120 12364 7160
rect 12404 7120 12439 7160
rect 13210 7120 13219 7160
rect 13259 7120 13268 7160
rect 13315 7120 13324 7160
rect 13364 7120 13373 7160
rect 13817 7120 13900 7160
rect 13940 7120 13948 7160
rect 13988 7120 13997 7160
rect 14083 7120 14092 7160
rect 14132 7120 14141 7160
rect 14731 7120 14764 7160
rect 14804 7120 14862 7160
rect 652 7036 980 7076
rect 0 6824 400 6844
rect 1036 6824 1076 7120
rect 1228 7076 1268 7120
rect 1612 7076 1652 7120
rect 2284 7076 2324 7120
rect 2668 7109 2904 7120
rect 1219 7036 1228 7076
rect 1268 7036 1313 7076
rect 1411 7036 1420 7076
rect 1460 7036 1652 7076
rect 2092 7036 2324 7076
rect 2092 6992 2132 7036
rect 2864 6992 2904 7109
rect 3628 7076 3668 7120
rect 4204 7076 4244 7120
rect 5644 7076 5684 7120
rect 3581 7036 3628 7076
rect 3668 7036 3677 7076
rect 3802 7036 3811 7076
rect 3851 7036 4244 7076
rect 4291 7036 4300 7076
rect 4340 7036 5684 7076
rect 5836 7076 5876 7120
rect 6700 7076 6740 7120
rect 7948 7076 7988 7120
rect 5836 7036 5972 7076
rect 6019 7036 6028 7076
rect 6068 7036 6740 7076
rect 7171 7036 7180 7076
rect 7220 7036 7988 7076
rect 5932 6992 5972 7036
rect 1481 6952 1603 6992
rect 1652 6952 1661 6992
rect 1786 6952 1795 6992
rect 1844 6952 1975 6992
rect 2083 6952 2092 6992
rect 2132 6952 2141 6992
rect 2441 6952 2572 6992
rect 2612 6952 2621 6992
rect 2668 6952 2707 6992
rect 2747 6952 2756 6992
rect 2864 6952 3820 6992
rect 3860 6952 3869 6992
rect 3994 6952 4003 6992
rect 4043 6952 4244 6992
rect 4291 6952 4300 6992
rect 4340 6952 4349 6992
rect 5609 6952 5740 6992
rect 5780 6952 5789 6992
rect 5923 6952 5932 6992
rect 5972 6952 6124 6992
rect 6164 6952 6173 6992
rect 6787 6952 6796 6992
rect 6836 6952 7276 6992
rect 7316 6952 7325 6992
rect 2668 6908 2708 6952
rect 2659 6868 2668 6908
rect 2708 6868 2717 6908
rect 0 6784 748 6824
rect 788 6784 797 6824
rect 1036 6784 4012 6824
rect 4052 6784 4061 6824
rect 0 6764 400 6784
rect 4204 6740 4244 6952
rect 4300 6908 4340 6952
rect 4300 6868 5836 6908
rect 5876 6868 5885 6908
rect 4343 6784 4352 6824
rect 4720 6784 4729 6824
rect 1132 6700 1516 6740
rect 1556 6700 1565 6740
rect 2860 6700 3916 6740
rect 3956 6700 3965 6740
rect 4204 6700 4780 6740
rect 4820 6700 4829 6740
rect 1132 6572 1172 6700
rect 1219 6616 1228 6656
rect 1268 6616 1996 6656
rect 2036 6616 2045 6656
rect 2153 6616 2284 6656
rect 2324 6616 2333 6656
rect 1132 6532 1267 6572
rect 1315 6532 1324 6572
rect 1364 6532 1612 6572
rect 1652 6532 1661 6572
rect 1708 6532 2764 6572
rect 2804 6532 2813 6572
rect 1227 6490 1267 6532
rect 1227 6488 1341 6490
rect 1708 6488 1748 6532
rect 2860 6488 2900 6700
rect 3401 6616 3436 6656
rect 3476 6616 3532 6656
rect 3572 6616 3581 6656
rect 6019 6616 6028 6656
rect 6068 6616 6604 6656
rect 6644 6616 6653 6656
rect 6874 6616 6883 6656
rect 6923 6616 7412 6656
rect 2947 6532 2956 6572
rect 2996 6532 6892 6572
rect 6932 6532 6941 6572
rect 4108 6488 4148 6532
rect 7372 6488 7412 6616
rect 7756 6488 7796 7036
rect 8140 6656 8180 7120
rect 9196 7076 9236 7120
rect 8707 7036 8716 7076
rect 8756 7036 9236 7076
rect 9484 7076 9524 7120
rect 9772 7076 9812 7120
rect 11788 7076 11828 7120
rect 12076 7076 12116 7120
rect 13324 7076 13364 7120
rect 14092 7076 14132 7120
rect 14862 7111 14902 7120
rect 14956 7120 15436 7160
rect 15476 7120 15485 7160
rect 15715 7120 15724 7160
rect 15764 7120 15773 7160
rect 15881 7120 16012 7160
rect 16052 7120 16061 7160
rect 16195 7120 16204 7160
rect 16244 7120 16636 7160
rect 16676 7120 16685 7160
rect 16771 7120 16780 7160
rect 16820 7120 16829 7160
rect 17347 7120 17356 7160
rect 17396 7120 17548 7160
rect 17588 7120 17597 7160
rect 17731 7120 17740 7160
rect 17780 7120 17789 7160
rect 17993 7120 18124 7160
rect 18164 7120 18173 7160
rect 18499 7120 18508 7160
rect 18548 7120 18700 7160
rect 18740 7120 18749 7160
rect 18874 7120 18883 7160
rect 18923 7120 18932 7160
rect 9484 7036 9812 7076
rect 10627 7036 10636 7076
rect 10676 7036 11828 7076
rect 11971 7036 11980 7076
rect 12020 7036 12116 7076
rect 13027 7036 13036 7076
rect 13076 7036 13364 7076
rect 13612 7036 14380 7076
rect 14420 7036 14429 7076
rect 14537 7036 14561 7076
rect 14601 7036 14668 7076
rect 14708 7036 14717 7076
rect 13612 6992 13652 7036
rect 14956 6992 14996 7120
rect 15532 7111 15572 7120
rect 15099 7036 15148 7076
rect 15188 7036 15230 7076
rect 15270 7036 15279 7076
rect 15724 6992 15764 7120
rect 16780 7076 16820 7120
rect 10330 6952 10339 6992
rect 10379 6952 10388 6992
rect 10627 6952 10636 6992
rect 10676 6952 10685 6992
rect 11299 6952 11308 6992
rect 11348 6952 11404 6992
rect 11444 6952 11479 6992
rect 12355 6952 12364 6992
rect 12404 6952 12413 6992
rect 13603 6952 13612 6992
rect 13652 6952 13661 6992
rect 14467 6952 14476 6992
rect 14516 6952 14764 6992
rect 14804 6952 14813 6992
rect 14860 6952 14996 6992
rect 15322 6952 15331 6992
rect 15371 6952 15380 6992
rect 15427 6952 15436 6992
rect 15476 6952 15764 6992
rect 16684 7036 16820 7076
rect 17740 7076 17780 7120
rect 18892 7076 18932 7120
rect 17740 7036 18316 7076
rect 18356 7036 18365 7076
rect 18595 7036 18604 7076
rect 18644 7036 18932 7076
rect 18988 7120 19001 7160
rect 19041 7120 19050 7160
rect 19158 7120 19167 7160
rect 19207 7120 19220 7160
rect 19262 7120 19271 7160
rect 19311 7120 19320 7160
rect 19363 7120 19372 7160
rect 19441 7120 19543 7160
rect 19603 7120 19612 7160
rect 19652 7120 19661 7160
rect 19843 7120 19852 7160
rect 19892 7120 19901 7160
rect 20105 7120 20236 7160
rect 20276 7120 20285 7160
rect 20410 7120 20419 7160
rect 20459 7120 20468 7160
rect 20515 7120 20524 7160
rect 20564 7120 20573 7160
rect 20620 7120 20663 7160
rect 20703 7120 20712 7160
rect 20794 7120 20803 7160
rect 20843 7120 20852 7160
rect 20899 7120 20908 7160
rect 20948 7120 20957 7160
rect 21187 7120 21196 7160
rect 21236 7120 21245 7160
rect 21298 7120 21318 7160
rect 21358 7120 21367 7160
rect 21435 7120 21444 7160
rect 21484 7120 22060 7160
rect 22100 7120 22109 7160
rect 22169 7120 22252 7160
rect 22292 7120 22300 7160
rect 22340 7120 22349 7160
rect 22409 7120 22531 7160
rect 22580 7120 22589 7160
rect 22697 7120 22828 7160
rect 22868 7120 22877 7160
rect 23008 7120 23017 7160
rect 23057 7120 23066 7160
rect 23128 7155 23191 7162
rect 23277 7193 23318 7202
rect 23317 7162 23318 7193
rect 23277 7144 23317 7153
rect 24154 7120 24163 7160
rect 24203 7120 24212 7160
rect 26947 7120 26956 7160
rect 26996 7120 27005 7160
rect 10348 6824 10388 6952
rect 10636 6908 10676 6952
rect 12364 6908 12404 6952
rect 14860 6908 14900 6952
rect 10636 6868 12404 6908
rect 14275 6868 14284 6908
rect 14324 6868 14900 6908
rect 15340 6908 15380 6952
rect 16684 6908 16724 7036
rect 18988 6992 19028 7120
rect 19271 7076 19311 7120
rect 19171 7036 19180 7076
rect 19220 7036 19311 7076
rect 19612 7076 19652 7120
rect 19852 7076 19892 7120
rect 19612 7036 19660 7076
rect 19700 7036 19709 7076
rect 19852 7036 20428 7076
rect 20468 7036 20477 7076
rect 17731 6952 17740 6992
rect 17780 6952 18988 6992
rect 19028 6952 19037 6992
rect 19354 6952 19363 6992
rect 19403 6952 19412 6992
rect 19913 6952 19939 6992
rect 19979 6952 20044 6992
rect 20084 6952 20093 6992
rect 15340 6868 16724 6908
rect 19372 6908 19412 6952
rect 20524 6908 20564 7120
rect 20620 7076 20660 7120
rect 20620 7036 20716 7076
rect 20756 7036 20765 7076
rect 20812 6908 20852 7120
rect 21196 7076 21236 7120
rect 23014 7076 23054 7120
rect 21196 7036 23500 7076
rect 23540 7036 23549 7076
rect 23657 7036 23779 7076
rect 23828 7036 23837 7076
rect 21283 6952 21292 6992
rect 21332 6952 21676 6992
rect 21716 6952 21725 6992
rect 22051 6952 22060 6992
rect 22100 6952 22732 6992
rect 22772 6952 22781 6992
rect 23177 6952 23308 6992
rect 23348 6952 23357 6992
rect 24172 6908 24212 7120
rect 24259 7036 24268 7076
rect 24308 7036 26275 7076
rect 26315 7036 26324 7076
rect 26956 6992 26996 7120
rect 26083 6952 26092 6992
rect 26132 6952 26996 6992
rect 19372 6868 20852 6908
rect 23020 6868 24212 6908
rect 23020 6824 23060 6868
rect 9292 6784 10388 6824
rect 12117 6784 12126 6824
rect 12494 6784 12503 6824
rect 16492 6784 19564 6824
rect 19604 6784 19613 6824
rect 19891 6784 19900 6824
rect 20268 6784 20277 6824
rect 22723 6784 22732 6824
rect 22772 6784 23060 6824
rect 27665 6784 27674 6824
rect 28042 6784 28051 6824
rect 8323 6700 8332 6740
rect 8372 6700 8468 6740
rect 8428 6656 8468 6700
rect 9292 6656 9332 6784
rect 10348 6740 10388 6784
rect 16492 6740 16532 6784
rect 10348 6700 11500 6740
rect 11540 6700 11549 6740
rect 13036 6700 16532 6740
rect 18499 6700 18508 6740
rect 18548 6700 18836 6740
rect 7843 6616 7852 6656
rect 7892 6616 8323 6656
rect 8363 6616 8372 6656
rect 8428 6616 8668 6656
rect 8708 6616 8717 6656
rect 9139 6616 9148 6656
rect 9188 6616 9332 6656
rect 9466 6616 9475 6656
rect 9515 6616 9772 6656
rect 9812 6616 9821 6656
rect 10121 6616 10243 6656
rect 10292 6616 10301 6656
rect 10531 6616 10540 6656
rect 10580 6616 10732 6656
rect 10772 6616 10781 6656
rect 7843 6532 7852 6572
rect 7892 6532 8372 6572
rect 8419 6532 8428 6572
rect 8468 6532 10484 6572
rect 8332 6488 8372 6532
rect 10444 6488 10484 6532
rect 11500 6488 11540 6700
rect 13036 6656 13076 6700
rect 11849 6616 11980 6656
rect 12020 6616 12029 6656
rect 12329 6616 12451 6656
rect 12500 6616 12509 6656
rect 13018 6616 13027 6656
rect 13067 6616 13076 6656
rect 13123 6616 13132 6656
rect 13172 6616 13507 6656
rect 13547 6616 14228 6656
rect 14659 6616 14668 6656
rect 14708 6616 14764 6656
rect 14804 6616 14839 6656
rect 15017 6616 15148 6656
rect 15188 6616 15197 6656
rect 16073 6616 16108 6656
rect 16148 6616 16204 6656
rect 16244 6616 16253 6656
rect 12556 6532 13748 6572
rect 12556 6488 12596 6532
rect 13708 6488 13748 6532
rect 14188 6488 14228 6616
rect 14371 6532 14380 6572
rect 14420 6532 15284 6572
rect 15244 6488 15284 6532
rect 16492 6488 16532 6700
rect 18796 6656 18836 6700
rect 19372 6700 19660 6740
rect 19700 6700 19709 6740
rect 19372 6656 19412 6700
rect 16666 6616 16675 6656
rect 16715 6616 16780 6656
rect 16820 6616 16855 6656
rect 16979 6616 17443 6656
rect 17483 6616 17492 6656
rect 17539 6616 17548 6656
rect 17588 6616 18211 6656
rect 18251 6616 18260 6656
rect 18473 6616 18508 6656
rect 18548 6616 18604 6656
rect 18644 6616 18653 6656
rect 18778 6616 18787 6656
rect 18827 6616 18836 6656
rect 18883 6616 18892 6656
rect 18932 6616 19063 6656
rect 19363 6616 19372 6656
rect 19412 6616 19421 6656
rect 19468 6616 20620 6656
rect 20660 6616 21388 6656
rect 21428 6616 21437 6656
rect 22243 6616 22252 6656
rect 22292 6616 22636 6656
rect 22676 6616 22685 6656
rect 23194 6616 23203 6656
rect 23243 6616 23596 6656
rect 23636 6616 23645 6656
rect 23779 6616 23788 6656
rect 23828 6616 24268 6656
rect 24308 6616 24317 6656
rect 16979 6498 17019 6616
rect 18604 6572 18644 6616
rect 18604 6532 18686 6572
rect 18726 6532 18735 6572
rect 1123 6448 1132 6488
rect 1172 6448 1181 6488
rect 1227 6450 1315 6488
rect 1301 6448 1315 6450
rect 1355 6448 1364 6488
rect 1514 6448 1523 6488
rect 1563 6448 1572 6488
rect 1690 6448 1699 6488
rect 1739 6448 1748 6488
rect 2057 6448 2188 6488
rect 2228 6448 2237 6488
rect 2362 6448 2371 6488
rect 2411 6448 2900 6488
rect 2947 6448 2956 6488
rect 2996 6448 3005 6488
rect 3209 6448 3340 6488
rect 3380 6448 3389 6488
rect 4090 6448 4099 6488
rect 4139 6448 4148 6488
rect 4195 6448 4204 6488
rect 4244 6448 6547 6488
rect 6587 6448 6596 6488
rect 6733 6448 6742 6488
rect 6782 6448 6796 6488
rect 6836 6448 6922 6488
rect 6979 6448 6988 6488
rect 7028 6448 7037 6488
rect 7241 6448 7372 6488
rect 7412 6448 7421 6488
rect 7651 6448 7660 6488
rect 7700 6448 7709 6488
rect 7756 6448 8227 6488
rect 8267 6448 8276 6488
rect 8332 6448 8535 6488
rect 8575 6448 8584 6488
rect 8803 6448 8812 6488
rect 8852 6448 8861 6488
rect 8986 6479 9004 6488
rect 0 6404 400 6424
rect 1132 6404 1172 6448
rect 0 6364 556 6404
rect 596 6364 605 6404
rect 1132 6364 1420 6404
rect 1460 6364 1469 6404
rect 0 6344 400 6364
rect 1516 6320 1556 6448
rect 2956 6404 2996 6448
rect 6988 6404 7028 6448
rect 7660 6404 7700 6448
rect 8812 6404 8852 6448
rect 8986 6439 8995 6479
rect 9044 6448 9175 6488
rect 9292 6448 9580 6488
rect 9620 6448 9628 6488
rect 9668 6448 9677 6488
rect 9763 6448 9772 6488
rect 9812 6448 9821 6488
rect 10051 6448 10060 6488
rect 10100 6448 10348 6488
rect 10388 6448 10397 6488
rect 10444 6448 10876 6488
rect 10916 6448 10964 6488
rect 11011 6448 11020 6488
rect 11060 6448 11308 6488
rect 11348 6448 11357 6488
rect 11491 6448 11500 6488
rect 11540 6448 11549 6488
rect 11779 6448 11788 6488
rect 11828 6448 11837 6488
rect 12547 6448 12556 6488
rect 12596 6448 12605 6488
rect 12920 6448 12929 6488
rect 12969 6448 12980 6488
rect 13123 6448 13132 6488
rect 13172 6479 13303 6488
rect 13172 6448 13228 6479
rect 9035 6439 9044 6448
rect 8986 6438 9044 6439
rect 1795 6364 1804 6404
rect 1844 6364 2996 6404
rect 3593 6364 3724 6404
rect 3764 6364 3773 6404
rect 4675 6364 4684 6404
rect 4724 6364 4733 6404
rect 6988 6364 7892 6404
rect 8515 6364 8524 6404
rect 8564 6364 8852 6404
rect 7852 6320 7892 6364
rect 9292 6320 9332 6448
rect 9772 6404 9812 6448
rect 10924 6404 10964 6448
rect 9641 6364 9772 6404
rect 9812 6364 10828 6404
rect 10868 6364 10877 6404
rect 10924 6364 11596 6404
rect 11636 6364 11645 6404
rect 11788 6320 11828 6448
rect 12940 6320 12980 6448
rect 13268 6448 13303 6479
rect 13577 6448 13708 6488
rect 13748 6448 13757 6488
rect 13865 6448 13996 6488
rect 14036 6448 14045 6488
rect 14179 6448 14188 6488
rect 14228 6448 14237 6488
rect 14467 6448 14476 6488
rect 14516 6448 14525 6488
rect 14572 6448 14947 6488
rect 14987 6448 14996 6488
rect 15235 6448 15244 6488
rect 15284 6448 15293 6488
rect 15497 6448 15628 6488
rect 15668 6448 15677 6488
rect 15881 6448 16012 6488
rect 16052 6448 16061 6488
rect 16492 6448 16828 6488
rect 16868 6448 16877 6488
rect 16961 6458 16970 6498
rect 17010 6458 17019 6498
rect 19468 6488 19508 6616
rect 20035 6532 20044 6572
rect 20084 6532 20323 6572
rect 20363 6532 20372 6572
rect 17731 6448 17740 6488
rect 17780 6448 18124 6488
rect 18164 6448 18173 6488
rect 18307 6448 18316 6488
rect 18356 6448 18487 6488
rect 18857 6448 18988 6488
rect 19028 6448 19037 6488
rect 19116 6448 19180 6488
rect 19220 6448 19276 6488
rect 19316 6448 19325 6488
rect 19450 6448 19459 6488
rect 19499 6448 19604 6488
rect 19834 6448 19843 6488
rect 19883 6448 19892 6488
rect 20009 6448 20140 6488
rect 20180 6448 20189 6488
rect 20698 6448 20707 6488
rect 20756 6448 20887 6488
rect 23177 6448 23308 6488
rect 23348 6448 23357 6488
rect 23596 6448 23644 6488
rect 23684 6448 23693 6488
rect 23753 6448 23884 6488
rect 23924 6448 23933 6488
rect 24067 6448 24076 6488
rect 24116 6448 24268 6488
rect 24308 6448 24317 6488
rect 24809 6448 24940 6488
rect 24980 6448 24989 6488
rect 25673 6448 25804 6488
rect 25844 6448 25853 6488
rect 13228 6404 13268 6439
rect 14476 6404 14516 6448
rect 13228 6364 14516 6404
rect 14572 6320 14612 6448
rect 1027 6280 1036 6320
rect 1076 6280 2188 6320
rect 2228 6280 2237 6320
rect 2441 6280 2476 6320
rect 2516 6280 2572 6320
rect 2612 6280 2621 6320
rect 7171 6280 7180 6320
rect 7220 6280 7756 6320
rect 7796 6280 7805 6320
rect 7852 6280 9332 6320
rect 10531 6280 10540 6320
rect 10580 6280 11788 6320
rect 11828 6280 11837 6320
rect 12739 6280 12748 6320
rect 12788 6280 12980 6320
rect 13891 6280 13900 6320
rect 13940 6280 14612 6320
rect 16012 6320 16052 6448
rect 18988 6430 19028 6439
rect 19276 6404 19316 6448
rect 17641 6364 17650 6404
rect 17690 6364 17699 6404
rect 19276 6364 19468 6404
rect 19508 6364 19517 6404
rect 17650 6320 17690 6364
rect 19564 6320 19604 6448
rect 16012 6280 19604 6320
rect 19852 6236 19892 6448
rect 23596 6404 23636 6448
rect 21571 6364 21580 6404
rect 21620 6364 21629 6404
rect 22243 6364 22252 6404
rect 22292 6364 22828 6404
rect 22868 6364 22877 6404
rect 23596 6364 25123 6404
rect 25163 6364 25172 6404
rect 24643 6280 24652 6320
rect 24692 6280 25996 6320
rect 26036 6280 26045 6320
rect 5635 6196 5644 6236
rect 5684 6196 5693 6236
rect 5897 6196 6028 6236
rect 6068 6196 6077 6236
rect 10627 6196 10636 6236
rect 10676 6196 10828 6236
rect 10868 6196 10877 6236
rect 19852 6196 20620 6236
rect 20660 6196 20669 6236
rect 20803 6196 20812 6236
rect 20852 6196 22636 6236
rect 22676 6196 22685 6236
rect 23875 6196 23884 6236
rect 23924 6196 24844 6236
rect 24884 6196 24893 6236
rect 5644 6152 5684 6196
rect 5644 6112 5932 6152
rect 5972 6112 8524 6152
rect 8564 6112 8573 6152
rect 18307 6112 18316 6152
rect 18356 6112 25324 6152
rect 25364 6112 25373 6152
rect 3103 6028 3112 6068
rect 3480 6028 3489 6068
rect 10877 6028 10886 6068
rect 11254 6028 11263 6068
rect 18651 6028 18660 6068
rect 19028 6028 19037 6068
rect 26425 6028 26434 6068
rect 26802 6028 26811 6068
rect 0 5984 400 6004
rect 0 5944 19372 5984
rect 19412 5944 19421 5984
rect 20419 5944 20428 5984
rect 20468 5944 21196 5984
rect 21236 5944 21245 5984
rect 0 5924 400 5944
rect 3523 5860 3532 5900
rect 3572 5860 3724 5900
rect 3764 5860 3773 5900
rect 4156 5860 4876 5900
rect 4916 5860 4925 5900
rect 7939 5860 7948 5900
rect 7988 5860 8428 5900
rect 8468 5860 8477 5900
rect 8803 5860 8812 5900
rect 8852 5860 9004 5900
rect 9044 5860 9053 5900
rect 11491 5860 11500 5900
rect 11540 5860 12172 5900
rect 12212 5860 12844 5900
rect 12884 5860 12893 5900
rect 13027 5860 13036 5900
rect 13076 5860 14284 5900
rect 14324 5860 14333 5900
rect 15331 5860 15340 5900
rect 15380 5860 15724 5900
rect 15764 5860 15773 5900
rect 16963 5860 16972 5900
rect 17012 5860 18124 5900
rect 18164 5860 18173 5900
rect 20131 5860 20140 5900
rect 20180 5860 20332 5900
rect 20372 5860 20381 5900
rect 20611 5860 20620 5900
rect 20660 5860 21484 5900
rect 21524 5860 21533 5900
rect 22627 5860 22636 5900
rect 22676 5860 24172 5900
rect 24212 5860 24268 5900
rect 24308 5860 24343 5900
rect 24931 5860 24940 5900
rect 24980 5860 25132 5900
rect 25172 5860 25181 5900
rect 3785 5776 3820 5816
rect 3860 5776 3916 5816
rect 3956 5776 3965 5816
rect 4156 5807 4196 5860
rect 4553 5776 4684 5816
rect 4724 5776 4733 5816
rect 5356 5776 6220 5816
rect 6260 5776 6269 5816
rect 12547 5776 12556 5816
rect 12596 5776 12605 5816
rect 17225 5776 17356 5816
rect 17396 5776 17405 5816
rect 21833 5776 21868 5816
rect 21908 5776 21964 5816
rect 22004 5776 22013 5816
rect 24643 5776 24652 5816
rect 24692 5776 25804 5816
rect 25844 5776 25853 5816
rect 4156 5758 4196 5767
rect 5356 5732 5396 5776
rect 12556 5732 12596 5776
rect 5347 5692 5356 5732
rect 5396 5692 5405 5732
rect 7555 5692 7564 5732
rect 7604 5692 7613 5732
rect 11203 5692 11212 5732
rect 11252 5692 11261 5732
rect 12556 5692 12940 5732
rect 12980 5692 12989 5732
rect 15043 5692 15052 5732
rect 15092 5692 15101 5732
rect 15619 5692 15628 5732
rect 15668 5692 16435 5732
rect 16475 5692 17548 5732
rect 17588 5692 17597 5732
rect 18211 5692 18220 5732
rect 18260 5692 18269 5732
rect 19180 5692 20716 5732
rect 20756 5692 22484 5732
rect 5836 5648 5876 5657
rect 3401 5608 3532 5648
rect 3572 5608 3581 5648
rect 3715 5608 3724 5648
rect 3764 5608 3773 5648
rect 4073 5608 4099 5648
rect 4139 5608 4204 5648
rect 4244 5608 4253 5648
rect 4771 5608 4780 5648
rect 4820 5608 5035 5648
rect 5075 5608 5097 5648
rect 5146 5608 5155 5648
rect 5195 5608 5204 5648
rect 5251 5608 5260 5648
rect 5300 5608 5684 5648
rect 5731 5608 5740 5648
rect 5780 5608 5836 5648
rect 5876 5608 5911 5648
rect 6007 5608 6016 5648
rect 6068 5608 6196 5648
rect 6874 5608 6883 5648
rect 6932 5608 8236 5648
rect 8276 5608 8285 5648
rect 8995 5608 9004 5648
rect 9044 5608 9196 5648
rect 9236 5608 9245 5648
rect 9292 5643 10388 5648
rect 10540 5643 10627 5648
rect 9292 5608 10627 5643
rect 10667 5608 10676 5648
rect 12940 5608 13036 5648
rect 13076 5608 13085 5648
rect 13171 5608 13180 5648
rect 13220 5608 13228 5648
rect 13268 5608 13351 5648
rect 14170 5608 14179 5648
rect 14219 5608 15916 5648
rect 15956 5608 15965 5648
rect 16621 5608 16630 5648
rect 16670 5608 16820 5648
rect 18874 5608 18883 5648
rect 18923 5643 19028 5648
rect 19180 5643 19220 5692
rect 18923 5608 19220 5643
rect 19337 5608 19468 5648
rect 19508 5608 19517 5648
rect 20323 5608 20332 5648
rect 20372 5608 21004 5648
rect 21044 5608 21053 5648
rect 21178 5608 21187 5648
rect 21227 5608 21236 5648
rect 21283 5608 21292 5648
rect 21332 5608 21463 5648
rect 22444 5643 22484 5692
rect 23980 5648 24020 5712
rect 22636 5643 22723 5648
rect 22444 5608 22723 5643
rect 22772 5608 22903 5648
rect 23980 5608 24652 5648
rect 24692 5608 24701 5648
rect 24826 5608 24835 5648
rect 24875 5608 24884 5648
rect 25001 5608 25132 5648
rect 25172 5608 25181 5648
rect 3724 5564 3764 5608
rect 3724 5524 4108 5564
rect 4148 5524 4157 5564
rect 5057 5312 5097 5608
rect 5164 5564 5204 5608
rect 5644 5564 5684 5608
rect 5836 5599 5876 5608
rect 8236 5564 8276 5608
rect 9292 5564 9332 5608
rect 10348 5603 10580 5608
rect 5164 5524 5276 5564
rect 5403 5524 5452 5564
rect 5492 5524 5534 5564
rect 5574 5524 5583 5564
rect 5626 5524 5635 5564
rect 5675 5524 5684 5564
rect 6377 5524 6499 5564
rect 6548 5524 6557 5564
rect 8236 5524 9332 5564
rect 9388 5524 10060 5564
rect 10100 5524 10109 5564
rect 10234 5524 10243 5564
rect 10283 5524 10292 5564
rect 12713 5524 12835 5564
rect 12884 5524 12893 5564
rect 5236 5396 5276 5524
rect 9388 5480 9428 5524
rect 5731 5440 5740 5480
rect 5780 5440 5972 5480
rect 6163 5440 6172 5480
rect 6212 5440 9428 5480
rect 9859 5440 9868 5480
rect 9908 5440 9917 5480
rect 5932 5396 5972 5440
rect 5236 5356 5740 5396
rect 5780 5356 5789 5396
rect 5932 5356 7372 5396
rect 7412 5356 7421 5396
rect 5932 5312 5972 5356
rect 4343 5272 4352 5312
rect 4720 5272 4729 5312
rect 5057 5272 5972 5312
rect 4099 5188 4108 5228
rect 4148 5188 5452 5228
rect 5492 5188 5501 5228
rect 5452 4892 5492 5188
rect 6355 5104 6364 5144
rect 6404 5104 6508 5144
rect 6548 5104 6557 5144
rect 7363 5104 7372 5144
rect 7412 5104 9139 5144
rect 9179 5104 9188 5144
rect 9868 5060 9908 5440
rect 10252 5144 10292 5524
rect 12117 5272 12126 5312
rect 12494 5272 12503 5312
rect 12940 5228 12980 5608
rect 13027 5524 13036 5564
rect 13076 5524 13795 5564
rect 13835 5524 13844 5564
rect 16108 5524 16492 5564
rect 16532 5524 16541 5564
rect 16108 5480 16148 5524
rect 13123 5440 13132 5480
rect 13172 5440 13996 5480
rect 14036 5440 14045 5480
rect 16099 5440 16108 5480
rect 16148 5440 16157 5480
rect 10339 5188 10348 5228
rect 10388 5188 13268 5228
rect 10051 5104 10060 5144
rect 10100 5104 10109 5144
rect 10252 5104 10828 5144
rect 10868 5104 10877 5144
rect 11770 5104 11779 5144
rect 11819 5104 13132 5144
rect 13172 5104 13181 5144
rect 9484 5020 9908 5060
rect 10060 5060 10100 5104
rect 13228 5060 13268 5188
rect 13516 5144 13556 5440
rect 16780 5144 16820 5608
rect 18988 5603 19220 5608
rect 19258 5524 19267 5564
rect 19316 5524 19447 5564
rect 20131 5524 20140 5564
rect 20180 5524 20908 5564
rect 20948 5524 20957 5564
rect 21196 5480 21236 5608
rect 22444 5603 22676 5608
rect 20419 5440 20428 5480
rect 20468 5440 21236 5480
rect 21484 5524 21495 5564
rect 21535 5524 21544 5564
rect 22330 5524 22339 5564
rect 22379 5524 22388 5564
rect 21484 5396 21524 5524
rect 22348 5480 22388 5524
rect 22348 5440 23636 5480
rect 20995 5356 21004 5396
rect 21044 5356 23060 5396
rect 23020 5312 23060 5356
rect 19891 5272 19900 5312
rect 20268 5272 20277 5312
rect 23020 5272 23540 5312
rect 20716 5188 22828 5228
rect 22868 5188 23308 5228
rect 23348 5188 23357 5228
rect 20716 5144 20756 5188
rect 13516 5104 13610 5144
rect 13786 5104 13795 5144
rect 13844 5104 13975 5144
rect 16780 5104 16972 5144
rect 17012 5104 17021 5144
rect 19459 5104 19468 5144
rect 19508 5104 20372 5144
rect 20707 5104 20716 5144
rect 20756 5104 20765 5144
rect 21065 5104 21196 5144
rect 21236 5104 21245 5144
rect 22339 5104 22348 5144
rect 22388 5104 23444 5144
rect 10060 5020 10772 5060
rect 9484 4976 9524 5020
rect 10732 4976 10772 5020
rect 10828 5020 11500 5060
rect 11540 5020 11549 5060
rect 11692 5020 12076 5060
rect 12116 5020 12125 5060
rect 12835 5020 12844 5060
rect 12884 5020 13076 5060
rect 6089 4936 6220 4976
rect 6260 4936 6269 4976
rect 9325 4936 9334 4976
rect 9374 4936 9524 4976
rect 9658 4936 9667 4976
rect 9707 4936 9716 4976
rect 9763 4936 9772 4976
rect 9812 4936 9943 4976
rect 10060 4936 10348 4976
rect 10388 4936 10397 4976
rect 10531 4936 10540 4976
rect 10580 4936 10589 4976
rect 10723 4936 10732 4976
rect 10772 4936 10781 4976
rect 9676 4892 9716 4936
rect 10060 4892 10100 4936
rect 10540 4892 10580 4936
rect 10828 4892 10868 5020
rect 11692 4976 11732 5020
rect 13036 4976 13076 5020
rect 13228 5020 13420 5060
rect 13460 5020 13469 5060
rect 13228 4976 13268 5020
rect 13570 5018 13610 5104
rect 20332 5060 20372 5104
rect 13769 5020 13900 5060
rect 13940 5020 13949 5060
rect 16003 5020 16012 5060
rect 16052 5020 16300 5060
rect 16340 5020 16349 5060
rect 19660 5020 20276 5060
rect 20332 5020 21236 5060
rect 22627 5020 22636 5060
rect 22676 5020 23054 5060
rect 23165 5020 23212 5060
rect 23252 5020 23261 5060
rect 13516 4978 13610 5018
rect 13516 4976 13556 4978
rect 19660 4976 19700 5020
rect 20236 4976 20276 5020
rect 21196 4976 21236 5020
rect 23014 4976 23054 5020
rect 23212 4976 23252 5020
rect 23404 4976 23444 5104
rect 23500 5060 23540 5272
rect 23596 5144 23636 5440
rect 24844 5144 24884 5608
rect 27665 5272 27674 5312
rect 28042 5272 28051 5312
rect 23587 5104 23596 5144
rect 23636 5104 23645 5144
rect 23962 5104 23971 5144
rect 24011 5104 24884 5144
rect 23500 5020 23870 5060
rect 23910 5020 23919 5060
rect 24067 5020 24076 5060
rect 24116 5020 24268 5060
rect 24308 5020 24317 5060
rect 23692 4976 23732 5020
rect 10915 4936 10924 4976
rect 10964 4936 10973 4976
rect 11299 4936 11308 4976
rect 11348 4936 11447 4976
rect 11487 4936 11496 4976
rect 11683 4936 11692 4976
rect 11732 4936 11741 4976
rect 11849 4936 11980 4976
rect 12020 4936 12029 4976
rect 12163 4936 12172 4976
rect 12212 4936 12221 4976
rect 12739 4936 12748 4976
rect 12788 4936 12797 4976
rect 12922 4936 12931 4976
rect 12971 4936 12980 4976
rect 13027 4936 13036 4976
rect 13076 4936 13085 4976
rect 13219 4936 13228 4976
rect 13268 4936 13277 4976
rect 13324 4936 13350 4976
rect 13390 4936 13399 4976
rect 13468 4936 13477 4976
rect 13517 4936 13556 4976
rect 13690 4936 13699 4976
rect 13748 4936 13879 4976
rect 13987 4936 13996 4976
rect 14047 4936 14167 4976
rect 14227 4936 14236 4976
rect 14276 4936 14284 4976
rect 14324 4936 14407 4976
rect 14851 4936 14860 4976
rect 14900 4936 15619 4976
rect 15659 4936 15668 4976
rect 16291 4936 16300 4976
rect 16340 4936 16492 4976
rect 16532 4936 16541 4976
rect 17347 4936 17356 4976
rect 17396 4936 19084 4976
rect 19124 4936 19133 4976
rect 19258 4936 19267 4976
rect 19307 4936 19651 4976
rect 19691 4936 19700 4976
rect 19747 4936 19756 4976
rect 19796 4936 19805 4976
rect 20227 4936 20236 4976
rect 20276 4936 20285 4976
rect 20396 4936 20405 4976
rect 20445 4936 20468 4976
rect 20515 4936 20524 4976
rect 20564 4936 20695 4976
rect 20899 4936 20908 4976
rect 20948 4936 21004 4976
rect 21044 4936 21079 4976
rect 21187 4936 21196 4976
rect 21236 4936 21245 4976
rect 21379 4936 21388 4976
rect 21428 4936 21559 4976
rect 22505 4936 22636 4976
rect 22676 4936 22685 4976
rect 22810 4936 22819 4976
rect 22859 4936 22868 4976
rect 23011 4936 23020 4976
rect 23060 4936 23069 4976
rect 23194 4936 23203 4976
rect 23243 4936 23252 4976
rect 23305 4936 23314 4976
rect 23354 4936 23444 4976
rect 23506 4936 23515 4976
rect 23555 4936 23636 4976
rect 23683 4936 23692 4976
rect 23732 4936 23741 4976
rect 24172 4967 24212 4976
rect 5452 4852 8852 4892
rect 8899 4852 8908 4892
rect 8948 4852 10100 4892
rect 10243 4852 10252 4892
rect 10292 4852 10444 4892
rect 10484 4852 10493 4892
rect 10540 4852 10868 4892
rect 10924 4892 10964 4936
rect 12172 4892 12212 4936
rect 10924 4852 11348 4892
rect 11465 4852 11587 4892
rect 11636 4852 11645 4892
rect 11779 4852 11788 4892
rect 11828 4852 12212 4892
rect 8812 4808 8852 4852
rect 10924 4808 10964 4852
rect 11308 4808 11348 4852
rect 12748 4808 12788 4936
rect 12940 4892 12980 4936
rect 12893 4852 12940 4892
rect 12980 4852 12989 4892
rect 7433 4768 7564 4808
rect 7604 4768 7613 4808
rect 8812 4768 10964 4808
rect 11081 4768 11123 4808
rect 11163 4768 11212 4808
rect 11252 4768 11261 4808
rect 11308 4768 12788 4808
rect 13027 4768 13036 4808
rect 13076 4768 13207 4808
rect 13324 4724 13364 4936
rect 19276 4892 19316 4936
rect 14764 4852 19316 4892
rect 19756 4892 19796 4936
rect 20428 4892 20468 4936
rect 22828 4892 22868 4936
rect 23596 4892 23636 4936
rect 19756 4852 20860 4892
rect 20900 4852 20909 4892
rect 22781 4852 22828 4892
rect 22868 4852 22877 4892
rect 23587 4852 23596 4892
rect 23636 4852 23645 4892
rect 14764 4808 14804 4852
rect 24172 4808 24212 4927
rect 13507 4768 13516 4808
rect 13556 4768 14804 4808
rect 14921 4768 15052 4808
rect 15092 4768 15101 4808
rect 18089 4768 18220 4808
rect 18260 4768 18269 4808
rect 19258 4768 19267 4808
rect 19307 4768 20428 4808
rect 20468 4768 20477 4808
rect 21449 4768 21580 4808
rect 21620 4768 21629 4808
rect 22810 4768 22819 4808
rect 22859 4768 23884 4808
rect 23924 4768 24212 4808
rect 9763 4684 9772 4724
rect 9812 4684 11980 4724
rect 12020 4684 15820 4724
rect 15860 4684 15869 4724
rect 19721 4684 19852 4724
rect 19892 4684 19901 4724
rect 23299 4684 23308 4724
rect 23348 4684 26188 4724
rect 26228 4684 26237 4724
rect 3103 4516 3112 4556
rect 3480 4516 3489 4556
rect 10877 4516 10886 4556
rect 11254 4516 11263 4556
rect 18651 4516 18660 4556
rect 19028 4516 19037 4556
rect 26425 4516 26434 4556
rect 26802 4516 26811 4556
rect 19267 4348 19276 4388
rect 19316 4348 19843 4388
rect 19883 4348 19892 4388
rect 20201 4348 20332 4388
rect 20372 4348 20381 4388
rect 20515 4348 20524 4388
rect 20564 4348 20668 4388
rect 20708 4348 20717 4388
rect 9091 4264 9100 4304
rect 9140 4264 10060 4304
rect 10100 4264 10109 4304
rect 9571 4180 9580 4220
rect 9620 4180 10196 4220
rect 20419 4180 20428 4220
rect 20468 4180 20477 4220
rect 20524 4180 21292 4220
rect 21332 4180 21341 4220
rect 10156 4136 10196 4180
rect 20428 4136 20468 4180
rect 20524 4136 20564 4180
rect 9763 4096 9772 4136
rect 9812 4096 9964 4136
rect 10004 4096 10013 4136
rect 10147 4096 10156 4136
rect 10196 4096 10205 4136
rect 19651 4096 19660 4136
rect 19700 4096 19709 4136
rect 19834 4096 19843 4136
rect 19892 4096 20023 4136
rect 20323 4096 20332 4136
rect 20372 4096 20468 4136
rect 20515 4096 20524 4136
rect 20564 4096 20573 4136
rect 20681 4096 20812 4136
rect 20852 4096 20861 4136
rect 19660 4052 19700 4096
rect 19660 4012 21004 4052
rect 21044 4012 21053 4052
rect 4343 3760 4352 3800
rect 4720 3760 4729 3800
rect 12117 3760 12126 3800
rect 12494 3760 12503 3800
rect 19891 3760 19900 3800
rect 20268 3760 20277 3800
rect 27665 3760 27674 3800
rect 28042 3760 28051 3800
rect 3103 3004 3112 3044
rect 3480 3004 3489 3044
rect 10877 3004 10886 3044
rect 11254 3004 11263 3044
rect 18651 3004 18660 3044
rect 19028 3004 19037 3044
rect 26425 3004 26434 3044
rect 26802 3004 26811 3044
rect 4343 2248 4352 2288
rect 4720 2248 4729 2288
rect 12117 2248 12126 2288
rect 12494 2248 12503 2288
rect 19891 2248 19900 2288
rect 20268 2248 20277 2288
rect 27665 2248 27674 2288
rect 28042 2248 28051 2288
rect 3103 1492 3112 1532
rect 3480 1492 3489 1532
rect 10877 1492 10886 1532
rect 11254 1492 11263 1532
rect 18651 1492 18660 1532
rect 19028 1492 19037 1532
rect 26425 1492 26434 1532
rect 26802 1492 26811 1532
rect 4343 736 4352 776
rect 4720 736 4729 776
rect 12117 736 12126 776
rect 12494 736 12503 776
rect 19891 736 19900 776
rect 20268 736 20277 776
rect 27665 736 27674 776
rect 28042 736 28051 776
<< via2 >>
rect 2092 28876 2132 28916
rect 13516 28876 13556 28916
rect 5644 28624 5684 28664
rect 12652 28624 12692 28664
rect 4876 28540 4916 28580
rect 14092 28540 14132 28580
rect 16492 28540 16532 28580
rect 30028 28540 30068 28580
rect 2380 28456 2420 28496
rect 4108 28456 4148 28496
rect 24652 28456 24692 28496
rect 27244 28456 27284 28496
rect 9196 28372 9236 28412
rect 13708 28372 13748 28412
rect 19468 28372 19508 28412
rect 28972 28372 29012 28412
rect 2476 28288 2516 28328
rect 12556 28288 12596 28328
rect 23884 28288 23924 28328
rect 26764 28288 26804 28328
rect 23116 28204 23156 28244
rect 30028 28204 30068 28244
rect 23788 28120 23828 28160
rect 28876 28120 28916 28160
rect 2092 28036 2132 28076
rect 13804 28036 13844 28076
rect 1900 27868 1940 27908
rect 1900 27700 1940 27740
rect 2092 27700 2132 27740
rect 4352 27952 4720 27992
rect 5356 27952 5396 27992
rect 11308 27952 11348 27992
rect 12126 27952 12494 27992
rect 13132 27952 13172 27992
rect 19900 27952 20268 27992
rect 27674 27952 28042 27992
rect 2284 27868 2324 27908
rect 3052 27868 3092 27908
rect 4972 27868 5012 27908
rect 8620 27868 8660 27908
rect 13900 27868 13940 27908
rect 26380 27868 26420 27908
rect 27052 27868 27092 27908
rect 2476 27784 2516 27824
rect 2956 27784 2987 27824
rect 2987 27784 2996 27824
rect 4108 27784 4139 27824
rect 4139 27784 4148 27824
rect 5548 27784 5588 27824
rect 9292 27784 9332 27824
rect 10732 27784 10772 27824
rect 19468 27784 19508 27824
rect 1516 27616 1556 27656
rect 2380 27700 2420 27740
rect 2860 27700 2900 27740
rect 6892 27700 6923 27740
rect 6923 27700 6932 27740
rect 3340 27616 3371 27656
rect 3371 27616 3380 27656
rect 2380 27532 2420 27572
rect 2572 27532 2612 27572
rect 2764 27532 2804 27572
rect 3052 27532 3092 27572
rect 3724 27532 3764 27572
rect 3628 27448 3668 27488
rect 10540 27700 10580 27740
rect 13900 27700 13940 27740
rect 18028 27700 18068 27740
rect 4492 27616 4532 27656
rect 5068 27616 5108 27656
rect 5260 27616 5291 27656
rect 5291 27616 5300 27656
rect 5740 27616 5752 27656
rect 5752 27616 5780 27656
rect 6220 27616 6232 27656
rect 6232 27616 6260 27656
rect 6700 27647 6740 27656
rect 6700 27616 6740 27647
rect 9676 27616 9688 27656
rect 9688 27616 9716 27656
rect 11500 27616 11540 27656
rect 13228 27616 13268 27656
rect 13516 27616 13556 27656
rect 14284 27616 14324 27656
rect 16684 27616 16715 27656
rect 16715 27616 16724 27656
rect 19660 27616 19700 27656
rect 4204 27532 4244 27572
rect 5356 27532 5396 27572
rect 5548 27532 5587 27572
rect 5587 27532 5588 27572
rect 6316 27532 6356 27572
rect 8428 27532 8468 27572
rect 9484 27532 9523 27572
rect 9523 27532 9524 27572
rect 10636 27523 10676 27563
rect 12364 27532 12404 27572
rect 25420 27784 25460 27824
rect 27724 27784 27764 27824
rect 23788 27700 23828 27740
rect 24172 27700 24212 27740
rect 25804 27700 25844 27740
rect 26188 27700 26228 27740
rect 28492 27700 28532 27740
rect 21868 27616 21899 27656
rect 21899 27616 21908 27656
rect 13804 27532 13844 27572
rect 14092 27532 14132 27572
rect 16876 27532 16916 27572
rect 24364 27616 24395 27656
rect 24395 27616 24404 27656
rect 25228 27616 25268 27656
rect 26380 27616 26420 27656
rect 26764 27647 26804 27656
rect 26764 27616 26795 27647
rect 26795 27616 26804 27647
rect 27244 27647 27284 27656
rect 27244 27616 27275 27647
rect 27275 27616 27284 27647
rect 27724 27647 27764 27656
rect 27724 27616 27755 27647
rect 27755 27616 27764 27647
rect 28684 27647 28724 27656
rect 28684 27616 28715 27647
rect 28715 27616 28724 27647
rect 22252 27532 22283 27572
rect 22283 27532 22292 27572
rect 24556 27532 24596 27572
rect 24748 27532 24779 27572
rect 24779 27532 24788 27572
rect 25900 27532 25940 27572
rect 26188 27532 26228 27572
rect 26476 27532 26516 27572
rect 26860 27532 26900 27572
rect 27436 27532 27476 27572
rect 28492 27532 28532 27572
rect 28780 27532 28820 27572
rect 29260 27532 29300 27572
rect 30796 27616 30836 27656
rect 30988 27532 31028 27572
rect 4396 27448 4436 27488
rect 4876 27448 4916 27488
rect 652 27364 692 27404
rect 6412 27364 6443 27404
rect 6443 27364 6452 27404
rect 11980 27448 12020 27488
rect 19564 27448 19604 27488
rect 27532 27448 27572 27488
rect 29932 27448 29972 27488
rect 30220 27448 30260 27488
rect 9196 27364 9236 27404
rect 18316 27364 18356 27404
rect 23692 27364 23732 27404
rect 25804 27364 25844 27404
rect 26380 27364 26420 27404
rect 2188 27280 2228 27320
rect 4012 27280 4052 27320
rect 4972 27280 5012 27320
rect 3112 27196 3480 27236
rect 4588 27196 4628 27236
rect 6316 27196 6356 27236
rect 8332 27196 8372 27236
rect 9484 27196 9524 27236
rect 10886 27196 11254 27236
rect 9868 27112 9908 27152
rect 16012 27280 16052 27320
rect 23116 27280 23156 27320
rect 18660 27196 19028 27236
rect 23404 27196 23444 27236
rect 25996 27196 26036 27236
rect 26434 27196 26802 27236
rect 26956 27196 26996 27236
rect 15244 27112 15284 27152
rect 19276 27112 19316 27152
rect 19756 27112 19796 27152
rect 3340 27028 3380 27068
rect 9676 27028 9716 27068
rect 10348 27028 10388 27068
rect 11980 27028 12020 27068
rect 14188 27028 14228 27068
rect 18412 27028 18452 27068
rect 22252 27028 22292 27068
rect 22444 27028 22484 27068
rect 23596 27028 23636 27068
rect 28108 27028 28148 27068
rect 29644 27028 29684 27068
rect 3628 26944 3668 26984
rect 1036 26860 1076 26900
rect 1516 26860 1556 26900
rect 2380 26860 2420 26900
rect 2764 26860 2804 26900
rect 3148 26860 3188 26900
rect 3340 26860 3380 26900
rect 4780 26860 4820 26900
rect 652 26776 692 26816
rect 1228 26776 1259 26816
rect 1259 26776 1268 26816
rect 1804 26776 1844 26816
rect 2092 26776 2132 26816
rect 4588 26776 4628 26816
rect 4876 26776 4916 26816
rect 2188 26692 2228 26732
rect 2668 26692 2708 26732
rect 1132 26608 1172 26648
rect 1996 26608 2036 26648
rect 2764 26608 2795 26648
rect 2795 26608 2804 26648
rect 6316 26860 6356 26900
rect 5548 26776 5588 26816
rect 2956 26692 2996 26732
rect 4972 26692 5003 26732
rect 5003 26692 5012 26732
rect 8908 26860 8948 26900
rect 10060 26860 10100 26900
rect 12268 26944 12308 26984
rect 13228 26860 13268 26900
rect 13516 26860 13556 26900
rect 13900 26944 13940 26984
rect 15436 26944 15476 26984
rect 15820 26944 15860 26984
rect 26764 26944 26804 26984
rect 27148 26944 27188 26984
rect 28780 26944 28820 26984
rect 29260 26944 29300 26984
rect 17260 26860 17300 26900
rect 8812 26776 8852 26816
rect 9196 26776 9236 26816
rect 9868 26776 9908 26816
rect 10252 26776 10283 26816
rect 10283 26776 10292 26816
rect 13324 26776 13364 26816
rect 18220 26860 18260 26900
rect 18796 26860 18836 26900
rect 19372 26860 19412 26900
rect 19660 26860 19700 26900
rect 15052 26776 15092 26816
rect 15340 26776 15380 26816
rect 16780 26776 16820 26816
rect 17548 26776 17549 26816
rect 17549 26776 17588 26816
rect 18028 26776 18040 26816
rect 18040 26776 18068 26816
rect 14092 26734 14132 26774
rect 8140 26692 8180 26732
rect 13516 26692 13556 26732
rect 13900 26692 13940 26732
rect 14284 26692 14324 26732
rect 14668 26692 14708 26732
rect 4108 26608 4148 26648
rect 8044 26608 8084 26648
rect 8332 26608 8372 26648
rect 12172 26608 12212 26648
rect 13420 26608 13460 26648
rect 13804 26608 13844 26648
rect 14572 26608 14612 26648
rect 6700 26524 6740 26564
rect 8620 26524 8660 26564
rect 11116 26524 11156 26564
rect 12940 26524 12980 26564
rect 14860 26692 14900 26732
rect 17644 26692 17684 26732
rect 18316 26692 18356 26732
rect 18604 26692 18644 26732
rect 15436 26608 15476 26648
rect 16588 26608 16628 26648
rect 17356 26608 17396 26648
rect 18892 26608 18932 26648
rect 19564 26776 19604 26816
rect 20236 26776 20276 26816
rect 4352 26440 4720 26480
rect 6796 26440 6836 26480
rect 7180 26440 7220 26480
rect 9484 26440 9524 26480
rect 9676 26440 9716 26480
rect 9964 26440 10004 26480
rect 12126 26440 12494 26480
rect 14764 26440 14804 26480
rect 20428 26692 20468 26732
rect 23020 26860 23060 26900
rect 23692 26860 23732 26900
rect 24940 26860 24980 26900
rect 26284 26860 26324 26900
rect 28396 26860 28436 26900
rect 29356 26860 29396 26900
rect 29548 26860 29588 26900
rect 29932 26860 29972 26900
rect 30316 26860 30356 26900
rect 20812 26776 20852 26816
rect 27724 26776 27764 26816
rect 27916 26776 27944 26816
rect 27944 26776 27956 26816
rect 28972 26776 29012 26816
rect 21964 26692 22004 26732
rect 26380 26692 26420 26732
rect 20236 26608 20276 26648
rect 21100 26608 21140 26648
rect 22444 26608 22484 26648
rect 22636 26608 22676 26648
rect 26764 26608 26804 26648
rect 19084 26524 19124 26564
rect 27244 26692 27284 26732
rect 27628 26692 27668 26732
rect 28300 26692 28340 26732
rect 28204 26608 28244 26648
rect 30124 26608 30164 26648
rect 18988 26440 19028 26480
rect 19900 26440 20268 26480
rect 20524 26440 20564 26480
rect 21676 26440 21716 26480
rect 27436 26440 27476 26480
rect 27674 26440 28042 26480
rect 28396 26440 28436 26480
rect 5644 26356 5684 26396
rect 14476 26356 14516 26396
rect 15340 26356 15380 26396
rect 16396 26356 16436 26396
rect 22924 26356 22964 26396
rect 3532 26272 3572 26312
rect 4876 26272 4916 26312
rect 6220 26272 6260 26312
rect 6892 26272 6932 26312
rect 7372 26272 7412 26312
rect 11884 26272 11924 26312
rect 13516 26272 13556 26312
rect 1132 26188 1172 26228
rect 3436 26188 3476 26228
rect 6028 26188 6068 26228
rect 6412 26188 6452 26228
rect 7180 26188 7220 26228
rect 12940 26188 12980 26228
rect 13132 26188 13172 26228
rect 652 26104 692 26144
rect 844 26104 875 26144
rect 875 26104 884 26144
rect 1420 26104 1460 26144
rect 1804 26104 1844 26144
rect 2860 26104 2900 26144
rect 4204 26104 4244 26144
rect 5740 26104 5780 26144
rect 6796 26104 6836 26144
rect 7756 26104 7796 26144
rect 8236 26104 8276 26144
rect 8524 26104 8564 26144
rect 9292 26104 9332 26144
rect 9772 26104 9812 26144
rect 10540 26104 10580 26144
rect 11116 26104 11156 26144
rect 11404 26104 11444 26144
rect 11692 26104 11723 26144
rect 11723 26104 11732 26144
rect 12268 26104 12308 26144
rect 12844 26104 12884 26144
rect 940 26020 980 26060
rect 1996 26020 2036 26060
rect 2476 26020 2516 26060
rect 3628 26020 3668 26060
rect 1612 25936 1652 25976
rect 2284 25936 2324 25976
rect 2668 25936 2699 25976
rect 2699 25936 2708 25976
rect 6412 26020 6452 26060
rect 8140 26020 8180 26060
rect 11212 25936 11252 25976
rect 11788 26020 11828 26060
rect 14188 26272 14228 26312
rect 14956 26272 14987 26312
rect 14987 26272 14996 26312
rect 16012 26272 16037 26312
rect 16037 26272 16052 26312
rect 13900 26188 13940 26228
rect 14476 26188 14516 26228
rect 15532 26188 15572 26228
rect 15724 26188 15764 26228
rect 29356 26524 29396 26564
rect 29164 26440 29204 26480
rect 30316 26440 30356 26480
rect 25132 26356 25172 26396
rect 18604 26272 18644 26312
rect 19084 26272 19124 26312
rect 19948 26272 19988 26312
rect 24460 26272 24500 26312
rect 17164 26188 17204 26228
rect 17740 26188 17780 26228
rect 18316 26188 18356 26228
rect 13420 26104 13439 26144
rect 13439 26104 13460 26144
rect 13804 26104 13844 26144
rect 14092 26104 14132 26144
rect 14860 26104 14891 26144
rect 14891 26104 14900 26144
rect 15340 26104 15380 26144
rect 15628 26104 15668 26144
rect 16204 26135 16244 26144
rect 16204 26104 16244 26135
rect 16876 26104 16907 26144
rect 16907 26104 16916 26144
rect 15436 26020 15476 26060
rect 12076 25936 12116 25976
rect 13228 25936 13268 25976
rect 17356 26104 17396 26144
rect 22156 26188 22196 26228
rect 22636 26188 22676 26228
rect 22828 26188 22868 26228
rect 23308 26188 23348 26228
rect 26476 26188 26516 26228
rect 26668 26188 26708 26228
rect 18028 26104 18059 26144
rect 18059 26104 18068 26144
rect 18988 26104 19028 26144
rect 19276 26104 19310 26144
rect 19310 26104 19316 26144
rect 20236 26104 20276 26144
rect 21292 26104 21299 26144
rect 21299 26104 21332 26144
rect 21676 26104 21699 26144
rect 21699 26104 21716 26144
rect 28108 26272 28148 26312
rect 29740 26272 29780 26312
rect 30604 26272 30644 26312
rect 30988 26272 31028 26312
rect 27532 26188 27572 26228
rect 27916 26188 27956 26228
rect 28780 26188 28820 26228
rect 28972 26188 29012 26228
rect 22444 26104 22484 26144
rect 23020 26104 23060 26144
rect 23596 26104 23636 26144
rect 26764 26104 26795 26144
rect 26795 26104 26804 26144
rect 27628 26104 27668 26144
rect 17644 26020 17684 26060
rect 17836 26020 17876 26060
rect 18316 26020 18356 26060
rect 18796 26020 18836 26060
rect 19756 26020 19796 26060
rect 20716 26020 20756 26060
rect 21388 26020 21428 26060
rect 24844 26020 24875 26060
rect 24875 26020 24884 26060
rect 18892 25936 18932 25976
rect 19660 25936 19700 25976
rect 20044 25936 20084 25976
rect 21484 25936 21524 25976
rect 21676 25936 21716 25976
rect 23116 25936 23156 25976
rect 23692 25936 23723 25976
rect 23723 25936 23732 25976
rect 6220 25852 6260 25892
rect 7276 25852 7316 25892
rect 8524 25852 8564 25892
rect 9196 25852 9236 25892
rect 11692 25852 11732 25892
rect 11980 25852 12020 25892
rect 29644 26104 29682 26144
rect 29682 26104 29684 26144
rect 30412 26104 30452 26144
rect 26956 26020 26996 26060
rect 27148 26020 27179 26060
rect 27179 26020 27188 26060
rect 27724 26020 27764 26060
rect 28012 26020 28052 26060
rect 28684 26020 28724 26060
rect 29356 26020 29396 26060
rect 30028 26020 30068 26060
rect 27916 25936 27956 25976
rect 13900 25852 13940 25892
rect 14188 25852 14228 25892
rect 14572 25852 14612 25892
rect 15340 25852 15380 25892
rect 16396 25852 16436 25892
rect 18508 25852 18548 25892
rect 20620 25852 20660 25892
rect 25132 25852 25172 25892
rect 28588 25936 28628 25976
rect 29452 25936 29492 25976
rect 28876 25852 28916 25892
rect 29548 25852 29588 25892
rect 30028 25852 30068 25892
rect 8812 25768 8852 25808
rect 14860 25768 14900 25808
rect 17740 25768 17780 25808
rect 24268 25768 24308 25808
rect 27916 25768 27956 25808
rect 28588 25768 28628 25808
rect 3112 25684 3480 25724
rect 6796 25684 6836 25724
rect 10886 25684 11254 25724
rect 6700 25600 6740 25640
rect 3532 25516 3572 25556
rect 4972 25516 5012 25556
rect 6412 25516 6452 25556
rect 1036 25348 1076 25388
rect 4108 25348 4148 25388
rect 5260 25348 5300 25388
rect 6988 25348 7028 25388
rect 844 25264 884 25304
rect 1132 25264 1172 25304
rect 9580 25348 9620 25388
rect 18660 25684 19028 25724
rect 20140 25684 20180 25724
rect 20908 25684 20948 25724
rect 26434 25684 26802 25724
rect 11404 25516 11444 25556
rect 11788 25432 11828 25472
rect 13516 25432 13556 25472
rect 14380 25516 14420 25556
rect 14764 25516 14804 25556
rect 19564 25516 19604 25556
rect 19948 25516 19988 25556
rect 21004 25516 21035 25556
rect 21035 25516 21044 25556
rect 24172 25516 24212 25556
rect 24748 25516 24788 25556
rect 28876 25516 28916 25556
rect 14092 25432 14132 25472
rect 14476 25432 14516 25472
rect 11116 25348 11156 25388
rect 13900 25348 13940 25388
rect 14380 25348 14420 25388
rect 14956 25432 14996 25472
rect 15724 25432 15764 25472
rect 3148 25264 3188 25304
rect 4492 25264 4532 25304
rect 6604 25264 6644 25304
rect 7180 25264 7220 25304
rect 7372 25264 7412 25304
rect 9100 25264 9140 25304
rect 11212 25264 11252 25304
rect 11692 25264 11732 25304
rect 11980 25264 12020 25304
rect 12748 25264 12757 25304
rect 12757 25264 12788 25304
rect 12940 25264 12980 25304
rect 4108 25180 4148 25220
rect 8908 25180 8948 25220
rect 9676 25180 9716 25220
rect 11404 25180 11444 25220
rect 6412 25096 6452 25136
rect 7084 25096 7124 25136
rect 7852 25096 7892 25136
rect 9964 25096 10004 25136
rect 10828 25096 10868 25136
rect 11308 25096 11339 25136
rect 11339 25096 11348 25136
rect 8140 25012 8180 25052
rect 4352 24928 4720 24968
rect 4876 24844 4916 24884
rect 8716 24844 8756 24884
rect 2092 24760 2132 24800
rect 3340 24760 3380 24800
rect 4492 24760 4532 24800
rect 7756 24760 7796 24800
rect 8140 24760 8180 24800
rect 4972 24676 5012 24716
rect 6796 24676 6836 24716
rect 14860 25264 14900 25304
rect 15916 25264 15956 25304
rect 16396 25264 16436 25304
rect 16780 25264 16820 25304
rect 16972 25264 17012 25304
rect 18988 25432 19028 25472
rect 20140 25432 20180 25472
rect 20908 25432 20948 25472
rect 23020 25432 23060 25472
rect 24940 25432 24980 25472
rect 28684 25432 28724 25472
rect 12844 25180 12884 25220
rect 13324 25180 13364 25220
rect 13708 25180 13748 25220
rect 14380 25180 14420 25220
rect 15436 25180 15476 25220
rect 16204 25180 16233 25220
rect 16233 25180 16244 25220
rect 12556 25096 12596 25136
rect 13420 25096 13460 25136
rect 13900 25096 13940 25136
rect 15724 25096 15764 25136
rect 16108 25096 16148 25136
rect 18604 25348 18644 25388
rect 19372 25348 19403 25388
rect 19403 25348 19412 25388
rect 19660 25348 19700 25388
rect 19852 25348 19892 25388
rect 20716 25348 20756 25388
rect 18508 25264 18548 25304
rect 19180 25264 19220 25304
rect 19468 25264 19506 25304
rect 19506 25264 19508 25304
rect 20140 25264 20180 25304
rect 20908 25264 20948 25304
rect 21292 25264 21332 25304
rect 21580 25264 21620 25304
rect 18028 25180 18068 25220
rect 18220 25180 18260 25220
rect 19564 25180 19595 25220
rect 19595 25180 19604 25220
rect 20044 25180 20084 25220
rect 16684 25096 16724 25136
rect 17644 25096 17684 25136
rect 18796 25096 18827 25136
rect 18827 25096 18836 25136
rect 14476 25012 14516 25052
rect 9100 24928 9140 24968
rect 11884 24928 11924 24968
rect 12126 24928 12494 24968
rect 9292 24844 9332 24884
rect 10732 24844 10772 24884
rect 11212 24844 11252 24884
rect 11980 24844 12020 24884
rect 16684 24928 16724 24968
rect 8620 24760 8660 24800
rect 9100 24760 9140 24800
rect 13228 24760 13268 24800
rect 14956 24760 14996 24800
rect 16108 24760 16148 24800
rect 18124 24760 18164 24800
rect 18316 24760 18356 24800
rect 18508 24760 18548 24800
rect 18796 24760 18827 24800
rect 18827 24760 18836 24800
rect 8812 24676 8841 24716
rect 8841 24676 8852 24716
rect 12844 24676 12884 24716
rect 1036 24592 1067 24632
rect 1067 24592 1076 24632
rect 4396 24592 4436 24632
rect 5068 24592 5108 24632
rect 5548 24592 5579 24632
rect 5579 24592 5588 24632
rect 6604 24592 6644 24632
rect 8908 24592 8948 24632
rect 19276 25012 19316 25052
rect 21388 25012 21428 25052
rect 19900 24928 20268 24968
rect 19276 24844 19316 24884
rect 21004 24844 21044 24884
rect 19468 24760 19508 24800
rect 21292 24760 21332 24800
rect 23308 25348 23348 25388
rect 25420 25348 25451 25388
rect 25451 25348 25460 25388
rect 28588 25348 28628 25388
rect 28876 25348 28916 25388
rect 22924 25264 22964 25304
rect 23212 25264 23252 25304
rect 24076 25264 24116 25304
rect 25228 25264 25268 25304
rect 27340 25264 27371 25304
rect 27371 25264 27380 25304
rect 23308 25180 23348 25220
rect 25996 25180 26036 25220
rect 28108 25180 28148 25220
rect 29644 25516 29684 25556
rect 29356 25432 29396 25472
rect 29452 25348 29492 25388
rect 30220 25180 30260 25220
rect 23212 25096 23252 25136
rect 24268 25096 24308 25136
rect 28396 25096 28436 25136
rect 28972 25012 29012 25052
rect 29164 25012 29204 25052
rect 27674 24928 28042 24968
rect 25324 24844 25364 24884
rect 22636 24760 22676 24800
rect 23020 24760 23051 24800
rect 23051 24760 23060 24800
rect 25036 24760 25076 24800
rect 14380 24676 14420 24716
rect 16012 24676 16052 24716
rect 19756 24676 19796 24716
rect 20140 24676 20180 24716
rect 21580 24676 21620 24716
rect 22348 24676 22388 24716
rect 25804 24676 25844 24716
rect 27436 24676 27476 24716
rect 11212 24592 11252 24632
rect 11500 24592 11540 24632
rect 11980 24592 12020 24632
rect 13324 24592 13364 24632
rect 13516 24592 13556 24632
rect 13900 24592 13940 24632
rect 1708 24508 1748 24548
rect 3340 24508 3380 24548
rect 3724 24508 3764 24548
rect 8236 24508 8276 24548
rect 8428 24508 8468 24548
rect 10348 24508 10388 24548
rect 11788 24508 11819 24548
rect 11819 24508 11828 24548
rect 29836 24676 29876 24716
rect 16108 24592 16148 24632
rect 16588 24623 16628 24632
rect 16588 24592 16619 24623
rect 16619 24592 16628 24623
rect 17164 24592 17195 24632
rect 17195 24592 17204 24632
rect 17740 24592 17780 24632
rect 18220 24592 18260 24632
rect 18508 24592 18548 24632
rect 18700 24592 18739 24632
rect 18739 24592 18740 24632
rect 18988 24592 19027 24632
rect 19027 24592 19028 24632
rect 19276 24592 19307 24632
rect 19307 24592 19316 24632
rect 21868 24592 21899 24632
rect 21899 24592 21908 24632
rect 22924 24592 22964 24632
rect 24364 24592 24404 24632
rect 27340 24592 27380 24632
rect 29644 24592 29684 24632
rect 30124 24592 30164 24632
rect 21580 24508 21620 24548
rect 23788 24508 23828 24548
rect 25324 24508 25364 24548
rect 28780 24508 28820 24548
rect 29068 24508 29108 24548
rect 2572 24424 2612 24464
rect 9580 24424 9620 24464
rect 11980 24424 12020 24464
rect 17356 24424 17396 24464
rect 18508 24424 18548 24464
rect 19564 24424 19604 24464
rect 22444 24424 22484 24464
rect 23212 24424 23252 24464
rect 460 24340 500 24380
rect 3532 24340 3572 24380
rect 29260 24424 29300 24464
rect 30988 24424 31028 24464
rect 4876 24340 4916 24380
rect 9196 24340 9236 24380
rect 12556 24340 12596 24380
rect 14860 24340 14900 24380
rect 15148 24340 15188 24380
rect 20332 24340 20372 24380
rect 20908 24340 20948 24380
rect 24460 24340 24500 24380
rect 25708 24340 25748 24380
rect 28396 24340 28436 24380
rect 28684 24340 28724 24380
rect 29452 24340 29492 24380
rect 30028 24340 30068 24380
rect 12844 24256 12884 24296
rect 14188 24256 14228 24296
rect 22060 24256 22100 24296
rect 25516 24256 25556 24296
rect 3112 24172 3480 24212
rect 9004 24172 9044 24212
rect 10636 24172 10676 24212
rect 10886 24172 11254 24212
rect 18660 24172 19028 24212
rect 24460 24172 24500 24212
rect 26434 24172 26802 24212
rect 10060 24088 10100 24128
rect 29740 24088 29780 24128
rect 4780 24004 4820 24044
rect 6796 24004 6827 24044
rect 6827 24004 6836 24044
rect 9964 24004 10004 24044
rect 10828 24004 10868 24044
rect 12748 24004 12788 24044
rect 13516 24004 13556 24044
rect 15820 24004 15860 24044
rect 16204 24004 16244 24044
rect 19852 24004 19892 24044
rect 22348 24004 22388 24044
rect 25900 24004 25931 24044
rect 25931 24004 25940 24044
rect 27436 24004 27476 24044
rect 28204 24004 28244 24044
rect 28876 24004 28916 24044
rect 29644 24004 29684 24044
rect 556 23920 596 23960
rect 5260 23836 5300 23876
rect 364 23752 404 23792
rect 940 23752 980 23792
rect 1420 23752 1460 23792
rect 2668 23752 2708 23792
rect 4204 23752 4244 23792
rect 4876 23752 4916 23792
rect 12364 23920 12404 23960
rect 18316 23920 18356 23960
rect 19660 23920 19700 23960
rect 24364 23920 24404 23960
rect 7084 23836 7124 23876
rect 8140 23836 8180 23876
rect 11308 23836 11348 23876
rect 11500 23836 11540 23876
rect 13516 23836 13556 23876
rect 15148 23836 15179 23876
rect 15179 23836 15188 23876
rect 15724 23836 15764 23876
rect 16300 23836 16340 23876
rect 16684 23836 16724 23876
rect 18124 23836 18164 23876
rect 30508 23920 30548 23960
rect 21292 23836 21332 23876
rect 8620 23752 8660 23792
rect 8908 23752 8948 23792
rect 9196 23752 9236 23792
rect 9964 23752 10004 23792
rect 10252 23752 10292 23792
rect 11116 23752 11156 23792
rect 12556 23752 12596 23792
rect 13036 23752 13076 23792
rect 15244 23752 15284 23792
rect 15628 23752 15668 23792
rect 15916 23752 15956 23792
rect 16876 23752 16916 23792
rect 17356 23752 17396 23792
rect 17644 23752 17684 23792
rect 18316 23752 18356 23792
rect 18892 23752 18932 23792
rect 19084 23752 19124 23792
rect 19852 23752 19892 23792
rect 20236 23752 20276 23792
rect 1228 23668 1268 23708
rect 3052 23668 3092 23708
rect 4780 23668 4820 23708
rect 6220 23668 6260 23708
rect 6988 23668 7028 23708
rect 9100 23668 9140 23708
rect 3532 23584 3572 23624
rect 5068 23584 5108 23624
rect 5836 23584 5876 23624
rect 6412 23584 6452 23624
rect 7660 23584 7700 23624
rect 7948 23584 7988 23624
rect 9196 23584 9236 23624
rect 10348 23668 10388 23708
rect 7180 23500 7220 23540
rect 10828 23668 10868 23708
rect 11404 23668 11444 23708
rect 12460 23668 12500 23708
rect 10636 23584 10676 23624
rect 16300 23668 16340 23708
rect 16972 23668 17012 23708
rect 16204 23584 16244 23624
rect 22636 23836 22667 23876
rect 22667 23836 22676 23876
rect 24076 23836 24116 23876
rect 25804 23836 25844 23876
rect 29164 23836 29204 23876
rect 21004 23752 21044 23792
rect 21772 23752 21812 23792
rect 22060 23752 22100 23792
rect 23116 23752 23156 23792
rect 24364 23752 24404 23792
rect 24940 23752 24980 23792
rect 25132 23752 25156 23792
rect 25156 23752 25172 23792
rect 25996 23752 26036 23792
rect 26188 23752 26228 23792
rect 27244 23752 27284 23792
rect 28204 23752 28244 23792
rect 17452 23668 17492 23708
rect 19756 23668 19796 23708
rect 18508 23584 18548 23624
rect 21388 23584 21428 23624
rect 22444 23584 22484 23624
rect 16876 23500 16916 23540
rect 19372 23500 19412 23540
rect 4352 23416 4720 23456
rect 9388 23416 9428 23456
rect 11884 23416 11924 23456
rect 12126 23416 12494 23456
rect 15916 23416 15956 23456
rect 16300 23416 16340 23456
rect 19900 23416 20268 23456
rect 556 23164 596 23204
rect 9004 23332 9044 23372
rect 10732 23332 10772 23372
rect 13420 23332 13460 23372
rect 2572 23248 2612 23288
rect 4300 23248 4340 23288
rect 4780 23248 4820 23288
rect 5644 23248 5684 23288
rect 6988 23248 7028 23288
rect 7372 23248 7412 23288
rect 8236 23248 8276 23288
rect 11692 23248 11732 23288
rect 5548 23164 5588 23204
rect 6604 23164 6644 23204
rect 7084 23164 7124 23204
rect 7468 23164 7508 23204
rect 7756 23164 7787 23204
rect 7787 23164 7796 23204
rect 172 23080 212 23120
rect 1036 23080 1067 23120
rect 1067 23080 1076 23120
rect 3340 23080 3380 23120
rect 3916 23080 3956 23120
rect 5068 23080 5108 23120
rect 6412 23080 6452 23120
rect 13228 23164 13268 23204
rect 14668 23248 14708 23288
rect 14476 23164 14516 23204
rect 23788 23668 23828 23708
rect 24556 23668 24596 23708
rect 25900 23668 25940 23708
rect 26284 23668 26324 23708
rect 25324 23584 25364 23624
rect 25516 23584 25547 23624
rect 25547 23584 25556 23624
rect 22732 23500 22772 23540
rect 17452 23332 17492 23372
rect 15628 23248 15668 23288
rect 16204 23248 16244 23288
rect 16684 23248 16724 23288
rect 17356 23248 17396 23288
rect 19468 23248 19508 23288
rect 20236 23248 20276 23288
rect 20812 23248 20852 23288
rect 21100 23248 21140 23288
rect 15244 23164 15284 23204
rect 8716 23080 8756 23120
rect 8908 23080 8948 23120
rect 9388 23080 9428 23120
rect 9868 23080 9899 23120
rect 9899 23080 9908 23120
rect 11788 23080 11828 23120
rect 13132 23080 13172 23120
rect 13516 23080 13556 23120
rect 1996 22996 2036 23036
rect 4684 22996 4724 23036
rect 5644 22996 5684 23036
rect 6220 22996 6260 23036
rect 7180 22996 7220 23036
rect 14572 23080 14612 23120
rect 7564 22996 7595 23036
rect 7595 22996 7604 23036
rect 7852 22996 7892 23036
rect 9100 22996 9131 23036
rect 9131 22996 9140 23036
rect 10348 22996 10388 23036
rect 11500 22996 11540 23036
rect 12844 22996 12884 23036
rect 13420 22996 13460 23036
rect 14188 22996 14228 23036
rect 15724 22996 15764 23036
rect 16108 22996 16148 23036
rect 17164 23164 17204 23204
rect 18892 23164 18932 23204
rect 19564 23164 19604 23204
rect 20524 23164 20564 23204
rect 21580 23164 21620 23204
rect 17452 23080 17492 23120
rect 17836 23080 17876 23120
rect 18604 23080 18605 23120
rect 18605 23080 18644 23120
rect 19660 23080 19691 23120
rect 19691 23080 19700 23120
rect 17164 22996 17187 23036
rect 17187 22996 17204 23036
rect 18316 22996 18356 23036
rect 7276 22912 7316 22952
rect 16396 22912 16436 22952
rect 5836 22828 5876 22868
rect 11212 22828 11252 22868
rect 11884 22828 11924 22868
rect 14572 22828 14612 22868
rect 16300 22828 16340 22868
rect 3112 22660 3480 22700
rect 21100 23080 21131 23120
rect 21131 23080 21140 23120
rect 21388 23080 21428 23120
rect 19564 22996 19604 23036
rect 20908 22996 20948 23036
rect 23308 23500 23348 23540
rect 28204 23500 28244 23540
rect 30220 23836 30260 23876
rect 29068 23752 29108 23792
rect 29644 23752 29684 23792
rect 28972 23668 29012 23708
rect 30316 23668 30356 23708
rect 29164 23584 29204 23624
rect 29548 23584 29588 23624
rect 29836 23584 29876 23624
rect 30988 23584 31028 23624
rect 28876 23500 28916 23540
rect 27674 23416 28042 23456
rect 28588 23416 28628 23456
rect 29548 23416 29588 23456
rect 25324 23332 25364 23372
rect 26572 23332 26612 23372
rect 27244 23248 27284 23288
rect 28204 23164 28244 23204
rect 29164 23164 29204 23204
rect 22732 23080 22772 23120
rect 24076 23080 24116 23120
rect 26284 23080 26324 23120
rect 26572 23080 26612 23120
rect 28588 23080 28628 23120
rect 28972 23080 29012 23120
rect 29452 23080 29492 23120
rect 29740 23080 29780 23120
rect 26380 22996 26420 23036
rect 26860 22996 26900 23036
rect 30028 22996 30068 23036
rect 22060 22912 22100 22952
rect 29164 22912 29204 22952
rect 29644 22912 29684 22952
rect 30412 22912 30452 22952
rect 17548 22828 17588 22868
rect 19084 22828 19124 22868
rect 19852 22828 19892 22868
rect 21580 22828 21620 22868
rect 24940 22828 24980 22868
rect 28780 22828 28820 22868
rect 9292 22744 9332 22784
rect 11500 22744 11540 22784
rect 21484 22744 21524 22784
rect 30124 22744 30164 22784
rect 8812 22660 8852 22700
rect 10886 22660 11254 22700
rect 16300 22660 16340 22700
rect 18660 22660 19028 22700
rect 26434 22660 26802 22700
rect 7276 22576 7316 22616
rect 9100 22576 9140 22616
rect 18316 22576 18356 22616
rect 1612 22408 1652 22448
rect 5644 22408 5684 22448
rect 4204 22324 4244 22364
rect 4684 22324 4724 22364
rect 6124 22324 6164 22364
rect 6508 22324 6548 22364
rect 6892 22492 6932 22532
rect 10732 22492 10772 22532
rect 11500 22492 11540 22532
rect 19468 22492 19508 22532
rect 21004 22492 21044 22532
rect 21676 22492 21716 22532
rect 8236 22408 8267 22448
rect 8267 22408 8276 22448
rect 9772 22408 9812 22448
rect 10252 22408 10292 22448
rect 7756 22324 7796 22364
rect 9100 22324 9140 22364
rect 10060 22324 10100 22364
rect 14764 22408 14804 22448
rect 17452 22408 17492 22448
rect 13132 22324 13172 22364
rect 556 22240 596 22280
rect 1804 22240 1844 22280
rect 2092 22240 2132 22280
rect 2572 22240 2612 22280
rect 3916 22240 3956 22280
rect 4972 22240 5003 22280
rect 5003 22240 5012 22280
rect 5644 22240 5669 22280
rect 5669 22240 5684 22280
rect 15724 22324 15764 22364
rect 16012 22324 16052 22364
rect 16300 22324 16340 22364
rect 16684 22324 16724 22364
rect 16972 22324 17012 22364
rect 17548 22324 17588 22364
rect 20812 22324 20852 22364
rect 21484 22324 21524 22364
rect 21772 22324 21812 22364
rect 22060 22324 22100 22364
rect 24460 22492 24500 22532
rect 26380 22492 26420 22532
rect 26860 22492 26900 22532
rect 27052 22492 27092 22532
rect 28972 22492 29012 22532
rect 30316 22408 30356 22448
rect 30604 22408 30644 22448
rect 30796 22408 30836 22448
rect 25804 22324 25844 22364
rect 27532 22324 27572 22364
rect 29356 22324 29396 22364
rect 7084 22240 7124 22280
rect 7564 22240 7595 22280
rect 7595 22240 7604 22280
rect 8236 22240 8276 22280
rect 8908 22240 8947 22280
rect 8947 22240 8948 22280
rect 9196 22240 9236 22280
rect 9868 22240 9908 22280
rect 11788 22240 11828 22280
rect 13516 22240 13556 22280
rect 14284 22240 14324 22280
rect 14860 22240 14900 22280
rect 16780 22240 16820 22280
rect 17164 22240 17195 22280
rect 17195 22240 17204 22280
rect 18412 22240 18452 22280
rect 19180 22240 19211 22280
rect 19211 22240 19220 22280
rect 19564 22240 19604 22280
rect 22156 22240 22196 22280
rect 22444 22240 22475 22280
rect 22475 22240 22484 22280
rect 24940 22240 24980 22280
rect 30124 22324 30164 22364
rect 25900 22240 25940 22280
rect 26764 22240 26804 22280
rect 27340 22240 27380 22280
rect 28780 22240 28820 22280
rect 30028 22240 30068 22280
rect 30508 22240 30548 22280
rect 30700 22240 30740 22280
rect 844 22156 884 22196
rect 4108 22156 4148 22196
rect 1228 22072 1267 22112
rect 1267 22072 1268 22112
rect 2860 22072 2900 22112
rect 3820 22072 3860 22112
rect 4396 22156 4427 22196
rect 4427 22156 4436 22196
rect 6124 22156 6164 22196
rect 6700 22156 6740 22196
rect 7372 22156 7412 22196
rect 8044 22156 8084 22196
rect 13228 22156 13268 22196
rect 4684 22072 4715 22112
rect 4715 22072 4724 22112
rect 6028 22072 6068 22112
rect 6604 22072 6644 22112
rect 14380 22156 14420 22196
rect 16012 22156 16052 22196
rect 16396 22156 16436 22196
rect 9676 22072 9716 22112
rect 10252 22072 10292 22112
rect 12940 22072 12980 22112
rect 19084 22156 19124 22196
rect 26956 22156 26996 22196
rect 27148 22156 27188 22196
rect 18412 22072 18451 22112
rect 18451 22072 18452 22112
rect 21676 22072 21716 22112
rect 24460 22072 24500 22112
rect 25516 22072 25556 22112
rect 30028 22072 30068 22112
rect 2380 21988 2420 22028
rect 6412 21988 6452 22028
rect 17260 21988 17300 22028
rect 18892 21988 18932 22028
rect 21484 21988 21524 22028
rect 25900 21988 25940 22028
rect 3340 21904 3380 21944
rect 4352 21904 4720 21944
rect 1516 21820 1556 21860
rect 5068 21820 5108 21860
rect 9676 21904 9716 21944
rect 12126 21904 12494 21944
rect 13516 21904 13556 21944
rect 16396 21904 16436 21944
rect 16972 21904 17012 21944
rect 19900 21904 20268 21944
rect 27674 21904 28042 21944
rect 6412 21820 6452 21860
rect 2572 21736 2612 21776
rect 3724 21652 3764 21692
rect 4492 21652 4532 21692
rect 4780 21652 4820 21692
rect 5740 21652 5780 21692
rect 6124 21736 6155 21776
rect 6155 21736 6164 21776
rect 6604 21736 6635 21776
rect 6635 21736 6644 21776
rect 7084 21736 7124 21776
rect 7756 21736 7796 21776
rect 6028 21652 6068 21692
rect 8236 21652 8267 21692
rect 8267 21652 8276 21692
rect 10060 21820 10100 21860
rect 17452 21820 17492 21860
rect 26188 21820 26228 21860
rect 8716 21736 8756 21776
rect 9580 21736 9620 21776
rect 13324 21736 13364 21776
rect 13708 21736 13748 21776
rect 15244 21736 15284 21776
rect 20140 21736 20180 21776
rect 24268 21736 24308 21776
rect 24940 21736 24980 21776
rect 25516 21736 25556 21776
rect 27532 21736 27572 21776
rect 8812 21652 8852 21692
rect 9676 21652 9716 21692
rect 10252 21652 10292 21692
rect 13420 21652 13460 21692
rect 16012 21652 16052 21692
rect 16204 21652 16244 21692
rect 16972 21652 17012 21692
rect 17356 21652 17396 21692
rect 18892 21652 18932 21692
rect 20428 21652 20468 21692
rect 21580 21652 21620 21692
rect 24556 21652 24596 21692
rect 26092 21652 26132 21692
rect 26380 21652 26420 21692
rect 2284 21568 2324 21608
rect 2668 21568 2708 21608
rect 3148 21568 3179 21608
rect 3179 21568 3188 21608
rect 3436 21568 3476 21608
rect 3820 21568 3860 21608
rect 4204 21568 4244 21608
rect 4588 21568 4628 21608
rect 5164 21568 5204 21608
rect 6316 21568 6356 21608
rect 6700 21568 6740 21608
rect 1036 21484 1076 21524
rect 940 21400 980 21440
rect 1324 21400 1364 21440
rect 1420 21316 1460 21356
rect 1228 21064 1268 21104
rect 2092 21484 2132 21524
rect 2860 21484 2900 21524
rect 4684 21484 4724 21524
rect 2572 21400 2612 21440
rect 8908 21568 8948 21608
rect 9580 21543 9620 21583
rect 5068 21484 5108 21524
rect 6124 21484 6164 21524
rect 6412 21484 6452 21524
rect 7468 21484 7508 21524
rect 7756 21484 7796 21524
rect 3340 21400 3380 21440
rect 4972 21400 5012 21440
rect 6028 21400 6068 21440
rect 8236 21484 8276 21524
rect 10540 21568 10580 21608
rect 11116 21568 11128 21608
rect 11128 21568 11156 21608
rect 11596 21568 11608 21608
rect 11608 21568 11636 21608
rect 11788 21568 11828 21608
rect 12844 21568 12884 21608
rect 13228 21568 13268 21608
rect 13516 21568 13556 21608
rect 13996 21568 14036 21608
rect 14380 21568 14411 21608
rect 14411 21568 14420 21608
rect 15628 21568 15668 21608
rect 16396 21568 16436 21608
rect 17068 21568 17108 21608
rect 17645 21568 17684 21608
rect 17684 21568 17685 21608
rect 10732 21484 10772 21524
rect 8812 21400 8852 21440
rect 9004 21400 9044 21440
rect 9964 21400 10004 21440
rect 19852 21568 19892 21608
rect 20716 21568 20756 21608
rect 21100 21568 21140 21608
rect 21868 21568 21908 21608
rect 22444 21568 22484 21608
rect 22636 21568 22676 21608
rect 24076 21568 24097 21608
rect 24097 21568 24116 21608
rect 13804 21484 13835 21524
rect 13835 21484 13844 21524
rect 14764 21484 14804 21524
rect 15532 21484 15563 21524
rect 15563 21484 15572 21524
rect 16108 21484 16148 21524
rect 16684 21484 16724 21524
rect 16876 21484 16916 21524
rect 17548 21484 17579 21524
rect 17579 21484 17588 21524
rect 17836 21484 17876 21524
rect 24652 21568 24692 21608
rect 25228 21568 25268 21608
rect 25804 21568 25844 21608
rect 27436 21568 27467 21608
rect 27467 21568 27476 21608
rect 28780 21568 28820 21608
rect 30988 21568 31028 21608
rect 18028 21484 18068 21524
rect 19084 21484 19124 21524
rect 20620 21484 20660 21524
rect 23500 21484 23540 21524
rect 23884 21484 23924 21524
rect 24460 21484 24500 21524
rect 15916 21400 15956 21440
rect 17932 21400 17972 21440
rect 19276 21400 19316 21440
rect 20716 21400 20756 21440
rect 22828 21400 22868 21440
rect 24172 21400 24212 21440
rect 25132 21400 25135 21440
rect 25135 21400 25172 21440
rect 2188 21316 2228 21356
rect 3436 21316 3476 21356
rect 5740 21316 5780 21356
rect 7084 21316 7124 21356
rect 7372 21316 7412 21356
rect 11692 21316 11732 21356
rect 11980 21316 12020 21356
rect 15724 21316 15764 21356
rect 16876 21316 16916 21356
rect 17068 21316 17108 21356
rect 4300 21232 4340 21272
rect 15148 21232 15188 21272
rect 17740 21232 17780 21272
rect 30796 21484 30836 21524
rect 30316 21400 30356 21440
rect 30892 21400 30932 21440
rect 21388 21316 21428 21356
rect 23788 21316 23819 21356
rect 23819 21316 23828 21356
rect 30604 21316 30644 21356
rect 30508 21232 30548 21272
rect 3112 21148 3480 21188
rect 3724 21148 3764 21188
rect 7852 21148 7892 21188
rect 8236 21148 8276 21188
rect 10886 21148 11254 21188
rect 18660 21148 19028 21188
rect 23308 21148 23348 21188
rect 26434 21148 26802 21188
rect 27244 21148 27284 21188
rect 30316 21148 30356 21188
rect 2956 21064 2996 21104
rect 6028 21064 6068 21104
rect 9100 21064 9140 21104
rect 19852 21064 19892 21104
rect 22924 21064 22964 21104
rect 1900 20980 1940 21020
rect 6124 20980 6164 21020
rect 7372 20980 7412 21020
rect 7564 20980 7604 21020
rect 7756 20980 7796 21020
rect 9196 20980 9236 21020
rect 13228 20980 13268 21020
rect 14764 20980 14804 21020
rect 16780 20980 16820 21020
rect 17836 20980 17876 21020
rect 18124 20980 18164 21020
rect 25228 20980 25268 21020
rect 30028 20980 30068 21020
rect 1804 20896 1844 20936
rect 3916 20896 3956 20936
rect 5164 20896 5204 20936
rect 748 20812 788 20852
rect 1132 20812 1172 20852
rect 2092 20812 2123 20852
rect 2123 20812 2132 20852
rect 2668 20812 2699 20852
rect 2699 20812 2708 20852
rect 3724 20812 3764 20852
rect 6412 20896 6452 20936
rect 6796 20896 6836 20936
rect 7084 20896 7124 20936
rect 10348 20896 10388 20936
rect 13132 20896 13172 20936
rect 13324 20896 13364 20936
rect 6220 20812 6260 20852
rect 7276 20812 7316 20852
rect 7948 20812 7988 20852
rect 8140 20812 8180 20852
rect 9388 20812 9428 20852
rect 9868 20812 9908 20852
rect 940 20728 980 20768
rect 1612 20728 1652 20768
rect 2188 20728 2228 20768
rect 2956 20728 2996 20768
rect 3340 20728 3380 20768
rect 5164 20728 5204 20768
rect 5644 20728 5684 20768
rect 7180 20728 7220 20768
rect 7564 20728 7604 20768
rect 748 20644 788 20684
rect 2860 20644 2900 20684
rect 3724 20644 3764 20684
rect 2380 20560 2420 20600
rect 3916 20560 3956 20600
rect 4780 20560 4820 20600
rect 268 20392 308 20432
rect 1132 20392 1172 20432
rect 1420 20476 1460 20516
rect 1708 20392 1748 20432
rect 2764 20392 2804 20432
rect 3436 20392 3476 20432
rect 4352 20392 4720 20432
rect 940 20308 980 20348
rect 2380 20308 2420 20348
rect 2956 20308 2996 20348
rect 1036 20140 1076 20180
rect 2188 20224 2228 20264
rect 6508 20644 6548 20684
rect 7852 20644 7892 20684
rect 9676 20728 9716 20768
rect 11020 20728 11060 20768
rect 8332 20644 8372 20684
rect 6988 20560 7028 20600
rect 7468 20560 7499 20600
rect 7499 20560 7508 20600
rect 9004 20644 9015 20684
rect 9015 20644 9044 20684
rect 10540 20644 10580 20684
rect 8812 20560 8843 20600
rect 8843 20560 8852 20600
rect 9100 20560 9140 20600
rect 9772 20560 9812 20600
rect 14860 20896 14900 20936
rect 15532 20896 15572 20936
rect 17452 20896 17492 20936
rect 13516 20812 13556 20852
rect 13708 20812 13748 20852
rect 15052 20812 15092 20852
rect 16396 20812 16436 20852
rect 16780 20812 16820 20852
rect 11596 20728 11636 20768
rect 13324 20728 13331 20768
rect 13331 20728 13364 20768
rect 18412 20896 18452 20936
rect 17260 20812 17291 20852
rect 17291 20812 17300 20852
rect 18604 20812 18635 20852
rect 18635 20812 18644 20852
rect 13996 20728 14036 20768
rect 14380 20728 14420 20768
rect 14860 20728 14900 20768
rect 15244 20728 15284 20768
rect 16012 20728 16052 20768
rect 16684 20728 16724 20768
rect 16972 20728 17012 20768
rect 17452 20728 17492 20768
rect 18028 20728 18068 20768
rect 18412 20728 18443 20768
rect 18443 20728 18452 20768
rect 20332 20896 20372 20936
rect 20428 20812 20468 20852
rect 24364 20896 24404 20936
rect 25132 20896 25172 20936
rect 25612 20896 25652 20936
rect 20620 20728 20660 20768
rect 12940 20644 12980 20684
rect 13228 20644 13268 20684
rect 13420 20644 13460 20684
rect 15916 20644 15955 20684
rect 15955 20644 15956 20684
rect 18316 20644 18356 20684
rect 22732 20812 22772 20852
rect 22924 20812 22964 20852
rect 24556 20812 24596 20852
rect 21292 20728 21332 20768
rect 21964 20728 22004 20768
rect 27244 20896 27284 20936
rect 29932 20896 29972 20936
rect 30604 20980 30644 21020
rect 30892 20896 30932 20936
rect 29548 20812 29588 20852
rect 22348 20728 22388 20768
rect 22636 20728 22676 20768
rect 23308 20728 23348 20768
rect 23596 20728 23635 20768
rect 23635 20728 23636 20768
rect 24172 20728 24212 20768
rect 24652 20728 24692 20768
rect 26092 20728 26132 20768
rect 27532 20728 27572 20768
rect 29164 20728 29195 20768
rect 29195 20728 29204 20768
rect 29932 20728 29972 20768
rect 30508 20728 30548 20768
rect 19564 20644 19604 20684
rect 19756 20644 19796 20684
rect 21580 20644 21620 20684
rect 22732 20644 22772 20684
rect 24364 20644 24404 20684
rect 25900 20644 25940 20684
rect 28108 20644 28148 20684
rect 28972 20644 29012 20684
rect 30220 20644 30260 20684
rect 11596 20560 11636 20600
rect 11884 20560 11924 20600
rect 12844 20560 12884 20600
rect 13900 20560 13940 20600
rect 15724 20560 15764 20600
rect 17164 20560 17204 20600
rect 17932 20560 17972 20600
rect 18124 20560 18155 20600
rect 18155 20560 18164 20600
rect 18988 20560 19028 20600
rect 19276 20560 19316 20600
rect 20236 20560 20276 20600
rect 21292 20560 21307 20600
rect 21307 20560 21332 20600
rect 21676 20560 21716 20600
rect 22636 20560 22676 20600
rect 25036 20560 25067 20600
rect 25067 20560 25076 20600
rect 25420 20560 25460 20600
rect 8140 20476 8180 20516
rect 9388 20476 9428 20516
rect 9676 20476 9716 20516
rect 21388 20476 21428 20516
rect 6220 20392 6260 20432
rect 8620 20392 8660 20432
rect 11884 20392 11924 20432
rect 12126 20392 12494 20432
rect 17068 20392 17108 20432
rect 18988 20392 19028 20432
rect 19660 20392 19700 20432
rect 19900 20392 20268 20432
rect 5068 20308 5108 20348
rect 5452 20308 5492 20348
rect 13420 20308 13460 20348
rect 13804 20308 13844 20348
rect 15148 20308 15188 20348
rect 20620 20308 20660 20348
rect 7660 20224 7700 20264
rect 8908 20224 8948 20264
rect 9580 20224 9611 20264
rect 9611 20224 9620 20264
rect 10636 20224 10676 20264
rect 11884 20224 11924 20264
rect 3244 20140 3284 20180
rect 5068 20140 5108 20180
rect 5452 20140 5492 20180
rect 9676 20140 9716 20180
rect 9964 20140 10004 20180
rect 1132 20056 1172 20096
rect 1804 20056 1811 20096
rect 1811 20056 1844 20096
rect 2092 20056 2132 20096
rect 2572 20056 2583 20096
rect 2583 20056 2612 20096
rect 3340 20056 3380 20096
rect 3724 20087 3764 20096
rect 3724 20056 3764 20087
rect 4492 20056 4532 20096
rect 1516 19972 1556 20012
rect 1708 19972 1748 20012
rect 2956 19972 2996 20012
rect 3820 19972 3860 20012
rect 4012 19972 4052 20012
rect 4396 19972 4436 20012
rect 4684 19972 4715 20012
rect 4715 19972 4724 20012
rect 2092 19888 2132 19928
rect 5164 19972 5204 20012
rect 5548 19972 5588 20012
rect 5740 19972 5780 20012
rect 12556 20140 12596 20180
rect 13036 20140 13076 20180
rect 13324 20140 13364 20180
rect 23500 20476 23540 20516
rect 30412 20476 30452 20516
rect 27674 20392 28042 20432
rect 21580 20308 21620 20348
rect 15724 20224 15764 20264
rect 16108 20224 16148 20264
rect 16876 20224 16916 20264
rect 17260 20224 17300 20264
rect 17836 20224 17876 20264
rect 18604 20224 18644 20264
rect 19564 20224 19604 20264
rect 19756 20224 19796 20264
rect 21388 20224 21428 20264
rect 14572 20140 14612 20180
rect 16204 20140 16244 20180
rect 6700 20056 6740 20096
rect 7180 20056 7220 20096
rect 7468 20056 7508 20096
rect 8332 20056 8372 20096
rect 8716 20056 8756 20096
rect 9004 20056 9044 20096
rect 10348 20056 10388 20096
rect 11596 20056 11636 20096
rect 11980 20056 12020 20096
rect 12364 20056 12395 20096
rect 12395 20056 12404 20096
rect 12844 20056 12884 20096
rect 14188 20056 14228 20096
rect 16972 20140 17012 20180
rect 5068 19888 5108 19928
rect 5836 19888 5876 19928
rect 1420 19804 1460 19844
rect 1708 19804 1748 19844
rect 2188 19804 2228 19844
rect 3340 19804 3380 19844
rect 5740 19804 5780 19844
rect 5356 19720 5396 19760
rect 3112 19636 3480 19676
rect 460 19384 500 19424
rect 2380 19384 2420 19424
rect 2572 19300 2612 19340
rect 5356 19384 5396 19424
rect 2860 19300 2900 19340
rect 6028 19804 6068 19844
rect 6028 19636 6068 19676
rect 6412 19972 6452 20012
rect 7084 19972 7115 20012
rect 7115 19972 7124 20012
rect 7372 19972 7412 20012
rect 6604 19888 6644 19928
rect 7948 19972 7988 20012
rect 8044 19888 8084 19928
rect 7276 19804 7316 19844
rect 8812 19804 8852 19844
rect 10060 19888 10100 19928
rect 10828 19972 10868 20012
rect 11116 19972 11156 20012
rect 13900 19972 13940 20012
rect 14380 19972 14420 20012
rect 15244 20056 15284 20096
rect 15532 20056 15572 20096
rect 15916 20056 15923 20096
rect 15923 20056 15956 20096
rect 15148 19972 15188 20012
rect 16012 19972 16043 20012
rect 16043 19972 16052 20012
rect 10444 19888 10484 19928
rect 15244 19888 15284 19928
rect 11596 19804 11627 19844
rect 11627 19804 11636 19844
rect 14572 19804 14612 19844
rect 18220 20140 18260 20180
rect 19276 20140 19316 20180
rect 20332 20140 20372 20180
rect 20524 20140 20564 20180
rect 17260 20056 17300 20096
rect 17932 20056 17972 20096
rect 18316 20056 18356 20096
rect 20428 20056 20468 20096
rect 21676 20056 21716 20096
rect 16684 19972 16724 20012
rect 18028 19972 18068 20012
rect 17356 19888 17396 19928
rect 16876 19804 16916 19844
rect 18700 19972 18740 20012
rect 12556 19720 12596 19760
rect 15820 19720 15860 19760
rect 17644 19720 17684 19760
rect 17932 19720 17972 19760
rect 19084 19972 19124 20012
rect 19564 19972 19604 20012
rect 30700 20308 30740 20348
rect 24364 20224 24404 20264
rect 27244 20224 27284 20264
rect 29932 20224 29972 20264
rect 22732 20140 22772 20180
rect 23884 20140 23924 20180
rect 25420 20140 25460 20180
rect 25612 20140 25652 20180
rect 29164 20140 29204 20180
rect 30220 20140 30260 20180
rect 23116 20056 23156 20096
rect 24076 20056 24116 20096
rect 24364 20056 24404 20096
rect 24748 20056 24788 20096
rect 26284 20056 26324 20096
rect 28204 20056 28244 20096
rect 29068 20087 29108 20096
rect 29068 20056 29099 20087
rect 29099 20056 29108 20087
rect 29836 20056 29876 20096
rect 22636 19972 22667 20012
rect 22667 19972 22676 20012
rect 19276 19888 19316 19928
rect 20332 19888 20372 19928
rect 21772 19888 21812 19928
rect 24172 19972 24212 20012
rect 27340 19972 27380 20012
rect 28108 19972 28148 20012
rect 25900 19888 25940 19928
rect 29548 19888 29588 19928
rect 29932 19888 29972 19928
rect 19084 19804 19124 19844
rect 22924 19804 22964 19844
rect 26092 19804 26132 19844
rect 26860 19804 26900 19844
rect 27148 19804 27188 19844
rect 21196 19720 21236 19760
rect 6508 19636 6548 19676
rect 8716 19636 8756 19676
rect 10886 19636 11254 19676
rect 13420 19636 13460 19676
rect 15436 19636 15476 19676
rect 18660 19636 19028 19676
rect 24460 19636 24500 19676
rect 7084 19552 7124 19592
rect 9004 19552 9044 19592
rect 15340 19552 15380 19592
rect 16012 19552 16052 19592
rect 23116 19552 23156 19592
rect 25324 19552 25364 19592
rect 25516 19552 25556 19592
rect 26434 19636 26802 19676
rect 25708 19552 25748 19592
rect 7948 19468 7988 19508
rect 8332 19468 8372 19508
rect 10444 19468 10484 19508
rect 5644 19300 5684 19340
rect 6700 19384 6740 19424
rect 7276 19384 7316 19424
rect 7756 19384 7796 19424
rect 8524 19384 8564 19424
rect 556 19216 596 19256
rect 1612 19216 1643 19256
rect 1643 19216 1652 19256
rect 2284 19216 2324 19256
rect 3820 19216 3860 19256
rect 4204 19216 4244 19256
rect 5452 19216 5492 19256
rect 5740 19216 5780 19256
rect 6028 19216 6068 19256
rect 1900 19132 1940 19172
rect 3148 19132 3177 19172
rect 3177 19132 3188 19172
rect 3532 19132 3572 19172
rect 4588 19132 4628 19172
rect 4780 19132 4820 19172
rect 2092 18880 2132 18920
rect 2476 18880 2516 18920
rect 6508 19300 6548 19340
rect 7084 19300 7124 19340
rect 9484 19384 9524 19424
rect 6412 19216 6452 19256
rect 8908 19300 8948 19340
rect 9580 19300 9620 19340
rect 8332 19216 8348 19256
rect 8348 19216 8372 19256
rect 9004 19216 9044 19256
rect 9388 19216 9428 19256
rect 9772 19216 9803 19256
rect 9803 19216 9812 19256
rect 10732 19384 10772 19424
rect 5836 19132 5876 19172
rect 6988 19132 7028 19172
rect 7372 19132 7412 19172
rect 7948 19132 7988 19172
rect 11788 19468 11828 19508
rect 12844 19468 12884 19508
rect 15052 19468 15092 19508
rect 16684 19468 16715 19508
rect 16715 19468 16724 19508
rect 16876 19468 16916 19508
rect 20716 19468 20756 19508
rect 22348 19468 22388 19508
rect 10924 19216 10964 19256
rect 11692 19384 11732 19424
rect 12748 19384 12788 19424
rect 13036 19300 13076 19340
rect 14956 19300 14996 19340
rect 20524 19384 20564 19424
rect 22156 19384 22196 19424
rect 23308 19384 23348 19424
rect 24076 19384 24116 19424
rect 26860 19384 26900 19424
rect 17260 19300 17300 19340
rect 17932 19300 17972 19340
rect 22924 19300 22964 19340
rect 23692 19300 23732 19340
rect 26380 19300 26420 19340
rect 11788 19216 11828 19256
rect 12652 19216 12692 19256
rect 13228 19216 13268 19256
rect 13804 19216 13844 19256
rect 14188 19216 14228 19256
rect 14572 19216 14574 19256
rect 14574 19216 14612 19256
rect 15532 19216 15572 19256
rect 16300 19216 16340 19256
rect 16588 19216 16628 19256
rect 16780 19216 16820 19256
rect 17836 19216 17876 19256
rect 18988 19247 19028 19256
rect 18988 19216 19028 19247
rect 21196 19216 21236 19256
rect 22156 19216 22196 19256
rect 22540 19216 22580 19256
rect 23116 19216 23156 19256
rect 24076 19216 24116 19256
rect 24460 19216 24500 19256
rect 8620 19132 8660 19172
rect 9676 19132 9716 19172
rect 11596 19132 11636 19172
rect 13132 19132 13172 19172
rect 15244 19132 15273 19172
rect 15273 19132 15284 19172
rect 15724 19132 15764 19172
rect 16684 19132 16713 19172
rect 16713 19132 16724 19172
rect 17068 19132 17108 19172
rect 17356 19132 17396 19172
rect 17644 19132 17684 19172
rect 18220 19132 18260 19172
rect 3820 19048 3860 19088
rect 4396 19048 4436 19088
rect 7084 19048 7124 19088
rect 7564 19048 7604 19088
rect 7756 19048 7796 19088
rect 4204 18964 4244 19004
rect 4352 18880 4720 18920
rect 2860 18796 2900 18836
rect 556 18628 596 18668
rect 1804 18712 1844 18752
rect 1420 18628 1460 18668
rect 3340 18712 3380 18752
rect 3724 18712 3764 18752
rect 4780 18712 4820 18752
rect 2380 18628 2420 18668
rect 3052 18628 3092 18668
rect 6508 18964 6548 19004
rect 8332 18964 8372 19004
rect 8524 18964 8564 19004
rect 8908 18964 8948 19004
rect 6412 18880 6452 18920
rect 5164 18712 5204 18752
rect 5452 18712 5492 18752
rect 5548 18628 5588 18668
rect 5740 18628 5780 18668
rect 6316 18712 6356 18752
rect 6796 18880 6836 18920
rect 7660 18880 7700 18920
rect 9772 19048 9812 19088
rect 10060 19048 10100 19088
rect 10732 19048 10763 19088
rect 10763 19048 10772 19088
rect 11404 19048 11444 19088
rect 11692 19048 11732 19088
rect 13516 19048 13556 19088
rect 14764 19048 14804 19088
rect 15052 19048 15083 19088
rect 15083 19048 15092 19088
rect 15340 19048 15380 19088
rect 15916 19048 15956 19088
rect 16396 19048 16436 19088
rect 9100 18964 9140 19004
rect 10828 18964 10868 19004
rect 11308 18964 11348 19004
rect 12940 18964 12980 19004
rect 15532 18964 15572 19004
rect 16684 18964 16724 19004
rect 18700 19132 18740 19172
rect 20428 19132 20468 19172
rect 20908 19132 20948 19172
rect 19468 18964 19508 19004
rect 9292 18880 9332 18920
rect 10540 18880 10580 18920
rect 11404 18880 11444 18920
rect 12126 18880 12494 18920
rect 15436 18880 15476 18920
rect 17548 18880 17588 18920
rect 19900 18880 20268 18920
rect 8044 18796 8084 18836
rect 10828 18796 10868 18836
rect 14956 18796 14996 18836
rect 7180 18712 7220 18752
rect 7948 18712 7988 18752
rect 9676 18712 9716 18752
rect 10444 18712 10484 18752
rect 10924 18712 10964 18752
rect 12556 18712 12596 18752
rect 13516 18712 13556 18752
rect 15244 18712 15284 18752
rect 6220 18628 6260 18668
rect 7276 18628 7316 18668
rect 1708 18544 1748 18584
rect 1900 18544 1925 18584
rect 1925 18544 1940 18584
rect 3148 18544 3188 18584
rect 1516 18460 1556 18500
rect 1804 18460 1827 18500
rect 1827 18460 1844 18500
rect 2092 18460 2132 18500
rect 2380 18460 2420 18500
rect 1228 18376 1268 18416
rect 2476 18376 2516 18416
rect 2668 18376 2708 18416
rect 3532 18544 3572 18584
rect 4012 18544 4052 18584
rect 5644 18544 5684 18584
rect 6604 18544 6644 18584
rect 9964 18628 10004 18668
rect 10348 18628 10388 18668
rect 13612 18628 13652 18668
rect 16204 18796 16244 18836
rect 16972 18712 17012 18752
rect 19564 18796 19604 18836
rect 22348 19132 22388 19172
rect 23404 19132 23444 19172
rect 23692 19132 23732 19172
rect 25324 19216 25364 19256
rect 26668 19216 26708 19256
rect 24844 19132 24884 19172
rect 22156 19048 22196 19088
rect 23020 19048 23060 19088
rect 23500 19048 23540 19088
rect 27436 19300 27476 19340
rect 27148 19216 27188 19256
rect 28684 19384 28724 19424
rect 24940 19048 24980 19088
rect 23788 18964 23828 19004
rect 24556 18964 24596 19004
rect 27532 18964 27572 19004
rect 20716 18880 20756 18920
rect 27674 18880 28042 18920
rect 29164 19048 29204 19088
rect 29548 19048 29588 19088
rect 25996 18796 26036 18836
rect 18604 18712 18644 18752
rect 18988 18712 19028 18752
rect 22540 18712 22580 18752
rect 24460 18712 24500 18752
rect 27436 18712 27476 18752
rect 16588 18628 16628 18668
rect 17260 18628 17300 18668
rect 18796 18628 18836 18668
rect 19180 18628 19220 18668
rect 24940 18628 24980 18668
rect 28684 18628 28724 18668
rect 2764 18292 2804 18332
rect 5164 18460 5204 18500
rect 5548 18460 5588 18500
rect 6796 18460 6836 18500
rect 5452 18376 5492 18416
rect 3112 18124 3480 18164
rect 2380 18040 2420 18080
rect 748 17956 779 17996
rect 779 17956 788 17996
rect 3724 17956 3764 17996
rect 1516 17872 1556 17912
rect 1996 17872 2036 17912
rect 2380 17872 2420 17912
rect 4876 17872 4916 17912
rect 1804 17788 1844 17828
rect 2284 17788 2324 17828
rect 940 17704 980 17744
rect 1132 17704 1172 17744
rect 1612 17704 1652 17744
rect 2860 17704 2900 17744
rect 3244 17704 3284 17744
rect 940 17452 980 17492
rect 1804 17452 1844 17492
rect 3724 17704 3764 17744
rect 4780 17788 4820 17828
rect 2668 17620 2708 17660
rect 2956 17620 2996 17660
rect 3148 17620 3188 17660
rect 6412 18208 6452 18248
rect 7660 18544 7700 18584
rect 8044 18544 8063 18584
rect 8063 18544 8084 18584
rect 8428 18544 8468 18584
rect 9100 18544 9140 18584
rect 9484 18544 9524 18584
rect 10732 18544 10772 18584
rect 13132 18544 13172 18584
rect 13516 18544 13547 18584
rect 13547 18544 13556 18584
rect 13804 18544 13844 18584
rect 14284 18544 14324 18584
rect 14764 18544 14804 18584
rect 8140 18460 8180 18500
rect 7660 18376 7700 18416
rect 7948 18376 7988 18416
rect 7564 18292 7604 18332
rect 8620 18460 8660 18500
rect 9388 18460 9428 18500
rect 10156 18460 10196 18500
rect 11020 18460 11060 18500
rect 14956 18544 14996 18584
rect 15436 18544 15476 18584
rect 16204 18544 16244 18584
rect 13324 18460 13364 18500
rect 14188 18460 14219 18500
rect 14219 18460 14228 18500
rect 14380 18460 14420 18500
rect 15244 18460 15284 18500
rect 15724 18460 15764 18500
rect 16684 18460 16724 18500
rect 16876 18460 16916 18500
rect 9196 18376 9236 18416
rect 10540 18376 10580 18416
rect 10732 18376 10772 18416
rect 11500 18376 11540 18416
rect 12076 18376 12116 18416
rect 18988 18544 19028 18584
rect 20620 18544 20660 18584
rect 20812 18544 20852 18584
rect 22156 18544 22196 18584
rect 22924 18544 22964 18584
rect 26284 18544 26324 18584
rect 17644 18460 17684 18500
rect 20332 18460 20372 18500
rect 21004 18460 21044 18500
rect 22444 18460 22484 18500
rect 20428 18376 20468 18416
rect 20812 18376 20852 18416
rect 27532 18544 27572 18584
rect 28588 18544 28628 18584
rect 28780 18544 28820 18584
rect 29260 18544 29300 18584
rect 25324 18460 25364 18500
rect 28108 18460 28148 18500
rect 28972 18460 29012 18500
rect 8524 18292 8564 18332
rect 9100 18292 9140 18332
rect 9292 18292 9332 18332
rect 9580 18292 9620 18332
rect 10636 18292 10676 18332
rect 11980 18292 12020 18332
rect 12172 18292 12212 18332
rect 14476 18292 14516 18332
rect 17068 18292 17108 18332
rect 17260 18292 17300 18332
rect 18700 18292 18740 18332
rect 20140 18292 20180 18332
rect 20716 18292 20756 18332
rect 21196 18292 21236 18332
rect 23212 18292 23252 18332
rect 23596 18292 23636 18332
rect 27340 18376 27380 18416
rect 28684 18376 28724 18416
rect 24844 18292 24884 18332
rect 27628 18292 27668 18332
rect 8044 18208 8084 18248
rect 8908 18208 8948 18248
rect 11500 18208 11540 18248
rect 16108 18208 16148 18248
rect 20524 18208 20564 18248
rect 6124 18040 6164 18080
rect 8140 18124 8180 18164
rect 9196 18124 9236 18164
rect 10732 18124 10772 18164
rect 10886 18124 11254 18164
rect 18660 18124 19028 18164
rect 26434 18124 26802 18164
rect 11692 18040 11732 18080
rect 15436 18040 15476 18080
rect 16780 18040 16820 18080
rect 17740 18040 17780 18080
rect 21004 18040 21044 18080
rect 10732 17956 10772 17996
rect 12076 17956 12116 17996
rect 13612 17956 13652 17996
rect 15532 17956 15572 17996
rect 17548 17956 17588 17996
rect 26092 17956 26132 17996
rect 5068 17872 5108 17912
rect 6604 17872 6644 17912
rect 7372 17872 7412 17912
rect 7564 17872 7604 17912
rect 8716 17872 8756 17912
rect 12844 17872 12884 17912
rect 14188 17872 14228 17912
rect 14764 17872 14804 17912
rect 20332 17872 20372 17912
rect 27436 17872 27476 17912
rect 28012 17872 28052 17912
rect 5452 17788 5492 17828
rect 5836 17788 5876 17828
rect 6508 17788 6548 17828
rect 6700 17788 6740 17828
rect 7756 17788 7796 17828
rect 2380 17536 2420 17576
rect 2860 17536 2900 17576
rect 2572 17452 2612 17492
rect 3628 17452 3668 17492
rect 12268 17788 12291 17828
rect 12291 17788 12308 17828
rect 12460 17788 12500 17828
rect 12652 17788 12692 17828
rect 6220 17704 6229 17744
rect 6229 17704 6260 17744
rect 6988 17704 7019 17744
rect 7019 17704 7028 17744
rect 7276 17704 7300 17744
rect 7300 17704 7316 17744
rect 8620 17704 8660 17744
rect 9196 17704 9236 17744
rect 5068 17620 5108 17660
rect 4780 17536 4820 17576
rect 5452 17620 5492 17660
rect 6412 17620 6452 17660
rect 7564 17620 7604 17660
rect 11308 17704 11348 17744
rect 11788 17704 11828 17744
rect 12076 17704 12116 17744
rect 13324 17704 13364 17744
rect 13612 17704 13652 17744
rect 8044 17620 8084 17660
rect 8908 17620 8948 17660
rect 9676 17620 9716 17660
rect 11212 17620 11252 17660
rect 11404 17620 11444 17660
rect 12172 17620 12212 17660
rect 12940 17620 12980 17660
rect 15820 17788 15860 17828
rect 18028 17788 18068 17828
rect 18892 17788 18932 17828
rect 20812 17788 20852 17828
rect 5548 17536 5588 17576
rect 5740 17536 5780 17576
rect 8524 17536 8564 17576
rect 9868 17536 9908 17576
rect 10156 17536 10196 17576
rect 10540 17536 10580 17576
rect 11500 17536 11540 17576
rect 11980 17536 12020 17576
rect 12268 17536 12308 17576
rect 8908 17452 8948 17492
rect 9772 17452 9812 17492
rect 14476 17704 14492 17744
rect 14492 17704 14516 17744
rect 14572 17620 14612 17660
rect 14764 17620 14804 17660
rect 15340 17620 15380 17660
rect 16204 17704 16244 17744
rect 16588 17704 16628 17744
rect 16780 17704 16811 17744
rect 16811 17704 16820 17744
rect 18988 17704 19028 17744
rect 19468 17704 19508 17744
rect 13036 17536 13076 17576
rect 13228 17536 13268 17576
rect 14284 17536 14315 17576
rect 14315 17536 14324 17576
rect 15244 17536 15284 17576
rect 13324 17452 13364 17492
rect 3052 17368 3092 17408
rect 3820 17368 3860 17408
rect 4352 17368 4720 17408
rect 1228 17284 1268 17324
rect 4876 17284 4916 17324
rect 5548 17368 5588 17408
rect 8524 17284 8564 17324
rect 844 17200 884 17240
rect 2380 17200 2420 17240
rect 3436 17200 3476 17240
rect 5644 17200 5684 17240
rect 6412 17200 6452 17240
rect 9772 17200 9812 17240
rect 940 17116 969 17156
rect 969 17116 980 17156
rect 1420 17116 1460 17156
rect 1612 17116 1652 17156
rect 1900 17116 1940 17156
rect 2476 17116 2516 17156
rect 3148 17116 3188 17156
rect 11884 17368 11924 17408
rect 12126 17368 12494 17408
rect 12556 17284 12596 17324
rect 15148 17284 15188 17324
rect 11788 17200 11828 17240
rect 13228 17200 13268 17240
rect 14092 17200 14123 17240
rect 14123 17200 14132 17240
rect 4780 17116 4820 17156
rect 5068 17116 5108 17156
rect 5836 17116 5876 17156
rect 6220 17116 6260 17156
rect 7372 17116 7412 17156
rect 8332 17116 8372 17156
rect 9292 17116 9332 17156
rect 10732 17116 10772 17156
rect 11404 17116 11444 17156
rect 11980 17116 12020 17156
rect 1516 17032 1556 17072
rect 1420 16948 1460 16988
rect 1996 17032 2036 17048
rect 1996 17008 2036 17032
rect 2572 17032 2612 17072
rect 5452 17032 5492 17072
rect 5740 17032 5747 17072
rect 5747 17032 5780 17072
rect 6316 17032 6356 17072
rect 6700 17032 6740 17072
rect 2092 16906 2132 16946
rect 1708 16864 1748 16904
rect 2668 16948 2708 16988
rect 3532 16948 3572 16988
rect 2476 16864 2516 16904
rect 2956 16864 2996 16904
rect 940 16780 971 16820
rect 971 16780 980 16820
rect 2380 16780 2420 16820
rect 1996 16444 2036 16484
rect 2764 16444 2804 16484
rect 1420 16360 1460 16400
rect 2668 16360 2708 16400
rect 1612 16276 1652 16316
rect 2092 16276 2132 16316
rect 1228 16192 1268 16232
rect 1708 16192 1739 16232
rect 1739 16192 1748 16232
rect 2380 16192 2418 16232
rect 2418 16192 2420 16232
rect 3112 16612 3480 16652
rect 3820 16360 3860 16400
rect 4012 16948 4052 16988
rect 5068 16948 5108 16988
rect 5836 16948 5876 16988
rect 6124 16948 6164 16988
rect 5740 16696 5780 16736
rect 5932 16696 5972 16736
rect 5932 16528 5972 16568
rect 4876 16444 4916 16484
rect 4396 16360 4436 16400
rect 3436 16276 3476 16316
rect 4108 16276 4148 16316
rect 4684 16276 4707 16316
rect 4707 16276 4724 16316
rect 7852 17032 7892 17072
rect 8236 17032 8276 17072
rect 9100 17032 9140 17072
rect 9484 17032 9524 17072
rect 10156 17032 10196 17072
rect 10828 17032 10868 17072
rect 11596 17032 11636 17072
rect 12460 17116 12500 17156
rect 12652 17116 12692 17156
rect 13036 17116 13047 17156
rect 13047 17116 13076 17156
rect 13996 17116 14036 17156
rect 14380 17116 14420 17156
rect 7084 16948 7124 16988
rect 7948 16948 7988 16988
rect 8524 16948 8564 16988
rect 8812 16948 8852 16988
rect 9676 16948 9716 16988
rect 9964 16948 10004 16988
rect 10348 16948 10388 16988
rect 7276 16864 7316 16904
rect 8428 16864 8468 16904
rect 9004 16864 9044 16904
rect 9868 16780 9908 16820
rect 13324 17032 13364 17072
rect 16012 17620 16052 17660
rect 17644 17620 17684 17660
rect 17932 17620 17972 17660
rect 16396 17536 16436 17576
rect 16684 17536 16724 17576
rect 16204 17452 16244 17492
rect 20332 17704 20372 17744
rect 20524 17704 20564 17744
rect 23500 17788 23540 17828
rect 24172 17788 24212 17828
rect 25900 17788 25940 17828
rect 27532 17788 27572 17828
rect 19180 17536 19220 17576
rect 21580 17735 21620 17744
rect 21580 17704 21620 17735
rect 21868 17704 21908 17744
rect 22060 17704 22100 17744
rect 23116 17704 23156 17744
rect 23788 17704 23828 17744
rect 24460 17704 24500 17744
rect 25708 17704 25720 17744
rect 25720 17704 25748 17744
rect 22636 17620 22676 17660
rect 23308 17620 23348 17660
rect 24940 17620 24980 17660
rect 27052 17620 27092 17660
rect 20140 17536 20180 17576
rect 20524 17536 20564 17576
rect 22156 17536 22196 17576
rect 22444 17536 22475 17576
rect 22475 17536 22484 17576
rect 23212 17536 23252 17576
rect 23500 17536 23540 17576
rect 27340 17536 27380 17576
rect 18700 17452 18740 17492
rect 20620 17452 20660 17492
rect 23596 17452 23636 17492
rect 19900 17368 20268 17408
rect 27674 17368 28042 17408
rect 21868 17284 21908 17324
rect 16876 17200 16916 17240
rect 19564 17200 19604 17240
rect 19852 17200 19892 17240
rect 15148 17116 15188 17156
rect 14284 17032 14324 17072
rect 11692 16948 11732 16988
rect 12364 16948 12404 16988
rect 11500 16864 11540 16904
rect 12556 16864 12596 16904
rect 13804 16780 13844 16820
rect 16012 17116 16052 17156
rect 16492 17116 16532 17156
rect 16780 17116 16820 17156
rect 17836 17116 17876 17156
rect 18220 17116 18260 17156
rect 20332 17200 20372 17240
rect 20428 17116 20468 17156
rect 22444 17116 22484 17156
rect 17740 17032 17780 17072
rect 18700 17032 18740 17072
rect 14380 16948 14420 16988
rect 15244 16948 15284 16988
rect 15532 16948 15572 16988
rect 14764 16864 14804 16904
rect 16300 16948 16340 16988
rect 16492 16948 16532 16988
rect 16972 16948 17012 16988
rect 17164 16948 17204 16988
rect 19180 17032 19220 17072
rect 19468 17032 19508 17072
rect 19948 17032 19988 17072
rect 20620 17032 20660 17072
rect 20908 17032 20939 17072
rect 20939 17032 20948 17072
rect 22156 17032 22196 17072
rect 23020 17032 23060 17072
rect 23500 17032 23540 17072
rect 19564 16948 19604 16988
rect 21868 16948 21908 16988
rect 25708 17200 25748 17240
rect 25900 17200 25940 17240
rect 28492 17200 28532 17240
rect 24460 17116 24500 17156
rect 27340 17116 27380 17156
rect 24556 17032 24596 17072
rect 25132 17032 25172 17072
rect 25324 17032 25364 17072
rect 27532 17032 27572 17072
rect 24364 16948 24404 16988
rect 24844 16948 24884 16988
rect 25036 16948 25076 16988
rect 26284 16948 26324 16988
rect 27436 16948 27476 16988
rect 17740 16864 17780 16904
rect 19756 16864 19796 16904
rect 21580 16864 21620 16904
rect 15628 16780 15668 16820
rect 16012 16780 16052 16820
rect 17932 16780 17972 16820
rect 20140 16780 20180 16820
rect 21868 16780 21908 16820
rect 24748 16780 24788 16820
rect 26188 16780 26228 16820
rect 28108 16780 28148 16820
rect 13036 16696 13076 16736
rect 13420 16696 13460 16736
rect 19948 16696 19988 16736
rect 8332 16612 8372 16652
rect 10444 16612 10484 16652
rect 8524 16528 8564 16568
rect 10156 16528 10196 16568
rect 5164 16360 5204 16400
rect 7372 16444 7412 16484
rect 7276 16360 7316 16400
rect 5548 16276 5588 16316
rect 5836 16276 5876 16316
rect 6316 16276 6339 16316
rect 6339 16276 6356 16316
rect 6700 16276 6740 16316
rect 10886 16612 11254 16652
rect 16108 16612 16148 16652
rect 18660 16612 19028 16652
rect 21292 16612 21332 16652
rect 25324 16612 25364 16652
rect 26434 16612 26802 16652
rect 11596 16528 11636 16568
rect 7660 16360 7700 16400
rect 8236 16360 8276 16400
rect 10444 16360 10484 16400
rect 10636 16391 10676 16400
rect 10636 16360 10644 16391
rect 10644 16360 10676 16391
rect 7180 16276 7220 16316
rect 8524 16276 8564 16316
rect 11692 16360 11732 16400
rect 11020 16276 11060 16316
rect 13324 16528 13364 16568
rect 16012 16528 16052 16568
rect 19756 16528 19796 16568
rect 23020 16528 23060 16568
rect 25420 16528 25460 16568
rect 15628 16444 15659 16484
rect 15659 16444 15668 16484
rect 17452 16444 17492 16484
rect 19372 16444 19412 16484
rect 22156 16444 22196 16484
rect 22348 16444 22388 16484
rect 23500 16444 23540 16484
rect 28300 16444 28340 16484
rect 13420 16360 13460 16400
rect 13804 16360 13844 16400
rect 14188 16360 14228 16400
rect 11884 16276 11924 16316
rect 4396 16192 4436 16232
rect 6604 16192 6644 16232
rect 8236 16192 8276 16232
rect 8812 16192 8843 16232
rect 8843 16192 8852 16232
rect 10444 16192 10484 16232
rect 10732 16192 10772 16232
rect 11212 16192 11252 16232
rect 11788 16192 11828 16232
rect 11980 16192 12005 16232
rect 12005 16192 12020 16232
rect 2572 16108 2601 16148
rect 2601 16108 2612 16148
rect 3628 16108 3668 16148
rect 4492 16108 4532 16148
rect 1420 16024 1451 16064
rect 1451 16024 1460 16064
rect 2764 16024 2804 16064
rect 3340 16024 3380 16064
rect 5068 16108 5108 16148
rect 6316 16108 6356 16148
rect 6988 16108 7028 16148
rect 6124 16024 6164 16064
rect 6796 16024 6836 16064
rect 2956 15940 2996 15980
rect 5164 15940 5204 15980
rect 6220 15940 6260 15980
rect 2476 15856 2516 15896
rect 4352 15856 4720 15896
rect 2572 15772 2612 15812
rect 1036 15688 1076 15728
rect 1708 15688 1748 15728
rect 3436 15688 3476 15728
rect 4012 15688 4043 15728
rect 4043 15688 4052 15728
rect 1420 15604 1460 15644
rect 2284 15604 2324 15644
rect 2668 15604 2708 15644
rect 2860 15604 2900 15644
rect 3340 15604 3380 15644
rect 7756 16108 7796 16148
rect 7948 16108 7988 16148
rect 9100 16108 9140 16148
rect 9676 16108 9716 16148
rect 9964 16108 10004 16148
rect 10252 16108 10292 16148
rect 12652 16276 12692 16316
rect 12460 16192 12500 16232
rect 12940 16192 12980 16232
rect 7564 16024 7604 16064
rect 9484 16024 9524 16064
rect 6988 15940 7028 15980
rect 11308 15940 11348 15980
rect 11596 15940 11636 15980
rect 13708 16276 13748 16316
rect 14092 16276 14132 16316
rect 15820 16360 15860 16400
rect 15532 16276 15572 16316
rect 16108 16276 16148 16316
rect 13324 16108 13364 16148
rect 13516 16108 13556 16148
rect 14476 16192 14516 16232
rect 14668 16192 14708 16232
rect 16684 16276 16724 16316
rect 17260 16276 17300 16316
rect 17644 16276 17684 16316
rect 20428 16360 20468 16400
rect 21484 16360 21524 16400
rect 22252 16360 22292 16400
rect 25420 16360 25460 16400
rect 26188 16360 26228 16400
rect 19372 16276 19412 16316
rect 20236 16276 20276 16316
rect 22348 16276 22388 16316
rect 22828 16276 22868 16316
rect 23596 16276 23636 16316
rect 25708 16276 25748 16316
rect 26860 16276 26900 16316
rect 16876 16192 16905 16232
rect 16905 16192 16916 16232
rect 17452 16192 17471 16232
rect 17471 16192 17492 16232
rect 17836 16192 17876 16232
rect 18508 16192 18520 16232
rect 18520 16192 18548 16232
rect 19852 16223 19892 16232
rect 19852 16192 19883 16223
rect 19883 16192 19892 16223
rect 20908 16192 20948 16232
rect 21196 16192 21227 16232
rect 21227 16192 21236 16232
rect 14380 16108 14420 16148
rect 15628 16108 15668 16148
rect 13612 16024 13643 16064
rect 13643 16024 13652 16064
rect 12940 15940 12980 15980
rect 13324 15940 13364 15980
rect 13708 15940 13748 15980
rect 14668 15940 14708 15980
rect 7852 15856 7892 15896
rect 8812 15856 8852 15896
rect 12126 15856 12494 15896
rect 14284 15856 14324 15896
rect 4876 15772 4916 15812
rect 5356 15688 5396 15728
rect 5740 15688 5780 15728
rect 7660 15772 7700 15812
rect 8524 15772 8564 15812
rect 5164 15604 5204 15644
rect 5452 15604 5492 15644
rect 6124 15604 6164 15644
rect 6412 15604 6452 15644
rect 7756 15688 7796 15728
rect 7372 15604 7412 15644
rect 7660 15604 7700 15644
rect 8044 15688 8084 15728
rect 8428 15688 8468 15728
rect 8620 15688 8660 15728
rect 10444 15688 10484 15728
rect 10636 15688 10676 15728
rect 16108 16108 16148 16148
rect 16492 16108 16532 16148
rect 15436 16024 15476 16064
rect 17548 16108 17588 16148
rect 20332 16108 20372 16148
rect 21292 16108 21332 16148
rect 21964 16108 22004 16148
rect 16972 16024 17012 16064
rect 18604 16024 18644 16064
rect 19756 16024 19796 16064
rect 22060 16024 22100 16064
rect 23500 16192 23531 16232
rect 23531 16192 23540 16232
rect 27628 16276 27668 16316
rect 28780 16360 28820 16400
rect 23692 16108 23732 16148
rect 25228 16192 25268 16232
rect 25900 16192 25940 16232
rect 26476 16192 26516 16232
rect 26764 16192 26804 16232
rect 28300 16192 28340 16232
rect 24556 16108 24596 16148
rect 23500 16024 23540 16064
rect 24268 16024 24308 16064
rect 25708 16024 25748 16064
rect 28108 16024 28148 16064
rect 28492 16024 28532 16064
rect 16012 15940 16052 15980
rect 16492 15940 16532 15980
rect 16876 15940 16916 15980
rect 18028 15940 18068 15980
rect 19564 15940 19604 15980
rect 21964 15940 22004 15980
rect 16204 15856 16244 15896
rect 19900 15856 20268 15896
rect 23788 15856 23828 15896
rect 13132 15772 13172 15812
rect 8524 15604 8564 15644
rect 8716 15604 8756 15644
rect 9388 15604 9428 15644
rect 9772 15604 9812 15644
rect 9964 15604 10004 15644
rect 652 15520 692 15560
rect 1228 15520 1268 15560
rect 1612 15520 1652 15560
rect 1516 15352 1556 15392
rect 3820 15520 3860 15560
rect 4396 15520 4436 15560
rect 5548 15520 5588 15560
rect 6220 15520 6251 15560
rect 6251 15520 6260 15560
rect 6796 15520 6836 15560
rect 7084 15520 7124 15560
rect 2380 15436 2420 15476
rect 2956 15436 2996 15476
rect 2572 15352 2612 15392
rect 4300 15436 4331 15476
rect 4331 15436 4340 15476
rect 3820 15268 3860 15308
rect 2476 15184 2516 15224
rect 4780 15184 4820 15224
rect 3112 15100 3480 15140
rect 4012 15100 4052 15140
rect 5932 15436 5955 15476
rect 5955 15436 5972 15476
rect 6412 15436 6452 15476
rect 8428 15436 8468 15476
rect 6316 15352 6356 15392
rect 7852 15352 7892 15392
rect 5548 15268 5588 15308
rect 5740 15268 5780 15308
rect 6700 15268 6740 15308
rect 8812 15268 8852 15308
rect 10924 15604 10964 15644
rect 11308 15604 11348 15644
rect 13228 15688 13268 15728
rect 13516 15688 13556 15728
rect 15436 15688 15476 15728
rect 9100 15520 9140 15560
rect 10252 15520 10277 15560
rect 10277 15520 10292 15560
rect 11116 15520 11132 15560
rect 11132 15520 11156 15560
rect 9676 15436 9716 15476
rect 8524 15184 8564 15224
rect 10348 15436 10388 15476
rect 10540 15436 10580 15476
rect 10732 15436 10772 15476
rect 14284 15604 14324 15644
rect 15148 15604 15188 15644
rect 15628 15604 15668 15644
rect 17836 15772 17876 15812
rect 18412 15772 18452 15812
rect 21676 15772 21716 15812
rect 24268 15772 24308 15812
rect 17260 15688 17300 15728
rect 18316 15688 18356 15728
rect 20428 15688 20468 15728
rect 21964 15688 22004 15728
rect 22348 15688 22379 15728
rect 22379 15688 22388 15728
rect 23020 15688 23060 15728
rect 23308 15688 23348 15728
rect 24940 15688 24980 15728
rect 25900 15688 25940 15728
rect 17932 15604 17972 15644
rect 18220 15604 18260 15644
rect 19180 15604 19220 15644
rect 19372 15604 19412 15644
rect 19852 15604 19892 15644
rect 22156 15604 22196 15644
rect 22636 15604 22676 15644
rect 22924 15604 22964 15644
rect 11884 15520 11907 15560
rect 11907 15520 11924 15560
rect 12172 15520 12212 15560
rect 11500 15352 11540 15392
rect 10348 15268 10388 15308
rect 9484 15184 9524 15224
rect 10540 15184 10580 15224
rect 9388 15100 9428 15140
rect 10444 15100 10484 15140
rect 10886 15100 11254 15140
rect 9484 15016 9524 15056
rect 11596 15016 11636 15056
rect 1804 14932 1844 14972
rect 4876 14932 4916 14972
rect 1036 14764 1067 14804
rect 1067 14764 1076 14804
rect 2092 14764 2132 14804
rect 4396 14764 4436 14804
rect 6700 14932 6740 14972
rect 7084 14932 7124 14972
rect 5836 14764 5876 14804
rect 6412 14764 6443 14804
rect 6443 14764 6452 14804
rect 6796 14764 6836 14804
rect 2668 14680 2708 14720
rect 3148 14680 3188 14720
rect 3628 14680 3668 14720
rect 4204 14680 4244 14720
rect 4588 14680 4628 14720
rect 5548 14680 5588 14720
rect 5932 14680 5972 14720
rect 3724 14596 3764 14636
rect 4108 14596 4148 14636
rect 652 14512 692 14552
rect 2668 14512 2708 14552
rect 3628 14512 3668 14552
rect 7180 14848 7220 14888
rect 8524 14848 8564 14888
rect 9196 14848 9236 14888
rect 11020 14848 11060 14888
rect 12364 15268 12395 15308
rect 12395 15268 12404 15308
rect 12940 15520 12980 15560
rect 14380 15520 14401 15560
rect 14401 15520 14420 15560
rect 14668 15520 14693 15560
rect 14693 15520 14708 15560
rect 15244 15520 15284 15560
rect 17260 15520 17300 15560
rect 13708 15436 13748 15476
rect 14284 15436 14324 15476
rect 12844 15352 12884 15392
rect 12940 15268 12980 15308
rect 13420 15268 13460 15308
rect 14188 15268 14228 15308
rect 13996 15184 14036 15224
rect 18700 15520 18740 15560
rect 19084 15520 19124 15560
rect 19948 15520 19988 15560
rect 20428 15520 20468 15560
rect 20908 15520 20948 15560
rect 21292 15520 21332 15560
rect 21868 15520 21908 15560
rect 22252 15520 22292 15560
rect 27674 15856 28042 15896
rect 28300 15772 28340 15812
rect 28780 15772 28820 15812
rect 26956 15688 26996 15728
rect 23692 15604 23732 15644
rect 27532 15604 27572 15644
rect 23788 15520 23828 15560
rect 24748 15520 24788 15560
rect 25420 15520 25460 15560
rect 25708 15520 25748 15560
rect 26764 15520 26804 15560
rect 27820 15520 27851 15560
rect 27851 15520 27860 15560
rect 28108 15520 28148 15560
rect 28396 15551 28436 15560
rect 17932 15436 17972 15476
rect 18412 15436 18452 15476
rect 18604 15436 18644 15476
rect 18892 15436 18923 15476
rect 18923 15436 18932 15476
rect 19756 15436 19796 15476
rect 20812 15436 20852 15476
rect 21484 15436 21524 15476
rect 21964 15436 22004 15476
rect 22540 15436 22580 15476
rect 23500 15436 23540 15476
rect 15244 15352 15284 15392
rect 16492 15352 16532 15392
rect 18028 15352 18068 15392
rect 28396 15520 28427 15551
rect 28427 15520 28436 15551
rect 28780 15520 28820 15560
rect 25228 15436 25268 15476
rect 28300 15436 28340 15476
rect 28492 15436 28532 15476
rect 19180 15352 19220 15392
rect 20044 15352 20084 15392
rect 20428 15352 20468 15392
rect 20716 15352 20756 15392
rect 22444 15352 22484 15392
rect 23884 15352 23924 15392
rect 24364 15352 24404 15392
rect 16396 15268 16436 15308
rect 19276 15268 19316 15308
rect 19564 15268 19604 15308
rect 19756 15268 19796 15308
rect 20524 15268 20564 15308
rect 23980 15268 24020 15308
rect 28972 15268 29012 15308
rect 17452 15184 17492 15224
rect 26284 15184 26324 15224
rect 15148 15100 15188 15140
rect 18660 15100 19028 15140
rect 20044 15100 20084 15140
rect 22252 15100 22292 15140
rect 26434 15100 26802 15140
rect 16300 15016 16340 15056
rect 19564 15016 19604 15056
rect 23308 15016 23348 15056
rect 23788 15016 23828 15056
rect 27148 15016 27188 15056
rect 13324 14932 13364 14972
rect 14956 14932 14996 14972
rect 17932 14932 17972 14972
rect 18124 14932 18164 14972
rect 19084 14932 19124 14972
rect 19756 14932 19796 14972
rect 20812 14932 20852 14972
rect 21964 14932 22004 14972
rect 14860 14848 14900 14888
rect 15628 14848 15668 14888
rect 7660 14764 7691 14804
rect 7691 14764 7700 14804
rect 9004 14764 9044 14804
rect 9292 14764 9332 14804
rect 9484 14764 9524 14804
rect 10060 14764 10100 14804
rect 10540 14764 10563 14804
rect 10563 14764 10580 14804
rect 11116 14764 11156 14804
rect 11980 14764 12020 14804
rect 12748 14764 12788 14804
rect 6700 14680 6740 14720
rect 8620 14680 8660 14720
rect 8908 14680 8948 14720
rect 13996 14764 14036 14804
rect 14764 14764 14804 14804
rect 15052 14764 15092 14804
rect 9676 14680 9716 14720
rect 10156 14680 10196 14720
rect 11692 14680 11732 14720
rect 12172 14680 12212 14720
rect 12844 14680 12884 14720
rect 6604 14596 6644 14636
rect 6988 14596 7028 14636
rect 7564 14596 7604 14636
rect 9580 14596 9620 14636
rect 9772 14596 9812 14636
rect 8236 14512 8276 14552
rect 8620 14512 8659 14552
rect 8659 14512 8660 14552
rect 10636 14596 10676 14636
rect 11116 14596 11156 14636
rect 9100 14512 9140 14552
rect 11020 14512 11060 14552
rect 13612 14680 13652 14720
rect 14188 14680 14228 14720
rect 14572 14680 14612 14720
rect 15148 14680 15188 14720
rect 19468 14848 19508 14888
rect 19948 14848 19988 14888
rect 21004 14848 21044 14888
rect 16684 14764 16724 14804
rect 18316 14764 18356 14804
rect 19756 14764 19796 14804
rect 21100 14764 21140 14804
rect 16108 14680 16137 14720
rect 16137 14680 16148 14720
rect 16396 14680 16436 14720
rect 17260 14680 17300 14720
rect 17452 14680 17483 14720
rect 17483 14680 17492 14720
rect 18604 14680 18644 14720
rect 21580 14764 21620 14804
rect 20524 14680 20535 14720
rect 20535 14680 20564 14720
rect 24076 14932 24116 14972
rect 25900 14932 25940 14972
rect 28396 14932 28436 14972
rect 22540 14764 22580 14804
rect 21676 14680 21716 14720
rect 22252 14680 22292 14720
rect 22444 14680 22469 14720
rect 22469 14680 22484 14720
rect 23308 14764 23348 14804
rect 11500 14596 11540 14636
rect 12460 14596 12500 14636
rect 14284 14596 14324 14636
rect 14764 14596 14804 14636
rect 15436 14596 15476 14636
rect 18220 14596 18260 14636
rect 18892 14596 18932 14636
rect 19084 14596 19124 14636
rect 19468 14596 19508 14636
rect 19852 14596 19892 14636
rect 20908 14596 20948 14636
rect 21580 14596 21620 14636
rect 11596 14512 11636 14552
rect 12748 14512 12788 14552
rect 13804 14512 13844 14552
rect 15244 14512 15284 14552
rect 16300 14512 16340 14552
rect 16684 14512 16724 14552
rect 17260 14512 17300 14552
rect 17644 14512 17684 14552
rect 18796 14512 18836 14552
rect 20140 14512 20180 14552
rect 20716 14512 20756 14552
rect 21196 14512 21227 14552
rect 21227 14512 21236 14552
rect 21676 14512 21716 14552
rect 1420 14428 1460 14468
rect 4780 14428 4820 14468
rect 14860 14428 14900 14468
rect 4352 14344 4720 14384
rect 9100 14344 9140 14384
rect 3244 14260 3284 14300
rect 3916 14260 3956 14300
rect 4204 14260 4244 14300
rect 4876 14260 4916 14300
rect 1228 14176 1268 14216
rect 4972 14176 5012 14216
rect 1612 14092 1652 14132
rect 556 14008 596 14048
rect 1036 14008 1076 14048
rect 1900 14008 1940 14048
rect 2572 14008 2612 14048
rect 2956 14008 2996 14048
rect 3244 14008 3284 14048
rect 5356 14092 5396 14132
rect 940 13924 980 13964
rect 2092 13840 2132 13880
rect 3148 13756 3188 13796
rect 3436 13756 3476 13796
rect 3112 13588 3480 13628
rect 844 13504 884 13544
rect 2572 13420 2603 13460
rect 2603 13420 2612 13460
rect 4684 14008 4724 14048
rect 4300 13924 4340 13964
rect 7468 14260 7508 14300
rect 10348 14260 10388 14300
rect 6508 14176 6548 14216
rect 12126 14344 12494 14384
rect 21964 14596 22004 14636
rect 22924 14680 22964 14720
rect 23692 14764 23732 14804
rect 28876 14848 28916 14888
rect 29836 14848 29876 14888
rect 23884 14680 23924 14720
rect 25132 14680 25172 14720
rect 27148 14764 27188 14804
rect 28684 14680 28724 14720
rect 29644 14680 29684 14720
rect 24652 14596 24683 14636
rect 24683 14596 24692 14636
rect 27820 14596 27860 14636
rect 22060 14512 22100 14552
rect 22348 14512 22388 14552
rect 23116 14512 23156 14552
rect 25516 14512 25556 14552
rect 21388 14428 21428 14468
rect 22540 14428 22580 14468
rect 23308 14428 23348 14468
rect 19900 14344 20268 14384
rect 23596 14344 23636 14384
rect 27674 14344 28042 14384
rect 10636 14260 10676 14300
rect 12748 14260 12788 14300
rect 9388 14176 9428 14216
rect 9676 14176 9716 14216
rect 5644 14092 5684 14132
rect 6124 14092 6164 14132
rect 9580 14092 9620 14132
rect 10156 14092 10196 14132
rect 10636 14092 10676 14132
rect 11308 14092 11348 14132
rect 14380 14176 14420 14216
rect 14668 14176 14708 14216
rect 16300 14176 16340 14216
rect 19180 14176 19220 14216
rect 20140 14176 20180 14216
rect 13516 14092 13556 14132
rect 13708 14092 13748 14132
rect 14764 14092 14804 14132
rect 15244 14092 15284 14132
rect 16012 14092 16052 14132
rect 5740 14008 5780 14048
rect 6604 14008 6644 14048
rect 4876 13924 4916 13964
rect 5836 13924 5876 13964
rect 4204 13840 4244 13880
rect 7756 14008 7760 14048
rect 7760 14008 7796 14048
rect 8044 14008 8084 14048
rect 8332 14008 8372 14048
rect 9292 14008 9332 14048
rect 10060 14008 10100 14048
rect 7180 13924 7220 13964
rect 9580 13924 9611 13964
rect 9611 13924 9620 13964
rect 10252 13924 10292 13964
rect 11404 14008 11444 14048
rect 11884 14008 11924 14048
rect 12268 14008 12308 14048
rect 12748 14008 12779 14048
rect 12779 14008 12788 14048
rect 23212 14260 23252 14300
rect 20620 14176 20660 14216
rect 23884 14176 23924 14216
rect 24172 14176 24203 14216
rect 24203 14176 24212 14216
rect 18700 14092 18740 14132
rect 13996 14008 14036 14048
rect 14476 14008 14516 14048
rect 12460 13924 12500 13964
rect 13324 13924 13364 13964
rect 14572 13924 14612 13964
rect 15052 13924 15083 13964
rect 15083 13924 15092 13964
rect 15628 13924 15651 13964
rect 15651 13924 15668 13964
rect 16396 14008 16436 14048
rect 17644 14008 17684 14048
rect 18220 14008 18260 14048
rect 18412 14008 18452 14048
rect 18796 14008 18836 14048
rect 16780 13924 16786 13964
rect 16786 13924 16820 13964
rect 17740 13924 17780 13964
rect 6508 13840 6548 13880
rect 7468 13840 7508 13880
rect 10156 13840 10196 13880
rect 12940 13840 12980 13880
rect 14284 13840 14324 13880
rect 16012 13840 16052 13880
rect 17644 13840 17684 13880
rect 5836 13756 5876 13796
rect 6220 13756 6260 13796
rect 8524 13756 8564 13796
rect 9772 13756 9812 13796
rect 10252 13756 10292 13796
rect 10540 13756 10580 13796
rect 10828 13756 10868 13796
rect 12364 13756 12404 13796
rect 13516 13756 13556 13796
rect 19468 13966 19508 14006
rect 20524 14092 20564 14132
rect 21580 14092 21620 14132
rect 25996 14176 26036 14216
rect 29644 14176 29684 14216
rect 21868 14092 21908 14132
rect 23596 14092 23636 14132
rect 25324 14092 25364 14132
rect 25900 14092 25940 14132
rect 20044 14008 20084 14048
rect 20812 14008 20852 14048
rect 21388 14008 21428 14048
rect 19756 13840 19796 13880
rect 18796 13756 18836 13796
rect 18988 13756 19028 13796
rect 20236 13924 20276 13964
rect 22060 14008 22100 14048
rect 22444 14008 22484 14048
rect 21196 13924 21236 13964
rect 22156 13924 22196 13964
rect 22732 13924 22772 13964
rect 22828 13840 22868 13880
rect 21196 13756 21236 13796
rect 7468 13672 7508 13712
rect 9868 13672 9908 13712
rect 10156 13672 10196 13712
rect 11884 13672 11924 13712
rect 13324 13672 13364 13712
rect 18412 13672 18452 13712
rect 19180 13672 19220 13712
rect 6412 13588 6452 13628
rect 10886 13588 11254 13628
rect 18660 13588 19028 13628
rect 5932 13420 5972 13460
rect 5068 13336 5108 13376
rect 5836 13252 5867 13292
rect 5867 13252 5876 13292
rect 652 13168 692 13208
rect 1804 13168 1844 13208
rect 2380 13168 2420 13208
rect 2956 13168 2987 13208
rect 2987 13168 2996 13208
rect 3916 13168 3956 13208
rect 4972 13168 5012 13208
rect 5452 13168 5492 13208
rect 6316 13504 6356 13544
rect 8620 13504 8660 13544
rect 14476 13504 14516 13544
rect 22636 13672 22676 13712
rect 19468 13588 19508 13628
rect 20716 13588 20756 13628
rect 20908 13588 20948 13628
rect 20332 13504 20372 13544
rect 20524 13504 20564 13544
rect 11308 13420 11348 13460
rect 12556 13420 12596 13460
rect 13612 13420 13652 13460
rect 14188 13420 14228 13460
rect 14572 13420 14612 13460
rect 15724 13420 15764 13460
rect 19468 13420 19508 13460
rect 19948 13420 19988 13460
rect 20620 13420 20660 13460
rect 20812 13420 20852 13460
rect 21676 13420 21716 13460
rect 6220 13252 6260 13292
rect 23404 14008 23444 14048
rect 23788 14008 23828 14048
rect 24364 14008 24404 14048
rect 24748 14008 24788 14048
rect 25708 14008 25748 14048
rect 27052 14008 27092 14048
rect 27532 14008 27563 14048
rect 27563 14008 27572 14048
rect 23692 13924 23732 13964
rect 26860 13924 26900 13964
rect 29836 13924 29876 13964
rect 28876 13840 28916 13880
rect 23500 13756 23540 13796
rect 24748 13756 24788 13796
rect 25324 13756 25364 13796
rect 29068 13756 29108 13796
rect 24172 13588 24212 13628
rect 26434 13588 26802 13628
rect 22828 13420 22868 13460
rect 23308 13420 23348 13460
rect 23692 13420 23732 13460
rect 24652 13420 24692 13460
rect 7276 13336 7316 13376
rect 18316 13336 18356 13376
rect 18700 13336 18740 13376
rect 20044 13336 20084 13376
rect 21196 13336 21236 13376
rect 22348 13336 22388 13376
rect 6508 13252 6548 13292
rect 7372 13252 7412 13292
rect 7948 13252 7988 13292
rect 8524 13252 8564 13292
rect 10060 13252 10100 13292
rect 10252 13252 10258 13292
rect 10258 13252 10292 13292
rect 11788 13252 11828 13292
rect 12364 13252 12404 13292
rect 13228 13252 13268 13292
rect 13516 13252 13556 13292
rect 13804 13252 13844 13292
rect 14764 13252 14804 13292
rect 15148 13252 15188 13292
rect 16204 13252 16244 13292
rect 16876 13252 16916 13292
rect 6796 13168 6836 13208
rect 7276 13168 7316 13208
rect 1132 13084 1172 13124
rect 4780 13084 4820 13124
rect 5932 13084 5972 13124
rect 6220 13084 6260 13124
rect 7084 13084 7124 13124
rect 7852 13168 7892 13208
rect 8908 13168 8916 13208
rect 8916 13168 8948 13208
rect 9772 13168 9803 13208
rect 9803 13168 9812 13208
rect 10540 13168 10580 13208
rect 11596 13168 11636 13208
rect 12460 13168 12500 13208
rect 14188 13168 14228 13208
rect 14476 13168 14516 13208
rect 15340 13168 15380 13208
rect 15724 13168 15764 13208
rect 1228 13000 1268 13040
rect 6028 13000 6059 13040
rect 6059 13000 6068 13040
rect 6316 13000 6356 13040
rect 7468 13000 7508 13040
rect 8044 13084 8084 13124
rect 10828 13084 10868 13124
rect 11212 13084 11252 13124
rect 11404 13084 11444 13124
rect 12556 13084 12596 13124
rect 13324 13084 13364 13124
rect 13804 13084 13844 13124
rect 14284 13084 14324 13124
rect 17068 13168 17108 13208
rect 17548 13168 17588 13208
rect 15244 13084 15284 13124
rect 15628 13084 15668 13124
rect 16012 13084 16052 13124
rect 18796 13168 18836 13208
rect 17356 13084 17396 13124
rect 17836 13084 17876 13124
rect 19852 13252 19892 13292
rect 20332 13252 20372 13292
rect 20812 13252 20852 13292
rect 22540 13252 22580 13292
rect 28684 13336 28724 13376
rect 23308 13252 23348 13292
rect 24556 13252 24596 13292
rect 24940 13252 24980 13292
rect 25900 13252 25940 13292
rect 28396 13252 28436 13292
rect 21868 13168 21908 13208
rect 22156 13168 22196 13208
rect 19756 13084 19796 13124
rect 20236 13084 20276 13124
rect 20716 13084 20756 13124
rect 10444 13000 10484 13040
rect 11788 13000 11828 13040
rect 12172 13000 12212 13040
rect 12940 13000 12980 13040
rect 13708 13000 13748 13040
rect 14188 13000 14228 13040
rect 15148 13000 15188 13040
rect 21004 13084 21044 13124
rect 23116 13168 23147 13208
rect 23147 13168 23156 13208
rect 23596 13168 23636 13208
rect 28780 13252 28820 13292
rect 24748 13168 24788 13208
rect 25324 13168 25364 13208
rect 27148 13168 27188 13208
rect 27532 13168 27563 13208
rect 27563 13168 27572 13208
rect 28972 13168 29012 13208
rect 21580 13084 21620 13124
rect 22060 13084 22100 13124
rect 22252 13084 22292 13124
rect 22732 13084 22772 13124
rect 23212 13084 23252 13124
rect 23788 13084 23828 13124
rect 23980 13084 24020 13124
rect 24268 13084 24308 13124
rect 24652 13084 24692 13124
rect 25036 13084 25076 13124
rect 25420 13084 25460 13124
rect 28204 13084 28244 13124
rect 21100 13000 21140 13040
rect 23404 13000 23444 13040
rect 27340 13000 27380 13040
rect 3916 12916 3956 12956
rect 7180 12916 7220 12956
rect 11212 12916 11252 12956
rect 19468 12916 19508 12956
rect 19756 12916 19796 12956
rect 22732 12916 22772 12956
rect 4352 12832 4720 12872
rect 652 12748 692 12788
rect 5932 12748 5972 12788
rect 460 12664 500 12704
rect 1804 12664 1844 12704
rect 2956 12664 2996 12704
rect 4780 12664 4820 12704
rect 2380 12580 2420 12620
rect 4492 12580 4532 12620
rect 4972 12580 5012 12620
rect 6796 12748 6836 12788
rect 7564 12748 7604 12788
rect 9676 12748 9716 12788
rect 5836 12664 5876 12704
rect 7084 12664 7124 12704
rect 5548 12580 5588 12620
rect 6796 12580 6836 12620
rect 6988 12580 7028 12620
rect 7180 12580 7220 12620
rect 940 12496 980 12536
rect 1708 12496 1748 12536
rect 2956 12496 2996 12536
rect 3916 12496 3956 12536
rect 4300 12496 4340 12536
rect 5164 12496 5204 12536
rect 6508 12527 6548 12536
rect 6508 12496 6548 12527
rect 28492 12916 28532 12956
rect 12126 12832 12494 12872
rect 13804 12832 13844 12872
rect 16588 12832 16628 12872
rect 19900 12832 20268 12872
rect 27674 12832 28042 12872
rect 16108 12748 16148 12788
rect 17068 12748 17108 12788
rect 21196 12748 21236 12788
rect 9100 12664 9140 12704
rect 9868 12664 9908 12704
rect 11500 12664 11540 12704
rect 8044 12580 8084 12620
rect 8332 12580 8372 12620
rect 8716 12580 8756 12620
rect 9004 12580 9044 12620
rect 11404 12580 11444 12620
rect 12076 12580 12116 12620
rect 12556 12664 12596 12704
rect 13420 12664 13460 12704
rect 13708 12664 13748 12704
rect 13804 12580 13844 12620
rect 14956 12664 14996 12704
rect 16012 12664 16052 12704
rect 16300 12664 16331 12704
rect 16331 12664 16340 12704
rect 16876 12664 16916 12704
rect 17644 12664 17684 12704
rect 19948 12664 19988 12704
rect 20524 12664 20564 12704
rect 21388 12664 21428 12704
rect 24940 12664 24980 12704
rect 14188 12611 14228 12620
rect 14188 12580 14219 12611
rect 14219 12580 14228 12611
rect 15532 12580 15572 12620
rect 15724 12580 15764 12620
rect 16396 12580 16436 12620
rect 17452 12580 17478 12620
rect 17478 12580 17492 12620
rect 19660 12580 19700 12620
rect 22540 12580 22580 12620
rect 3052 12412 3092 12452
rect 4780 12412 4820 12452
rect 7468 12496 7508 12536
rect 9100 12496 9140 12536
rect 9580 12496 9620 12536
rect 11212 12496 11252 12536
rect 6412 12412 6452 12452
rect 6604 12412 6644 12452
rect 7084 12412 7124 12452
rect 8140 12412 8180 12452
rect 8620 12412 8660 12452
rect 10156 12412 10196 12452
rect 11884 12496 11924 12536
rect 12940 12496 12980 12536
rect 12748 12412 12788 12452
rect 10348 12328 10388 12368
rect 13804 12328 13844 12368
rect 7852 12244 7892 12284
rect 8044 12244 8084 12284
rect 9196 12244 9236 12284
rect 9676 12244 9716 12284
rect 10732 12244 10772 12284
rect 13900 12244 13931 12284
rect 13931 12244 13940 12284
rect 3112 12076 3480 12116
rect 6316 12076 6356 12116
rect 12652 12160 12692 12200
rect 5548 11992 5588 12032
rect 1420 11908 1460 11948
rect 6988 11908 7028 11948
rect 7468 11908 7508 11948
rect 1132 11824 1172 11864
rect 3052 11824 3092 11864
rect 1420 11740 1460 11780
rect 2380 11740 2420 11780
rect 3148 11740 3188 11780
rect 4204 11824 4244 11864
rect 6220 11740 6260 11780
rect 6796 11740 6836 11780
rect 7468 11740 7508 11780
rect 8428 11740 8468 11780
rect 10886 12076 11254 12116
rect 12940 11992 12980 12032
rect 9580 11908 9620 11948
rect 12460 11908 12500 11948
rect 12748 11908 12788 11948
rect 10060 11824 10100 11864
rect 10156 11740 10196 11780
rect 12460 11740 12500 11780
rect 13324 12076 13364 12116
rect 15340 12496 15380 12536
rect 16588 12496 16628 12536
rect 16972 12496 17012 12536
rect 17260 12496 17300 12536
rect 25516 12664 25547 12704
rect 25547 12664 25556 12704
rect 18700 12496 18740 12536
rect 18892 12496 18932 12536
rect 19372 12496 19412 12536
rect 19756 12496 19796 12536
rect 20524 12496 20564 12536
rect 20716 12496 20756 12536
rect 21868 12496 21899 12536
rect 21899 12496 21908 12536
rect 25900 12664 25940 12704
rect 26860 12664 26900 12704
rect 27340 12664 27380 12704
rect 28204 12664 28244 12704
rect 25804 12580 25844 12620
rect 26956 12580 26967 12620
rect 26967 12580 26996 12620
rect 27244 12580 27284 12620
rect 27436 12580 27476 12620
rect 17068 12412 17091 12452
rect 17091 12412 17108 12452
rect 19084 12412 19124 12452
rect 18124 12328 18164 12368
rect 26188 12496 26228 12536
rect 26764 12496 26804 12536
rect 27052 12496 27092 12536
rect 27820 12496 27860 12536
rect 23116 12403 23156 12443
rect 23404 12412 23444 12452
rect 25036 12412 25076 12452
rect 25804 12412 25844 12452
rect 27436 12412 27476 12452
rect 27916 12412 27956 12452
rect 28108 12412 28148 12452
rect 19756 12244 19796 12284
rect 21100 12244 21140 12284
rect 21772 12244 21812 12284
rect 23596 12244 23636 12284
rect 15820 12160 15860 12200
rect 17068 12160 17108 12200
rect 27244 12328 27284 12368
rect 28396 12328 28436 12368
rect 28876 12328 28916 12368
rect 25420 12244 25460 12284
rect 27532 12244 27572 12284
rect 20236 12160 20276 12200
rect 27724 12160 27764 12200
rect 18660 12076 19028 12116
rect 19660 12076 19700 12116
rect 22828 12076 22868 12116
rect 16684 11824 16724 11864
rect 26434 12076 26802 12116
rect 26284 11992 26324 12032
rect 27916 11992 27956 12032
rect 17548 11908 17588 11948
rect 19276 11908 19316 11948
rect 21292 11908 21332 11948
rect 28876 11908 28916 11948
rect 17452 11824 17492 11864
rect 22732 11824 22772 11864
rect 15148 11740 15188 11780
rect 15436 11740 15476 11780
rect 15820 11740 15826 11780
rect 15826 11740 15860 11780
rect 17164 11740 17204 11780
rect 1228 11656 1268 11696
rect 1708 11656 1748 11696
rect 3340 11656 3351 11696
rect 3351 11656 3380 11696
rect 4204 11656 4244 11696
rect 4396 11656 4436 11696
rect 4972 11656 5012 11696
rect 5164 11656 5204 11696
rect 5452 11656 5492 11696
rect 5740 11656 5780 11696
rect 6316 11656 6356 11696
rect 6604 11656 6644 11696
rect 7756 11656 7796 11696
rect 8044 11656 8084 11696
rect 9004 11656 9044 11696
rect 11500 11656 11540 11696
rect 11980 11656 12020 11696
rect 12172 11656 12212 11696
rect 13228 11656 13268 11696
rect 1612 11572 1652 11612
rect 3052 11572 3092 11612
rect 5068 11572 5108 11612
rect 6124 11572 6164 11612
rect 4108 11488 4148 11528
rect 5260 11488 5300 11528
rect 9004 11488 9044 11528
rect 1804 11404 1844 11444
rect 5164 11404 5204 11444
rect 3724 11320 3764 11360
rect 4352 11320 4720 11360
rect 4108 11236 4148 11276
rect 1612 11152 1652 11192
rect 2380 11152 2420 11192
rect 2764 11152 2804 11192
rect 3052 11152 3092 11192
rect 5452 11152 5492 11192
rect 6604 11152 6644 11192
rect 748 11068 788 11108
rect 940 11068 980 11108
rect 3148 11068 3188 11108
rect 4588 11068 4628 11108
rect 5260 11068 5300 11108
rect 1132 10984 1172 11024
rect 1612 10984 1652 11024
rect 1804 10984 1844 11024
rect 2092 10984 2132 11024
rect 3340 10984 3380 11024
rect 10348 11572 10388 11612
rect 12844 11572 12884 11612
rect 11020 11488 11051 11528
rect 11051 11488 11060 11528
rect 12652 11488 12692 11528
rect 13036 11488 13076 11528
rect 11980 11404 12020 11444
rect 14764 11656 14804 11696
rect 16300 11656 16340 11696
rect 14188 11572 14228 11612
rect 14380 11488 14411 11528
rect 14411 11488 14420 11528
rect 13804 11404 13844 11444
rect 14956 11572 14996 11612
rect 15244 11572 15284 11612
rect 18892 11740 18923 11780
rect 18923 11740 18932 11780
rect 20236 11740 20276 11780
rect 21964 11740 22004 11780
rect 22540 11740 22580 11780
rect 23596 11740 23636 11780
rect 23884 11740 23924 11780
rect 27628 11824 27668 11864
rect 27916 11824 27956 11864
rect 28204 11824 28244 11864
rect 27724 11740 27764 11780
rect 17740 11656 17780 11696
rect 18508 11656 18548 11696
rect 18700 11656 18740 11696
rect 19468 11656 19508 11696
rect 20812 11656 20852 11696
rect 21868 11656 21908 11696
rect 17452 11572 17492 11612
rect 17932 11572 17972 11612
rect 21580 11572 21620 11612
rect 21772 11572 21812 11612
rect 24172 11656 24212 11696
rect 26956 11656 26996 11696
rect 27148 11656 27188 11696
rect 24364 11572 24404 11612
rect 27436 11656 27476 11696
rect 20908 11488 20948 11528
rect 24940 11488 24980 11528
rect 27532 11488 27572 11528
rect 17260 11404 17300 11444
rect 19372 11404 19412 11444
rect 23308 11404 23348 11444
rect 24460 11404 24500 11444
rect 10060 11320 10100 11360
rect 10252 11320 10292 11360
rect 10732 11320 10772 11360
rect 12126 11320 12494 11360
rect 19900 11320 20268 11360
rect 21292 11320 21332 11360
rect 27674 11320 28042 11360
rect 8428 11236 8468 11276
rect 9772 11236 9812 11276
rect 10636 11236 10676 11276
rect 7372 11152 7412 11192
rect 8524 11152 8564 11192
rect 7852 11068 7892 11108
rect 8716 11068 8756 11108
rect 9580 11152 9620 11192
rect 9196 11068 9236 11108
rect 10156 11068 10196 11108
rect 11500 11152 11540 11192
rect 12556 11152 12596 11192
rect 2188 10900 2228 10940
rect 4396 10984 4427 11024
rect 4427 10984 4436 11024
rect 4684 10984 4695 11024
rect 4695 10984 4724 11024
rect 5164 10984 5204 11024
rect 5548 10984 5588 11024
rect 6028 10984 6051 11024
rect 6051 10984 6068 11024
rect 6988 10984 7028 11024
rect 7468 10984 7499 11024
rect 7499 10984 7508 11024
rect 8620 10984 8631 11024
rect 8631 10984 8660 11024
rect 9004 10984 9044 11024
rect 11020 10984 11060 11024
rect 1996 10816 2036 10856
rect 3112 10564 3480 10604
rect 3820 10900 3860 10940
rect 5836 10816 5876 10856
rect 6700 10900 6740 10940
rect 14380 11236 14420 11276
rect 17740 11236 17780 11276
rect 13228 11152 13259 11192
rect 13259 11152 13268 11192
rect 14188 11152 14228 11192
rect 15052 11152 15092 11192
rect 16780 11152 16820 11192
rect 17452 11152 17492 11192
rect 18700 11152 18740 11192
rect 20524 11152 20564 11192
rect 12652 11068 12692 11108
rect 16204 11068 16244 11108
rect 18796 11068 18836 11108
rect 25804 11236 25844 11276
rect 27436 11236 27476 11276
rect 23788 11152 23828 11192
rect 24364 11152 24404 11192
rect 25324 11152 25364 11192
rect 26188 11152 26228 11192
rect 21868 11068 21908 11108
rect 22444 11068 22484 11108
rect 12268 10984 12269 11024
rect 12269 10984 12308 11024
rect 12844 10984 12884 11024
rect 13708 10984 13748 11024
rect 16396 10984 16436 11024
rect 16780 10984 16820 11024
rect 16972 10984 17012 11024
rect 17548 10984 17588 11024
rect 18124 10984 18164 11024
rect 19180 10984 19220 11024
rect 19564 11015 19604 11024
rect 19564 10984 19595 11015
rect 19595 10984 19604 11015
rect 20332 10984 20372 11024
rect 20908 10984 20948 11024
rect 21484 10984 21524 11024
rect 9196 10900 9236 10940
rect 9772 10900 9812 10940
rect 11308 10900 11348 10940
rect 12172 10900 12203 10940
rect 12203 10900 12212 10940
rect 12748 10900 12779 10940
rect 12779 10900 12788 10940
rect 13900 10900 13940 10940
rect 10156 10816 10196 10856
rect 13804 10816 13844 10856
rect 15244 10900 15284 10940
rect 15052 10816 15092 10856
rect 9964 10732 10004 10772
rect 10636 10732 10676 10772
rect 18124 10732 18164 10772
rect 9100 10648 9140 10688
rect 9580 10564 9620 10604
rect 10252 10564 10292 10604
rect 10886 10564 11254 10604
rect 13228 10564 13268 10604
rect 7948 10480 7988 10520
rect 10444 10480 10484 10520
rect 11884 10480 11924 10520
rect 1996 10396 2036 10436
rect 2956 10396 2996 10436
rect 3532 10396 3572 10436
rect 4780 10396 4820 10436
rect 8716 10396 8756 10436
rect 9196 10396 9236 10436
rect 3340 10312 3380 10352
rect 3628 10312 3668 10352
rect 5068 10312 5108 10352
rect 5740 10312 5780 10352
rect 940 10228 980 10268
rect 1612 10228 1652 10268
rect 1996 10228 2027 10268
rect 2027 10228 2036 10268
rect 2764 10228 2804 10268
rect 4204 10228 4244 10268
rect 4492 10228 4532 10268
rect 4876 10228 4916 10268
rect 5260 10228 5300 10268
rect 5548 10228 5588 10268
rect 6700 10228 6740 10268
rect 6988 10228 7028 10268
rect 7852 10228 7892 10268
rect 11308 10228 11348 10268
rect 1804 10144 1844 10184
rect 2572 10144 2612 10184
rect 2956 10144 2996 10184
rect 3436 10144 3476 10184
rect 4972 10144 5012 10184
rect 5164 10144 5171 10184
rect 5171 10144 5204 10184
rect 5932 10144 5937 10184
rect 5937 10144 5972 10184
rect 6220 10144 6260 10184
rect 7372 10144 7397 10184
rect 7397 10144 7412 10184
rect 7948 10144 7988 10184
rect 9100 10144 9140 10184
rect 10156 10144 10196 10184
rect 16396 10480 16436 10520
rect 14764 10396 14804 10436
rect 16300 10396 16340 10436
rect 18316 10396 18356 10436
rect 11692 10228 11723 10268
rect 11723 10228 11732 10268
rect 12652 10228 12683 10268
rect 12683 10228 12692 10268
rect 13324 10312 13364 10352
rect 13996 10312 14036 10352
rect 14188 10312 14228 10352
rect 14380 10312 14420 10352
rect 13324 10144 13364 10184
rect 13900 10144 13940 10184
rect 1612 10060 1652 10100
rect 2476 10060 2516 10100
rect 4396 10060 4436 10100
rect 4780 10060 4820 10100
rect 3820 9976 3860 10016
rect 4204 9976 4244 10016
rect 5452 9976 5492 10016
rect 3436 9892 3476 9932
rect 7564 10018 7604 10058
rect 9676 10060 9716 10100
rect 10252 10060 10292 10100
rect 7756 9976 7796 10016
rect 8524 9976 8564 10016
rect 9772 9976 9812 10016
rect 10732 10060 10772 10100
rect 13036 10060 13076 10100
rect 13804 10060 13844 10100
rect 14764 10144 14804 10184
rect 15148 10144 15179 10184
rect 15179 10144 15188 10184
rect 15724 10144 15764 10184
rect 16204 10144 16244 10184
rect 16492 10144 16532 10184
rect 16972 10144 17012 10184
rect 17260 10144 17300 10184
rect 17548 10144 17588 10184
rect 21100 10900 21140 10940
rect 21676 10900 21716 10940
rect 22348 10900 22388 10940
rect 18660 10564 19028 10604
rect 22732 10816 22763 10856
rect 22763 10816 22772 10856
rect 18988 10396 19028 10436
rect 14668 10060 14708 10100
rect 16012 10060 16052 10100
rect 11020 9976 11060 10016
rect 11980 9976 12020 10016
rect 12556 9976 12596 10016
rect 13420 9976 13460 10016
rect 13708 9976 13748 10016
rect 8332 9892 8372 9932
rect 10060 9892 10100 9932
rect 10444 9892 10484 9932
rect 13516 9892 13556 9932
rect 15244 9976 15284 10016
rect 16300 9976 16340 10016
rect 18892 10228 18932 10268
rect 21772 10732 21812 10772
rect 20140 10480 20180 10520
rect 21292 10480 21332 10520
rect 21484 10396 21524 10436
rect 24172 10984 24212 11024
rect 24460 11015 24500 11024
rect 24460 10984 24491 11015
rect 24491 10984 24500 11015
rect 26956 10984 26987 11024
rect 26987 10984 26996 11024
rect 28492 10984 28532 11024
rect 25612 10900 25652 10940
rect 27148 10900 27188 10940
rect 27340 10900 27371 10940
rect 27371 10900 27380 10940
rect 25228 10732 25268 10772
rect 26434 10564 26802 10604
rect 27148 10312 27188 10352
rect 24172 10228 24178 10268
rect 24178 10228 24212 10268
rect 27052 10228 27092 10268
rect 19084 10144 19124 10184
rect 21868 10144 21908 10184
rect 23308 10144 23348 10184
rect 24940 10144 24980 10184
rect 25228 10144 25268 10184
rect 25996 10144 26036 10184
rect 18892 10060 18932 10100
rect 22732 10060 22772 10100
rect 19468 9976 19508 10016
rect 20332 9976 20372 10016
rect 21484 9976 21524 10016
rect 22540 9976 22580 10016
rect 23884 9976 23924 10016
rect 26092 9976 26132 10016
rect 26284 9976 26324 10016
rect 20524 9892 20564 9932
rect 21868 9892 21908 9932
rect 2284 9808 2324 9848
rect 2956 9808 2996 9848
rect 4352 9808 4720 9848
rect 6316 9808 6356 9848
rect 8812 9808 8852 9848
rect 10348 9808 10388 9848
rect 12126 9808 12494 9848
rect 12556 9808 12596 9848
rect 16108 9808 16148 9848
rect 19900 9808 20268 9848
rect 27674 9808 28042 9848
rect 1708 9724 1748 9764
rect 5836 9724 5876 9764
rect 6604 9724 6644 9764
rect 8524 9724 8564 9764
rect 9388 9724 9428 9764
rect 11788 9724 11828 9764
rect 2668 9640 2708 9680
rect 2956 9640 2996 9680
rect 4780 9640 4820 9680
rect 5260 9640 5300 9680
rect 940 9556 980 9596
rect 7660 9640 7700 9680
rect 8332 9640 8363 9680
rect 8363 9640 8372 9680
rect 8620 9640 8660 9680
rect 12556 9640 12596 9680
rect 13324 9640 13364 9680
rect 13900 9640 13940 9680
rect 9004 9556 9044 9596
rect 10060 9556 10100 9596
rect 11692 9556 11732 9596
rect 12076 9556 12116 9596
rect 12940 9556 12980 9596
rect 844 9472 884 9512
rect 3436 9472 3476 9512
rect 3724 9472 3764 9512
rect 5836 9472 5876 9512
rect 6220 9472 6260 9512
rect 7564 9472 7604 9512
rect 7852 9472 7892 9512
rect 8428 9472 8468 9512
rect 9388 9472 9428 9512
rect 9772 9472 9779 9512
rect 9779 9472 9812 9512
rect 9964 9472 10004 9512
rect 10444 9472 10475 9512
rect 10475 9472 10484 9512
rect 10636 9472 10676 9512
rect 11212 9472 11252 9512
rect 11500 9472 11540 9512
rect 12460 9472 12500 9512
rect 14764 9556 14804 9596
rect 19756 9724 19796 9764
rect 20428 9724 20468 9764
rect 24268 9724 24308 9764
rect 15628 9640 15668 9680
rect 17932 9640 17972 9680
rect 18412 9640 18452 9680
rect 19276 9640 19316 9680
rect 22828 9640 22859 9680
rect 22859 9640 22868 9680
rect 16204 9556 16244 9596
rect 17260 9556 17300 9596
rect 21484 9556 21524 9596
rect 1516 9388 1556 9428
rect 460 8884 500 8924
rect 3340 9388 3380 9428
rect 4204 9388 4244 9428
rect 4876 9388 4916 9428
rect 5164 9388 5170 9428
rect 5170 9388 5204 9428
rect 6124 9388 6164 9428
rect 6796 9388 6836 9428
rect 8812 9388 8852 9428
rect 5356 9304 5396 9344
rect 5548 9304 5588 9344
rect 7276 9304 7316 9344
rect 5068 9220 5108 9260
rect 7084 9220 7115 9260
rect 7115 9220 7124 9260
rect 8044 9220 8084 9260
rect 13132 9472 13172 9512
rect 13516 9472 13556 9512
rect 13996 9503 14036 9512
rect 13996 9472 14036 9503
rect 14668 9472 14708 9512
rect 15724 9472 15764 9512
rect 16012 9472 16052 9512
rect 16396 9472 16436 9512
rect 17836 9472 17876 9512
rect 19660 9472 19700 9512
rect 9196 9388 9236 9428
rect 9676 9388 9716 9428
rect 11884 9388 11924 9428
rect 13228 9388 13268 9428
rect 9100 9304 9140 9344
rect 14668 9304 14708 9344
rect 17356 9388 17396 9428
rect 17644 9388 17684 9428
rect 18700 9388 18740 9428
rect 18988 9388 19028 9428
rect 17548 9304 17588 9344
rect 18892 9304 18932 9344
rect 9868 9220 9908 9260
rect 17260 9220 17300 9260
rect 18508 9220 18548 9260
rect 9292 9136 9332 9176
rect 3112 9052 3480 9092
rect 6316 9052 6356 9092
rect 10886 9052 11254 9092
rect 14572 9052 14612 9092
rect 18660 9052 19028 9092
rect 7372 8968 7412 9008
rect 9676 8968 9716 9008
rect 3724 8884 3764 8924
rect 4972 8884 5012 8924
rect 8140 8884 8180 8924
rect 9772 8884 9812 8924
rect 10828 8884 10868 8924
rect 5164 8800 5204 8840
rect 6220 8800 6260 8840
rect 2476 8716 2516 8756
rect 4780 8716 4820 8756
rect 172 8632 212 8672
rect 2956 8632 2996 8672
rect 4204 8632 4244 8672
rect 4684 8632 4724 8672
rect 5068 8632 5108 8672
rect 5356 8632 5396 8672
rect 5644 8632 5684 8672
rect 2092 8548 2132 8588
rect 4876 8548 4916 8588
rect 2572 8380 2612 8420
rect 3724 8380 3764 8420
rect 460 8044 500 8084
rect 8716 8800 8756 8840
rect 9388 8800 9428 8840
rect 10252 8800 10292 8840
rect 7276 8716 7307 8756
rect 7307 8716 7316 8756
rect 8428 8716 8468 8756
rect 9100 8747 9140 8756
rect 9100 8716 9139 8747
rect 9139 8716 9140 8747
rect 9772 8716 9812 8756
rect 10732 8716 10772 8756
rect 13036 8884 13076 8924
rect 12844 8800 12884 8840
rect 15052 8800 15092 8840
rect 20332 9472 20372 9512
rect 22540 9472 22580 9512
rect 23308 9472 23348 9512
rect 20140 9388 20180 9428
rect 21196 9388 21236 9428
rect 24172 9640 24212 9680
rect 25996 9640 26036 9680
rect 27340 9640 27380 9680
rect 25900 9556 25940 9596
rect 25228 9472 25268 9512
rect 25996 9472 26036 9512
rect 26284 9472 26315 9512
rect 26315 9472 26324 9512
rect 24844 9388 24884 9428
rect 26092 9388 26132 9428
rect 24460 9304 24500 9344
rect 25708 9304 25748 9344
rect 26434 9052 26802 9092
rect 20140 8884 20171 8924
rect 20171 8884 20180 8924
rect 21580 8884 21620 8924
rect 24076 8884 24116 8924
rect 18412 8800 18452 8840
rect 19564 8800 19604 8840
rect 12940 8716 12980 8756
rect 13228 8716 13268 8756
rect 16492 8716 16532 8756
rect 17260 8716 17300 8756
rect 17548 8716 17588 8756
rect 6316 8632 6347 8672
rect 6347 8632 6356 8672
rect 6604 8632 6644 8672
rect 7084 8632 7124 8672
rect 7372 8632 7412 8672
rect 8044 8632 8084 8672
rect 8524 8632 8564 8672
rect 9292 8632 9332 8672
rect 9676 8632 9716 8672
rect 10060 8632 10100 8672
rect 10252 8632 10292 8672
rect 10540 8632 10580 8672
rect 11500 8632 11540 8672
rect 13420 8632 13460 8672
rect 13612 8632 13652 8672
rect 16204 8632 16244 8672
rect 18028 8632 18068 8672
rect 18604 8716 18644 8756
rect 20812 8716 20852 8756
rect 21100 8716 21140 8756
rect 21292 8716 21332 8756
rect 21868 8716 21908 8756
rect 23596 8716 23636 8756
rect 23884 8716 23924 8756
rect 24364 8716 24404 8756
rect 26572 8716 26595 8756
rect 26595 8716 26612 8756
rect 5932 8548 5972 8588
rect 6796 8548 6836 8588
rect 7564 8548 7604 8588
rect 11692 8548 11732 8588
rect 13324 8548 13364 8588
rect 20428 8632 20468 8672
rect 21388 8632 21428 8672
rect 21580 8632 21620 8672
rect 21772 8632 21812 8672
rect 23116 8632 23156 8672
rect 23980 8632 24020 8672
rect 24556 8632 24596 8672
rect 24844 8632 24884 8672
rect 25708 8632 25748 8672
rect 25900 8632 25940 8672
rect 26476 8632 26516 8672
rect 27052 8632 27092 8672
rect 20908 8548 20948 8588
rect 24076 8548 24116 8588
rect 8140 8464 8171 8504
rect 8171 8464 8180 8504
rect 9196 8464 9236 8504
rect 9964 8464 10004 8504
rect 11404 8464 11444 8504
rect 11788 8464 11828 8504
rect 12748 8464 12788 8504
rect 14476 8464 14516 8504
rect 15532 8464 15572 8504
rect 18124 8464 18164 8504
rect 8428 8380 8468 8420
rect 20812 8464 20852 8504
rect 22732 8464 22772 8504
rect 23404 8464 23444 8504
rect 26476 8464 26516 8504
rect 4352 8296 4720 8336
rect 5068 8296 5108 8336
rect 11788 8296 11828 8336
rect 12126 8296 12494 8336
rect 19900 8296 20268 8336
rect 27674 8296 28042 8336
rect 5548 8212 5588 8252
rect 6892 8212 6932 8252
rect 10636 8212 10676 8252
rect 1420 8128 1460 8168
rect 2092 8128 2132 8168
rect 3820 8128 3860 8168
rect 4204 8128 4244 8168
rect 5740 8128 5780 8168
rect 7564 8128 7604 8168
rect 9484 8128 9524 8168
rect 9772 8128 9803 8168
rect 9803 8128 9812 8168
rect 940 8044 980 8084
rect 1516 8044 1556 8084
rect 5068 8044 5097 8084
rect 5097 8044 5108 8084
rect 5452 8044 5492 8084
rect 11980 8212 12020 8252
rect 14956 8212 14996 8252
rect 18028 8212 18068 8252
rect 22444 8212 22484 8252
rect 23212 8212 23252 8252
rect 11500 8128 11540 8168
rect 11884 8128 11924 8168
rect 12268 8128 12308 8168
rect 13804 8128 13844 8168
rect 14092 8128 14132 8168
rect 15436 8128 15476 8168
rect 16396 8128 16436 8168
rect 19660 8128 19700 8168
rect 21196 8128 21236 8168
rect 12076 8044 12116 8084
rect 12556 8044 12596 8084
rect 14476 8044 14516 8084
rect 14860 8044 14900 8084
rect 18028 8044 18068 8084
rect 19180 8044 19220 8084
rect 20620 8044 20660 8084
rect 21100 8044 21140 8084
rect 21388 8128 21428 8168
rect 23308 8128 23339 8168
rect 23339 8128 23348 8168
rect 23596 8128 23636 8168
rect 25900 8128 25940 8168
rect 26284 8128 26315 8168
rect 26315 8128 26324 8168
rect 22444 8044 22484 8084
rect 25996 8044 26036 8084
rect 26380 8044 26420 8084
rect 1804 7960 1844 8000
rect 2092 7960 2132 8000
rect 2284 7960 2324 8000
rect 3724 7991 3764 8000
rect 3724 7960 3755 7991
rect 3755 7960 3764 7991
rect 4684 7960 4724 8000
rect 5356 7991 5396 8000
rect 5356 7960 5396 7991
rect 6028 7960 6068 8000
rect 6316 7960 6356 8000
rect 7948 7960 7988 8000
rect 8140 7960 8180 8000
rect 8428 7960 8468 8000
rect 9964 7960 10004 8000
rect 10252 7960 10292 8000
rect 10636 7960 10676 8000
rect 1228 7876 1268 7916
rect 2188 7876 2228 7916
rect 2764 7876 2804 7916
rect 2572 7792 2612 7832
rect 10828 7960 10868 8000
rect 11692 7960 11732 8000
rect 11980 7960 12020 8000
rect 12364 7991 12404 8000
rect 12364 7960 12404 7991
rect 12748 7960 12788 8000
rect 13324 7960 13364 8000
rect 14380 7960 14420 8000
rect 14668 7960 14697 8000
rect 14697 7960 14708 8000
rect 14956 7991 14996 8000
rect 14956 7960 14996 7991
rect 15532 7960 15572 8000
rect 17356 7960 17396 8000
rect 17740 7960 17780 8000
rect 18124 7960 18164 8000
rect 18604 7960 18644 8000
rect 20908 7960 20948 8000
rect 6220 7876 6260 7916
rect 8812 7876 8852 7916
rect 12076 7876 12116 7916
rect 4780 7792 4820 7832
rect 14764 7876 14804 7916
rect 13612 7792 13652 7832
rect 2188 7708 2228 7748
rect 6220 7708 6260 7748
rect 7660 7708 7700 7748
rect 13900 7708 13940 7748
rect 652 7624 692 7664
rect 3724 7624 3764 7664
rect 8908 7624 8948 7664
rect 11692 7624 11732 7664
rect 3112 7540 3480 7580
rect 10886 7540 11254 7580
rect 2380 7456 2420 7496
rect 7180 7456 7220 7496
rect 10252 7456 10292 7496
rect 1708 7372 1748 7412
rect 2284 7372 2324 7412
rect 5356 7372 5387 7412
rect 5387 7372 5396 7412
rect 1036 7288 1076 7328
rect 844 7204 884 7244
rect 1228 7204 1268 7244
rect 1516 7204 1556 7244
rect 2188 7288 2228 7328
rect 3340 7288 3380 7328
rect 4300 7288 4340 7328
rect 5260 7288 5300 7328
rect 5644 7288 5684 7328
rect 3052 7204 3092 7244
rect 4876 7204 4916 7244
rect 5740 7204 5780 7244
rect 1900 7120 1940 7160
rect 22348 7960 22388 8000
rect 22636 7960 22676 8000
rect 23404 7960 23444 8000
rect 19180 7876 19220 7916
rect 19372 7876 19412 7916
rect 20812 7876 20852 7916
rect 20236 7708 20276 7748
rect 20524 7708 20564 7748
rect 18660 7540 19028 7580
rect 8812 7372 8852 7412
rect 9292 7372 9332 7412
rect 12652 7372 12692 7412
rect 13996 7372 14027 7412
rect 14027 7372 14036 7412
rect 14380 7372 14420 7412
rect 18124 7372 18164 7412
rect 18892 7372 18932 7412
rect 20908 7372 20948 7412
rect 15052 7288 15092 7328
rect 15244 7288 15284 7328
rect 19564 7288 19604 7328
rect 20236 7288 20276 7328
rect 20716 7288 20756 7328
rect 6508 7204 6548 7244
rect 7564 7204 7595 7244
rect 7595 7204 7604 7244
rect 11596 7204 11636 7244
rect 11788 7204 11828 7244
rect 13324 7204 13364 7244
rect 15148 7204 15188 7244
rect 23596 7960 23636 8000
rect 23788 7960 23828 8000
rect 24076 7960 24116 8000
rect 24556 7960 24596 8000
rect 24844 7960 24884 8000
rect 25612 7960 25652 8000
rect 22828 7876 22868 7916
rect 24460 7876 24500 7916
rect 26188 7876 26228 7916
rect 26860 7960 26900 8000
rect 26764 7876 26795 7916
rect 26795 7876 26804 7916
rect 22540 7792 22580 7832
rect 23116 7792 23156 7832
rect 23308 7792 23348 7832
rect 25900 7792 25940 7832
rect 23020 7708 23060 7748
rect 25132 7708 25172 7748
rect 23500 7624 23540 7664
rect 25996 7624 26036 7664
rect 26434 7540 26802 7580
rect 25612 7456 25652 7496
rect 23788 7372 23828 7412
rect 24364 7372 24404 7412
rect 23116 7288 23156 7328
rect 20044 7204 20084 7244
rect 20332 7204 20372 7244
rect 20524 7204 20564 7244
rect 23020 7204 23060 7244
rect 3436 7120 3476 7160
rect 3724 7120 3764 7160
rect 5164 7120 5204 7160
rect 6220 7120 6260 7160
rect 6604 7120 6644 7160
rect 7660 7120 7700 7160
rect 9100 7120 9140 7160
rect 9772 7120 9812 7160
rect 10540 7120 10580 7160
rect 11116 7120 11156 7160
rect 11308 7120 11348 7160
rect 11692 7120 11732 7160
rect 12268 7120 12308 7160
rect 13900 7120 13940 7160
rect 14764 7120 14804 7160
rect 1228 7036 1268 7076
rect 1420 7036 1460 7076
rect 3628 7036 3668 7076
rect 4300 7036 4340 7076
rect 6028 7036 6068 7076
rect 7180 7036 7220 7076
rect 1612 6952 1643 6992
rect 1643 6952 1652 6992
rect 1804 6952 1835 6992
rect 1835 6952 1844 6992
rect 2572 6952 2612 6992
rect 3820 6952 3860 6992
rect 5740 6952 5780 6992
rect 5932 6952 5972 6992
rect 6124 6952 6164 6992
rect 6796 6952 6836 6992
rect 2668 6868 2708 6908
rect 748 6784 788 6824
rect 4012 6784 4052 6824
rect 5836 6868 5876 6908
rect 4352 6784 4720 6824
rect 1516 6700 1556 6740
rect 3916 6700 3956 6740
rect 4780 6700 4820 6740
rect 1996 6616 2036 6656
rect 2284 6616 2324 6656
rect 1324 6532 1364 6572
rect 2764 6532 2804 6572
rect 3532 6616 3572 6656
rect 6604 6616 6644 6656
rect 2956 6532 2996 6572
rect 6892 6532 6932 6572
rect 8716 7036 8756 7076
rect 16012 7120 16052 7160
rect 16204 7120 16244 7160
rect 17548 7120 17588 7160
rect 18124 7120 18164 7160
rect 18700 7120 18740 7160
rect 10636 7036 10676 7076
rect 11980 7036 12020 7076
rect 13036 7036 13076 7076
rect 14380 7036 14420 7076
rect 14668 7036 14708 7076
rect 15148 7036 15188 7076
rect 11308 6952 11348 6992
rect 12364 6952 12404 6992
rect 14476 6952 14516 6992
rect 18316 7036 18356 7076
rect 18604 7036 18644 7076
rect 19372 7120 19401 7160
rect 19401 7120 19412 7160
rect 20236 7120 20276 7160
rect 22060 7120 22100 7160
rect 22252 7120 22292 7160
rect 22540 7120 22571 7160
rect 22571 7120 22580 7160
rect 22828 7120 22868 7160
rect 14284 6868 14324 6908
rect 19180 7036 19220 7076
rect 19660 7036 19700 7076
rect 20428 7036 20468 7076
rect 17740 6952 17780 6992
rect 18988 6952 19028 6992
rect 20044 6952 20084 6992
rect 20716 7036 20756 7076
rect 23500 7036 23540 7076
rect 23788 7036 23819 7076
rect 23819 7036 23828 7076
rect 21292 6952 21332 6992
rect 22060 6952 22100 6992
rect 23308 6952 23348 6992
rect 24268 7036 24308 7076
rect 12126 6784 12494 6824
rect 19564 6784 19604 6824
rect 19900 6784 20268 6824
rect 22732 6784 22772 6824
rect 27674 6784 28042 6824
rect 8332 6700 8372 6740
rect 11500 6700 11540 6740
rect 18508 6700 18548 6740
rect 9772 6616 9812 6656
rect 10252 6616 10283 6656
rect 10283 6616 10292 6656
rect 10732 6616 10772 6656
rect 7852 6532 7892 6572
rect 11980 6616 12020 6656
rect 12460 6616 12491 6656
rect 12491 6616 12500 6656
rect 14764 6616 14804 6656
rect 15148 6616 15188 6656
rect 16204 6616 16244 6656
rect 14380 6532 14420 6572
rect 19660 6700 19700 6740
rect 16780 6616 16820 6656
rect 17548 6616 17588 6656
rect 18604 6616 18644 6656
rect 18892 6616 18932 6656
rect 20620 6616 20660 6656
rect 21388 6616 21428 6656
rect 22252 6616 22292 6656
rect 23596 6616 23636 6656
rect 23788 6616 23828 6656
rect 2188 6448 2228 6488
rect 3340 6448 3380 6488
rect 4204 6448 4244 6488
rect 6796 6448 6836 6488
rect 7372 6448 7412 6488
rect 9004 6479 9044 6488
rect 556 6364 596 6404
rect 1420 6364 1460 6404
rect 9004 6448 9035 6479
rect 9035 6448 9044 6479
rect 9580 6448 9620 6488
rect 10060 6448 10100 6488
rect 11308 6448 11348 6488
rect 13132 6448 13172 6488
rect 1804 6364 1844 6404
rect 3724 6364 3764 6404
rect 4684 6364 4724 6404
rect 8524 6364 8564 6404
rect 9772 6364 9812 6404
rect 10828 6364 10868 6404
rect 11596 6364 11636 6404
rect 13708 6448 13748 6488
rect 13996 6448 14036 6488
rect 15628 6448 15668 6488
rect 16012 6448 16052 6488
rect 18124 6448 18164 6488
rect 18316 6448 18356 6488
rect 18988 6479 19028 6488
rect 18988 6448 19028 6479
rect 19180 6448 19220 6488
rect 20140 6448 20180 6488
rect 20716 6448 20747 6488
rect 20747 6448 20756 6488
rect 23308 6448 23348 6488
rect 23884 6448 23924 6488
rect 24268 6448 24308 6488
rect 24940 6448 24980 6488
rect 25804 6448 25844 6488
rect 1036 6280 1076 6320
rect 2188 6280 2228 6320
rect 2476 6280 2516 6320
rect 7756 6280 7796 6320
rect 10540 6280 10580 6320
rect 11788 6280 11828 6320
rect 13900 6280 13940 6320
rect 19468 6364 19508 6404
rect 21580 6364 21620 6404
rect 22828 6364 22868 6404
rect 24652 6280 24692 6320
rect 6028 6196 6068 6236
rect 10636 6196 10676 6236
rect 20620 6196 20660 6236
rect 20812 6196 20852 6236
rect 24844 6196 24884 6236
rect 5932 6112 5972 6152
rect 8524 6112 8564 6152
rect 18316 6112 18356 6152
rect 25324 6112 25364 6152
rect 3112 6028 3480 6068
rect 10886 6028 11254 6068
rect 18660 6028 19028 6068
rect 26434 6028 26802 6068
rect 19372 5944 19412 5984
rect 20428 5944 20468 5984
rect 21196 5944 21236 5984
rect 3724 5860 3764 5900
rect 4876 5860 4916 5900
rect 7948 5860 7988 5900
rect 9004 5860 9044 5900
rect 11500 5860 11540 5900
rect 12844 5860 12884 5900
rect 13036 5860 13076 5900
rect 14284 5860 14324 5900
rect 15340 5860 15380 5900
rect 18124 5860 18164 5900
rect 20140 5860 20180 5900
rect 20620 5860 20660 5900
rect 22636 5860 22676 5900
rect 24172 5860 24212 5900
rect 24940 5860 24980 5900
rect 3820 5776 3860 5816
rect 4684 5776 4724 5816
rect 6220 5776 6260 5816
rect 17356 5776 17396 5816
rect 21964 5776 22004 5816
rect 25804 5776 25844 5816
rect 7564 5692 7604 5732
rect 11212 5692 11252 5732
rect 12940 5692 12980 5732
rect 15052 5692 15092 5732
rect 15628 5692 15668 5732
rect 17548 5692 17588 5732
rect 18220 5692 18260 5732
rect 20716 5692 20756 5732
rect 3532 5608 3572 5648
rect 4204 5608 4244 5648
rect 4780 5608 4820 5648
rect 5740 5608 5780 5648
rect 6028 5608 6056 5648
rect 6056 5608 6068 5648
rect 6892 5608 6923 5648
rect 6923 5608 6932 5648
rect 8236 5608 8276 5648
rect 9004 5608 9044 5648
rect 13228 5608 13268 5648
rect 15916 5608 15956 5648
rect 19468 5608 19508 5648
rect 20332 5608 20372 5648
rect 21292 5608 21332 5648
rect 22732 5608 22763 5648
rect 22763 5608 22772 5648
rect 24652 5608 24692 5648
rect 25132 5608 25172 5648
rect 4108 5524 4148 5564
rect 5452 5524 5492 5564
rect 6508 5524 6539 5564
rect 6539 5524 6548 5564
rect 10060 5524 10100 5564
rect 12844 5524 12875 5564
rect 12875 5524 12884 5564
rect 5740 5356 5780 5396
rect 7372 5356 7412 5396
rect 4352 5272 4720 5312
rect 4108 5188 4148 5228
rect 5452 5188 5492 5228
rect 6508 5104 6548 5144
rect 7372 5104 7412 5144
rect 12126 5272 12494 5312
rect 13036 5524 13076 5564
rect 16492 5524 16532 5564
rect 13996 5440 14036 5480
rect 10348 5188 10388 5228
rect 13132 5104 13172 5144
rect 19276 5524 19307 5564
rect 19307 5524 19316 5564
rect 20908 5524 20948 5564
rect 20428 5440 20468 5480
rect 21004 5356 21044 5396
rect 19900 5272 20268 5312
rect 22828 5188 22868 5228
rect 23308 5188 23348 5228
rect 13804 5104 13835 5144
rect 13835 5104 13844 5144
rect 19468 5104 19508 5144
rect 21196 5104 21236 5144
rect 22348 5104 22388 5144
rect 11500 5020 11540 5060
rect 12844 5020 12884 5060
rect 6220 4936 6260 4976
rect 9772 4936 9812 4976
rect 10348 4936 10388 4976
rect 13420 5020 13460 5060
rect 13900 5020 13940 5060
rect 16300 5020 16340 5060
rect 22636 5020 22676 5060
rect 23212 5020 23252 5060
rect 27674 5272 28042 5312
rect 24268 5020 24308 5060
rect 11308 4936 11348 4976
rect 11980 4936 12020 4976
rect 13708 4936 13739 4976
rect 13739 4936 13748 4976
rect 13996 4936 14007 4976
rect 14007 4936 14036 4976
rect 14284 4936 14324 4976
rect 16492 4936 16532 4976
rect 17356 4936 17396 4976
rect 20524 4936 20564 4976
rect 20908 4936 20948 4976
rect 21388 4936 21428 4976
rect 22636 4936 22676 4976
rect 8908 4852 8948 4892
rect 10252 4852 10292 4892
rect 11596 4852 11627 4892
rect 11627 4852 11636 4892
rect 11788 4852 11828 4892
rect 12940 4852 12980 4892
rect 7564 4768 7604 4808
rect 11212 4768 11252 4808
rect 13036 4768 13076 4808
rect 22828 4852 22868 4892
rect 23596 4852 23636 4892
rect 15052 4768 15092 4808
rect 18220 4768 18260 4808
rect 20428 4768 20468 4808
rect 21580 4768 21620 4808
rect 23884 4768 23924 4808
rect 9772 4684 9812 4724
rect 11980 4684 12020 4724
rect 19852 4684 19892 4724
rect 26188 4684 26228 4724
rect 3112 4516 3480 4556
rect 10886 4516 11254 4556
rect 18660 4516 19028 4556
rect 26434 4516 26802 4556
rect 19276 4348 19316 4388
rect 20332 4348 20372 4388
rect 20524 4348 20564 4388
rect 9100 4264 9140 4304
rect 9580 4180 9620 4220
rect 20428 4180 20468 4220
rect 21292 4180 21332 4220
rect 9772 4096 9812 4136
rect 19852 4096 19883 4136
rect 19883 4096 19892 4136
rect 20812 4096 20852 4136
rect 21004 4012 21044 4052
rect 4352 3760 4720 3800
rect 12126 3760 12494 3800
rect 19900 3760 20268 3800
rect 27674 3760 28042 3800
rect 3112 3004 3480 3044
rect 10886 3004 11254 3044
rect 18660 3004 19028 3044
rect 26434 3004 26802 3044
rect 4352 2248 4720 2288
rect 12126 2248 12494 2288
rect 19900 2248 20268 2288
rect 27674 2248 28042 2288
rect 3112 1492 3480 1532
rect 10886 1492 11254 1532
rect 18660 1492 19028 1532
rect 26434 1492 26802 1532
rect 4352 736 4720 776
rect 12126 736 12494 776
rect 19900 736 20268 776
rect 27674 736 28042 776
<< metal3 >>
rect 2092 28916 2132 28925
rect 2092 28076 2132 28876
rect 3128 28600 3208 29000
rect 3896 28600 3976 29000
rect 4664 28600 4744 29000
rect 5432 28600 5512 29000
rect 5644 28664 5684 28673
rect 2092 28027 2132 28036
rect 2380 28496 2420 28505
rect 1900 27908 1940 27917
rect 2284 27908 2324 27917
rect 1940 27868 2284 27908
rect 1900 27859 1940 27868
rect 2284 27859 2324 27868
rect 1900 27740 1940 27749
rect 1516 27656 1556 27665
rect 652 27404 692 27413
rect 652 26816 692 27364
rect 652 26144 692 26776
rect 1036 26900 1076 26909
rect 1036 26396 1076 26860
rect 1516 26900 1556 27616
rect 1228 26816 1268 26825
rect 1132 26648 1172 26657
rect 1132 26513 1172 26608
rect 1036 26347 1076 26356
rect 1228 26312 1268 26776
rect 1228 26263 1268 26272
rect 1132 26228 1172 26237
rect 652 25640 692 26104
rect 844 26144 884 26153
rect 844 26009 884 26104
rect 940 26060 980 26069
rect 652 25591 692 25600
rect 844 25304 884 25313
rect 940 25304 980 26020
rect 884 25264 980 25304
rect 844 25255 884 25264
rect 460 24380 500 24389
rect 364 23792 404 23801
rect 172 23120 212 23129
rect 76 20516 116 20525
rect 76 13880 116 20476
rect 76 13831 116 13840
rect 172 8672 212 23080
rect 172 8623 212 8632
rect 268 20432 308 20441
rect 268 7328 308 20392
rect 364 17996 404 23752
rect 460 19424 500 24340
rect 556 23960 596 23969
rect 556 23204 596 23920
rect 940 23876 980 25264
rect 1036 25388 1076 25397
rect 1036 24800 1076 25348
rect 1132 25304 1172 26188
rect 1420 26144 1460 26153
rect 1420 26060 1460 26104
rect 1420 26009 1460 26020
rect 1132 25255 1172 25264
rect 1036 24760 1172 24800
rect 940 23792 980 23836
rect 940 23741 980 23752
rect 1036 24632 1076 24641
rect 556 23155 596 23164
rect 1036 23120 1076 24592
rect 1036 23071 1076 23080
rect 556 22280 596 22289
rect 556 20600 596 22240
rect 844 22196 884 22205
rect 748 20852 788 20947
rect 748 20803 788 20812
rect 556 20551 596 20560
rect 748 20684 788 20693
rect 556 20348 596 20357
rect 556 19928 596 20308
rect 556 19888 692 19928
rect 460 19375 500 19384
rect 556 19256 596 19265
rect 556 18668 596 19216
rect 556 18619 596 18628
rect 652 18248 692 19888
rect 652 18199 692 18208
rect 364 17947 404 17956
rect 460 18164 500 18173
rect 364 17324 404 17333
rect 364 8924 404 17284
rect 460 12704 500 18124
rect 652 17996 692 18005
rect 652 17828 692 17956
rect 748 17996 788 20644
rect 748 17947 788 17956
rect 652 17788 788 17828
rect 652 17408 692 17417
rect 652 15560 692 17368
rect 556 15520 652 15560
rect 556 14048 596 15520
rect 652 15511 692 15520
rect 556 13999 596 14008
rect 652 14552 692 14561
rect 460 12655 500 12664
rect 556 13880 596 13889
rect 460 8924 500 8933
rect 364 8884 460 8924
rect 460 8875 500 8884
rect 460 8084 500 8093
rect 460 7949 500 8044
rect 268 7279 308 7288
rect 556 6404 596 13840
rect 652 13208 692 14512
rect 652 12788 692 13168
rect 652 12739 692 12748
rect 748 11108 788 17788
rect 844 17408 884 22156
rect 1036 21524 1076 21533
rect 940 21440 980 21449
rect 940 20768 980 21400
rect 1036 21389 1076 21484
rect 1132 21020 1172 24760
rect 1420 24128 1460 24137
rect 1420 23792 1460 24088
rect 1420 23743 1460 23752
rect 1228 23708 1268 23717
rect 1228 22112 1268 23668
rect 1228 22063 1268 22072
rect 1516 21860 1556 26860
rect 1804 26816 1844 26825
rect 1804 26564 1844 26776
rect 1804 26515 1844 26524
rect 1804 26144 1844 26153
rect 1612 25976 1652 25985
rect 1612 22448 1652 25936
rect 1708 24548 1748 24557
rect 1708 24413 1748 24508
rect 1612 22399 1652 22408
rect 1804 24128 1844 26104
rect 1804 22280 1844 24088
rect 1900 23960 1940 27700
rect 2092 27740 2132 27749
rect 2092 27605 2132 27700
rect 2380 27740 2420 28456
rect 2476 28328 2516 28337
rect 2476 27824 2516 28288
rect 3148 28076 3188 28600
rect 3148 28027 3188 28036
rect 3052 27908 3092 27917
rect 2476 27775 2516 27784
rect 2956 27824 2996 27833
rect 2860 27740 2900 27749
rect 2380 27691 2420 27700
rect 2668 27700 2860 27740
rect 2380 27572 2420 27581
rect 2380 27404 2420 27532
rect 2572 27572 2612 27667
rect 2572 27523 2612 27532
rect 2380 27355 2420 27364
rect 2188 27320 2228 27329
rect 2092 26816 2132 26825
rect 1996 26648 2036 26657
rect 1996 26060 2036 26608
rect 1996 26011 2036 26020
rect 2092 25892 2132 26776
rect 2188 26732 2228 27280
rect 2188 26683 2228 26692
rect 2284 27068 2324 27077
rect 2284 25976 2324 27028
rect 2284 25927 2324 25936
rect 2380 26900 2420 26909
rect 2092 25843 2132 25852
rect 2380 24884 2420 26860
rect 2476 26900 2516 26909
rect 2476 26060 2516 26860
rect 2668 26732 2708 27700
rect 2860 27691 2900 27700
rect 2956 27689 2996 27784
rect 2764 27572 2804 27581
rect 2764 26900 2804 27532
rect 3052 27572 3092 27868
rect 3052 27523 3092 27532
rect 3340 27656 3380 27665
rect 3340 27488 3380 27616
rect 3724 27572 3764 27581
rect 3764 27532 3860 27572
rect 3724 27523 3764 27532
rect 3340 27439 3380 27448
rect 3628 27488 3668 27497
rect 3112 27236 3480 27245
rect 3112 27187 3480 27196
rect 3628 27236 3668 27448
rect 3628 27187 3668 27196
rect 3724 27404 3764 27413
rect 3340 27068 3380 27077
rect 2764 26851 2804 26860
rect 3148 26900 3188 26909
rect 2668 26228 2708 26692
rect 2956 26732 2996 26741
rect 2668 26179 2708 26188
rect 2764 26648 2804 26657
rect 2476 26011 2516 26020
rect 2668 25976 2708 25985
rect 2668 25841 2708 25936
rect 2572 25220 2612 25229
rect 2380 24844 2516 24884
rect 1900 23911 1940 23920
rect 2092 24800 2132 24809
rect 1804 22231 1844 22240
rect 1996 23036 2036 23045
rect 1516 21811 1556 21820
rect 1708 21524 1748 21533
rect 1324 21440 1364 21449
rect 1132 20971 1172 20980
rect 1228 21104 1268 21113
rect 940 20719 980 20728
rect 1132 20852 1172 20861
rect 1132 20432 1172 20812
rect 1132 20383 1172 20392
rect 940 20348 980 20357
rect 940 18500 980 20308
rect 1228 20264 1268 21064
rect 1228 20215 1268 20224
rect 940 18451 980 18460
rect 1036 20180 1076 20189
rect 940 17912 980 17921
rect 940 17744 980 17872
rect 940 17695 980 17704
rect 844 17359 884 17368
rect 940 17492 980 17501
rect 844 17240 884 17249
rect 844 13544 884 17200
rect 940 17156 980 17452
rect 940 17107 980 17116
rect 940 16820 980 16829
rect 940 13964 980 16780
rect 1036 15728 1076 20140
rect 1132 20096 1172 20105
rect 1132 19592 1172 20056
rect 1132 19543 1172 19552
rect 1228 18416 1268 18425
rect 1132 17996 1172 18005
rect 1132 17744 1172 17956
rect 1132 17695 1172 17704
rect 1228 17324 1268 18376
rect 1228 17275 1268 17284
rect 1036 15679 1076 15688
rect 1132 17240 1172 17249
rect 1036 14804 1076 14813
rect 1036 14048 1076 14764
rect 1036 13999 1076 14008
rect 940 13915 980 13924
rect 844 13495 884 13504
rect 1132 13124 1172 17200
rect 1228 16988 1268 16997
rect 1228 16232 1268 16948
rect 1228 16183 1268 16192
rect 1228 15560 1268 15569
rect 1228 14216 1268 15520
rect 1228 14167 1268 14176
rect 1132 13075 1172 13084
rect 1228 13040 1268 13049
rect 940 12536 980 12547
rect 940 12452 980 12496
rect 940 12403 980 12412
rect 1132 11864 1172 11873
rect 748 11059 788 11068
rect 940 11108 980 11117
rect 940 10268 980 11068
rect 844 9764 884 9773
rect 844 9512 884 9724
rect 940 9596 980 10228
rect 1132 11024 1172 11824
rect 1228 11696 1268 13000
rect 1228 11647 1268 11656
rect 1132 10100 1172 10984
rect 1228 10184 1268 10193
rect 1228 10100 1268 10144
rect 1132 10060 1268 10100
rect 940 9547 980 9556
rect 652 7664 692 7673
rect 652 7529 692 7624
rect 844 7244 884 9472
rect 940 8168 980 8179
rect 940 8084 980 8128
rect 940 8035 980 8044
rect 1228 7916 1268 10060
rect 844 7195 884 7204
rect 1036 7328 1076 7337
rect 748 6824 788 6833
rect 748 6689 788 6784
rect 556 6355 596 6364
rect 1036 6320 1076 7288
rect 1228 7244 1268 7876
rect 1228 7195 1268 7204
rect 1228 7076 1268 7085
rect 1228 6941 1268 7036
rect 1324 6572 1364 21400
rect 1420 21356 1460 21365
rect 1420 20852 1460 21316
rect 1516 20852 1556 20861
rect 1420 20812 1516 20852
rect 1420 20516 1460 20525
rect 1420 19844 1460 20476
rect 1516 20096 1556 20812
rect 1516 20012 1556 20056
rect 1516 19932 1556 19972
rect 1612 20768 1652 20777
rect 1420 19795 1460 19804
rect 1612 19256 1652 20728
rect 1708 20432 1748 21484
rect 1900 21020 1940 21029
rect 1804 20936 1844 20945
rect 1804 20801 1844 20896
rect 1708 20383 1748 20392
rect 1900 20180 1940 20980
rect 1900 20131 1940 20140
rect 1708 20012 1748 20107
rect 1708 19963 1748 19972
rect 1804 20096 1844 20105
rect 1420 18668 1460 18677
rect 1420 17156 1460 18628
rect 1516 18500 1556 18509
rect 1516 17912 1556 18460
rect 1516 17863 1556 17872
rect 1612 17744 1652 19216
rect 1708 19844 1748 19853
rect 1708 18752 1748 19804
rect 1708 18703 1748 18712
rect 1804 18752 1844 20056
rect 1996 19844 2036 22996
rect 2092 22280 2132 24760
rect 2092 22231 2132 22240
rect 2380 22028 2420 22037
rect 2284 21608 2324 21617
rect 2092 21524 2132 21533
rect 2092 20852 2132 21484
rect 2092 20803 2132 20812
rect 2188 21356 2228 21365
rect 2188 20768 2228 21316
rect 2188 20264 2228 20728
rect 2188 20215 2228 20224
rect 1996 19795 2036 19804
rect 2092 20096 2132 20105
rect 2092 19928 2132 20056
rect 1900 19172 1940 19181
rect 1900 19037 1940 19132
rect 2092 18920 2132 19888
rect 2092 18871 2132 18880
rect 2188 19844 2228 19853
rect 1804 18703 1844 18712
rect 1708 18584 1748 18593
rect 1708 18332 1748 18544
rect 1900 18584 1940 18593
rect 1708 18283 1748 18292
rect 1804 18500 1844 18509
rect 1804 18248 1844 18460
rect 1804 18199 1844 18208
rect 1420 17107 1460 17116
rect 1516 17704 1612 17744
rect 1516 17072 1556 17704
rect 1612 17695 1652 17704
rect 1708 17828 1748 17837
rect 1516 17023 1556 17032
rect 1612 17156 1652 17165
rect 1420 16988 1460 16997
rect 1420 16400 1460 16948
rect 1420 16351 1460 16360
rect 1612 16316 1652 17116
rect 1708 17072 1748 17788
rect 1804 17828 1844 17837
rect 1804 17492 1844 17788
rect 1804 17357 1844 17452
rect 1900 17300 1940 18544
rect 2092 18500 2132 18509
rect 2092 18332 2132 18460
rect 2092 18283 2132 18292
rect 1996 17912 2036 17921
rect 1996 17660 2036 17872
rect 2188 17828 2228 19804
rect 2188 17779 2228 17788
rect 2284 19256 2324 21568
rect 2380 21104 2420 21988
rect 2380 21055 2420 21064
rect 2284 17828 2324 19216
rect 2380 20600 2420 20609
rect 2380 20348 2420 20560
rect 2380 19424 2420 20308
rect 2380 18668 2420 19384
rect 2476 19088 2516 24844
rect 2572 24464 2612 25180
rect 2572 24415 2612 24424
rect 2668 23876 2708 23885
rect 2668 23792 2708 23836
rect 2668 23741 2708 23752
rect 2764 23792 2804 26608
rect 2956 26396 2996 26692
rect 3148 26732 3188 26860
rect 3340 26900 3380 27028
rect 3340 26851 3380 26860
rect 3628 26984 3668 26993
rect 3628 26849 3668 26944
rect 3148 26683 3188 26692
rect 2860 26356 2996 26396
rect 2860 26144 2900 26356
rect 3532 26312 3572 26321
rect 2860 26095 2900 26104
rect 3436 26228 3476 26237
rect 3436 26060 3476 26188
rect 3436 26011 3476 26020
rect 3112 25724 3480 25733
rect 3112 25675 3480 25684
rect 3532 25556 3572 26272
rect 3628 26060 3668 26069
rect 3628 25925 3668 26020
rect 3532 25507 3572 25516
rect 3148 25304 3188 25313
rect 3148 25169 3188 25264
rect 3340 24800 3380 24809
rect 3340 24548 3380 24760
rect 3340 24413 3380 24508
rect 3724 24548 3764 27364
rect 3820 27236 3860 27532
rect 3916 27404 3956 28600
rect 4108 28496 4148 28505
rect 4108 27824 4148 28456
rect 4684 28160 4724 28600
rect 4684 28111 4724 28120
rect 4876 28580 4916 28589
rect 4352 27992 4720 28001
rect 4352 27943 4720 27952
rect 4108 27775 4148 27784
rect 4396 27656 4436 27665
rect 3916 27355 3956 27364
rect 4204 27572 4244 27581
rect 4012 27320 4052 27329
rect 3820 27196 3956 27236
rect 3724 24499 3764 24508
rect 3820 26228 3860 26237
rect 3532 24380 3572 24389
rect 3112 24212 3480 24221
rect 3112 24163 3480 24172
rect 2764 23743 2804 23752
rect 3052 23708 3092 23717
rect 2572 23288 2612 23297
rect 2572 22280 2612 23248
rect 2860 23204 2900 23213
rect 2860 22784 2900 23164
rect 3052 23204 3092 23668
rect 3532 23624 3572 24340
rect 3532 23575 3572 23584
rect 3724 24380 3764 24389
rect 3052 23155 3092 23164
rect 3340 23120 3380 23129
rect 3340 23036 3380 23080
rect 3340 22985 3380 22996
rect 2572 22231 2612 22240
rect 2764 22744 2900 22784
rect 3532 22952 3572 22961
rect 2764 21860 2804 22744
rect 3112 22700 3480 22709
rect 3112 22651 3480 22660
rect 2860 22112 2900 22121
rect 2860 21977 2900 22072
rect 3436 22028 3476 22037
rect 3340 21944 3380 21953
rect 2764 21820 2996 21860
rect 2572 21776 2612 21785
rect 2572 21440 2612 21736
rect 2668 21608 2708 21617
rect 2668 21473 2708 21568
rect 2860 21524 2900 21533
rect 2572 21305 2612 21400
rect 2860 21272 2900 21484
rect 2956 21524 2996 21820
rect 2956 21475 2996 21484
rect 3148 21608 3188 21617
rect 3148 21356 3188 21568
rect 3340 21440 3380 21904
rect 3436 21608 3476 21988
rect 3436 21559 3476 21568
rect 3340 21391 3380 21400
rect 2860 21223 2900 21232
rect 2956 21316 3188 21356
rect 3436 21356 3476 21451
rect 2956 21104 2996 21316
rect 3436 21307 3476 21316
rect 3112 21188 3480 21197
rect 3112 21139 3480 21148
rect 2956 21055 2996 21064
rect 2668 20852 2708 20861
rect 2572 20096 2612 20105
rect 2572 19340 2612 20056
rect 2572 19291 2612 19300
rect 2476 19048 2612 19088
rect 2476 18920 2516 18929
rect 2476 18785 2516 18880
rect 2380 18619 2420 18628
rect 2380 18500 2420 18509
rect 2380 18080 2420 18460
rect 2476 18416 2516 18425
rect 2476 18281 2516 18376
rect 2380 18031 2420 18040
rect 2284 17744 2324 17788
rect 2380 17912 2420 17921
rect 2380 17777 2420 17872
rect 2284 17664 2324 17704
rect 1996 17620 2228 17660
rect 1900 17260 2036 17300
rect 1900 17156 1940 17165
rect 1708 17032 1844 17072
rect 1420 16064 1460 16073
rect 1420 15929 1460 16024
rect 1420 15644 1460 15653
rect 1420 15476 1460 15604
rect 1612 15560 1652 16276
rect 1708 16904 1748 16913
rect 1708 16232 1748 16864
rect 1708 16183 1748 16192
rect 1708 15728 1748 15737
rect 1708 15593 1748 15688
rect 1612 15511 1652 15520
rect 1420 15427 1460 15436
rect 1516 15392 1556 15401
rect 1420 14468 1460 14477
rect 1420 11948 1460 14428
rect 1420 11899 1460 11908
rect 1420 11780 1460 11789
rect 1420 8168 1460 11740
rect 1516 9428 1556 15352
rect 1804 14972 1844 17032
rect 1900 16988 1940 17116
rect 1900 16939 1940 16948
rect 1996 17156 2036 17260
rect 1996 17048 2036 17116
rect 1996 16484 2036 17008
rect 1996 15644 2036 16444
rect 2092 16946 2132 16955
rect 2092 16316 2132 16906
rect 2092 16267 2132 16276
rect 1996 15595 2036 15604
rect 1804 14923 1844 14932
rect 2092 14804 2132 14813
rect 1612 14132 1652 14141
rect 1612 13997 1652 14092
rect 1900 14048 1940 14057
rect 1804 13208 1844 13217
rect 1804 12704 1844 13168
rect 1804 12655 1844 12664
rect 1708 12536 1748 12547
rect 1708 12452 1748 12496
rect 1708 12403 1748 12412
rect 1708 11696 1748 11705
rect 1612 11612 1652 11621
rect 1612 11192 1652 11572
rect 1612 11143 1652 11152
rect 1612 11024 1652 11033
rect 1612 10268 1652 10984
rect 1612 10219 1652 10228
rect 1516 9379 1556 9388
rect 1612 10100 1652 10109
rect 1420 8119 1460 8128
rect 1516 8084 1556 8093
rect 1516 7244 1556 8044
rect 1324 6523 1364 6532
rect 1420 7076 1460 7085
rect 1420 6404 1460 7036
rect 1516 6740 1556 7204
rect 1612 6992 1652 10060
rect 1708 9764 1748 11656
rect 1900 11696 1940 14008
rect 2092 13880 2132 14764
rect 2092 13831 2132 13840
rect 2188 12980 2228 17620
rect 2380 17576 2420 17585
rect 2380 17240 2420 17536
rect 2572 17492 2612 19048
rect 2668 18740 2708 20812
rect 2860 20768 2900 20777
rect 2860 20684 2900 20728
rect 2764 20432 2804 20441
rect 2764 18836 2804 20392
rect 2860 19340 2900 20644
rect 2956 20768 2996 20777
rect 2956 20348 2996 20728
rect 2956 20299 2996 20308
rect 3340 20768 3380 20777
rect 3148 20264 3188 20273
rect 2860 19004 2900 19300
rect 2860 18955 2900 18964
rect 2956 20012 2996 20021
rect 2956 18920 2996 19972
rect 3148 19844 3188 20224
rect 3244 20180 3284 20189
rect 3244 20045 3284 20140
rect 3340 20096 3380 20728
rect 3436 20432 3476 20441
rect 3436 20297 3476 20392
rect 3340 20047 3380 20056
rect 3340 19844 3380 19853
rect 3148 19804 3340 19844
rect 3340 19795 3380 19804
rect 3112 19676 3480 19685
rect 3112 19627 3480 19636
rect 3532 19340 3572 22912
rect 3724 21692 3764 24340
rect 3820 23120 3860 26188
rect 3916 24464 3956 27196
rect 3916 24415 3956 24424
rect 3820 23071 3860 23080
rect 3916 23204 3956 23213
rect 3916 23120 3956 23164
rect 3916 23069 3956 23080
rect 3916 22280 3956 22289
rect 3724 21557 3764 21652
rect 3820 22112 3860 22121
rect 3820 21608 3860 22072
rect 3820 21559 3860 21568
rect 3436 19300 3572 19340
rect 3628 21524 3668 21533
rect 3148 19172 3188 19181
rect 3148 19037 3188 19132
rect 3340 18920 3380 18929
rect 2956 18880 3188 18920
rect 2860 18836 2900 18845
rect 2764 18796 2860 18836
rect 2860 18787 2900 18796
rect 2668 18691 2708 18700
rect 2860 18668 2900 18677
rect 2668 18416 2708 18425
rect 2668 17996 2708 18376
rect 2860 18416 2900 18628
rect 3052 18668 3092 18677
rect 3052 18500 3092 18628
rect 3148 18584 3188 18880
rect 3340 18752 3380 18880
rect 3340 18703 3380 18712
rect 3148 18535 3188 18544
rect 3052 18451 3092 18460
rect 2860 18367 2900 18376
rect 2764 18332 2804 18341
rect 2764 18197 2804 18292
rect 2956 18332 2996 18341
rect 2668 17947 2708 17956
rect 2860 17744 2900 17839
rect 2860 17695 2900 17704
rect 2668 17660 2708 17669
rect 2668 17525 2708 17620
rect 2956 17660 2996 18292
rect 3436 18332 3476 19300
rect 3436 18283 3476 18292
rect 3532 19172 3572 19181
rect 3532 18584 3572 19132
rect 3112 18164 3480 18173
rect 3112 18115 3480 18124
rect 3532 17996 3572 18544
rect 3436 17956 3572 17996
rect 3244 17744 3284 17753
rect 2860 17576 2900 17585
rect 2572 17443 2612 17452
rect 2860 17492 2900 17536
rect 2860 17441 2900 17452
rect 2380 17191 2420 17200
rect 2476 17156 2516 17165
rect 2476 17021 2516 17116
rect 2572 17072 2612 17083
rect 2956 17072 2996 17620
rect 3148 17660 3188 17669
rect 2284 16988 2324 16997
rect 2284 15980 2324 16948
rect 2572 16988 2612 17032
rect 2860 17032 2996 17072
rect 3052 17408 3092 17417
rect 2572 16939 2612 16948
rect 2668 16988 2708 16997
rect 2476 16904 2516 16913
rect 2380 16820 2420 16829
rect 2380 16685 2420 16780
rect 2380 16232 2420 16241
rect 2380 16097 2420 16192
rect 2284 15940 2420 15980
rect 2284 15644 2324 15653
rect 2284 15509 2324 15604
rect 2380 15476 2420 15940
rect 2476 15896 2516 16864
rect 2668 16400 2708 16948
rect 2668 16351 2708 16360
rect 2764 16484 2804 16493
rect 2764 16232 2804 16444
rect 2668 16192 2804 16232
rect 2476 15847 2516 15856
rect 2572 16148 2612 16157
rect 2572 15812 2612 16108
rect 2572 15763 2612 15772
rect 2668 15644 2708 16192
rect 2764 16064 2804 16073
rect 2764 15929 2804 16024
rect 2668 15595 2708 15604
rect 2860 15644 2900 17032
rect 2860 15595 2900 15604
rect 2956 16904 2996 16913
rect 3052 16904 3092 17368
rect 3148 17156 3188 17620
rect 3244 17609 3284 17704
rect 3436 17240 3476 17956
rect 3628 17744 3668 21484
rect 3820 21272 3860 21281
rect 3724 21188 3764 21197
rect 3724 20852 3764 21148
rect 3724 20803 3764 20812
rect 3724 20684 3764 20693
rect 3724 20549 3764 20644
rect 3724 20180 3764 20189
rect 3724 20096 3764 20140
rect 3724 20045 3764 20056
rect 3820 20012 3860 21232
rect 3916 20936 3956 22240
rect 3916 20887 3956 20896
rect 3820 19963 3860 19972
rect 3916 20600 3956 20609
rect 3724 19760 3764 19769
rect 3724 18752 3764 19720
rect 3820 19256 3860 19351
rect 3820 19207 3860 19216
rect 3724 18703 3764 18712
rect 3820 19088 3860 19097
rect 3724 18248 3764 18257
rect 3724 17996 3764 18208
rect 3724 17947 3764 17956
rect 3628 17695 3668 17704
rect 3724 17828 3764 17839
rect 3724 17744 3764 17788
rect 3724 17695 3764 17704
rect 3436 17191 3476 17200
rect 3532 17660 3572 17669
rect 3148 17107 3188 17116
rect 3532 16988 3572 17620
rect 3532 16939 3572 16948
rect 3628 17492 3668 17501
rect 2996 16864 3092 16904
rect 2956 15980 2996 16864
rect 3112 16652 3480 16661
rect 3112 16603 3480 16612
rect 3436 16316 3476 16325
rect 2380 15427 2420 15436
rect 2956 15476 2996 15940
rect 3340 16064 3380 16073
rect 3340 15644 3380 16024
rect 3436 15728 3476 16276
rect 3628 16148 3668 17452
rect 3820 17408 3860 19048
rect 3820 17359 3860 17368
rect 3820 16400 3860 16409
rect 3820 16265 3860 16360
rect 3628 16099 3668 16108
rect 3820 16148 3860 16157
rect 3436 15679 3476 15688
rect 3724 15812 3764 15821
rect 3340 15595 3380 15604
rect 2956 15427 2996 15436
rect 2572 15392 2612 15401
rect 2476 15224 2516 15233
rect 2476 15089 2516 15184
rect 2572 15056 2612 15352
rect 2572 15007 2612 15016
rect 2668 15224 2708 15233
rect 2668 14720 2708 15184
rect 3112 15140 3480 15149
rect 3112 15091 3480 15100
rect 3724 15056 3764 15772
rect 3820 15560 3860 16108
rect 3820 15511 3860 15520
rect 3628 15016 3764 15056
rect 3820 15308 3860 15317
rect 2668 14671 2708 14680
rect 3148 14720 3188 14729
rect 2668 14552 2708 14561
rect 2380 14132 2420 14141
rect 2380 13208 2420 14092
rect 2572 14048 2612 14057
rect 2572 13460 2612 14008
rect 2572 13411 2612 13420
rect 2188 12940 2324 12980
rect 1900 11647 1940 11656
rect 1804 11444 1844 11453
rect 1804 11024 1844 11404
rect 2092 11024 2132 11033
rect 1804 10975 1844 10984
rect 1900 10984 2092 11024
rect 1708 9715 1748 9724
rect 1804 10184 1844 10193
rect 1900 10184 1940 10984
rect 2092 10975 2132 10984
rect 2188 10940 2228 10949
rect 1996 10856 2036 10865
rect 1996 10436 2036 10816
rect 1996 10387 2036 10396
rect 1844 10144 1940 10184
rect 1996 10268 2036 10277
rect 1804 9512 1844 10144
rect 1708 9472 1844 9512
rect 1708 7412 1748 9472
rect 1708 7363 1748 7372
rect 1804 8000 1844 8009
rect 1612 6943 1652 6952
rect 1804 6992 1844 7960
rect 1900 7160 1940 7169
rect 1900 7025 1940 7120
rect 1516 6691 1556 6700
rect 1420 6355 1460 6364
rect 1804 6404 1844 6952
rect 1996 6656 2036 10228
rect 2092 10268 2132 10277
rect 2092 8588 2132 10228
rect 2092 8168 2132 8548
rect 2092 8119 2132 8128
rect 2092 8000 2132 8009
rect 2092 7916 2132 7960
rect 2092 7865 2132 7876
rect 2188 7916 2228 10900
rect 2284 10184 2324 12940
rect 2380 12620 2420 13168
rect 2380 12571 2420 12580
rect 2380 11780 2420 11789
rect 2380 11645 2420 11740
rect 2380 11192 2420 11201
rect 2380 11024 2420 11152
rect 2380 10975 2420 10984
rect 2476 10352 2516 10361
rect 2284 10144 2420 10184
rect 2188 7867 2228 7876
rect 2284 9848 2324 9857
rect 2284 8000 2324 9808
rect 2188 7748 2228 7757
rect 2188 7328 2228 7708
rect 2284 7412 2324 7960
rect 2380 7496 2420 10144
rect 2476 10100 2516 10312
rect 2476 10051 2516 10060
rect 2572 10184 2612 10193
rect 2380 7447 2420 7456
rect 2476 8756 2516 8765
rect 2284 7363 2324 7372
rect 2188 7279 2228 7288
rect 1996 6607 2036 6616
rect 2284 6656 2324 6665
rect 2284 6521 2324 6616
rect 1804 6355 1844 6364
rect 2188 6488 2228 6497
rect 1036 6271 1076 6280
rect 2188 6320 2228 6448
rect 2188 6271 2228 6280
rect 2476 6320 2516 8716
rect 2572 8420 2612 10144
rect 2668 9680 2708 14512
rect 2956 14048 2996 14057
rect 2956 13208 2996 14008
rect 3148 13796 3188 14680
rect 3628 14720 3668 15016
rect 3628 14552 3668 14680
rect 3628 14503 3668 14512
rect 3724 14636 3764 14645
rect 3244 14300 3284 14309
rect 3244 14048 3284 14260
rect 3244 13999 3284 14008
rect 3148 13747 3188 13756
rect 3436 13796 3476 13891
rect 3436 13747 3476 13756
rect 3628 13796 3668 13805
rect 3112 13628 3480 13637
rect 3112 13579 3480 13588
rect 2956 12704 2996 13168
rect 2956 12655 2996 12664
rect 2956 12536 2996 12545
rect 2956 12368 2996 12496
rect 2764 12328 2996 12368
rect 3052 12452 3092 12461
rect 2764 11192 2804 12328
rect 3052 12284 3092 12412
rect 2764 11143 2804 11152
rect 2956 12244 3092 12284
rect 2956 10436 2996 12244
rect 3112 12116 3480 12125
rect 3112 12067 3480 12076
rect 3052 11864 3092 11873
rect 3052 11612 3092 11824
rect 3052 11192 3092 11572
rect 3052 11143 3092 11152
rect 3148 11780 3188 11789
rect 3148 11108 3188 11740
rect 3340 11696 3380 11705
rect 3340 11192 3380 11656
rect 3340 11143 3380 11152
rect 3148 11059 3188 11068
rect 3628 11108 3668 13756
rect 3724 11360 3764 14596
rect 3724 11311 3764 11320
rect 3820 11108 3860 15268
rect 3916 14300 3956 20560
rect 4012 20180 4052 27280
rect 4108 26648 4148 26657
rect 4108 25388 4148 26608
rect 4204 26312 4244 27532
rect 4396 27488 4436 27616
rect 4396 27439 4436 27448
rect 4492 27656 4532 27665
rect 4492 26816 4532 27616
rect 4876 27488 4916 28540
rect 5356 27992 5396 28001
rect 4972 27908 5012 27917
rect 4972 27824 5012 27868
rect 4972 27784 5204 27824
rect 4876 27439 4916 27448
rect 5068 27656 5108 27665
rect 4972 27320 5012 27329
rect 4492 26767 4532 26776
rect 4588 27236 4628 27245
rect 4588 26816 4628 27196
rect 4972 27185 5012 27280
rect 4588 26767 4628 26776
rect 4780 26900 4820 26909
rect 4352 26480 4720 26489
rect 4352 26431 4720 26440
rect 4204 26272 4532 26312
rect 4108 25339 4148 25348
rect 4204 26144 4244 26153
rect 4108 25220 4148 25229
rect 4108 25085 4148 25180
rect 4204 24632 4244 26104
rect 4492 25304 4532 26272
rect 4492 25255 4532 25264
rect 4352 24968 4720 24977
rect 4352 24919 4720 24928
rect 4492 24800 4532 24809
rect 4492 24665 4532 24760
rect 4396 24632 4436 24641
rect 4204 23792 4244 24592
rect 4204 23743 4244 23752
rect 4300 24592 4396 24632
rect 4300 23624 4340 24592
rect 4396 24497 4436 24592
rect 4780 24044 4820 26860
rect 4876 26816 4916 26825
rect 4876 26312 4916 26776
rect 4876 24884 4916 26272
rect 4972 26732 5012 26741
rect 4972 25556 5012 26692
rect 4972 25507 5012 25516
rect 4876 24380 4916 24844
rect 4972 24968 5012 24977
rect 4972 24716 5012 24928
rect 4972 24667 5012 24676
rect 5068 24884 5108 27616
rect 5068 24632 5108 24844
rect 5068 24583 5108 24592
rect 4876 24331 4916 24340
rect 4780 23995 4820 24004
rect 4876 23792 4916 23801
rect 4300 23575 4340 23584
rect 4780 23708 4820 23717
rect 4352 23456 4720 23465
rect 4352 23407 4720 23416
rect 4108 23288 4148 23297
rect 4108 23036 4148 23248
rect 4300 23288 4340 23297
rect 4300 23120 4340 23248
rect 4780 23288 4820 23668
rect 4780 23239 4820 23248
rect 4300 23071 4340 23080
rect 4108 22987 4148 22996
rect 4684 23036 4724 23045
rect 4588 22700 4628 22709
rect 4204 22364 4244 22373
rect 4108 22196 4148 22205
rect 4108 22061 4148 22156
rect 4204 21944 4244 22324
rect 4396 22280 4436 22291
rect 4396 22196 4436 22240
rect 4396 22147 4436 22156
rect 4588 22112 4628 22660
rect 4684 22364 4724 22996
rect 4876 22700 4916 23752
rect 5068 23624 5108 23633
rect 5068 23120 5108 23584
rect 5068 23036 5108 23080
rect 5068 22987 5108 22996
rect 4876 22651 4916 22660
rect 5164 22616 5204 27784
rect 5260 27656 5300 27665
rect 5260 26480 5300 27616
rect 5356 27572 5396 27952
rect 5356 27523 5396 27532
rect 5260 26431 5300 26440
rect 5452 26312 5492 28600
rect 5452 26263 5492 26272
rect 5548 27824 5588 27833
rect 5548 27572 5588 27784
rect 5644 27656 5684 28624
rect 6200 28600 6280 29000
rect 6968 28600 7048 29000
rect 7736 28600 7816 29000
rect 8504 28600 8584 29000
rect 9272 28600 9352 29000
rect 10040 28600 10120 29000
rect 10808 28600 10888 29000
rect 11576 28600 11656 29000
rect 12344 28600 12424 29000
rect 12652 28664 12692 28673
rect 6220 27908 6260 28600
rect 6220 27859 6260 27868
rect 6892 27740 6932 27749
rect 5644 27607 5684 27616
rect 5740 27656 5780 27665
rect 5548 26816 5588 27532
rect 5356 26144 5396 26153
rect 5260 25808 5300 25817
rect 5260 25388 5300 25768
rect 5260 24632 5300 25348
rect 5260 24583 5300 24592
rect 4724 22324 4916 22364
rect 4684 22315 4724 22324
rect 4698 22121 4738 22193
rect 4588 22063 4628 22072
rect 4684 22112 4738 22121
rect 4684 22063 4738 22072
rect 4012 20131 4052 20140
rect 4108 21904 4244 21944
rect 4352 21944 4720 21953
rect 4012 20012 4052 20021
rect 4012 18584 4052 19972
rect 4012 16988 4052 18544
rect 4012 16939 4052 16948
rect 4108 16484 4148 21904
rect 4352 21895 4720 21904
rect 4780 21860 4820 21869
rect 4492 21776 4532 21785
rect 4492 21692 4532 21736
rect 4492 21641 4532 21652
rect 4780 21692 4820 21820
rect 4780 21643 4820 21652
rect 4204 21608 4244 21617
rect 4204 21272 4244 21568
rect 4588 21608 4628 21619
rect 4588 21524 4628 21568
rect 4876 21608 4916 22324
rect 4588 21475 4628 21484
rect 4684 21524 4724 21533
rect 4876 21524 4916 21568
rect 4724 21484 4916 21524
rect 4684 21475 4724 21484
rect 4876 21473 4916 21484
rect 4972 22280 5012 22289
rect 4972 21440 5012 22240
rect 5068 21944 5108 21955
rect 5068 21860 5108 21904
rect 5068 21811 5108 21820
rect 5164 21776 5204 22576
rect 5164 21727 5204 21736
rect 5260 23876 5300 23885
rect 5164 21608 5204 21617
rect 4972 21391 5012 21400
rect 5068 21524 5108 21533
rect 4204 21223 4244 21232
rect 4300 21272 4340 21281
rect 4300 21188 4340 21232
rect 4300 21137 4340 21148
rect 4876 21188 4916 21197
rect 4204 21104 4244 21113
rect 4204 19760 4244 21064
rect 4780 20600 4820 20609
rect 4352 20432 4720 20441
rect 4352 20383 4720 20392
rect 4492 20264 4532 20273
rect 4492 20096 4532 20224
rect 4396 20012 4436 20021
rect 4396 19877 4436 19972
rect 4492 19844 4532 20056
rect 4684 20012 4724 20021
rect 4780 20012 4820 20560
rect 4724 19972 4820 20012
rect 4684 19963 4724 19972
rect 4492 19795 4532 19804
rect 4204 19256 4244 19720
rect 4876 19424 4916 21148
rect 4876 19375 4916 19384
rect 4972 20600 5012 20609
rect 4972 19508 5012 20560
rect 5068 20348 5108 21484
rect 5164 21473 5204 21568
rect 5164 21104 5204 21113
rect 5164 20936 5204 21064
rect 5164 20887 5204 20896
rect 5164 20768 5204 20777
rect 5164 20600 5204 20728
rect 5164 20551 5204 20560
rect 5068 20299 5108 20308
rect 5068 20180 5108 20189
rect 5068 20045 5108 20140
rect 5164 20012 5204 20021
rect 4204 19207 4244 19216
rect 4396 19256 4436 19265
rect 4396 19088 4436 19216
rect 4588 19172 4628 19267
rect 4588 19123 4628 19132
rect 4780 19172 4820 19181
rect 4972 19172 5012 19468
rect 4396 19039 4436 19048
rect 4204 19004 4244 19013
rect 4204 18836 4244 18964
rect 4352 18920 4720 18929
rect 4352 18871 4720 18880
rect 4204 17744 4244 18796
rect 4780 18752 4820 19132
rect 4780 18703 4820 18712
rect 4876 19132 5012 19172
rect 5068 19928 5108 19937
rect 4876 18080 4916 19132
rect 4780 18040 4916 18080
rect 4972 19004 5012 19013
rect 4780 17828 4820 18040
rect 4780 17779 4820 17788
rect 4876 17912 4916 17921
rect 4876 17777 4916 17872
rect 4204 17695 4244 17704
rect 4780 17576 4820 17587
rect 4780 17492 4820 17536
rect 4780 17443 4820 17452
rect 4876 17576 4916 17585
rect 4352 17408 4720 17417
rect 4352 17359 4720 17368
rect 4876 17324 4916 17536
rect 4876 17275 4916 17284
rect 4780 17156 4820 17165
rect 4780 17021 4820 17116
rect 4876 16568 4916 16577
rect 4876 16484 4916 16528
rect 4108 16444 4244 16484
rect 4108 16316 4148 16325
rect 4012 15728 4052 15737
rect 4012 15593 4052 15688
rect 4108 15644 4148 16276
rect 4108 15595 4148 15604
rect 3916 13208 3956 14260
rect 3916 13159 3956 13168
rect 4012 15140 4052 15149
rect 3916 12956 3956 12965
rect 3916 12536 3956 12916
rect 3916 12487 3956 12496
rect 3820 11068 3956 11108
rect 3628 11059 3668 11068
rect 3340 11024 3380 11033
rect 3340 10772 3380 10984
rect 3820 10940 3860 10949
rect 3532 10900 3820 10940
rect 3532 10772 3572 10900
rect 3820 10891 3860 10900
rect 3340 10732 3572 10772
rect 3112 10604 3480 10613
rect 3112 10555 3480 10564
rect 2956 10387 2996 10396
rect 3532 10436 3572 10732
rect 3532 10387 3572 10396
rect 3820 10772 3860 10781
rect 3340 10352 3380 10361
rect 2668 9631 2708 9640
rect 2764 10268 2804 10277
rect 2572 8371 2612 8380
rect 2764 7916 2804 10228
rect 2956 10268 2996 10277
rect 2956 10184 2996 10228
rect 2668 7876 2764 7916
rect 2572 7832 2612 7841
rect 2572 6992 2612 7792
rect 2572 6943 2612 6952
rect 2668 6908 2708 7876
rect 2764 7867 2804 7876
rect 2860 10016 2900 10025
rect 2668 6859 2708 6868
rect 2764 6572 2804 6581
rect 2860 6572 2900 9976
rect 2956 9848 2996 10144
rect 2956 9799 2996 9808
rect 2956 9680 2996 9689
rect 2956 8840 2996 9640
rect 3340 9428 3380 10312
rect 3628 10352 3668 10361
rect 3436 10184 3476 10279
rect 3628 10217 3668 10312
rect 3436 10135 3476 10144
rect 3820 10184 3860 10732
rect 3820 10135 3860 10144
rect 3820 10016 3860 10025
rect 3436 9932 3476 9941
rect 3436 9512 3476 9892
rect 3724 9512 3764 9521
rect 3476 9472 3572 9512
rect 3436 9463 3476 9472
rect 3340 9379 3380 9388
rect 3112 9092 3480 9101
rect 3112 9043 3480 9052
rect 2956 8800 3092 8840
rect 2804 6532 2900 6572
rect 2956 8672 2996 8681
rect 2956 6572 2996 8632
rect 3052 7748 3092 8800
rect 3052 7699 3092 7708
rect 3112 7580 3480 7589
rect 3112 7531 3480 7540
rect 3340 7328 3380 7337
rect 3052 7244 3092 7253
rect 3052 7160 3092 7204
rect 3052 7109 3092 7120
rect 2764 6523 2804 6532
rect 2956 6523 2996 6532
rect 3340 6488 3380 7288
rect 3436 7160 3476 7169
rect 3532 7160 3572 9472
rect 3724 8924 3764 9472
rect 3476 7120 3572 7160
rect 3628 8884 3724 8924
rect 3436 7111 3476 7120
rect 3628 7076 3668 8884
rect 3724 8875 3764 8884
rect 3820 9512 3860 9976
rect 3724 8420 3764 8429
rect 3724 8000 3764 8380
rect 3820 8168 3860 9472
rect 3820 8033 3860 8128
rect 3724 7951 3764 7960
rect 3724 7664 3764 7673
rect 3724 7160 3764 7624
rect 3724 7111 3764 7120
rect 3628 7027 3668 7036
rect 3820 6992 3860 7001
rect 3340 6439 3380 6448
rect 3532 6656 3572 6665
rect 2476 6271 2516 6280
rect 3112 6068 3480 6077
rect 3112 6019 3480 6028
rect 3532 5648 3572 6616
rect 3724 6404 3764 6413
rect 3724 5900 3764 6364
rect 3724 5851 3764 5860
rect 3820 5816 3860 6952
rect 3916 6740 3956 11068
rect 4012 6824 4052 15100
rect 4204 14972 4244 16444
rect 4876 16433 4916 16444
rect 4396 16400 4436 16409
rect 4396 16232 4436 16360
rect 4396 16183 4436 16192
rect 4492 16316 4532 16325
rect 4492 16148 4532 16276
rect 4492 16099 4532 16108
rect 4684 16316 4724 16325
rect 4684 16148 4724 16276
rect 4684 16099 4724 16108
rect 4352 15896 4720 15905
rect 4352 15847 4720 15856
rect 4876 15812 4916 15821
rect 4396 15560 4436 15569
rect 4204 14923 4244 14932
rect 4300 15476 4340 15485
rect 4204 14804 4244 14815
rect 4204 14720 4244 14764
rect 4204 14671 4244 14680
rect 4108 14636 4148 14645
rect 4108 14468 4148 14596
rect 4300 14552 4340 15436
rect 4396 14804 4436 15520
rect 4780 15224 4820 15233
rect 4396 14755 4436 14764
rect 4588 15140 4628 15149
rect 4108 14419 4148 14428
rect 4204 14512 4340 14552
rect 4588 14720 4628 15100
rect 4588 14552 4628 14680
rect 4108 14300 4148 14309
rect 4108 11528 4148 14260
rect 4204 14300 4244 14512
rect 4588 14503 4628 14512
rect 4780 14468 4820 15184
rect 4780 14419 4820 14428
rect 4876 14972 4916 15772
rect 4352 14384 4720 14393
rect 4352 14335 4720 14344
rect 4204 14251 4244 14260
rect 4876 14300 4916 14932
rect 4876 14251 4916 14260
rect 4972 14216 5012 18964
rect 5068 17912 5108 19888
rect 5164 19760 5204 19972
rect 5164 19711 5204 19720
rect 5164 18752 5204 18761
rect 5164 18617 5204 18712
rect 5068 17863 5108 17872
rect 5164 18500 5204 18509
rect 5068 17660 5108 17669
rect 5068 17525 5108 17620
rect 5068 17324 5108 17333
rect 5068 17156 5108 17284
rect 5068 17107 5108 17116
rect 5068 16988 5108 16997
rect 5068 16484 5108 16948
rect 5068 16435 5108 16444
rect 5164 16400 5204 18460
rect 5164 16351 5204 16360
rect 4972 14167 5012 14176
rect 5068 16148 5108 16157
rect 4684 14048 4724 14057
rect 4300 13964 4340 13975
rect 4204 13880 4244 13889
rect 4204 11864 4244 13840
rect 4300 13880 4340 13924
rect 4300 13831 4340 13840
rect 4684 13124 4724 14008
rect 4876 13964 4916 13973
rect 4684 13075 4724 13084
rect 4780 13124 4820 13133
rect 4352 12872 4720 12881
rect 4352 12823 4720 12832
rect 4396 12704 4436 12713
rect 4300 12536 4340 12545
rect 4300 12401 4340 12496
rect 4204 11815 4244 11824
rect 4108 11276 4148 11488
rect 4108 11227 4148 11236
rect 4204 11696 4244 11705
rect 4108 11108 4148 11117
rect 4108 7916 4148 11068
rect 4204 10268 4244 11656
rect 4396 11696 4436 12664
rect 4780 12704 4820 13084
rect 4780 12655 4820 12664
rect 4492 12620 4532 12629
rect 4492 12485 4532 12580
rect 4396 11647 4436 11656
rect 4780 12452 4820 12461
rect 4352 11360 4720 11369
rect 4352 11311 4720 11320
rect 4684 11192 4724 11201
rect 4588 11108 4628 11117
rect 4396 11024 4436 11033
rect 4396 10889 4436 10984
rect 4588 10973 4628 11068
rect 4684 11024 4724 11152
rect 4204 10219 4244 10228
rect 4492 10268 4532 10277
rect 4396 10184 4436 10195
rect 4396 10100 4436 10144
rect 4492 10133 4532 10228
rect 4396 10051 4436 10060
rect 4204 10016 4244 10025
rect 4204 9428 4244 9976
rect 4684 10016 4724 10984
rect 4780 10436 4820 12412
rect 4780 10387 4820 10396
rect 4876 10268 4916 13924
rect 5068 13376 5108 16108
rect 5164 15980 5204 16020
rect 5164 15896 5204 15940
rect 5164 15644 5204 15856
rect 5164 15595 5204 15604
rect 5068 13327 5108 13336
rect 5164 15308 5204 15317
rect 4972 13208 5012 13217
rect 5164 13208 5204 15268
rect 4972 12620 5012 13168
rect 4972 12571 5012 12580
rect 5068 13168 5204 13208
rect 5068 12452 5108 13168
rect 5260 12980 5300 23836
rect 5356 19760 5396 26104
rect 5452 26060 5492 26069
rect 5452 20348 5492 26020
rect 5548 24632 5588 26776
rect 5548 23204 5588 24592
rect 5644 26396 5684 26405
rect 5644 23288 5684 26356
rect 5740 26144 5780 27616
rect 6220 27656 6260 27665
rect 6220 27521 6260 27616
rect 6700 27656 6740 27665
rect 6316 27572 6356 27581
rect 5740 26095 5780 26104
rect 5932 27488 5972 27497
rect 5644 23239 5684 23248
rect 5740 25640 5780 25649
rect 5548 23155 5588 23164
rect 5644 23036 5684 23045
rect 5548 22700 5588 22709
rect 5548 20600 5588 22660
rect 5644 22448 5684 22996
rect 5644 22399 5684 22408
rect 5644 22280 5684 22289
rect 5644 21440 5684 22240
rect 5644 20768 5684 21400
rect 5740 21692 5780 25600
rect 5836 23708 5876 23719
rect 5836 23624 5876 23668
rect 5836 23575 5876 23584
rect 5740 21356 5780 21652
rect 5740 21307 5780 21316
rect 5836 22868 5876 22877
rect 5644 20719 5684 20728
rect 5740 21188 5780 21197
rect 5548 20560 5684 20600
rect 5452 20299 5492 20308
rect 5452 20180 5492 20189
rect 5452 20012 5492 20140
rect 5644 20180 5684 20560
rect 5740 20348 5780 21148
rect 5740 20299 5780 20308
rect 5644 20131 5684 20140
rect 5836 20180 5876 22828
rect 5836 20131 5876 20140
rect 5452 19963 5492 19972
rect 5548 20012 5588 20021
rect 5356 19711 5396 19720
rect 5356 19424 5396 19433
rect 5356 15728 5396 19384
rect 5452 19424 5492 19433
rect 5452 19256 5492 19384
rect 5452 19207 5492 19216
rect 5452 18752 5492 18761
rect 5452 18617 5492 18712
rect 5548 18668 5588 19972
rect 5740 20012 5780 20021
rect 5740 19844 5780 19972
rect 5740 19760 5780 19804
rect 5740 19709 5780 19720
rect 5836 19928 5876 19937
rect 5644 19340 5684 19349
rect 5644 19205 5684 19300
rect 5740 19256 5780 19265
rect 5740 19004 5780 19216
rect 5740 18955 5780 18964
rect 5836 19172 5876 19888
rect 5548 18619 5588 18628
rect 5740 18668 5780 18677
rect 5644 18584 5684 18593
rect 5548 18500 5588 18509
rect 5452 18416 5492 18425
rect 5452 17828 5492 18376
rect 5452 17779 5492 17788
rect 5452 17660 5492 17669
rect 5452 17492 5492 17620
rect 5548 17576 5588 18460
rect 5548 17527 5588 17536
rect 5452 17072 5492 17452
rect 5548 17408 5588 17417
rect 5548 17273 5588 17368
rect 5644 17240 5684 18544
rect 5740 17576 5780 18628
rect 5740 17527 5780 17536
rect 5836 17828 5876 19132
rect 5836 17324 5876 17788
rect 5644 17191 5684 17200
rect 5740 17240 5780 17249
rect 5452 16988 5492 17032
rect 5452 16939 5492 16948
rect 5740 17072 5780 17200
rect 5836 17156 5876 17284
rect 5836 17107 5876 17116
rect 5548 16904 5588 16913
rect 5548 16316 5588 16864
rect 5740 16904 5780 17032
rect 5740 16855 5780 16864
rect 5836 16988 5876 16997
rect 5740 16736 5780 16745
rect 5548 16267 5588 16276
rect 5644 16484 5684 16493
rect 5356 15679 5396 15688
rect 5548 15728 5588 15737
rect 5452 15644 5492 15653
rect 5452 15392 5492 15604
rect 5548 15560 5588 15688
rect 5548 15511 5588 15520
rect 5452 15343 5492 15352
rect 5548 15308 5588 15317
rect 5452 14972 5492 14981
rect 5356 14132 5396 14141
rect 5356 13880 5396 14092
rect 5356 13831 5396 13840
rect 5452 13376 5492 14932
rect 5548 14720 5588 15268
rect 5548 14671 5588 14680
rect 5644 14132 5684 16444
rect 5740 15728 5780 16696
rect 5740 15679 5780 15688
rect 5836 16316 5876 16948
rect 5932 16736 5972 27448
rect 6316 27236 6356 27532
rect 6700 27488 6740 27616
rect 6700 27439 6740 27448
rect 6316 27187 6356 27196
rect 6412 27404 6452 27413
rect 6316 26900 6356 26909
rect 6124 26648 6164 26657
rect 6028 26228 6068 26237
rect 6028 26093 6068 26188
rect 6124 22364 6164 26608
rect 6220 26312 6260 26321
rect 6220 25892 6260 26272
rect 6220 25843 6260 25852
rect 6220 24548 6260 24557
rect 6220 23708 6260 24508
rect 6220 23540 6260 23668
rect 6220 23491 6260 23500
rect 6124 22315 6164 22324
rect 6220 23036 6260 23045
rect 6124 22196 6164 22205
rect 6028 22112 6068 22121
rect 6028 21860 6068 22072
rect 6028 21811 6068 21820
rect 6124 21776 6164 22156
rect 6124 21727 6164 21736
rect 6028 21692 6068 21701
rect 6028 21557 6068 21652
rect 6124 21608 6164 21648
rect 6124 21524 6164 21568
rect 6028 21440 6068 21449
rect 6028 21305 6068 21400
rect 6028 21104 6068 21113
rect 6028 20852 6068 21064
rect 6124 21020 6164 21484
rect 6124 20971 6164 20980
rect 6220 20852 6260 22996
rect 6316 21776 6356 26860
rect 6412 26228 6452 27364
rect 6412 26179 6452 26188
rect 6700 26564 6740 26573
rect 6604 26144 6644 26153
rect 6412 26060 6452 26069
rect 6412 25556 6452 26020
rect 6412 25507 6452 25516
rect 6604 25304 6644 26104
rect 6700 25640 6740 26524
rect 6796 26480 6836 26489
rect 6796 26144 6836 26440
rect 6892 26312 6932 27700
rect 6892 26263 6932 26272
rect 6796 26095 6836 26104
rect 6700 25591 6740 25600
rect 6796 25724 6836 25733
rect 6412 25136 6452 25145
rect 6412 23624 6452 25096
rect 6604 24632 6644 25264
rect 6796 24884 6836 25684
rect 6988 25556 7028 28600
rect 7756 27404 7796 28600
rect 7756 27355 7796 27364
rect 8044 27656 8084 27665
rect 7180 27320 7220 27329
rect 7180 26480 7220 27280
rect 7180 26431 7220 26440
rect 8044 26648 8084 27616
rect 8428 27572 8468 27581
rect 8332 27236 8372 27245
rect 7276 26396 7316 26405
rect 6604 24583 6644 24592
rect 6700 24844 6836 24884
rect 6892 25516 7028 25556
rect 7084 26228 7124 26237
rect 6700 23876 6740 24844
rect 6796 24716 6836 24725
rect 6796 24044 6836 24676
rect 6796 23995 6836 24004
rect 6700 23836 6836 23876
rect 6412 23489 6452 23584
rect 6604 23204 6644 23213
rect 6412 23120 6452 23129
rect 6412 22784 6452 23080
rect 6412 22735 6452 22744
rect 6508 22448 6548 22459
rect 6508 22364 6548 22408
rect 6508 22315 6548 22324
rect 6604 22280 6644 23164
rect 6412 22112 6452 22123
rect 6412 22028 6452 22072
rect 6604 22112 6644 22240
rect 6604 22063 6644 22072
rect 6700 22196 6740 22205
rect 6412 21979 6452 21988
rect 6604 21944 6644 21953
rect 6316 21727 6356 21736
rect 6412 21860 6452 21869
rect 6028 20812 6164 20852
rect 6028 19844 6068 19939
rect 6028 19795 6068 19804
rect 6028 19676 6068 19685
rect 6028 19541 6068 19636
rect 5932 16687 5972 16696
rect 6028 19256 6068 19265
rect 5836 15560 5876 16276
rect 5836 15511 5876 15520
rect 5932 16568 5972 16577
rect 5932 15728 5972 16528
rect 5932 15476 5972 15688
rect 5932 15427 5972 15436
rect 5644 13964 5684 14092
rect 5740 15308 5780 15317
rect 5740 14048 5780 15268
rect 5836 15140 5876 15149
rect 5836 14804 5876 15100
rect 5836 14132 5876 14764
rect 5932 14720 5972 14731
rect 5932 14636 5972 14680
rect 5932 14587 5972 14596
rect 5836 14083 5876 14092
rect 5932 14468 5972 14477
rect 5740 13999 5780 14008
rect 5644 13915 5684 13924
rect 5836 13964 5876 13973
rect 5836 13796 5876 13924
rect 5836 13747 5876 13756
rect 5836 13460 5876 13469
rect 5452 13336 5588 13376
rect 5548 13292 5588 13336
rect 5452 13208 5492 13217
rect 5452 13073 5492 13168
rect 5260 12940 5396 12980
rect 4972 12412 5108 12452
rect 5164 12536 5204 12545
rect 4972 11696 5012 12412
rect 4972 11561 5012 11656
rect 5164 11696 5204 12496
rect 5164 11647 5204 11656
rect 5068 11612 5108 11621
rect 5068 11024 5108 11572
rect 5260 11528 5300 11537
rect 5068 10975 5108 10984
rect 5164 11444 5204 11453
rect 5164 11024 5204 11404
rect 5260 11108 5300 11488
rect 5260 11059 5300 11068
rect 5164 10975 5204 10984
rect 5164 10604 5204 10613
rect 4876 10219 4916 10228
rect 5068 10352 5108 10361
rect 4972 10184 5012 10193
rect 4684 9967 4724 9976
rect 4780 10100 4820 10109
rect 4352 9848 4720 9857
rect 4352 9799 4720 9808
rect 4780 9680 4820 10060
rect 4780 9631 4820 9640
rect 4204 9379 4244 9388
rect 4876 9428 4916 9437
rect 4684 8840 4724 8849
rect 4108 7867 4148 7876
rect 4204 8672 4244 8681
rect 4204 8168 4244 8632
rect 4684 8672 4724 8800
rect 4684 8504 4724 8632
rect 4684 8455 4724 8464
rect 4780 8756 4820 8765
rect 4352 8336 4720 8345
rect 4352 8287 4720 8296
rect 4204 8000 4244 8128
rect 4780 8084 4820 8716
rect 4876 8588 4916 9388
rect 4972 8924 5012 10144
rect 4972 8875 5012 8884
rect 5068 9260 5108 10312
rect 5164 10184 5204 10564
rect 5164 9428 5204 10144
rect 5260 10268 5300 10277
rect 5260 9680 5300 10228
rect 5260 9631 5300 9640
rect 5356 9512 5396 12940
rect 5548 12620 5588 13252
rect 5836 13292 5876 13420
rect 5932 13460 5972 14428
rect 5932 13411 5972 13420
rect 5836 12704 5876 13252
rect 5932 13124 5972 13133
rect 5932 12788 5972 13084
rect 6028 13040 6068 19216
rect 6124 18080 6164 20812
rect 6220 20803 6260 20812
rect 6316 21608 6356 21617
rect 6220 20432 6260 20443
rect 6220 20348 6260 20392
rect 6220 20299 6260 20308
rect 6220 19508 6260 19517
rect 6220 18668 6260 19468
rect 6316 19256 6356 21568
rect 6412 21524 6452 21820
rect 6604 21776 6644 21904
rect 6604 21727 6644 21736
rect 6412 21475 6452 21484
rect 6508 21608 6548 21617
rect 6412 20936 6452 20945
rect 6412 20432 6452 20896
rect 6508 20936 6548 21568
rect 6700 21608 6740 22156
rect 6796 22196 6836 23836
rect 6892 23060 6932 25516
rect 6988 25388 7028 25397
rect 6988 25253 7028 25348
rect 7084 25136 7124 26188
rect 7180 26228 7220 26237
rect 7180 25304 7220 26188
rect 7276 25892 7316 26356
rect 7372 26312 7412 26321
rect 7372 26228 7412 26272
rect 7372 26177 7412 26188
rect 7276 25843 7316 25852
rect 7756 26144 7796 26153
rect 7180 25255 7220 25264
rect 7372 25304 7412 25313
rect 7372 25169 7412 25264
rect 7084 25087 7124 25096
rect 7756 24800 7796 26104
rect 7852 25136 7892 25145
rect 7852 25001 7892 25096
rect 7756 24751 7796 24760
rect 7084 23876 7124 23971
rect 7084 23827 7124 23836
rect 7468 23960 7508 23969
rect 6988 23708 7028 23717
rect 7028 23668 7412 23708
rect 6988 23659 7028 23668
rect 7180 23540 7220 23549
rect 6988 23372 7028 23383
rect 6988 23288 7028 23332
rect 6988 23239 7028 23248
rect 7084 23204 7124 23213
rect 6892 23020 7028 23060
rect 6796 22147 6836 22156
rect 6892 22532 6932 22541
rect 6740 21568 6836 21608
rect 6700 21559 6740 21568
rect 6508 20887 6548 20896
rect 6796 20936 6836 21568
rect 6892 21104 6932 22492
rect 6892 21055 6932 21064
rect 6796 20887 6836 20896
rect 6604 20852 6644 20861
rect 6412 20383 6452 20392
rect 6508 20684 6548 20693
rect 6412 20012 6452 20021
rect 6412 19877 6452 19972
rect 6508 19676 6548 20644
rect 6508 19340 6548 19636
rect 6508 19291 6548 19300
rect 6604 19928 6644 20812
rect 6988 20768 7028 23020
rect 7084 22532 7124 23164
rect 7180 23036 7220 23500
rect 7180 22987 7220 22996
rect 7276 23288 7316 23297
rect 7276 22952 7316 23248
rect 7372 23288 7412 23668
rect 7372 23239 7412 23248
rect 7468 23204 7508 23920
rect 7468 23155 7508 23164
rect 7660 23624 7700 23633
rect 7276 22903 7316 22912
rect 7564 23036 7604 23045
rect 7084 22483 7124 22492
rect 7276 22616 7316 22625
rect 7084 22280 7124 22289
rect 7084 21776 7124 22240
rect 7124 21736 7220 21776
rect 7084 21727 7124 21736
rect 7084 21356 7124 21365
rect 7084 20936 7124 21316
rect 7084 20887 7124 20896
rect 6892 20728 7028 20768
rect 7180 20768 7220 21736
rect 7276 20852 7316 22576
rect 7564 22280 7604 22996
rect 7372 22196 7412 22205
rect 7372 21356 7412 22156
rect 7564 22145 7604 22240
rect 7660 21776 7700 23584
rect 7948 23624 7988 23633
rect 7756 23204 7796 23213
rect 7756 22448 7796 23164
rect 7756 22364 7796 22408
rect 7756 22313 7796 22324
rect 7852 23036 7892 23045
rect 7564 21736 7700 21776
rect 7756 21776 7796 21785
rect 7372 21307 7412 21316
rect 7468 21524 7508 21533
rect 7276 20803 7316 20812
rect 7372 21020 7412 21029
rect 6604 19340 6644 19888
rect 6700 20096 6740 20105
rect 6700 19676 6740 20056
rect 6700 19627 6740 19636
rect 6604 19291 6644 19300
rect 6700 19424 6740 19433
rect 6316 19207 6356 19216
rect 6412 19256 6452 19265
rect 6412 19088 6452 19216
rect 6412 19048 6548 19088
rect 6508 19004 6548 19048
rect 6508 18955 6548 18964
rect 6412 18920 6452 18929
rect 6412 18785 6452 18880
rect 6604 18920 6644 18929
rect 6220 18619 6260 18628
rect 6316 18752 6356 18763
rect 6316 18668 6356 18712
rect 6316 18619 6356 18628
rect 6604 18584 6644 18880
rect 6604 18500 6644 18544
rect 6604 18449 6644 18460
rect 6412 18248 6452 18257
rect 6124 18031 6164 18040
rect 6220 18080 6260 18089
rect 6220 17744 6260 18040
rect 6220 17695 6260 17704
rect 6412 17660 6452 18208
rect 6700 18164 6740 19384
rect 6796 18920 6836 18929
rect 6796 18785 6836 18880
rect 6796 18500 6836 18509
rect 6796 18365 6836 18460
rect 6700 18124 6836 18164
rect 6700 17996 6740 18005
rect 6412 17492 6452 17620
rect 6412 17443 6452 17452
rect 6508 17912 6548 17952
rect 6508 17828 6548 17872
rect 6412 17240 6452 17249
rect 6220 17156 6260 17165
rect 6124 16988 6164 16997
rect 6124 16568 6164 16948
rect 6124 16519 6164 16528
rect 6124 16064 6164 16073
rect 6124 15644 6164 16024
rect 6220 15980 6260 17116
rect 6316 17072 6356 17081
rect 6316 16937 6356 17032
rect 6316 16484 6356 16493
rect 6316 16316 6356 16444
rect 6412 16400 6452 17200
rect 6412 16351 6452 16360
rect 6316 16267 6356 16276
rect 6220 15931 6260 15940
rect 6316 16148 6356 16157
rect 6124 15595 6164 15604
rect 6220 15560 6260 15569
rect 6124 14132 6164 14141
rect 6124 13997 6164 14092
rect 6220 13796 6260 15520
rect 6316 15560 6356 16108
rect 6316 15511 6356 15520
rect 6412 15644 6452 15653
rect 6412 15476 6452 15604
rect 6412 15427 6452 15436
rect 6220 13747 6260 13756
rect 6316 15392 6356 15401
rect 6316 13544 6356 15352
rect 6412 14804 6452 14899
rect 6412 14755 6452 14764
rect 6412 14636 6452 14645
rect 6412 13628 6452 14596
rect 6508 14216 6548 17788
rect 6604 17912 6644 17921
rect 6604 17576 6644 17872
rect 6700 17828 6740 17956
rect 6700 17779 6740 17788
rect 6604 17527 6644 17536
rect 6700 17492 6740 17501
rect 6700 17072 6740 17452
rect 6700 17023 6740 17032
rect 6796 16484 6836 18124
rect 6604 16444 6836 16484
rect 6604 16232 6644 16444
rect 6604 16183 6644 16192
rect 6700 16316 6740 16325
rect 6700 16064 6740 16276
rect 6604 16024 6740 16064
rect 6796 16316 6836 16325
rect 6796 16064 6836 16276
rect 6604 15308 6644 16024
rect 6796 16015 6836 16024
rect 6796 15560 6836 15569
rect 6604 15259 6644 15268
rect 6700 15308 6740 15317
rect 6700 14972 6740 15268
rect 6700 14923 6740 14932
rect 6796 14804 6836 15520
rect 6700 14720 6740 14729
rect 6604 14636 6644 14645
rect 6604 14501 6644 14596
rect 6508 14167 6548 14176
rect 6604 14048 6644 14057
rect 6412 13579 6452 13588
rect 6508 13880 6548 13889
rect 6316 13495 6356 13504
rect 6220 13460 6260 13469
rect 6028 12991 6068 13000
rect 6124 13376 6164 13385
rect 5932 12739 5972 12748
rect 5836 12655 5876 12664
rect 5548 12032 5588 12580
rect 5548 11983 5588 11992
rect 5644 12452 5684 12461
rect 5452 11696 5492 11705
rect 5452 11192 5492 11656
rect 5452 11143 5492 11152
rect 5548 11696 5588 11705
rect 5548 11024 5588 11656
rect 5548 10604 5588 10984
rect 5548 10555 5588 10564
rect 5548 10352 5588 10363
rect 5548 10268 5588 10312
rect 5548 10219 5588 10228
rect 5164 9379 5204 9388
rect 5260 9472 5396 9512
rect 5452 10016 5492 10025
rect 5068 8672 5108 9220
rect 5068 8623 5108 8632
rect 5164 8840 5204 8849
rect 4876 8539 4916 8548
rect 4012 6775 4052 6784
rect 4108 7748 4148 7757
rect 3916 6691 3956 6700
rect 3820 5767 3860 5776
rect 3532 5599 3572 5608
rect 4108 5564 4148 7708
rect 4204 6488 4244 7960
rect 4684 8000 4724 8011
rect 4684 7916 4724 7960
rect 4684 7867 4724 7876
rect 4780 7832 4820 8044
rect 4300 7328 4340 7337
rect 4300 7076 4340 7288
rect 4300 7027 4340 7036
rect 4352 6824 4720 6833
rect 4352 6775 4720 6784
rect 4204 5648 4244 6448
rect 4780 6740 4820 7792
rect 4684 6404 4724 6413
rect 4684 5816 4724 6364
rect 4684 5767 4724 5776
rect 4204 5599 4244 5608
rect 4780 5648 4820 6700
rect 4876 8420 4916 8429
rect 4876 7244 4916 8380
rect 5068 8336 5108 8345
rect 5068 8084 5108 8296
rect 5068 8035 5108 8044
rect 4876 5900 4916 7204
rect 5164 7160 5204 8800
rect 5260 7328 5300 9472
rect 5356 9344 5396 9353
rect 5356 8672 5396 9304
rect 5356 8623 5396 8632
rect 5452 8084 5492 9976
rect 5644 9932 5684 12412
rect 5932 12368 5972 12377
rect 5740 11696 5780 11705
rect 5740 11108 5780 11656
rect 5740 11059 5780 11068
rect 5836 10856 5876 10865
rect 5548 9344 5588 9353
rect 5548 8252 5588 9304
rect 5644 8840 5684 9892
rect 5644 8791 5684 8800
rect 5740 10352 5780 10361
rect 5740 8756 5780 10312
rect 5836 9764 5876 10816
rect 5836 9715 5876 9724
rect 5932 10184 5972 12328
rect 6124 11612 6164 13336
rect 6220 13292 6260 13420
rect 6220 13243 6260 13252
rect 6508 13292 6548 13840
rect 6604 13376 6644 14008
rect 6604 13327 6644 13336
rect 6508 13243 6548 13252
rect 6316 13208 6356 13217
rect 6220 13124 6260 13133
rect 6220 11780 6260 13084
rect 6316 13040 6356 13168
rect 6316 12991 6356 13000
rect 6412 12452 6452 12547
rect 6412 12403 6452 12412
rect 6508 12536 6548 12545
rect 6220 11731 6260 11740
rect 6316 12116 6356 12125
rect 6316 11696 6356 12076
rect 6316 11647 6356 11656
rect 6124 11563 6164 11572
rect 6028 11024 6068 11033
rect 6028 10772 6068 10984
rect 6028 10723 6068 10732
rect 5932 9764 5972 10144
rect 5932 9715 5972 9724
rect 6220 10184 6260 10193
rect 5836 9512 5876 9521
rect 5836 9377 5876 9472
rect 6220 9512 6260 10144
rect 6124 9428 6164 9437
rect 5740 8716 6068 8756
rect 5548 8203 5588 8212
rect 5644 8672 5684 8681
rect 5452 8035 5492 8044
rect 5356 8000 5396 8009
rect 5356 7412 5396 7960
rect 5356 7363 5396 7372
rect 5260 7279 5300 7288
rect 5644 7328 5684 8632
rect 5932 8588 5972 8597
rect 5644 7279 5684 7288
rect 5740 8168 5780 8177
rect 5740 7244 5780 8128
rect 5740 7195 5780 7204
rect 5932 7160 5972 8548
rect 5164 7111 5204 7120
rect 5836 7120 5972 7160
rect 6028 8000 6068 8716
rect 4876 5851 4916 5860
rect 5740 6992 5780 7001
rect 4780 5599 4820 5608
rect 5740 5648 5780 6952
rect 5836 6908 5876 7120
rect 6028 7076 6068 7960
rect 6028 7027 6068 7036
rect 5836 6859 5876 6868
rect 5932 6992 5972 7001
rect 5932 6152 5972 6952
rect 6124 6992 6164 9388
rect 6220 8840 6260 9472
rect 6220 7916 6260 8800
rect 6316 9848 6356 9857
rect 6316 9092 6356 9808
rect 6316 8672 6356 9052
rect 6316 8623 6356 8632
rect 6316 8084 6356 8093
rect 6316 8000 6356 8044
rect 6316 7949 6356 7960
rect 6220 7867 6260 7876
rect 6220 7748 6260 7757
rect 6220 7160 6260 7708
rect 6508 7244 6548 12496
rect 6604 12452 6644 12461
rect 6604 11696 6644 12412
rect 6604 11192 6644 11656
rect 6604 11143 6644 11152
rect 6700 10940 6740 14680
rect 6796 13208 6836 14764
rect 6796 12788 6836 13168
rect 6796 12739 6836 12748
rect 6796 12620 6836 12629
rect 6796 11948 6836 12580
rect 6796 11899 6836 11908
rect 6796 11780 6836 11789
rect 6796 11645 6836 11740
rect 6700 10268 6740 10900
rect 6700 10219 6740 10228
rect 6604 9764 6644 9773
rect 6604 8672 6644 9724
rect 6604 8623 6644 8632
rect 6796 9428 6836 9437
rect 6796 8588 6836 9388
rect 6796 8539 6836 8548
rect 6892 8252 6932 20728
rect 7180 20719 7220 20728
rect 6988 20600 7028 20609
rect 6988 19172 7028 20560
rect 7084 20432 7124 20441
rect 7084 20012 7124 20392
rect 7372 20180 7412 20980
rect 7468 20768 7508 21484
rect 7564 21020 7604 21736
rect 7756 21692 7796 21736
rect 7564 20971 7604 20980
rect 7660 21652 7796 21692
rect 7468 20719 7508 20728
rect 7564 20768 7604 20777
rect 7468 20600 7508 20609
rect 7468 20465 7508 20560
rect 7372 20131 7412 20140
rect 7564 20180 7604 20728
rect 7660 20264 7700 21652
rect 7852 21608 7892 22996
rect 7852 21559 7892 21568
rect 7756 21524 7796 21533
rect 7756 21020 7796 21484
rect 7756 20971 7796 20980
rect 7852 21188 7892 21197
rect 7852 20684 7892 21148
rect 7948 20852 7988 23584
rect 8044 23060 8084 26608
rect 8140 26732 8180 26741
rect 8140 26060 8180 26692
rect 8332 26648 8372 27196
rect 8332 26599 8372 26608
rect 8140 26011 8180 26020
rect 8236 26144 8276 26153
rect 8140 25052 8180 25061
rect 8140 24917 8180 25012
rect 8140 24800 8180 24809
rect 8140 23876 8180 24760
rect 8236 24548 8276 26104
rect 8428 25640 8468 27532
rect 8524 26396 8564 28600
rect 9196 28412 9236 28421
rect 8620 27908 8660 27917
rect 8620 27773 8660 27868
rect 8908 27488 8948 27497
rect 8908 26900 8948 27448
rect 9196 27404 9236 28372
rect 9292 27824 9332 28600
rect 10060 28244 10100 28600
rect 10060 28195 10100 28204
rect 9292 27775 9332 27784
rect 9388 27824 9428 27833
rect 8948 26860 9044 26900
rect 8908 26851 8948 26860
rect 8812 26816 8852 26825
rect 8524 26347 8564 26356
rect 8620 26564 8660 26573
rect 8524 26144 8564 26153
rect 8524 26009 8564 26104
rect 8236 24499 8276 24508
rect 8332 25600 8468 25640
rect 8524 25892 8564 25901
rect 8332 24464 8372 25600
rect 8332 24415 8372 24424
rect 8428 24548 8468 24557
rect 8140 23827 8180 23836
rect 8236 23960 8276 23969
rect 8236 23288 8276 23920
rect 8236 23239 8276 23248
rect 8332 23372 8372 23381
rect 8044 23020 8180 23060
rect 8044 22784 8084 22793
rect 8044 22196 8084 22744
rect 8044 22147 8084 22156
rect 8140 22028 8180 23020
rect 8236 22448 8276 22543
rect 8236 22399 8276 22408
rect 7948 20717 7988 20812
rect 8044 21988 8180 22028
rect 8236 22280 8276 22289
rect 7660 20215 7700 20224
rect 7756 20348 7796 20357
rect 7564 20131 7604 20140
rect 7084 19592 7124 19972
rect 7084 19508 7124 19552
rect 7084 19459 7124 19468
rect 7180 20096 7220 20105
rect 7084 19340 7124 19349
rect 7084 19205 7124 19300
rect 6988 19123 7028 19132
rect 7084 19088 7124 19097
rect 7084 18248 7124 19048
rect 7180 18920 7220 20056
rect 7468 20096 7508 20105
rect 7372 20012 7412 20021
rect 7372 19877 7412 19972
rect 7276 19844 7316 19853
rect 7276 19424 7316 19804
rect 7276 19375 7316 19384
rect 7180 18871 7220 18880
rect 7276 19256 7316 19296
rect 7276 19172 7316 19216
rect 7372 19172 7412 19181
rect 7276 19132 7372 19172
rect 7084 18199 7124 18208
rect 7180 18752 7220 18761
rect 6988 17744 7028 17753
rect 6988 17576 7028 17704
rect 6988 17527 7028 17536
rect 7084 16988 7124 16997
rect 7084 16484 7124 16948
rect 7084 16435 7124 16444
rect 7180 16316 7220 18712
rect 7276 18668 7316 19132
rect 7372 19123 7412 19132
rect 7276 17912 7316 18628
rect 7372 18752 7412 18761
rect 7372 18080 7412 18712
rect 7372 18031 7412 18040
rect 7276 17863 7316 17872
rect 7372 17912 7412 17921
rect 7276 17744 7316 17753
rect 7276 16904 7316 17704
rect 7372 17744 7412 17872
rect 7372 17695 7412 17704
rect 7372 17408 7412 17417
rect 7372 17156 7412 17368
rect 7372 17107 7412 17116
rect 7276 16736 7316 16864
rect 7276 16696 7412 16736
rect 7276 16568 7316 16577
rect 7276 16400 7316 16528
rect 7372 16484 7412 16696
rect 7372 16435 7412 16444
rect 7276 16351 7316 16360
rect 7180 16267 7220 16276
rect 6988 16148 7028 16243
rect 6988 16099 7028 16108
rect 6988 15980 7028 15989
rect 6988 14636 7028 15940
rect 7372 15644 7412 15653
rect 7084 15560 7124 15569
rect 7084 14972 7124 15520
rect 7084 14923 7124 14932
rect 7180 15560 7220 15569
rect 7180 14888 7220 15520
rect 7180 14839 7220 14848
rect 7276 15392 7316 15401
rect 6988 14587 7028 14596
rect 7180 13964 7220 13973
rect 7084 13124 7124 13133
rect 7084 12704 7124 13084
rect 7180 12956 7220 13924
rect 7276 13376 7316 15352
rect 7372 15308 7412 15604
rect 7372 15259 7412 15268
rect 7468 14300 7508 20056
rect 7756 19424 7796 20308
rect 7852 19760 7892 20644
rect 8044 20096 8084 21988
rect 8140 21860 8180 21869
rect 8140 21188 8180 21820
rect 8236 21692 8276 22240
rect 8236 21643 8276 21652
rect 8140 21139 8180 21148
rect 8236 21524 8276 21533
rect 8236 21188 8276 21484
rect 8236 21139 8276 21148
rect 8332 21020 8372 23332
rect 8236 20980 8372 21020
rect 8140 20852 8180 20861
rect 8140 20717 8180 20812
rect 8140 20516 8180 20525
rect 8140 20432 8180 20476
rect 8140 20381 8180 20392
rect 8044 20056 8180 20096
rect 7852 19711 7892 19720
rect 7948 20012 7988 20021
rect 7948 19508 7988 19972
rect 8044 19928 8084 19937
rect 8044 19844 8084 19888
rect 8044 19793 8084 19804
rect 7948 19459 7988 19468
rect 7756 19375 7796 19384
rect 8044 19424 8084 19433
rect 7948 19172 7988 19181
rect 7564 19088 7604 19097
rect 7564 18500 7604 19048
rect 7756 19088 7796 19097
rect 7660 18920 7700 18929
rect 7660 18668 7700 18880
rect 7660 18584 7700 18628
rect 7660 18535 7700 18544
rect 7564 18451 7604 18460
rect 7660 18416 7700 18425
rect 7564 18332 7604 18341
rect 7564 17912 7604 18292
rect 7564 17863 7604 17872
rect 7660 18248 7700 18376
rect 7564 17744 7604 17755
rect 7564 17660 7604 17704
rect 7564 17611 7604 17620
rect 7660 17156 7700 18208
rect 7756 17828 7796 19048
rect 7852 18920 7892 18929
rect 7852 18584 7892 18880
rect 7948 18752 7988 19132
rect 8044 18836 8084 19384
rect 8140 18920 8180 20056
rect 8140 18871 8180 18880
rect 8044 18787 8084 18796
rect 7948 18703 7988 18712
rect 8044 18584 8084 18593
rect 7852 18544 7988 18584
rect 7948 18416 7988 18544
rect 7948 18367 7988 18376
rect 8044 18248 8084 18544
rect 8044 18199 8084 18208
rect 8140 18500 8180 18509
rect 8140 18164 8180 18460
rect 8140 18115 8180 18124
rect 7756 17779 7796 17788
rect 8140 17996 8180 18005
rect 7948 17744 7988 17753
rect 7948 17240 7988 17704
rect 7948 17191 7988 17200
rect 8044 17660 8084 17669
rect 7660 17107 7700 17116
rect 7852 17072 7892 17081
rect 7660 16400 7700 16409
rect 7564 16148 7604 16159
rect 7564 16064 7604 16108
rect 7564 16015 7604 16024
rect 7660 15812 7700 16360
rect 7660 15763 7700 15772
rect 7756 16148 7796 16157
rect 7756 15728 7796 16108
rect 7852 15896 7892 17032
rect 7852 15847 7892 15856
rect 7948 16988 7988 16997
rect 7948 16148 7988 16948
rect 7756 15679 7796 15688
rect 7660 15644 7700 15653
rect 7660 15509 7700 15604
rect 7852 15392 7892 15401
rect 7660 14804 7700 14813
rect 7468 14251 7508 14260
rect 7564 14636 7604 14645
rect 7468 13880 7508 13975
rect 7468 13831 7508 13840
rect 7276 13327 7316 13336
rect 7468 13712 7508 13721
rect 7372 13292 7412 13301
rect 7180 12907 7220 12916
rect 7276 13208 7316 13217
rect 7084 12655 7124 12664
rect 6988 12620 7028 12629
rect 6988 11948 7028 12580
rect 7180 12620 7220 12629
rect 7180 12485 7220 12580
rect 7084 12452 7124 12461
rect 7084 12317 7124 12412
rect 7276 12368 7316 13168
rect 7276 12319 7316 12328
rect 6988 11899 7028 11908
rect 7084 11696 7124 11705
rect 6988 11024 7028 11033
rect 6988 10268 7028 10984
rect 6988 10219 7028 10228
rect 7084 9512 7124 11656
rect 7372 11192 7412 13252
rect 7468 13040 7508 13672
rect 7468 12991 7508 13000
rect 7564 12788 7604 14596
rect 7564 12739 7604 12748
rect 7468 12536 7508 12545
rect 7468 11948 7508 12496
rect 7468 11899 7508 11908
rect 7372 10184 7412 11152
rect 7468 11780 7508 11789
rect 7468 11024 7508 11740
rect 7468 10975 7508 10984
rect 7372 10135 7412 10144
rect 7564 10058 7604 10067
rect 7564 10016 7604 10018
rect 7564 9923 7604 9976
rect 7660 9680 7700 14764
rect 7756 14048 7796 14057
rect 7756 13880 7796 14008
rect 7756 13831 7796 13840
rect 7852 13208 7892 15352
rect 7948 13292 7988 16108
rect 8044 15728 8084 17620
rect 8044 15679 8084 15688
rect 7948 13243 7988 13252
rect 8044 14048 8084 14057
rect 7852 13159 7892 13168
rect 8044 13124 8084 14008
rect 8044 12788 8084 13084
rect 8044 12739 8084 12748
rect 8044 12620 8084 12629
rect 7852 12284 7892 12293
rect 7756 11696 7796 11705
rect 7756 10016 7796 11656
rect 7852 11108 7892 12244
rect 8044 12284 8084 12580
rect 8140 12452 8180 17956
rect 8236 17072 8276 20980
rect 8332 20684 8372 20693
rect 8332 20096 8372 20644
rect 8332 19508 8372 20056
rect 8332 19459 8372 19468
rect 8332 19256 8372 19265
rect 8332 19004 8372 19216
rect 8332 18955 8372 18964
rect 8428 18752 8468 24508
rect 8524 20096 8564 25852
rect 8620 24800 8660 26524
rect 8716 26480 8756 26489
rect 8716 24884 8756 26440
rect 8812 26144 8852 26776
rect 8812 25808 8852 26104
rect 8812 25759 8852 25768
rect 8908 25304 8948 25315
rect 8908 25220 8948 25264
rect 8908 25171 8948 25180
rect 8716 24835 8756 24844
rect 8908 25052 8948 25061
rect 8620 24751 8660 24760
rect 8812 24716 8852 24725
rect 8812 24581 8852 24676
rect 8908 24632 8948 25012
rect 8908 24583 8948 24592
rect 9004 24212 9044 26860
rect 9196 26816 9236 27364
rect 9196 26767 9236 26776
rect 9100 26732 9140 26741
rect 9100 25304 9140 26692
rect 9292 26480 9332 26489
rect 9292 26144 9332 26440
rect 9292 26095 9332 26104
rect 9196 25892 9236 25901
rect 9196 25757 9236 25852
rect 9100 25169 9140 25264
rect 9100 24968 9140 25063
rect 9100 24919 9140 24928
rect 9292 24884 9332 24893
rect 9100 24800 9140 24809
rect 9100 24665 9140 24760
rect 9292 24716 9332 24844
rect 9292 24667 9332 24676
rect 8620 23792 8660 23801
rect 8620 23540 8660 23752
rect 8620 21524 8660 23500
rect 8812 23792 8852 23801
rect 8716 23120 8756 23129
rect 8716 22448 8756 23080
rect 8812 22868 8852 23752
rect 8908 23792 8948 23803
rect 8908 23708 8948 23752
rect 8908 23659 8948 23668
rect 9004 23624 9044 24172
rect 9196 24380 9236 24389
rect 9196 23792 9236 24340
rect 9196 23743 9236 23752
rect 9004 23575 9044 23584
rect 9100 23708 9140 23717
rect 8908 23372 8948 23381
rect 8908 23120 8948 23332
rect 8908 23071 8948 23080
rect 9004 23372 9044 23381
rect 8812 22828 8948 22868
rect 8812 22700 8852 22709
rect 8812 22616 8852 22660
rect 8812 22565 8852 22576
rect 8716 22408 8852 22448
rect 8812 22112 8852 22408
rect 8908 22280 8948 22828
rect 8908 22231 8948 22240
rect 8812 22072 8948 22112
rect 8812 21944 8852 21953
rect 8620 20432 8660 21484
rect 8716 21776 8756 21785
rect 8716 20516 8756 21736
rect 8812 21692 8852 21904
rect 8812 21643 8852 21652
rect 8908 21608 8948 22072
rect 8908 21559 8948 21568
rect 8812 21440 8852 21451
rect 8812 21356 8852 21400
rect 9004 21440 9044 23332
rect 9100 23036 9140 23668
rect 9100 22987 9140 22996
rect 9196 23624 9236 23633
rect 9100 22616 9140 22625
rect 9100 22364 9140 22576
rect 9100 22315 9140 22324
rect 9196 22280 9236 23584
rect 9388 23456 9428 27784
rect 10732 27824 10772 27833
rect 9772 27740 9812 27749
rect 9676 27656 9716 27665
rect 9484 27572 9524 27581
rect 9484 27236 9524 27532
rect 9524 27196 9620 27236
rect 9484 27187 9524 27196
rect 9388 23120 9428 23416
rect 9388 23071 9428 23080
rect 9484 26480 9524 26489
rect 9292 22784 9332 22793
rect 9292 22364 9332 22744
rect 9292 22315 9332 22324
rect 9196 22231 9236 22240
rect 9004 21391 9044 21400
rect 9292 22028 9332 22037
rect 8812 21307 8852 21316
rect 9004 21188 9044 21197
rect 9004 20684 9044 21148
rect 9100 21104 9140 21113
rect 9100 20969 9140 21064
rect 9196 21020 9236 21029
rect 8716 20467 8756 20476
rect 8812 20600 8852 20609
rect 8812 20465 8852 20560
rect 8620 20383 8660 20392
rect 8908 20264 8948 20273
rect 8716 20096 8756 20105
rect 8524 20056 8716 20096
rect 8524 19424 8564 20056
rect 8716 20047 8756 20056
rect 8812 19844 8852 19853
rect 8524 19375 8564 19384
rect 8716 19676 8756 19685
rect 8620 19256 8660 19267
rect 8620 19172 8660 19216
rect 8620 19123 8660 19132
rect 8332 18712 8468 18752
rect 8524 19004 8564 19013
rect 8332 17996 8372 18712
rect 8524 18668 8564 18964
rect 8524 18619 8564 18628
rect 8332 17947 8372 17956
rect 8428 18584 8468 18593
rect 8236 16400 8276 17032
rect 8332 17156 8372 17165
rect 8332 16652 8372 17116
rect 8428 16904 8468 18544
rect 8620 18500 8660 18509
rect 8620 18365 8660 18460
rect 8524 18332 8564 18341
rect 8524 17744 8564 18292
rect 8716 17912 8756 19636
rect 8812 18164 8852 19804
rect 8908 19760 8948 20224
rect 9004 20264 9044 20644
rect 9004 20215 9044 20224
rect 9100 20600 9140 20609
rect 8908 19340 8948 19720
rect 9004 20096 9044 20105
rect 9004 19592 9044 20056
rect 9004 19543 9044 19552
rect 8908 19291 8948 19300
rect 9004 19256 9044 19265
rect 8908 19004 8948 19013
rect 8908 18248 8948 18964
rect 8908 18199 8948 18208
rect 8812 18115 8852 18124
rect 8716 17863 8756 17872
rect 8524 17695 8564 17704
rect 8620 17744 8660 17753
rect 8524 17576 8564 17585
rect 8524 17324 8564 17536
rect 8524 17275 8564 17284
rect 8524 17072 8564 17081
rect 8524 16988 8564 17032
rect 8524 16937 8564 16948
rect 8428 16855 8468 16864
rect 8332 16484 8372 16612
rect 8524 16568 8564 16577
rect 8332 16444 8468 16484
rect 8276 16360 8372 16400
rect 8236 16351 8276 16360
rect 8236 16232 8276 16241
rect 8236 16148 8276 16192
rect 8236 16097 8276 16108
rect 8332 15644 8372 16360
rect 8332 15595 8372 15604
rect 8428 15728 8468 16444
rect 8524 16433 8564 16528
rect 8524 16316 8564 16325
rect 8524 15812 8564 16276
rect 8524 15763 8564 15772
rect 8428 15476 8468 15688
rect 8620 15728 8660 17704
rect 8908 17744 8948 17753
rect 8908 17660 8948 17704
rect 8908 17609 8948 17620
rect 8908 17492 8948 17501
rect 8908 17324 8948 17452
rect 8812 16988 8852 16997
rect 8524 15644 8564 15653
rect 8524 15509 8564 15604
rect 8428 15427 8468 15436
rect 8524 15224 8564 15233
rect 8524 14888 8564 15184
rect 8524 14839 8564 14848
rect 8620 14720 8660 15688
rect 8620 14671 8660 14680
rect 8716 16948 8812 16988
rect 8716 15644 8756 16948
rect 8812 16939 8852 16948
rect 8812 16820 8852 16829
rect 8812 16232 8852 16780
rect 8812 15896 8852 16192
rect 8812 15847 8852 15856
rect 8140 12403 8180 12412
rect 8236 14552 8276 14561
rect 8044 12235 8084 12244
rect 8044 11696 8084 11705
rect 8044 11561 8084 11656
rect 7852 11059 7892 11068
rect 7948 10520 7988 10529
rect 7756 9932 7796 9976
rect 7756 9852 7796 9892
rect 7852 10268 7892 10277
rect 7660 9631 7700 9640
rect 7084 9463 7124 9472
rect 7564 9512 7604 9521
rect 7276 9344 7316 9353
rect 7084 9260 7124 9269
rect 7084 8672 7124 9220
rect 7276 8756 7316 9304
rect 7276 8707 7316 8716
rect 7372 9008 7412 9017
rect 7084 8623 7124 8632
rect 7372 8672 7412 8968
rect 7372 8623 7412 8632
rect 7564 8588 7604 9472
rect 7852 9512 7892 10228
rect 7852 9463 7892 9472
rect 7948 10184 7988 10480
rect 7564 8539 7604 8548
rect 6892 8203 6932 8212
rect 7564 8168 7604 8177
rect 6508 7195 6548 7204
rect 7180 7496 7220 7505
rect 6220 7111 6260 7120
rect 6604 7160 6644 7169
rect 6124 6943 6164 6952
rect 6604 6656 6644 7120
rect 7180 7076 7220 7456
rect 7564 7244 7604 8128
rect 7948 8000 7988 10144
rect 8044 9260 8084 9269
rect 8044 8672 8084 9220
rect 8140 8924 8180 8933
rect 8140 8789 8180 8884
rect 8044 8623 8084 8632
rect 7564 7195 7604 7204
rect 7660 7748 7700 7757
rect 7660 7160 7700 7708
rect 7660 7111 7700 7120
rect 7180 7027 7220 7036
rect 6604 6607 6644 6616
rect 6796 6992 6836 7001
rect 6796 6488 6836 6952
rect 6796 6439 6836 6448
rect 6892 6572 6932 6581
rect 7852 6572 7892 6581
rect 5932 6103 5972 6112
rect 6028 6236 6068 6245
rect 4108 5228 4148 5524
rect 5452 5564 5492 5573
rect 4352 5312 4720 5321
rect 4352 5263 4720 5272
rect 4108 5179 4148 5188
rect 5452 5228 5492 5524
rect 5740 5396 5780 5608
rect 6028 5648 6068 6196
rect 6028 5599 6068 5608
rect 6220 5816 6260 5825
rect 5740 5347 5780 5356
rect 5452 5179 5492 5188
rect 6220 4976 6260 5776
rect 6892 5648 6932 6532
rect 7756 6532 7852 6572
rect 6892 5599 6932 5608
rect 7372 6488 7412 6497
rect 6508 5564 6548 5573
rect 6508 5144 6548 5524
rect 6508 5095 6548 5104
rect 7372 5396 7412 6448
rect 7756 6320 7796 6532
rect 7852 6523 7892 6532
rect 7756 6271 7796 6280
rect 7948 5900 7988 7960
rect 8140 8504 8180 8513
rect 8140 8000 8180 8464
rect 8140 7951 8180 7960
rect 7948 5851 7988 5860
rect 7372 5144 7412 5356
rect 7372 5095 7412 5104
rect 7564 5732 7604 5741
rect 6220 4927 6260 4936
rect 7564 4808 7604 5692
rect 8236 5648 8276 14512
rect 8620 14552 8660 14561
rect 8332 14048 8372 14057
rect 8332 13913 8372 14008
rect 8524 13796 8564 13805
rect 8524 13661 8564 13756
rect 8620 13544 8660 14512
rect 8716 13964 8756 15604
rect 8812 15308 8852 15317
rect 8812 14132 8852 15268
rect 8908 15224 8948 17284
rect 9004 16904 9044 19216
rect 9100 19256 9140 20560
rect 9100 19207 9140 19216
rect 9100 19004 9140 19013
rect 9100 18869 9140 18964
rect 9196 18752 9236 20980
rect 9292 19088 9332 21988
rect 9388 20852 9428 20861
rect 9388 20717 9428 20812
rect 9388 20516 9428 20525
rect 9388 19256 9428 20476
rect 9388 19207 9428 19216
rect 9484 19424 9524 26440
rect 9580 25640 9620 27196
rect 9676 27068 9716 27616
rect 9676 27019 9716 27028
rect 9676 26816 9716 26825
rect 9676 26480 9716 26776
rect 9676 26431 9716 26440
rect 9772 26144 9812 27700
rect 10540 27740 10580 27749
rect 10060 27236 10100 27245
rect 9868 27152 9908 27161
rect 9868 26816 9908 27112
rect 10060 26900 10100 27196
rect 10348 27068 10388 27077
rect 10060 26851 10100 26860
rect 10156 26984 10196 26993
rect 9868 26767 9908 26776
rect 9772 26095 9812 26104
rect 9964 26480 10004 26489
rect 9580 25388 9620 25600
rect 9580 25339 9620 25348
rect 9580 25220 9620 25229
rect 9580 24464 9620 25180
rect 9676 25220 9716 25231
rect 9676 25136 9716 25180
rect 9676 25087 9716 25096
rect 9964 25136 10004 26440
rect 9580 24415 9620 24424
rect 9964 24044 10004 25096
rect 9964 23995 10004 24004
rect 10060 24128 10100 24137
rect 10060 23993 10100 24088
rect 9964 23792 10004 23801
rect 9868 23752 9964 23792
rect 9868 23120 9908 23752
rect 9964 23743 10004 23752
rect 10156 23540 10196 26944
rect 10252 26816 10292 26825
rect 10252 23792 10292 26776
rect 10348 24548 10388 27028
rect 10540 26144 10580 27700
rect 10636 27563 10676 27572
rect 10636 27068 10676 27523
rect 10636 27019 10676 27028
rect 10540 26095 10580 26104
rect 10732 25052 10772 27784
rect 10828 27404 10868 28600
rect 10828 27355 10868 27364
rect 11308 27992 11348 28001
rect 10886 27236 11254 27245
rect 10886 27187 11254 27196
rect 11116 26564 11156 26573
rect 11116 26144 11156 26524
rect 11308 26228 11348 27952
rect 11116 26095 11156 26104
rect 11212 26144 11252 26153
rect 11212 25976 11252 26104
rect 11212 25927 11252 25936
rect 10886 25724 11254 25733
rect 10886 25675 11254 25684
rect 11116 25556 11156 25565
rect 11116 25388 11156 25516
rect 11116 25339 11156 25348
rect 11212 25304 11252 25313
rect 10828 25220 10868 25231
rect 10828 25136 10868 25180
rect 10828 25087 10868 25096
rect 10732 25003 10772 25012
rect 10348 24499 10388 24508
rect 10732 24884 10772 24893
rect 10636 24296 10676 24305
rect 10636 24212 10676 24256
rect 10636 24161 10676 24172
rect 10252 23743 10292 23752
rect 10348 24128 10388 24137
rect 10348 23708 10388 24088
rect 10348 23659 10388 23668
rect 10636 23624 10676 23633
rect 10156 23500 10388 23540
rect 9868 23036 9908 23080
rect 9868 22987 9908 22996
rect 10252 23288 10292 23297
rect 9772 22448 9812 22457
rect 9676 22112 9716 22121
rect 9676 21944 9716 22072
rect 9580 21776 9620 21871
rect 9580 21727 9620 21736
rect 9676 21692 9716 21904
rect 9676 21643 9716 21652
rect 9580 21583 9620 21592
rect 9580 21104 9620 21543
rect 9580 21055 9620 21064
rect 9676 20768 9716 20777
rect 9676 20684 9716 20728
rect 9676 20633 9716 20644
rect 9772 20600 9812 22408
rect 10252 22448 10292 23248
rect 10348 23036 10388 23500
rect 10348 22987 10388 22996
rect 10252 22399 10292 22408
rect 10060 22364 10100 22373
rect 9868 22280 9908 22289
rect 9868 20852 9908 22240
rect 10060 22229 10100 22324
rect 10252 22112 10292 22121
rect 10060 21860 10100 21869
rect 10060 21725 10100 21820
rect 10252 21692 10292 22072
rect 9964 21440 10004 21449
rect 9964 21188 10004 21400
rect 9964 21139 10004 21148
rect 10060 21104 10100 21113
rect 10060 21020 10100 21064
rect 9868 20803 9908 20812
rect 9964 20980 10100 21020
rect 9964 20852 10004 20980
rect 9964 20803 10004 20812
rect 9676 20516 9716 20525
rect 9292 19048 9428 19088
rect 9196 18703 9236 18712
rect 9292 18920 9332 18929
rect 9004 16855 9044 16864
rect 9100 18584 9140 18593
rect 9100 18332 9140 18544
rect 9196 18416 9236 18511
rect 9292 18500 9332 18880
rect 9388 18920 9428 19048
rect 9388 18871 9428 18880
rect 9484 18584 9524 19384
rect 9580 20264 9620 20273
rect 9580 19844 9620 20224
rect 9676 20180 9716 20476
rect 9676 20131 9716 20140
rect 9580 19424 9620 19804
rect 9772 19508 9812 20560
rect 10252 20516 10292 21652
rect 10540 21608 10580 21617
rect 9772 19459 9812 19468
rect 9868 20348 9908 20357
rect 9580 19340 9620 19384
rect 9580 19289 9620 19300
rect 9772 19256 9812 19351
rect 9772 19207 9812 19216
rect 9676 19172 9716 19181
rect 9676 18752 9716 19132
rect 9676 18703 9716 18712
rect 9772 19088 9812 19097
rect 9388 18500 9428 18509
rect 9292 18460 9388 18500
rect 9196 18367 9236 18376
rect 9100 17072 9140 18292
rect 9292 18332 9332 18341
rect 8908 15175 8948 15184
rect 9004 16400 9044 16409
rect 9004 16148 9044 16360
rect 9004 14804 9044 16108
rect 9100 16148 9140 17032
rect 9196 18164 9236 18173
rect 9292 18164 9332 18292
rect 9236 18124 9332 18164
rect 9196 17744 9236 18124
rect 9196 17576 9236 17704
rect 9196 16820 9236 17536
rect 9196 16771 9236 16780
rect 9292 17156 9332 17165
rect 9292 16988 9332 17116
rect 9100 16099 9140 16108
rect 9100 15728 9140 15737
rect 9100 15560 9140 15688
rect 9100 14888 9140 15520
rect 9196 14888 9236 14897
rect 9100 14848 9196 14888
rect 9196 14839 9236 14848
rect 9004 14755 9044 14764
rect 9292 14804 9332 16948
rect 9388 15644 9428 18460
rect 9484 17744 9524 18544
rect 9484 17695 9524 17704
rect 9580 18332 9620 18341
rect 9484 17072 9524 17081
rect 9484 16820 9524 17032
rect 9484 16771 9524 16780
rect 9484 16064 9524 16073
rect 9484 15812 9524 16024
rect 9484 15763 9524 15772
rect 9388 15595 9428 15604
rect 9484 15644 9524 15653
rect 9484 15224 9524 15604
rect 9484 15175 9524 15184
rect 9388 15140 9428 15149
rect 9388 15005 9428 15100
rect 9484 15056 9524 15065
rect 9484 14921 9524 15016
rect 8908 14720 8948 14729
rect 8908 14636 8948 14680
rect 8908 14585 8948 14596
rect 9100 14552 9140 14561
rect 9100 14384 9140 14512
rect 9100 14335 9140 14344
rect 8812 14083 8852 14092
rect 9292 14048 9332 14764
rect 9484 14804 9524 14813
rect 9388 14216 9428 14225
rect 9388 14081 9428 14176
rect 9292 13999 9332 14008
rect 8716 13924 8852 13964
rect 8620 13495 8660 13504
rect 8524 13292 8564 13301
rect 8332 12620 8372 12629
rect 8332 12485 8372 12580
rect 8428 11780 8468 11789
rect 8428 11276 8468 11740
rect 8332 9932 8372 9941
rect 8332 9680 8372 9892
rect 8332 6740 8372 9640
rect 8428 9512 8468 11236
rect 8524 11192 8564 13252
rect 8716 12620 8756 12629
rect 8716 12485 8756 12580
rect 8620 12452 8660 12461
rect 8620 12317 8660 12412
rect 8524 11143 8564 11152
rect 8716 11108 8756 11117
rect 8620 11024 8660 11033
rect 8524 10016 8564 10025
rect 8524 9881 8564 9976
rect 8428 8756 8468 9472
rect 8428 8707 8468 8716
rect 8524 9764 8564 9773
rect 8524 8672 8564 9724
rect 8620 9680 8660 10984
rect 8716 10436 8756 11068
rect 8716 9680 8756 10396
rect 8812 9848 8852 13924
rect 9100 13712 9140 13721
rect 8908 13292 8948 13301
rect 8908 13208 8948 13252
rect 8908 13157 8948 13168
rect 9100 12704 9140 13672
rect 9100 12655 9140 12664
rect 9004 12620 9044 12629
rect 9004 12485 9044 12580
rect 9100 12536 9140 12545
rect 9004 11696 9044 11791
rect 9100 11696 9140 12496
rect 9044 11656 9140 11696
rect 9196 12284 9236 12293
rect 9004 11647 9044 11656
rect 9004 11528 9044 11537
rect 9004 11024 9044 11488
rect 9196 11108 9236 12244
rect 9196 11059 9236 11068
rect 9004 10975 9044 10984
rect 9196 10940 9236 10949
rect 9100 10688 9140 10697
rect 9100 10184 9140 10648
rect 9100 10135 9140 10144
rect 9196 10436 9236 10900
rect 8812 9799 8852 9808
rect 8716 9640 9044 9680
rect 8620 9631 8660 9640
rect 9004 9596 9044 9640
rect 9004 9547 9044 9556
rect 8812 9428 8852 9437
rect 8428 8420 8468 8429
rect 8428 8000 8468 8380
rect 8428 7951 8468 7960
rect 8332 6691 8372 6700
rect 8524 6404 8564 8632
rect 8716 8840 8756 8849
rect 8716 7076 8756 8800
rect 8812 8756 8852 9388
rect 9196 9428 9236 10396
rect 9196 9379 9236 9388
rect 9388 9764 9428 9773
rect 9388 9512 9428 9724
rect 9100 9344 9140 9353
rect 9100 8924 9140 9304
rect 9292 9176 9332 9185
rect 9100 8884 9236 8924
rect 9100 8756 9140 8765
rect 8812 8716 9100 8756
rect 9100 8707 9140 8716
rect 9196 8504 9236 8884
rect 9196 8455 9236 8464
rect 9292 8672 9332 9136
rect 9388 8840 9428 9472
rect 9388 8791 9428 8800
rect 8812 7916 8852 7925
rect 8812 7412 8852 7876
rect 8812 7363 8852 7372
rect 8908 7664 8948 7673
rect 8716 7027 8756 7036
rect 8524 6152 8564 6364
rect 8524 6103 8564 6112
rect 8236 5599 8276 5608
rect 8908 4892 8948 7624
rect 9292 7412 9332 8632
rect 9484 8168 9524 14764
rect 9580 14636 9620 18292
rect 9676 17996 9716 18005
rect 9676 17660 9716 17956
rect 9676 17072 9716 17620
rect 9772 17492 9812 19048
rect 9868 17744 9908 20308
rect 9964 20180 10004 20189
rect 9964 19592 10004 20140
rect 10060 19928 10100 19937
rect 10060 19760 10100 19888
rect 10060 19711 10100 19720
rect 9964 19543 10004 19552
rect 10156 19508 10196 19517
rect 10060 19088 10100 19097
rect 9868 17695 9908 17704
rect 9964 18668 10004 18677
rect 9772 17408 9812 17452
rect 9868 17576 9908 17585
rect 9868 17441 9908 17536
rect 9772 17359 9812 17368
rect 9772 17240 9812 17249
rect 9772 17105 9812 17200
rect 9676 16988 9716 17032
rect 9676 16736 9716 16948
rect 9964 16988 10004 18628
rect 9964 16939 10004 16948
rect 9676 16687 9716 16696
rect 9868 16820 9908 16829
rect 9868 16685 9908 16780
rect 9676 16148 9716 16157
rect 9676 15476 9716 16108
rect 9964 16148 10004 16157
rect 9772 15644 9812 15653
rect 9964 15644 10004 16108
rect 9812 15604 9908 15644
rect 9772 15595 9812 15604
rect 9676 15427 9716 15436
rect 9580 14587 9620 14596
rect 9676 14720 9716 14729
rect 9580 14132 9620 14227
rect 9676 14216 9716 14680
rect 9676 14167 9716 14176
rect 9772 14636 9812 14645
rect 9580 14083 9620 14092
rect 9580 13964 9620 13973
rect 9580 13829 9620 13924
rect 9772 13964 9812 14596
rect 9772 13915 9812 13924
rect 9772 13796 9812 13805
rect 9772 13208 9812 13756
rect 9868 13712 9908 15604
rect 9964 15595 10004 15604
rect 9868 13663 9908 13672
rect 9964 15476 10004 15485
rect 9772 13073 9812 13168
rect 9868 13292 9908 13301
rect 9676 12788 9716 12797
rect 9580 12536 9620 12545
rect 9580 11948 9620 12496
rect 9676 12284 9716 12748
rect 9868 12704 9908 13252
rect 9868 12655 9908 12664
rect 9676 12235 9716 12244
rect 9580 11192 9620 11908
rect 9580 11143 9620 11152
rect 9772 11276 9812 11285
rect 9772 10940 9812 11236
rect 9964 10940 10004 15436
rect 10060 14804 10100 19048
rect 10156 18500 10196 19468
rect 10252 18920 10292 20476
rect 10348 20936 10388 20945
rect 10348 20096 10388 20896
rect 10540 20684 10580 21568
rect 10540 20635 10580 20644
rect 10636 20600 10676 23584
rect 10732 23372 10772 24844
rect 11212 24884 11252 25264
rect 11212 24632 11252 24844
rect 11212 24583 11252 24592
rect 11308 25136 11348 26188
rect 11500 27656 11540 27665
rect 11404 26144 11444 26155
rect 11404 26060 11444 26104
rect 11404 26011 11444 26020
rect 11404 25892 11444 25901
rect 11404 25556 11444 25852
rect 11404 25507 11444 25516
rect 10886 24212 11254 24221
rect 10886 24163 11254 24172
rect 10828 24044 10868 24053
rect 11308 24044 11348 25096
rect 11404 25220 11444 25229
rect 11404 25136 11444 25180
rect 11404 25085 11444 25096
rect 10828 23708 10868 24004
rect 11116 24004 11348 24044
rect 11500 24632 11540 27616
rect 11116 23792 11156 24004
rect 11116 23743 11156 23752
rect 11212 23876 11252 23885
rect 10828 23659 10868 23668
rect 10732 23323 10772 23332
rect 11212 22868 11252 23836
rect 11212 22819 11252 22828
rect 11308 23876 11348 23885
rect 10886 22700 11254 22709
rect 10886 22651 11254 22660
rect 10732 22532 10772 22541
rect 10732 22397 10772 22492
rect 11116 22532 11156 22541
rect 11116 21608 11156 22492
rect 11116 21559 11156 21568
rect 10732 21524 10772 21533
rect 10732 20852 10772 21484
rect 10886 21188 11254 21197
rect 10886 21139 11254 21148
rect 10732 20803 10772 20812
rect 11020 20768 11060 20777
rect 11060 20728 11156 20768
rect 11020 20633 11060 20728
rect 10636 20560 10868 20600
rect 10348 20047 10388 20056
rect 10636 20264 10676 20273
rect 10444 19928 10484 19937
rect 10252 18871 10292 18880
rect 10348 19508 10388 19517
rect 10348 18668 10388 19468
rect 10444 19508 10484 19888
rect 10636 19760 10676 20224
rect 10828 20180 10868 20560
rect 10924 20180 10964 20189
rect 10828 20140 10924 20180
rect 10924 20131 10964 20140
rect 11116 20180 11156 20728
rect 11116 20131 11156 20140
rect 10828 20012 10868 20021
rect 10636 19711 10676 19720
rect 10732 19972 10828 20012
rect 10444 19459 10484 19468
rect 10732 19424 10772 19972
rect 10828 19963 10868 19972
rect 11116 20012 11156 20021
rect 11116 19877 11156 19972
rect 10886 19676 11254 19685
rect 10886 19627 11254 19636
rect 10732 19375 10772 19384
rect 10540 19256 10580 19265
rect 10540 18920 10580 19216
rect 10924 19256 10964 19265
rect 11308 19256 11348 23836
rect 11500 23876 11540 24592
rect 11500 23827 11540 23836
rect 10964 19216 11348 19256
rect 11404 23708 11444 23717
rect 11404 19256 11444 23668
rect 11500 23288 11540 23297
rect 11500 23036 11540 23248
rect 11500 22987 11540 22996
rect 11500 22784 11540 22793
rect 11500 22532 11540 22744
rect 11500 22483 11540 22492
rect 11596 21608 11636 28600
rect 12364 28328 12404 28600
rect 12364 28279 12404 28288
rect 12556 28328 12596 28337
rect 12126 27992 12494 28001
rect 12126 27943 12494 27952
rect 11788 27572 11828 27581
rect 11788 26816 11828 27532
rect 12364 27572 12404 27581
rect 11980 27488 12020 27497
rect 11980 27068 12020 27448
rect 11980 27019 12020 27028
rect 12364 27152 12404 27532
rect 11692 26228 11732 26237
rect 11692 26144 11732 26188
rect 11692 26093 11732 26104
rect 11788 26060 11828 26776
rect 12268 26984 12308 26993
rect 12172 26648 12212 26657
rect 12268 26648 12308 26944
rect 12364 26900 12404 27112
rect 12364 26851 12404 26860
rect 12556 26900 12596 28288
rect 12556 26851 12596 26860
rect 12212 26608 12308 26648
rect 12172 26599 12212 26608
rect 12126 26480 12494 26489
rect 12126 26431 12494 26440
rect 11788 26011 11828 26020
rect 11884 26312 11924 26321
rect 11692 25892 11732 25901
rect 11692 25640 11732 25852
rect 11884 25640 11924 26272
rect 12268 26144 12308 26153
rect 12076 25976 12116 25985
rect 11692 25600 11924 25640
rect 11980 25892 12020 25901
rect 11692 25304 11732 25600
rect 11692 25255 11732 25264
rect 11788 25472 11828 25481
rect 11788 24548 11828 25432
rect 11980 25304 12020 25852
rect 12076 25472 12116 25936
rect 12076 25423 12116 25432
rect 11980 25255 12020 25264
rect 11884 25220 11924 25229
rect 11884 24968 11924 25180
rect 12268 25136 12308 26104
rect 11884 24919 11924 24928
rect 11980 25096 12308 25136
rect 12556 25136 12596 25145
rect 11980 24884 12020 25096
rect 12126 24968 12494 24977
rect 12126 24919 12494 24928
rect 11980 24632 12020 24844
rect 11980 24583 12020 24592
rect 12556 24548 12596 25096
rect 11788 24499 11828 24508
rect 12460 24508 12596 24548
rect 11980 24464 12020 24473
rect 11884 23456 11924 23465
rect 11692 23288 11732 23297
rect 11692 21608 11732 23248
rect 11884 23288 11924 23416
rect 11884 23239 11924 23248
rect 11788 23120 11828 23129
rect 11788 22280 11828 23080
rect 11980 23120 12020 24424
rect 12364 24380 12404 24389
rect 12364 23960 12404 24340
rect 12364 23911 12404 23920
rect 12460 23708 12500 24508
rect 12556 24380 12596 24389
rect 12556 23792 12596 24340
rect 12556 23743 12596 23752
rect 12460 23659 12500 23668
rect 12652 23708 12692 28624
rect 13112 28600 13192 29000
rect 13516 28916 13556 28925
rect 13036 28328 13076 28337
rect 12940 26564 12980 26573
rect 12844 26228 12884 26237
rect 12844 26144 12884 26188
rect 12940 26228 12980 26524
rect 12940 26179 12980 26188
rect 12844 26093 12884 26104
rect 12748 25304 12788 25313
rect 12748 24044 12788 25264
rect 12940 25304 12980 25313
rect 12844 25220 12884 25229
rect 12844 24716 12884 25180
rect 12844 24667 12884 24676
rect 12844 24296 12884 24305
rect 12844 24161 12884 24256
rect 12748 23995 12788 24004
rect 12652 23659 12692 23668
rect 12126 23456 12494 23465
rect 12126 23407 12494 23416
rect 12940 23372 12980 25264
rect 13036 23960 13076 28288
rect 13132 28160 13172 28600
rect 13132 28111 13172 28120
rect 13132 27992 13172 28001
rect 13132 26396 13172 27952
rect 13228 27656 13268 27665
rect 13228 26900 13268 27616
rect 13516 27656 13556 28876
rect 13880 28600 13960 29000
rect 14648 28600 14728 29000
rect 15416 28600 15496 29000
rect 16184 28600 16264 29000
rect 23096 28600 23176 29000
rect 23864 28600 23944 29000
rect 24632 28600 24712 29000
rect 25400 28600 25480 29000
rect 26168 28600 26248 29000
rect 26936 28600 27016 29000
rect 27704 28600 27784 29000
rect 28472 28600 28552 29000
rect 29240 28600 29320 29000
rect 30008 28600 30088 29000
rect 30776 28600 30856 29000
rect 13708 28412 13748 28421
rect 13516 27607 13556 27616
rect 13612 28160 13652 28169
rect 13228 26851 13268 26860
rect 13516 26984 13556 26995
rect 13516 26900 13556 26944
rect 13516 26851 13556 26860
rect 13324 26816 13364 26825
rect 13132 26356 13268 26396
rect 13132 26228 13172 26237
rect 13132 25976 13172 26188
rect 13132 25927 13172 25936
rect 13228 25976 13268 26356
rect 13228 25927 13268 25936
rect 13324 26060 13364 26776
rect 13516 26732 13556 26741
rect 13420 26648 13460 26657
rect 13420 26144 13460 26608
rect 13516 26597 13556 26692
rect 13420 26095 13460 26104
rect 13516 26312 13556 26321
rect 13324 25388 13364 26020
rect 13516 25472 13556 26272
rect 13516 25423 13556 25432
rect 13324 25348 13460 25388
rect 13324 25220 13364 25229
rect 13228 24800 13268 24809
rect 13228 24632 13268 24760
rect 13228 24583 13268 24592
rect 13324 24632 13364 25180
rect 13036 23911 13076 23920
rect 13228 24296 13268 24305
rect 12940 23323 12980 23332
rect 13036 23792 13076 23801
rect 11980 23071 12020 23080
rect 12844 23036 12884 23045
rect 11884 22868 11924 22877
rect 11884 22733 11924 22828
rect 11788 22231 11828 22240
rect 12126 21944 12494 21953
rect 12126 21895 12494 21904
rect 11788 21608 11828 21617
rect 11692 21568 11788 21608
rect 11596 21559 11636 21568
rect 11692 21356 11732 21365
rect 11596 21272 11636 21281
rect 11596 20768 11636 21232
rect 11692 21221 11732 21316
rect 11788 21104 11828 21568
rect 12844 21608 12884 22996
rect 12844 21559 12884 21568
rect 12940 22112 12980 22121
rect 11788 21055 11828 21064
rect 11980 21356 12020 21365
rect 11596 20719 11636 20728
rect 11596 20600 11636 20609
rect 11596 20096 11636 20560
rect 10540 18871 10580 18880
rect 10732 19088 10772 19097
rect 10732 18920 10772 19048
rect 10348 18619 10388 18628
rect 10444 18752 10484 18761
rect 10156 18451 10196 18460
rect 10156 17576 10196 17585
rect 10156 17072 10196 17536
rect 10444 17156 10484 18712
rect 10732 18584 10772 18880
rect 10828 19004 10868 19013
rect 10828 18836 10868 18964
rect 10828 18787 10868 18796
rect 10924 18752 10964 19216
rect 11404 19088 11444 19216
rect 11404 19039 11444 19048
rect 11500 20056 11596 20096
rect 11308 19004 11348 19013
rect 10924 18703 10964 18712
rect 11020 18920 11060 18929
rect 10540 18416 10580 18427
rect 10540 18332 10580 18376
rect 10732 18416 10772 18544
rect 11020 18500 11060 18880
rect 11020 18451 11060 18460
rect 10732 18367 10772 18376
rect 10540 18283 10580 18292
rect 10636 18332 10676 18341
rect 10156 17023 10196 17032
rect 10252 17116 10484 17156
rect 10540 17576 10580 17585
rect 10060 14755 10100 14764
rect 10156 16568 10196 16577
rect 10156 15560 10196 16528
rect 10252 16148 10292 17116
rect 10348 16988 10388 16997
rect 10348 16652 10388 16948
rect 10348 16603 10388 16612
rect 10444 16652 10484 16661
rect 10444 16484 10484 16612
rect 10444 16400 10484 16444
rect 10444 16349 10484 16360
rect 10252 15896 10292 16108
rect 10252 15847 10292 15856
rect 10444 16232 10484 16241
rect 10444 15896 10484 16192
rect 10444 15847 10484 15856
rect 10444 15728 10484 15739
rect 10444 15644 10484 15688
rect 10444 15595 10484 15604
rect 10156 14720 10196 15520
rect 10156 14671 10196 14680
rect 10252 15560 10292 15569
rect 10156 14384 10196 14393
rect 10156 14132 10196 14344
rect 10060 14048 10100 14057
rect 10060 13913 10100 14008
rect 10156 13880 10196 14092
rect 10156 13831 10196 13840
rect 10252 13964 10292 15520
rect 10348 15476 10388 15571
rect 10348 15427 10388 15436
rect 10540 15476 10580 17536
rect 10636 16568 10676 18292
rect 10732 18164 10772 18173
rect 10732 17996 10772 18124
rect 10886 18164 11254 18173
rect 10886 18115 11254 18124
rect 10732 17947 10772 17956
rect 11308 17744 11348 18964
rect 11404 18920 11444 18929
rect 11500 18920 11540 20056
rect 11596 20047 11636 20056
rect 11884 20600 11924 20609
rect 11884 20432 11924 20560
rect 11884 20264 11924 20392
rect 11596 19844 11636 19853
rect 11596 19709 11636 19804
rect 11692 19508 11732 19517
rect 11692 19424 11732 19468
rect 11692 19373 11732 19384
rect 11788 19508 11828 19517
rect 11788 19256 11828 19468
rect 11788 19207 11828 19216
rect 11444 18880 11540 18920
rect 11404 18871 11444 18880
rect 11500 18416 11540 18880
rect 11500 18367 11540 18376
rect 11596 19172 11636 19181
rect 11500 18248 11540 18259
rect 11500 18164 11540 18208
rect 11500 18115 11540 18124
rect 11308 17695 11348 17704
rect 11212 17660 11252 17669
rect 10636 16519 10676 16528
rect 10732 17156 10772 17165
rect 11212 17156 11252 17620
rect 11404 17660 11444 17669
rect 11404 17576 11444 17620
rect 11404 17525 11444 17536
rect 11500 17576 11540 17585
rect 11596 17576 11636 19132
rect 11692 19088 11732 19097
rect 11692 18920 11732 19048
rect 11692 18871 11732 18880
rect 11540 17536 11636 17576
rect 11692 18080 11732 18089
rect 11692 17744 11732 18040
rect 11500 17408 11540 17536
rect 11500 17359 11540 17368
rect 11404 17156 11444 17165
rect 11212 17116 11404 17156
rect 10732 16484 10772 17116
rect 10828 17072 10868 17081
rect 10828 16937 10868 17032
rect 10886 16652 11254 16661
rect 10886 16603 11254 16612
rect 10732 16444 10964 16484
rect 10636 16400 10676 16409
rect 10636 15728 10676 16360
rect 10636 15679 10676 15688
rect 10732 16232 10772 16241
rect 10540 15427 10580 15436
rect 10732 15476 10772 16192
rect 10924 15644 10964 16444
rect 11020 16400 11060 16409
rect 11020 16316 11060 16360
rect 11020 16265 11060 16276
rect 10924 15595 10964 15604
rect 11212 16232 11252 16243
rect 11212 16148 11252 16192
rect 11116 15560 11156 15569
rect 11212 15560 11252 16108
rect 11308 15980 11348 15989
rect 11308 15812 11348 15940
rect 11308 15763 11348 15772
rect 11404 15896 11444 17116
rect 11596 17072 11636 17081
rect 11156 15520 11252 15560
rect 11116 15511 11156 15520
rect 10348 15308 10388 15317
rect 10348 14300 10388 15268
rect 10540 15224 10580 15233
rect 10444 15140 10484 15149
rect 10444 15005 10484 15100
rect 10540 14804 10580 15184
rect 10348 14165 10388 14260
rect 10444 14764 10540 14804
rect 10252 13796 10292 13924
rect 10252 13747 10292 13756
rect 10156 13712 10196 13721
rect 10060 13292 10100 13301
rect 10156 13292 10196 13672
rect 10252 13292 10292 13301
rect 10156 13252 10252 13292
rect 10060 13157 10100 13252
rect 10156 12452 10196 12461
rect 10060 11864 10100 11959
rect 10060 11815 10100 11824
rect 10156 11780 10196 12412
rect 9772 10891 9812 10900
rect 9868 10900 10004 10940
rect 10060 11696 10100 11705
rect 10060 11360 10100 11656
rect 9484 8119 9524 8128
rect 9580 10604 9620 10613
rect 9292 7363 9332 7372
rect 9100 7160 9140 7169
rect 9004 6488 9044 6497
rect 9004 5900 9044 6448
rect 9004 5648 9044 5860
rect 9004 5599 9044 5608
rect 8908 4843 8948 4852
rect 7564 4759 7604 4768
rect 3112 4556 3480 4565
rect 3112 4507 3480 4516
rect 9100 4304 9140 7120
rect 9100 4255 9140 4264
rect 9580 6488 9620 10564
rect 9676 10100 9716 10109
rect 9676 9428 9716 10060
rect 9772 10016 9812 10025
rect 9772 9512 9812 9976
rect 9772 9463 9812 9472
rect 9676 9379 9716 9388
rect 9868 9260 9908 10900
rect 10060 10856 10100 11320
rect 10156 11108 10196 11740
rect 10252 11360 10292 13252
rect 10444 13040 10484 14764
rect 10540 14755 10580 14764
rect 10636 14636 10676 14645
rect 10636 14468 10676 14596
rect 10636 14300 10676 14428
rect 10636 14251 10676 14260
rect 10636 14132 10676 14141
rect 10540 13796 10580 13805
rect 10540 13208 10580 13756
rect 10636 13376 10676 14092
rect 10636 13327 10676 13336
rect 10540 13159 10580 13168
rect 10444 12991 10484 13000
rect 10732 12872 10772 15436
rect 11212 15308 11252 15520
rect 11308 15644 11348 15653
rect 11308 15392 11348 15604
rect 11308 15343 11348 15352
rect 11212 15259 11252 15268
rect 10886 15140 11254 15149
rect 10886 15091 11254 15100
rect 11116 14972 11156 14981
rect 11020 14888 11060 14897
rect 10828 14804 10868 14813
rect 10828 13796 10868 14764
rect 11020 14552 11060 14848
rect 11116 14804 11156 14932
rect 11116 14755 11156 14764
rect 11308 14972 11348 14981
rect 11020 14503 11060 14512
rect 11116 14636 11156 14647
rect 11116 14552 11156 14596
rect 11116 14503 11156 14512
rect 11308 14132 11348 14932
rect 11404 14216 11444 15856
rect 11500 16904 11540 16913
rect 11500 15392 11540 16864
rect 11596 16568 11636 17032
rect 11692 16988 11732 17704
rect 11788 17744 11828 17753
rect 11884 17744 11924 20224
rect 11980 20096 12020 21316
rect 12940 20684 12980 22072
rect 12940 20635 12980 20644
rect 12844 20600 12884 20609
rect 12126 20432 12494 20441
rect 12126 20383 12494 20392
rect 12844 20348 12884 20560
rect 12844 20299 12884 20308
rect 12556 20180 12596 20189
rect 11980 20047 12020 20056
rect 12364 20096 12404 20105
rect 12364 19760 12404 20056
rect 12364 19711 12404 19720
rect 12556 19760 12596 20140
rect 12126 18920 12494 18929
rect 12126 18871 12494 18880
rect 12556 18752 12596 19720
rect 12652 20180 12692 20189
rect 12652 19256 12692 20140
rect 13036 20180 13076 23752
rect 13228 23204 13268 24256
rect 13132 23120 13172 23129
rect 13132 22364 13172 23080
rect 13132 22315 13172 22324
rect 13228 22196 13268 23164
rect 13228 21608 13268 22156
rect 13324 21776 13364 24592
rect 13420 25136 13460 25348
rect 13420 23372 13460 25096
rect 13516 24632 13556 24641
rect 13516 24044 13556 24592
rect 13516 23995 13556 24004
rect 13516 23876 13556 23885
rect 13516 23741 13556 23836
rect 13420 23323 13460 23332
rect 13420 23120 13460 23129
rect 13420 23036 13460 23080
rect 13420 22985 13460 22996
rect 13516 23120 13556 23129
rect 13324 21727 13364 21736
rect 13420 22364 13460 22373
rect 13420 21692 13460 22324
rect 13516 22280 13556 23080
rect 13612 23060 13652 28120
rect 13708 26144 13748 28372
rect 13804 28076 13844 28085
rect 13804 27740 13844 28036
rect 13900 27908 13940 28600
rect 13900 27859 13940 27868
rect 14092 28580 14132 28589
rect 13900 27740 13940 27749
rect 13804 27700 13900 27740
rect 13900 27691 13940 27700
rect 13804 27572 13844 27581
rect 13804 26648 13844 27532
rect 14092 27572 14132 28540
rect 14092 27523 14132 27532
rect 14284 27656 14324 27665
rect 14188 27068 14228 27077
rect 13900 26984 13940 26995
rect 13900 26900 13940 26944
rect 13900 26851 13940 26860
rect 14092 26774 14132 26783
rect 13804 26599 13844 26608
rect 13900 26732 13940 26741
rect 13900 26396 13940 26692
rect 13900 26347 13940 26356
rect 14092 26564 14132 26734
rect 14188 26564 14228 27028
rect 14284 26732 14324 27616
rect 14668 27068 14708 28600
rect 15340 27908 15380 27917
rect 14668 27019 14708 27028
rect 15244 27152 15284 27161
rect 15244 26984 15284 27112
rect 15244 26935 15284 26944
rect 15052 26816 15092 26825
rect 14284 26683 14324 26692
rect 14668 26732 14708 26741
rect 14092 26524 14228 26564
rect 14572 26648 14612 26657
rect 14572 26564 14612 26608
rect 13900 26228 13940 26237
rect 13804 26144 13844 26153
rect 13708 26104 13804 26144
rect 13804 26095 13844 26104
rect 13900 26060 13940 26188
rect 13900 26011 13940 26020
rect 13996 26144 14036 26153
rect 13900 25892 13940 25901
rect 13996 25892 14036 26104
rect 13940 25852 14036 25892
rect 14092 26144 14132 26524
rect 14572 26513 14612 26524
rect 14476 26396 14516 26405
rect 14516 26356 14612 26396
rect 14476 26347 14516 26356
rect 13900 25843 13940 25852
rect 14092 25724 14132 26104
rect 13804 25684 14132 25724
rect 14188 26312 14228 26321
rect 14188 25892 14228 26272
rect 14476 26228 14516 26237
rect 13708 25220 13748 25229
rect 13708 25085 13748 25180
rect 13804 25136 13844 25684
rect 14188 25640 14228 25852
rect 14092 25472 14132 25481
rect 13900 25432 14092 25472
rect 13900 25388 13940 25432
rect 14092 25423 14132 25432
rect 14188 25388 14228 25600
rect 14380 26188 14476 26228
rect 14380 25556 14420 26188
rect 14476 26179 14516 26188
rect 14380 25507 14420 25516
rect 14476 25892 14516 25901
rect 14476 25472 14516 25852
rect 14572 25892 14612 26356
rect 14572 25843 14612 25852
rect 14476 25423 14516 25432
rect 14380 25388 14420 25397
rect 14188 25348 14380 25388
rect 13900 25339 13940 25348
rect 14380 25339 14420 25348
rect 14380 25220 14420 25229
rect 13900 25136 13940 25145
rect 13804 25096 13900 25136
rect 13900 24884 13940 25096
rect 13900 24632 13940 24844
rect 14380 24716 14420 25180
rect 14668 25220 14708 26692
rect 14860 26732 14900 26741
rect 14860 26597 14900 26692
rect 14764 26480 14804 26489
rect 14764 25556 14804 26440
rect 14956 26396 14996 26407
rect 14956 26312 14996 26356
rect 14956 26263 14996 26272
rect 14860 26144 14900 26153
rect 14860 26009 14900 26104
rect 14764 25507 14804 25516
rect 14860 25808 14900 25817
rect 14860 25304 14900 25768
rect 14860 25255 14900 25264
rect 14956 25472 14996 25481
rect 14668 25171 14708 25180
rect 14380 24667 14420 24676
rect 14476 25052 14516 25061
rect 13900 24583 13940 24592
rect 14188 24296 14228 24305
rect 13612 23020 13748 23060
rect 13516 21944 13556 22240
rect 13516 21895 13556 21904
rect 13708 21776 13748 23020
rect 14188 23036 14228 24256
rect 14188 22987 14228 22996
rect 14284 23960 14324 23969
rect 14284 22280 14324 23920
rect 14476 23204 14516 25012
rect 14764 25052 14804 25061
rect 14476 23120 14516 23164
rect 14668 23624 14708 23633
rect 14668 23288 14708 23584
rect 14476 23040 14516 23080
rect 14572 23120 14612 23129
rect 14572 22868 14612 23080
rect 14572 22819 14612 22828
rect 14284 22231 14324 22240
rect 13708 21727 13748 21736
rect 14380 22196 14420 22205
rect 13132 21568 13228 21608
rect 13132 20936 13172 21568
rect 13228 21559 13268 21568
rect 13324 21608 13364 21617
rect 13324 21188 13364 21568
rect 13132 20887 13172 20896
rect 13228 21020 13268 21029
rect 13228 20684 13268 20980
rect 13324 20936 13364 21148
rect 13324 20887 13364 20896
rect 13228 20635 13268 20644
rect 13324 20768 13364 20777
rect 13324 20600 13364 20728
rect 13324 20551 13364 20560
rect 13420 20684 13460 21652
rect 13516 21608 13556 21617
rect 13516 20852 13556 21568
rect 13996 21608 14036 21617
rect 13804 21524 13844 21533
rect 13516 20717 13556 20812
rect 13708 21356 13748 21365
rect 13708 20852 13748 21316
rect 13708 20768 13748 20812
rect 13708 20688 13748 20728
rect 13420 20348 13460 20644
rect 13420 20299 13460 20308
rect 13804 20348 13844 21484
rect 13996 20768 14036 21568
rect 13900 20600 13940 20628
rect 13996 20600 14036 20728
rect 14380 21608 14420 22156
rect 14380 20768 14420 21568
rect 14380 20719 14420 20728
rect 13940 20560 13996 20600
rect 13900 20551 13940 20560
rect 13996 20551 14036 20560
rect 14572 20684 14612 20693
rect 13804 20299 13844 20308
rect 14380 20348 14420 20357
rect 12844 20096 12884 20105
rect 12844 19508 12884 20056
rect 12844 19459 12884 19468
rect 12652 19207 12692 19216
rect 12748 19424 12788 19433
rect 12556 18703 12596 18712
rect 12076 18416 12116 18425
rect 11980 18332 12020 18341
rect 11980 18197 12020 18292
rect 11828 17704 11924 17744
rect 11788 17695 11828 17704
rect 11788 17576 11828 17585
rect 11788 17240 11828 17536
rect 11884 17408 11924 17704
rect 12076 17996 12116 18376
rect 12076 17744 12116 17956
rect 12076 17695 12116 17704
rect 12172 18332 12212 18341
rect 12172 17660 12212 18292
rect 12268 17996 12308 18005
rect 12268 17828 12308 17956
rect 12556 17996 12596 18005
rect 12268 17779 12308 17788
rect 12460 17912 12500 17923
rect 12460 17828 12500 17872
rect 12460 17779 12500 17788
rect 12172 17611 12212 17620
rect 11884 17359 11924 17368
rect 11980 17576 12020 17585
rect 11788 17191 11828 17200
rect 11980 17156 12020 17536
rect 12268 17576 12308 17671
rect 12268 17527 12308 17536
rect 12126 17408 12494 17417
rect 12126 17359 12494 17368
rect 12556 17324 12596 17956
rect 12556 17240 12596 17284
rect 11980 17107 12020 17116
rect 12460 17200 12596 17240
rect 12460 17156 12500 17200
rect 12556 17189 12596 17200
rect 12652 17828 12692 17837
rect 12652 17240 12692 17788
rect 12460 17107 12500 17116
rect 12652 17156 12692 17200
rect 12652 17105 12692 17116
rect 11692 16939 11732 16948
rect 12364 16988 12404 16997
rect 11980 16820 12020 16829
rect 11884 16736 11924 16745
rect 11596 16519 11636 16528
rect 11692 16652 11732 16661
rect 11692 16400 11732 16612
rect 11692 16351 11732 16360
rect 11884 16316 11924 16696
rect 11884 16267 11924 16276
rect 11788 16232 11828 16243
rect 11788 16148 11828 16192
rect 11788 16099 11828 16108
rect 11980 16232 12020 16780
rect 12364 16820 12404 16948
rect 12364 16771 12404 16780
rect 12556 16904 12596 16913
rect 11500 15343 11540 15352
rect 11596 15980 11636 15989
rect 11596 15056 11636 15940
rect 11596 15007 11636 15016
rect 11884 15560 11924 15569
rect 11884 14972 11924 15520
rect 11980 15476 12020 16192
rect 12460 16400 12500 16409
rect 12460 16232 12500 16360
rect 12460 16183 12500 16192
rect 12126 15896 12494 15905
rect 12126 15847 12494 15856
rect 12460 15728 12500 15737
rect 11980 15427 12020 15436
rect 12172 15560 12212 15569
rect 12172 15425 12212 15520
rect 11884 14923 11924 14932
rect 12172 15308 12212 15317
rect 11980 14804 12020 14813
rect 11692 14720 11732 14729
rect 11404 14167 11444 14176
rect 11500 14636 11540 14645
rect 11500 14552 11540 14596
rect 11308 14083 11348 14092
rect 11500 14132 11540 14512
rect 11596 14552 11636 14561
rect 11596 14384 11636 14512
rect 11596 14335 11636 14344
rect 10828 13747 10868 13756
rect 11404 14048 11444 14057
rect 10886 13628 11254 13637
rect 10886 13579 11254 13588
rect 11404 13544 11444 14008
rect 11404 13495 11444 13504
rect 11308 13460 11348 13469
rect 11212 13292 11252 13301
rect 10444 12832 10772 12872
rect 10828 13124 10868 13133
rect 10348 12368 10388 12377
rect 10348 11612 10388 12328
rect 10348 11563 10388 11572
rect 10444 11444 10484 12832
rect 10828 12620 10868 13084
rect 11212 13124 11252 13252
rect 11212 13075 11252 13084
rect 10828 12571 10868 12580
rect 11212 12956 11252 12965
rect 11212 12536 11252 12916
rect 11212 12487 11252 12496
rect 10636 12284 10676 12293
rect 10252 11311 10292 11320
rect 10348 11404 10484 11444
rect 10540 11864 10580 11873
rect 10156 11059 10196 11068
rect 10156 10856 10196 10865
rect 10060 10816 10156 10856
rect 9964 10772 10004 10781
rect 9964 9512 10004 10732
rect 10156 10184 10196 10816
rect 10060 9932 10100 9941
rect 10060 9797 10100 9892
rect 9964 9463 10004 9472
rect 10060 9596 10100 9605
rect 9868 9211 9908 9220
rect 9676 9008 9716 9017
rect 9676 8672 9716 8968
rect 9772 8924 9812 9019
rect 9772 8875 9812 8884
rect 9676 8623 9716 8632
rect 9772 8756 9812 8765
rect 9772 8168 9812 8716
rect 10060 8672 10100 9556
rect 9772 8119 9812 8128
rect 9964 8504 10004 8513
rect 9964 8000 10004 8464
rect 9964 7951 10004 7960
rect 9772 7160 9812 7169
rect 9772 6656 9812 7120
rect 9772 6607 9812 6616
rect 9580 4220 9620 6448
rect 10060 6488 10100 8632
rect 10060 6439 10100 6448
rect 10156 8840 10196 10144
rect 10252 10604 10292 10613
rect 10252 10100 10292 10564
rect 10252 10051 10292 10060
rect 10348 9848 10388 11404
rect 10348 9799 10388 9808
rect 10444 10520 10484 10529
rect 10444 9932 10484 10480
rect 10444 9512 10484 9892
rect 10444 9463 10484 9472
rect 10252 8840 10292 8868
rect 10156 8800 10252 8840
rect 9580 4171 9620 4180
rect 9772 6404 9812 6413
rect 9772 4976 9812 6364
rect 10060 5564 10100 5573
rect 10156 5564 10196 8800
rect 10252 8791 10292 8800
rect 10252 8672 10292 8681
rect 10252 8000 10292 8632
rect 10252 7496 10292 7960
rect 10252 7447 10292 7456
rect 10540 8672 10580 11824
rect 10636 11276 10676 12244
rect 10732 12284 10772 12293
rect 10732 12032 10772 12244
rect 10886 12116 11254 12125
rect 10886 12067 11254 12076
rect 10732 11983 10772 11992
rect 11020 11528 11060 11537
rect 10636 11227 10676 11236
rect 10732 11360 10772 11369
rect 10636 10772 10676 10781
rect 10636 9512 10676 10732
rect 10732 10100 10772 11320
rect 11020 11024 11060 11488
rect 11020 10975 11060 10984
rect 11308 10940 11348 13420
rect 11404 13376 11444 13385
rect 11404 13124 11444 13336
rect 11404 12620 11444 13084
rect 11500 12704 11540 14092
rect 11596 13208 11636 13219
rect 11596 13124 11636 13168
rect 11596 13075 11636 13084
rect 11692 12980 11732 14680
rect 11980 14636 12020 14764
rect 12172 14720 12212 15268
rect 12364 15308 12404 15317
rect 12364 15173 12404 15268
rect 12172 14671 12212 14680
rect 11980 14587 12020 14596
rect 12460 14636 12500 15688
rect 12460 14587 12500 14596
rect 12126 14384 12494 14393
rect 12126 14335 12494 14344
rect 11788 14300 11828 14309
rect 11788 13292 11828 14260
rect 12268 14216 12308 14225
rect 11884 14048 11924 14057
rect 11884 13712 11924 14008
rect 12268 14048 12308 14176
rect 12268 13999 12308 14008
rect 12460 13964 12500 13973
rect 12460 13829 12500 13924
rect 12364 13796 12404 13805
rect 11924 13672 12020 13712
rect 11884 13663 11924 13672
rect 11788 13243 11828 13252
rect 11500 12655 11540 12664
rect 11596 12940 11732 12980
rect 11788 13040 11828 13049
rect 11404 12571 11444 12580
rect 11500 11696 11540 11705
rect 11500 11192 11540 11656
rect 10886 10604 11254 10613
rect 10886 10555 11254 10564
rect 10732 10051 10772 10060
rect 11020 10436 11060 10445
rect 10636 9463 10676 9472
rect 11020 10016 11060 10396
rect 11308 10268 11348 10900
rect 11308 10219 11348 10228
rect 11404 11024 11444 11033
rect 11020 9260 11060 9976
rect 11212 9512 11252 9521
rect 11252 9472 11348 9512
rect 11212 9463 11252 9472
rect 10540 7160 10580 8632
rect 10636 9220 11060 9260
rect 10636 8252 10676 9220
rect 10886 9092 11254 9101
rect 10886 9043 11254 9052
rect 10828 8924 10868 8933
rect 10636 8203 10676 8212
rect 10732 8756 10772 8765
rect 10100 5524 10196 5564
rect 10252 6656 10292 6665
rect 10252 5648 10292 6616
rect 10540 6320 10580 7120
rect 10540 6271 10580 6280
rect 10636 8000 10676 8009
rect 10636 7076 10676 7960
rect 10636 6236 10676 7036
rect 10732 6656 10772 8716
rect 10828 8000 10868 8884
rect 10828 7951 10868 7960
rect 10886 7580 11254 7589
rect 10886 7531 11254 7540
rect 10732 6607 10772 6616
rect 11116 7160 11156 7169
rect 10828 6404 10868 6413
rect 11116 6404 11156 7120
rect 11308 7160 11348 9472
rect 11404 8504 11444 10984
rect 11500 9512 11540 11152
rect 11500 9377 11540 9472
rect 11404 8455 11444 8464
rect 11500 8672 11540 8681
rect 11500 8168 11540 8632
rect 11500 8119 11540 8128
rect 11308 7111 11348 7120
rect 11500 8000 11540 8009
rect 10868 6364 11156 6404
rect 11308 6992 11348 7001
rect 11308 6488 11348 6952
rect 11500 6740 11540 7960
rect 11596 7244 11636 12940
rect 11692 10268 11732 10277
rect 11692 9596 11732 10228
rect 11788 9764 11828 13000
rect 11884 12536 11924 12545
rect 11884 10520 11924 12496
rect 11980 11864 12020 13672
rect 12364 13292 12404 13756
rect 12556 13460 12596 16864
rect 12652 16316 12692 16325
rect 12652 15308 12692 16276
rect 12652 15259 12692 15268
rect 12748 14804 12788 19384
rect 13036 19340 13076 20140
rect 13324 20180 13364 20189
rect 13036 19291 13076 19300
rect 13132 19760 13172 19769
rect 13132 19172 13172 19720
rect 13324 19676 13364 20140
rect 14188 20096 14228 20105
rect 13900 20012 13940 20021
rect 13324 19627 13364 19636
rect 13420 19676 13460 19685
rect 12940 19004 12980 19013
rect 12940 18869 12980 18964
rect 13132 19004 13172 19132
rect 13132 18955 13172 18964
rect 13228 19424 13268 19433
rect 13228 19256 13268 19384
rect 13132 18584 13172 18593
rect 13132 17996 13172 18544
rect 13132 17947 13172 17956
rect 12844 17912 12884 17921
rect 12844 17576 12884 17872
rect 12844 17527 12884 17536
rect 12940 17660 12980 17669
rect 12940 17525 12980 17620
rect 13036 17576 13076 17585
rect 13036 17156 13076 17536
rect 13228 17576 13268 19216
rect 13228 17240 13268 17536
rect 13324 18500 13364 18509
rect 13324 17744 13364 18460
rect 13420 18080 13460 19636
rect 13804 19256 13844 19265
rect 13516 19088 13556 19097
rect 13516 18752 13556 19048
rect 13516 18584 13556 18712
rect 13516 18535 13556 18544
rect 13612 18668 13652 18677
rect 13420 18031 13460 18040
rect 13324 17492 13364 17704
rect 13612 17996 13652 18628
rect 13804 18584 13844 19216
rect 13804 18500 13844 18544
rect 13804 18451 13844 18460
rect 13612 17744 13652 17956
rect 13612 17695 13652 17704
rect 13324 17443 13364 17452
rect 13228 17191 13268 17200
rect 13036 17107 13076 17116
rect 12940 17072 12980 17081
rect 12844 16400 12884 16409
rect 12844 15980 12884 16360
rect 12940 16232 12980 17032
rect 13228 17072 13268 17081
rect 12940 16183 12980 16192
rect 13036 16736 13076 16745
rect 12844 15931 12884 15940
rect 12940 15980 12980 16020
rect 12940 15896 12980 15940
rect 12844 15728 12884 15737
rect 12844 15476 12884 15688
rect 12940 15560 12980 15856
rect 12940 15511 12980 15520
rect 12844 15392 12884 15436
rect 12844 15341 12884 15352
rect 12940 15308 12980 15317
rect 12940 15173 12980 15268
rect 12556 13411 12596 13420
rect 12652 14764 12748 14804
rect 12652 13292 12692 14764
rect 12748 14755 12788 14764
rect 12844 14972 12884 14981
rect 12844 14720 12884 14932
rect 12844 14671 12884 14680
rect 12748 14552 12788 14561
rect 12748 14300 12788 14512
rect 12748 14251 12788 14260
rect 12940 14132 12980 14141
rect 12748 14048 12788 14057
rect 12748 13628 12788 14008
rect 12940 13880 12980 14092
rect 12940 13831 12980 13840
rect 12748 13579 12788 13588
rect 12364 13243 12404 13252
rect 12460 13252 12692 13292
rect 12172 13208 12212 13217
rect 12172 13040 12212 13168
rect 12460 13208 12500 13252
rect 13036 13208 13076 16696
rect 13132 16232 13172 16241
rect 13132 15812 13172 16192
rect 13228 16148 13268 17032
rect 13324 17072 13364 17081
rect 13324 16568 13364 17032
rect 13804 16820 13844 16829
rect 13324 16519 13364 16528
rect 13420 16736 13460 16745
rect 13420 16400 13460 16696
rect 13324 16148 13364 16157
rect 13228 16108 13324 16148
rect 13324 16099 13364 16108
rect 13132 15763 13172 15772
rect 13324 15980 13364 15989
rect 13228 15728 13268 15737
rect 12460 13159 12500 13168
rect 12940 13168 13076 13208
rect 13132 15308 13172 15317
rect 12172 12991 12212 13000
rect 12556 13124 12596 13133
rect 12126 12872 12494 12881
rect 12126 12823 12494 12832
rect 12556 12704 12596 13084
rect 12940 13040 12980 13168
rect 13132 13124 13172 15268
rect 13228 14720 13268 15688
rect 13324 14972 13364 15940
rect 13324 14923 13364 14932
rect 13420 15308 13460 16360
rect 13708 16484 13748 16493
rect 13708 16316 13748 16444
rect 13804 16400 13844 16780
rect 13804 16351 13844 16360
rect 13708 16267 13748 16276
rect 13516 16148 13556 16157
rect 13516 15728 13556 16108
rect 13516 15679 13556 15688
rect 13612 16064 13652 16073
rect 13420 14804 13460 15268
rect 13420 14764 13556 14804
rect 13228 14680 13460 14720
rect 13228 14552 13268 14561
rect 13228 13292 13268 14512
rect 13324 14384 13364 14393
rect 13324 13964 13364 14344
rect 13324 13712 13364 13924
rect 13324 13663 13364 13672
rect 13228 13243 13268 13252
rect 12940 12991 12980 13000
rect 13036 13084 13172 13124
rect 13324 13124 13364 13219
rect 12556 12655 12596 12664
rect 12076 12620 12116 12629
rect 12076 12485 12116 12580
rect 12940 12536 12980 12545
rect 12748 12452 12788 12461
rect 12652 12200 12692 12209
rect 11980 11696 12020 11824
rect 12460 11948 12500 11957
rect 12460 11780 12500 11908
rect 12500 11740 12596 11780
rect 12460 11731 12500 11740
rect 11980 11647 12020 11656
rect 12172 11696 12212 11705
rect 12172 11561 12212 11656
rect 11980 11444 12020 11453
rect 11980 10940 12020 11404
rect 12126 11360 12494 11369
rect 12126 11311 12494 11320
rect 12556 11192 12596 11740
rect 12652 11528 12692 12160
rect 12652 11479 12692 11488
rect 12748 11948 12788 12412
rect 12556 11143 12596 11152
rect 12652 11108 12692 11117
rect 12268 11024 12308 11033
rect 12172 10940 12212 10949
rect 11980 10900 12172 10940
rect 12172 10891 12212 10900
rect 12268 10889 12308 10984
rect 12652 10973 12692 11068
rect 12748 10940 12788 11908
rect 12940 12032 12980 12496
rect 12844 11612 12884 11621
rect 12844 11024 12884 11572
rect 12940 11108 12980 11992
rect 13036 11528 13076 13084
rect 13324 13075 13364 13084
rect 13420 12872 13460 14680
rect 13516 14132 13556 14764
rect 13612 14720 13652 16024
rect 13708 15980 13748 15989
rect 13708 15812 13748 15940
rect 13708 15476 13748 15772
rect 13708 15427 13748 15436
rect 13612 14671 13652 14680
rect 13804 14552 13844 14561
rect 13516 14083 13556 14092
rect 13708 14132 13748 14141
rect 13516 13796 13556 13805
rect 13516 13544 13556 13756
rect 13516 13292 13556 13504
rect 13516 13243 13556 13252
rect 13612 13460 13652 13469
rect 13420 12832 13556 12872
rect 13420 12704 13460 12713
rect 13420 12569 13460 12664
rect 13324 12116 13364 12125
rect 13036 11479 13076 11488
rect 13228 11696 13268 11705
rect 13228 11192 13268 11656
rect 13228 11143 13268 11152
rect 12940 11059 12980 11068
rect 12844 10975 12884 10984
rect 12748 10891 12788 10900
rect 11884 10471 11924 10480
rect 13228 10604 13268 10613
rect 12652 10268 12692 10277
rect 11788 9715 11828 9724
rect 11980 10016 12020 10025
rect 11980 9596 12020 9976
rect 12556 10016 12596 10025
rect 12126 9848 12494 9857
rect 12126 9799 12494 9808
rect 12556 9848 12596 9976
rect 12556 9799 12596 9808
rect 12556 9680 12596 9689
rect 12076 9596 12116 9605
rect 11980 9556 12076 9596
rect 11692 9547 11732 9556
rect 12076 9547 12116 9556
rect 12460 9512 12500 9521
rect 11884 9428 11924 9437
rect 11692 8588 11732 8597
rect 11692 8000 11732 8548
rect 11692 7865 11732 7960
rect 11788 8504 11828 8513
rect 11788 8336 11828 8464
rect 11596 7195 11636 7204
rect 11692 7664 11732 7673
rect 11692 7160 11732 7624
rect 11788 7244 11828 8296
rect 11884 8168 11924 9388
rect 11980 9428 12020 9437
rect 11980 8252 12020 9388
rect 12460 9377 12500 9472
rect 12126 8336 12494 8345
rect 12126 8287 12494 8296
rect 11980 8203 12020 8212
rect 11884 8119 11924 8128
rect 12268 8168 12308 8177
rect 12076 8084 12116 8093
rect 11788 7195 11828 7204
rect 11980 8000 12020 8009
rect 11692 7111 11732 7120
rect 11500 6691 11540 6700
rect 11980 7076 12020 7960
rect 12076 7916 12116 8044
rect 12076 7867 12116 7876
rect 12268 7160 12308 8128
rect 12556 8084 12596 9640
rect 12556 8035 12596 8044
rect 12268 7111 12308 7120
rect 12364 8000 12404 8009
rect 11980 6656 12020 7036
rect 12364 6992 12404 7960
rect 12652 7412 12692 10228
rect 13036 10100 13076 10109
rect 12940 9596 12980 9605
rect 12844 8840 12884 8849
rect 12748 8504 12788 8513
rect 12748 8000 12788 8464
rect 12748 7951 12788 7960
rect 12652 7363 12692 7372
rect 12364 6943 12404 6952
rect 12126 6824 12494 6833
rect 12126 6775 12494 6784
rect 11980 6607 12020 6616
rect 12460 6656 12500 6665
rect 10828 6355 10868 6364
rect 10636 6187 10676 6196
rect 10886 6068 11254 6077
rect 10886 6019 11254 6028
rect 10060 5496 10100 5524
rect 9772 4724 9812 4936
rect 10252 4892 10292 5608
rect 11212 5732 11252 5741
rect 10348 5228 10388 5237
rect 10348 4976 10388 5188
rect 10348 4927 10388 4936
rect 10252 4843 10292 4852
rect 11212 4808 11252 5692
rect 11308 4976 11348 6448
rect 12460 6488 12500 6616
rect 12460 6439 12500 6448
rect 11596 6404 11636 6413
rect 11500 5900 11540 5909
rect 11500 5060 11540 5860
rect 11500 5011 11540 5020
rect 11308 4927 11348 4936
rect 11596 4892 11636 6364
rect 11596 4843 11636 4852
rect 11788 6320 11828 6329
rect 11788 4892 11828 6280
rect 12844 5900 12884 8800
rect 12940 8756 12980 9556
rect 13036 8924 13076 10060
rect 13132 9512 13172 9521
rect 13132 9377 13172 9472
rect 13228 9428 13268 10564
rect 13324 10352 13364 12076
rect 13324 10303 13364 10312
rect 13324 10184 13364 10193
rect 13324 9680 13364 10144
rect 13324 9631 13364 9640
rect 13420 10016 13460 10025
rect 13228 9379 13268 9388
rect 13036 8875 13076 8884
rect 12940 8707 12980 8716
rect 13228 8756 13268 8765
rect 12844 5851 12884 5860
rect 13036 7076 13076 7085
rect 13036 5900 13076 7036
rect 12940 5732 12980 5741
rect 13036 5732 13076 5860
rect 12980 5692 13076 5732
rect 13132 6488 13172 6497
rect 12940 5664 12980 5692
rect 12844 5564 12884 5573
rect 12126 5312 12494 5321
rect 12126 5263 12494 5272
rect 12844 5060 12884 5524
rect 13036 5564 13076 5573
rect 12844 5011 12884 5020
rect 12940 5060 12980 5069
rect 11788 4843 11828 4852
rect 11980 4976 12020 4985
rect 11212 4759 11252 4768
rect 9772 4136 9812 4684
rect 11980 4724 12020 4936
rect 12940 4892 12980 5020
rect 12940 4843 12980 4852
rect 13036 4808 13076 5524
rect 13132 5144 13172 6448
rect 13228 5648 13268 8716
rect 13420 8672 13460 9976
rect 13516 9932 13556 12832
rect 13612 12536 13652 13420
rect 13708 13040 13748 14092
rect 13804 13292 13844 14512
rect 13804 13243 13844 13252
rect 13708 12704 13748 13000
rect 13804 13124 13844 13133
rect 13804 12989 13844 13084
rect 13804 12872 13844 12881
rect 13804 12737 13844 12832
rect 13708 12655 13748 12664
rect 13804 12620 13844 12629
rect 13804 12536 13844 12580
rect 13612 12496 13844 12536
rect 13804 12368 13844 12377
rect 13804 12233 13844 12328
rect 13900 12284 13940 19972
rect 14188 19256 14228 20056
rect 14380 20012 14420 20308
rect 14572 20180 14612 20644
rect 14572 20131 14612 20140
rect 14380 19963 14420 19972
rect 14188 19207 14228 19216
rect 14572 19844 14612 19853
rect 14572 19256 14612 19804
rect 14572 19207 14612 19216
rect 14284 18920 14324 18929
rect 14284 18668 14324 18880
rect 14284 18584 14324 18628
rect 14284 18533 14324 18544
rect 14188 18500 14228 18509
rect 14188 17912 14228 18460
rect 14188 17863 14228 17872
rect 14380 18500 14420 18509
rect 14284 17576 14324 17585
rect 14092 17240 14132 17251
rect 13996 17156 14036 17165
rect 13996 15224 14036 17116
rect 14092 17156 14132 17200
rect 14132 17116 14228 17156
rect 14092 17107 14132 17116
rect 14092 16484 14132 16493
rect 14092 16316 14132 16444
rect 14188 16400 14228 17116
rect 14284 17072 14324 17536
rect 14380 17156 14420 18460
rect 14476 18332 14516 18341
rect 14476 17744 14516 18292
rect 14476 17695 14516 17704
rect 14380 17107 14420 17116
rect 14572 17660 14612 17669
rect 14284 17023 14324 17032
rect 14188 16351 14228 16360
rect 14380 16988 14420 16997
rect 14092 15812 14132 16276
rect 14380 16148 14420 16948
rect 14380 16099 14420 16108
rect 14476 16820 14516 16829
rect 14476 16232 14516 16780
rect 14284 16064 14324 16073
rect 14284 15896 14324 16024
rect 14092 15772 14228 15812
rect 13996 15175 14036 15184
rect 14188 15308 14228 15772
rect 14284 15644 14324 15856
rect 14476 15728 14516 16192
rect 14476 15679 14516 15688
rect 14284 15595 14324 15604
rect 14380 15560 14420 15569
rect 14188 15173 14228 15268
rect 14284 15476 14324 15485
rect 14284 14972 14324 15436
rect 14284 14923 14324 14932
rect 13996 14804 14036 14813
rect 13996 14636 14036 14764
rect 13996 14300 14036 14596
rect 14188 14720 14228 14729
rect 14188 14552 14228 14680
rect 14188 14503 14228 14512
rect 14284 14636 14324 14645
rect 13996 14251 14036 14260
rect 13996 14048 14036 14057
rect 14036 14008 14132 14048
rect 13996 13999 14036 14008
rect 13900 12235 13940 12244
rect 13804 11444 13844 11453
rect 13708 11024 13748 11033
rect 13708 10016 13748 10984
rect 13804 10856 13844 11404
rect 13804 10807 13844 10816
rect 13900 10940 13940 10949
rect 13900 10688 13940 10900
rect 13708 9967 13748 9976
rect 13804 10648 13940 10688
rect 13804 10100 13844 10648
rect 13996 10352 14036 10361
rect 13516 9512 13556 9892
rect 13516 9463 13556 9472
rect 13420 8623 13460 8632
rect 13612 8672 13652 8681
rect 13324 8588 13364 8597
rect 13324 8000 13364 8548
rect 13324 7244 13364 7960
rect 13612 7832 13652 8632
rect 13804 8168 13844 10060
rect 13900 10184 13940 10193
rect 13900 9680 13940 10144
rect 13900 9631 13940 9640
rect 13804 8119 13844 8128
rect 13996 9512 14036 10312
rect 13612 7783 13652 7792
rect 13900 7748 13940 7757
rect 13324 7109 13364 7204
rect 13708 7244 13748 7253
rect 13708 6488 13748 7204
rect 13708 6439 13748 6448
rect 13900 7160 13940 7708
rect 13996 7412 14036 9472
rect 14092 8168 14132 14008
rect 14284 13880 14324 14596
rect 14380 14216 14420 15520
rect 14572 14888 14612 17620
rect 14668 16736 14708 23248
rect 14764 22448 14804 25012
rect 14956 24800 14996 25432
rect 14956 24751 14996 24760
rect 15052 24632 15092 26776
rect 15340 26816 15380 27868
rect 15436 27236 15476 28600
rect 15436 27187 15476 27196
rect 16012 27320 16052 27329
rect 15436 26984 15476 26993
rect 15436 26849 15476 26944
rect 15820 26984 15860 26993
rect 15340 26396 15380 26776
rect 15340 26347 15380 26356
rect 15436 26648 15476 26657
rect 15340 26144 15380 26239
rect 15340 26095 15380 26104
rect 15436 26060 15476 26608
rect 15436 26011 15476 26020
rect 15532 26228 15572 26237
rect 15340 25892 15380 25901
rect 14956 24592 15092 24632
rect 15244 25220 15284 25229
rect 14860 24380 14900 24389
rect 14860 23792 14900 24340
rect 14860 23743 14900 23752
rect 14764 22399 14804 22408
rect 14860 22280 14900 22289
rect 14764 21524 14804 21533
rect 14764 21020 14804 21484
rect 14764 20971 14804 20980
rect 14860 20936 14900 22240
rect 14860 20887 14900 20896
rect 14860 20768 14900 20777
rect 14860 20633 14900 20728
rect 14956 19592 14996 24592
rect 15148 24380 15188 24389
rect 15148 23876 15188 24340
rect 15148 23827 15188 23836
rect 15244 23792 15284 25180
rect 15244 23204 15284 23752
rect 15244 23155 15284 23164
rect 15244 21776 15284 21785
rect 15052 21524 15092 21533
rect 15052 21356 15092 21484
rect 15244 21524 15284 21736
rect 15244 21475 15284 21484
rect 15052 21307 15092 21316
rect 15148 21272 15188 21281
rect 14956 19543 14996 19552
rect 15052 20852 15092 20861
rect 15052 19508 15092 20812
rect 15148 20348 15188 21232
rect 15340 21272 15380 25852
rect 15436 25220 15476 25315
rect 15436 25171 15476 25180
rect 15532 21860 15572 26188
rect 15724 26228 15764 26237
rect 15628 26144 15668 26153
rect 15628 24128 15668 26104
rect 15724 25472 15764 26188
rect 15820 25892 15860 26944
rect 16012 26312 16052 27280
rect 16204 26732 16244 28600
rect 16204 26683 16244 26692
rect 16492 28580 16532 28589
rect 16396 26564 16436 26573
rect 16396 26396 16436 26524
rect 16396 26347 16436 26356
rect 16012 26263 16052 26272
rect 16204 26144 16244 26153
rect 16204 26060 16244 26104
rect 16204 26009 16244 26020
rect 15820 25843 15860 25852
rect 16396 25892 16436 25901
rect 15724 25423 15764 25432
rect 15916 25304 15956 25313
rect 15628 24079 15668 24088
rect 15724 25136 15764 25145
rect 15724 23876 15764 25096
rect 15820 24128 15860 24139
rect 15820 24044 15860 24088
rect 15820 23995 15860 24004
rect 15628 23792 15668 23803
rect 15628 23708 15668 23752
rect 15628 23288 15668 23668
rect 15628 23239 15668 23248
rect 15724 23036 15764 23836
rect 15916 23792 15956 25264
rect 16396 25304 16436 25852
rect 16396 25255 16436 25264
rect 16204 25220 16244 25229
rect 16108 25136 16148 25145
rect 16108 24800 16148 25096
rect 16108 24751 16148 24760
rect 15916 23456 15956 23752
rect 15916 23407 15956 23416
rect 16012 24716 16052 24725
rect 15724 22987 15764 22996
rect 15724 22364 15764 22373
rect 16012 22364 16052 24676
rect 15764 22324 15860 22364
rect 15724 22315 15764 22324
rect 15532 21811 15572 21820
rect 15628 21608 15668 21617
rect 15340 21223 15380 21232
rect 15532 21524 15572 21533
rect 15532 20936 15572 21484
rect 15532 20887 15572 20896
rect 15244 20768 15284 20777
rect 15244 20600 15284 20728
rect 15244 20551 15284 20560
rect 15148 20299 15188 20308
rect 15244 20096 15284 20105
rect 15052 19459 15092 19468
rect 15148 20012 15188 20021
rect 14956 19340 14996 19349
rect 14764 19088 14804 19097
rect 14804 19048 14900 19088
rect 14764 19039 14804 19048
rect 14764 18584 14804 18593
rect 14764 17912 14804 18544
rect 14764 17828 14804 17872
rect 14764 17748 14804 17788
rect 14764 17660 14804 17669
rect 14764 16904 14804 17620
rect 14764 16855 14804 16864
rect 14668 16696 14804 16736
rect 14668 16484 14708 16493
rect 14668 16232 14708 16444
rect 14668 16183 14708 16192
rect 14668 15980 14708 15989
rect 14668 15560 14708 15940
rect 14668 15511 14708 15520
rect 14572 14848 14708 14888
rect 14380 14167 14420 14176
rect 14572 14720 14612 14729
rect 14188 13460 14228 13469
rect 14188 13208 14228 13420
rect 14188 13159 14228 13168
rect 14284 13124 14324 13840
rect 14476 14048 14516 14057
rect 14476 13544 14516 14008
rect 14476 13208 14516 13504
rect 14572 13964 14612 14680
rect 14668 14216 14708 14848
rect 14764 14804 14804 16696
rect 14860 14888 14900 19048
rect 14956 18836 14996 19300
rect 14956 18787 14996 18796
rect 15052 19088 15092 19097
rect 14956 18584 14996 18593
rect 14956 14972 14996 18544
rect 14956 14923 14996 14932
rect 14860 14839 14900 14848
rect 14764 14755 14804 14764
rect 15052 14804 15092 19048
rect 15148 19004 15188 19972
rect 15148 17324 15188 18964
rect 15244 19928 15284 20056
rect 15244 19172 15284 19888
rect 15532 20096 15572 20105
rect 15436 19676 15476 19685
rect 15340 19592 15380 19601
rect 15340 19424 15380 19552
rect 15340 19375 15380 19384
rect 15244 18920 15284 19132
rect 15244 18871 15284 18880
rect 15340 19088 15380 19097
rect 15244 18752 15284 18761
rect 15244 18500 15284 18712
rect 15244 18080 15284 18460
rect 15340 18248 15380 19048
rect 15436 18920 15476 19636
rect 15436 18871 15476 18880
rect 15532 19256 15572 20056
rect 15532 19004 15572 19216
rect 15340 18199 15380 18208
rect 15436 18584 15476 18593
rect 15436 18500 15476 18544
rect 15244 18031 15284 18040
rect 15436 18080 15476 18460
rect 15436 18031 15476 18040
rect 15532 17996 15572 18964
rect 15532 17947 15572 17956
rect 15340 17660 15380 17669
rect 15244 17576 15284 17585
rect 15244 17441 15284 17536
rect 15148 17275 15188 17284
rect 15340 17240 15380 17620
rect 15340 17200 15572 17240
rect 15148 17156 15188 17165
rect 15340 17156 15380 17200
rect 15188 17116 15380 17156
rect 15148 17107 15188 17116
rect 15244 16988 15284 16997
rect 15148 16904 15188 16913
rect 15148 16568 15188 16864
rect 15148 15644 15188 16528
rect 15244 16820 15284 16948
rect 15244 16148 15284 16780
rect 15244 16099 15284 16108
rect 15148 15595 15188 15604
rect 15244 15560 15284 15569
rect 15244 15392 15284 15520
rect 15052 14755 15092 14764
rect 15148 15140 15188 15149
rect 15148 14720 15188 15100
rect 15148 14671 15188 14680
rect 14668 14167 14708 14176
rect 14764 14636 14804 14645
rect 14764 14132 14804 14596
rect 15244 14552 15284 15352
rect 15244 14503 15284 14512
rect 14764 14083 14804 14092
rect 14860 14468 14900 14477
rect 14572 13460 14612 13924
rect 14572 13411 14612 13420
rect 14668 14048 14708 14057
rect 14476 13159 14516 13168
rect 14668 13124 14708 14008
rect 14284 13075 14324 13084
rect 14572 13084 14708 13124
rect 14764 13292 14804 13301
rect 14188 13040 14228 13049
rect 14188 12620 14228 13000
rect 14188 12571 14228 12580
rect 14188 11612 14228 11621
rect 14188 11192 14228 11572
rect 14188 10352 14228 11152
rect 14188 10303 14228 10312
rect 14380 11528 14420 11537
rect 14380 11276 14420 11488
rect 14380 10352 14420 11236
rect 14380 10303 14420 10312
rect 14572 9092 14612 13084
rect 14764 11864 14804 13252
rect 14764 11815 14804 11824
rect 14764 11696 14804 11705
rect 14764 10436 14804 11656
rect 14764 10387 14804 10396
rect 14764 10184 14804 10193
rect 14668 10100 14708 10109
rect 14668 9512 14708 10060
rect 14764 9596 14804 10144
rect 14764 9547 14804 9556
rect 14668 9463 14708 9472
rect 14572 9043 14612 9052
rect 14668 9344 14708 9353
rect 14092 8119 14132 8128
rect 14476 8504 14516 8513
rect 14476 8084 14516 8464
rect 13996 7363 14036 7372
rect 14380 8000 14420 8009
rect 14380 7412 14420 7960
rect 14380 7363 14420 7372
rect 13900 6320 13940 7120
rect 14380 7076 14420 7085
rect 14284 6908 14324 6917
rect 13900 6271 13940 6280
rect 13996 6488 14036 6497
rect 13228 5513 13268 5608
rect 13804 5648 13844 5657
rect 13132 5095 13172 5104
rect 13804 5144 13844 5608
rect 13804 5095 13844 5104
rect 13996 5480 14036 6448
rect 13420 5060 13460 5069
rect 13900 5060 13940 5069
rect 13460 5020 13748 5060
rect 13420 5011 13460 5020
rect 13708 4976 13748 5020
rect 13708 4927 13748 4936
rect 13900 4925 13940 5020
rect 13996 4976 14036 5440
rect 13996 4927 14036 4936
rect 14284 5900 14324 6868
rect 14380 6572 14420 7036
rect 14476 6992 14516 8044
rect 14668 8000 14708 9304
rect 14860 8084 14900 14428
rect 14956 14384 14996 14393
rect 14956 12704 14996 14344
rect 15244 14132 15284 14141
rect 14956 12116 14996 12664
rect 14956 12067 14996 12076
rect 15052 13964 15092 13973
rect 14956 11864 14996 11873
rect 14956 11612 14996 11824
rect 14956 11563 14996 11572
rect 15052 11192 15092 13924
rect 15148 13292 15188 13303
rect 15148 13208 15188 13252
rect 15244 13292 15284 14092
rect 15340 14048 15380 17116
rect 15436 17072 15476 17081
rect 15436 16064 15476 17032
rect 15532 16988 15572 17200
rect 15532 16939 15572 16948
rect 15628 16820 15668 21568
rect 15724 21356 15764 21365
rect 15724 20600 15764 21316
rect 15724 20551 15764 20560
rect 15724 20264 15764 20273
rect 15820 20264 15860 22324
rect 16012 22315 16052 22324
rect 16108 24632 16148 24641
rect 16108 23036 16148 24592
rect 16204 24044 16244 25180
rect 16396 25136 16436 25145
rect 16204 23995 16244 24004
rect 16300 24044 16340 24053
rect 16300 23876 16340 24004
rect 16300 23827 16340 23836
rect 16300 23708 16340 23719
rect 16204 23624 16244 23633
rect 16204 23288 16244 23584
rect 16300 23624 16340 23668
rect 16300 23575 16340 23584
rect 16204 23239 16244 23248
rect 16300 23456 16340 23465
rect 16012 22196 16052 22205
rect 16012 21692 16052 22156
rect 16108 21692 16148 22996
rect 16300 22868 16340 23416
rect 16300 22819 16340 22828
rect 16396 22952 16436 25096
rect 16300 22700 16340 22709
rect 16300 22364 16340 22660
rect 16300 22280 16340 22324
rect 16300 22200 16340 22240
rect 16396 22196 16436 22912
rect 16396 22112 16436 22156
rect 16396 22063 16436 22072
rect 16396 21944 16436 21953
rect 16204 21692 16244 21701
rect 16108 21652 16204 21692
rect 16012 21643 16052 21652
rect 16204 21643 16244 21652
rect 16396 21608 16436 21904
rect 16396 21559 16436 21568
rect 16108 21524 16148 21533
rect 15764 20224 15860 20264
rect 15916 21440 15956 21449
rect 15916 20684 15956 21400
rect 15724 19172 15764 20224
rect 15916 20096 15956 20644
rect 16012 20768 16052 20777
rect 16012 20633 16052 20728
rect 15916 20047 15956 20056
rect 16108 20264 16148 21484
rect 15820 20012 15860 20021
rect 15820 19760 15860 19972
rect 15820 19711 15860 19720
rect 16012 20012 16052 20021
rect 15724 19123 15764 19132
rect 15820 19592 15860 19601
rect 15628 16771 15668 16780
rect 15724 18500 15764 18509
rect 15628 16568 15668 16579
rect 15628 16484 15668 16528
rect 15628 16435 15668 16444
rect 15436 15980 15476 16024
rect 15436 15931 15476 15940
rect 15532 16316 15572 16325
rect 15436 15812 15476 15823
rect 15436 15728 15476 15772
rect 15436 15679 15476 15688
rect 15340 13999 15380 14008
rect 15436 14636 15476 14645
rect 15244 13243 15284 13252
rect 15148 13159 15188 13168
rect 15340 13208 15380 13217
rect 15244 13124 15284 13133
rect 15148 13040 15188 13049
rect 15148 12452 15188 13000
rect 15148 12403 15188 12412
rect 15148 11780 15188 11789
rect 15148 11645 15188 11740
rect 15244 11612 15284 13084
rect 15340 12704 15380 13168
rect 15340 12655 15380 12664
rect 15244 11563 15284 11572
rect 15340 12536 15380 12545
rect 15052 11143 15092 11152
rect 15244 10940 15284 10949
rect 15052 10856 15092 10865
rect 15052 8840 15092 10816
rect 15148 10268 15188 10277
rect 15148 10184 15188 10228
rect 15148 10133 15188 10144
rect 15052 8791 15092 8800
rect 15244 10016 15284 10900
rect 14860 8035 14900 8044
rect 14956 8252 14996 8261
rect 14668 7076 14708 7960
rect 14956 8000 14996 8212
rect 14956 7951 14996 7960
rect 15052 8000 15092 8009
rect 14668 7027 14708 7036
rect 14764 7916 14804 7925
rect 14764 7160 14804 7876
rect 15052 7328 15092 7960
rect 15052 7279 15092 7288
rect 15148 7244 15188 7339
rect 15244 7328 15284 9976
rect 15244 7279 15284 7288
rect 15148 7195 15188 7204
rect 14476 6943 14516 6952
rect 14764 6656 14804 7120
rect 14764 6607 14804 6616
rect 15148 7076 15188 7085
rect 15148 6656 15188 7036
rect 15148 6607 15188 6616
rect 14380 6523 14420 6532
rect 14284 4976 14324 5860
rect 15340 5900 15380 12496
rect 15436 11780 15476 14596
rect 15532 12620 15572 16276
rect 15628 16148 15668 16157
rect 15628 15644 15668 16108
rect 15628 15595 15668 15604
rect 15628 14888 15668 14897
rect 15628 13964 15668 14848
rect 15628 13915 15668 13924
rect 15724 13460 15764 18460
rect 15820 17996 15860 19552
rect 16012 19592 16052 19972
rect 16012 19543 16052 19552
rect 15820 17947 15860 17956
rect 15916 19088 15956 19097
rect 15916 18920 15956 19048
rect 15820 17828 15860 17837
rect 15820 16820 15860 17788
rect 15820 16771 15860 16780
rect 15820 16400 15860 16409
rect 15820 14384 15860 16360
rect 15820 14335 15860 14344
rect 15724 13411 15764 13420
rect 15724 13292 15764 13332
rect 15724 13208 15764 13252
rect 15628 13124 15668 13135
rect 15628 13040 15668 13084
rect 15628 12991 15668 13000
rect 15532 12571 15572 12580
rect 15628 12704 15668 12713
rect 15436 11731 15476 11740
rect 15628 9680 15668 12664
rect 15724 12620 15764 13168
rect 15724 12571 15764 12580
rect 15820 12452 15860 12461
rect 15820 12200 15860 12412
rect 15820 11780 15860 12160
rect 15820 11731 15860 11740
rect 15628 9631 15668 9640
rect 15724 10184 15764 10279
rect 15724 9512 15764 10144
rect 15724 9463 15764 9472
rect 15532 8504 15572 8513
rect 15436 8168 15476 8196
rect 15532 8168 15572 8464
rect 15476 8128 15572 8168
rect 15436 8119 15476 8128
rect 15532 8000 15572 8128
rect 15532 7951 15572 7960
rect 15340 5851 15380 5860
rect 15628 6488 15668 6497
rect 14284 4927 14324 4936
rect 15052 5732 15092 5741
rect 13036 4759 13076 4768
rect 15052 4808 15092 5692
rect 15628 5732 15668 6448
rect 15628 5683 15668 5692
rect 15916 5648 15956 18880
rect 16108 18668 16148 20224
rect 16396 20852 16436 20861
rect 16204 20180 16244 20189
rect 16204 20045 16244 20140
rect 16300 19592 16340 19601
rect 16108 18619 16148 18628
rect 16204 19256 16244 19265
rect 16204 18836 16244 19216
rect 16204 18584 16244 18796
rect 16204 18535 16244 18544
rect 16300 19256 16340 19552
rect 16396 19340 16436 20812
rect 16396 19291 16436 19300
rect 16108 18248 16148 18257
rect 16108 18164 16148 18208
rect 16108 18113 16148 18124
rect 16204 17744 16244 17839
rect 16204 17695 16244 17704
rect 16012 17660 16052 17669
rect 16052 17620 16148 17660
rect 16012 17611 16052 17620
rect 16012 17156 16052 17167
rect 16012 17072 16052 17116
rect 16012 17023 16052 17032
rect 16012 16820 16052 16831
rect 16012 16736 16052 16780
rect 16012 16687 16052 16696
rect 16108 16652 16148 17620
rect 16012 16568 16052 16577
rect 16012 15980 16052 16528
rect 16108 16316 16148 16612
rect 16108 16267 16148 16276
rect 16204 17492 16244 17501
rect 16108 16148 16148 16157
rect 16108 16013 16148 16108
rect 16012 15931 16052 15940
rect 16204 15896 16244 17452
rect 16204 15847 16244 15856
rect 16300 16988 16340 19216
rect 16396 19088 16436 19099
rect 16396 19004 16436 19048
rect 16396 18955 16436 18964
rect 16300 15644 16340 16948
rect 16396 17576 16436 17585
rect 16396 16232 16436 17536
rect 16492 17156 16532 28540
rect 19468 28412 19508 28421
rect 17164 28244 17204 28253
rect 16684 27656 16724 27665
rect 16588 26648 16628 26657
rect 16588 26513 16628 26608
rect 16588 26228 16628 26237
rect 16588 24632 16628 26188
rect 16684 25136 16724 27616
rect 16876 27572 16916 27581
rect 16876 27437 16916 27532
rect 16876 27152 16916 27161
rect 16780 26900 16820 26909
rect 16780 26816 16820 26860
rect 16780 26765 16820 26776
rect 16876 26144 16916 27112
rect 16876 26095 16916 26104
rect 17164 26228 17204 28204
rect 19468 27824 19508 28372
rect 23116 28244 23156 28600
rect 23884 28328 23924 28600
rect 24652 28496 24692 28600
rect 24652 28447 24692 28456
rect 23884 28279 23924 28288
rect 23116 28195 23156 28204
rect 23788 28160 23828 28169
rect 19900 27992 20268 28001
rect 19900 27943 20268 27952
rect 19468 27775 19508 27784
rect 18028 27740 18068 27749
rect 17932 27236 17972 27245
rect 17260 26900 17300 26909
rect 17260 26816 17300 26860
rect 17548 26816 17588 26825
rect 17260 26776 17548 26816
rect 17548 26767 17588 26776
rect 17644 26732 17684 26741
rect 17356 26648 17396 26657
rect 16780 25892 16820 25901
rect 16780 25472 16820 25852
rect 16780 25304 16820 25432
rect 16780 25255 16820 25264
rect 16972 25304 17012 25313
rect 16684 25087 16724 25096
rect 16972 25136 17012 25264
rect 16972 25087 17012 25096
rect 16588 19592 16628 24592
rect 16684 24968 16724 24977
rect 16684 23876 16724 24928
rect 16684 23288 16724 23836
rect 16684 23239 16724 23248
rect 16780 24884 16820 24893
rect 16780 23060 16820 24844
rect 17164 24884 17204 26188
rect 17260 26564 17300 26573
rect 17260 25388 17300 26524
rect 17356 26144 17396 26608
rect 17356 26095 17396 26104
rect 17644 26060 17684 26692
rect 17260 25348 17396 25388
rect 17164 24835 17204 24844
rect 17164 24716 17204 24725
rect 17164 24632 17204 24676
rect 17356 24632 17396 25348
rect 17644 25136 17684 26020
rect 17740 26228 17780 26237
rect 17740 25808 17780 26188
rect 17740 25759 17780 25768
rect 17836 26060 17876 26069
rect 17836 25556 17876 26020
rect 17836 25507 17876 25516
rect 17644 25087 17684 25096
rect 17740 24632 17780 24643
rect 17356 24592 17492 24632
rect 17164 24581 17204 24592
rect 17356 24464 17396 24473
rect 17356 24128 17396 24424
rect 16876 23876 16916 23887
rect 16876 23792 16916 23836
rect 16876 23743 16916 23752
rect 17356 23792 17396 24088
rect 17356 23743 17396 23752
rect 16972 23708 17012 23717
rect 16972 23573 17012 23668
rect 17452 23708 17492 24592
rect 17740 24548 17780 24592
rect 17740 24499 17780 24508
rect 17452 23659 17492 23668
rect 17644 23792 17684 23801
rect 16684 23020 16820 23060
rect 16876 23540 16916 23549
rect 16684 22364 16724 23020
rect 16684 22315 16724 22324
rect 16780 22280 16820 22289
rect 16684 21524 16724 21533
rect 16684 20852 16724 21484
rect 16780 21020 16820 22240
rect 16876 21776 16916 23500
rect 17452 23372 17492 23381
rect 17356 23288 17396 23297
rect 17164 23204 17204 23213
rect 17164 23060 17204 23164
rect 17356 23153 17396 23248
rect 17452 23120 17492 23332
rect 17452 23071 17492 23080
rect 16972 23036 17204 23060
rect 16972 23020 17164 23036
rect 16972 22364 17012 23020
rect 17164 22987 17204 22996
rect 17548 22868 17588 22877
rect 16972 21944 17012 22324
rect 17452 22448 17492 22457
rect 17164 22280 17204 22289
rect 17164 22145 17204 22240
rect 16972 21895 17012 21904
rect 17260 22028 17300 22037
rect 17068 21860 17108 21869
rect 16876 21524 16916 21736
rect 16972 21692 17012 21787
rect 16972 21643 17012 21652
rect 17068 21608 17108 21820
rect 17068 21559 17108 21568
rect 16876 21475 16916 21484
rect 16780 20971 16820 20980
rect 16876 21356 16916 21365
rect 16684 20768 16724 20812
rect 16684 20717 16724 20728
rect 16780 20852 16820 20861
rect 16588 19543 16628 19552
rect 16684 20012 16724 20021
rect 16684 19508 16724 19972
rect 16684 19459 16724 19468
rect 16588 19256 16628 19265
rect 16588 18668 16628 19216
rect 16780 19256 16820 20812
rect 16876 20264 16916 21316
rect 17068 21356 17108 21365
rect 16972 21188 17012 21197
rect 16972 20768 17012 21148
rect 16972 20719 17012 20728
rect 17068 20432 17108 21316
rect 17260 21188 17300 21988
rect 17452 21860 17492 22408
rect 17548 22364 17588 22828
rect 17548 22315 17588 22324
rect 17644 22196 17684 23752
rect 17836 23540 17876 23549
rect 17836 23120 17876 23500
rect 17836 22985 17876 23080
rect 17644 22156 17780 22196
rect 17452 21811 17492 21820
rect 17260 21139 17300 21148
rect 17356 21692 17396 21701
rect 17260 20852 17300 20861
rect 17068 20383 17108 20392
rect 17164 20600 17204 20609
rect 16876 20215 16916 20224
rect 16972 20180 17012 20189
rect 16876 19844 16916 19853
rect 16876 19709 16916 19804
rect 16780 19207 16820 19216
rect 16876 19508 16916 19517
rect 16684 19172 16724 19181
rect 16684 19004 16724 19132
rect 16684 18955 16724 18964
rect 16876 18752 16916 19468
rect 16588 18500 16628 18628
rect 16780 18712 16916 18752
rect 16972 18752 17012 20140
rect 16588 18451 16628 18460
rect 16684 18500 16724 18509
rect 16684 18248 16724 18460
rect 16492 17107 16532 17116
rect 16588 17744 16628 17753
rect 16492 16988 16532 16999
rect 16492 16904 16532 16948
rect 16492 16855 16532 16864
rect 16396 16192 16532 16232
rect 16492 16148 16532 16192
rect 16492 16099 16532 16108
rect 16300 15056 16340 15604
rect 16492 15980 16532 15989
rect 16492 15392 16532 15940
rect 16492 15343 16532 15352
rect 16396 15308 16436 15317
rect 16396 15224 16436 15268
rect 16396 15173 16436 15184
rect 16300 15007 16340 15016
rect 16108 14720 16148 14729
rect 16012 14132 16052 14141
rect 16012 13997 16052 14092
rect 16012 13880 16052 13889
rect 16012 13628 16052 13840
rect 16012 13579 16052 13588
rect 16012 13124 16052 13133
rect 16012 12704 16052 13084
rect 16108 12788 16148 14680
rect 16396 14720 16436 14729
rect 16300 14552 16340 14561
rect 16204 14512 16300 14552
rect 16204 13292 16244 14512
rect 16300 14503 16340 14512
rect 16204 13243 16244 13252
rect 16300 14216 16340 14225
rect 16300 13292 16340 14176
rect 16396 14048 16436 14680
rect 16588 14636 16628 17704
rect 16684 17576 16724 18208
rect 16780 18080 16820 18712
rect 16972 18703 17012 18712
rect 17068 19172 17108 19181
rect 17068 18584 17108 19132
rect 17164 18668 17204 20560
rect 17260 20516 17300 20812
rect 17260 20467 17300 20476
rect 17260 20264 17300 20273
rect 17260 20096 17300 20224
rect 17260 19340 17300 20056
rect 17356 19928 17396 21652
rect 17645 21608 17685 21617
rect 17644 21568 17645 21608
rect 17644 21559 17685 21568
rect 17548 21524 17588 21533
rect 17452 20936 17492 20945
rect 17452 20768 17492 20896
rect 17452 20684 17492 20728
rect 17452 20604 17492 20644
rect 17356 19879 17396 19888
rect 17452 20180 17492 20189
rect 17260 19291 17300 19300
rect 17356 19172 17396 19181
rect 17260 18668 17300 18677
rect 17164 18628 17260 18668
rect 17260 18619 17300 18628
rect 17068 18544 17204 18584
rect 16780 17744 16820 18040
rect 16780 17695 16820 17704
rect 16876 18500 16916 18509
rect 16684 17527 16724 17536
rect 16876 17240 16916 18460
rect 16876 17191 16916 17200
rect 16972 18500 17012 18509
rect 16780 17156 16820 17165
rect 16684 16484 16724 16493
rect 16684 16316 16724 16444
rect 16684 14804 16724 16276
rect 16780 15560 16820 17116
rect 16972 16988 17012 18460
rect 16876 16820 16916 16829
rect 16876 16232 16916 16780
rect 16876 16183 16916 16192
rect 16972 16064 17012 16948
rect 16972 16015 17012 16024
rect 17068 18332 17108 18341
rect 17164 18332 17204 18544
rect 17260 18332 17300 18341
rect 17164 18292 17260 18332
rect 16780 15511 16820 15520
rect 16876 15980 16916 15989
rect 16684 14755 16724 14764
rect 16588 14587 16628 14596
rect 16396 13999 16436 14008
rect 16684 14552 16724 14561
rect 16300 13243 16340 13252
rect 16108 12739 16148 12748
rect 16300 13124 16340 13133
rect 16012 12655 16052 12664
rect 16300 12704 16340 13084
rect 16300 12655 16340 12664
rect 16396 13040 16436 13049
rect 16396 12620 16436 13000
rect 16396 12571 16436 12580
rect 16588 12872 16628 12881
rect 16588 12536 16628 12832
rect 16588 12487 16628 12496
rect 16108 12368 16148 12377
rect 16012 10100 16052 10109
rect 16012 9512 16052 10060
rect 16108 9848 16148 12328
rect 16684 11864 16724 14512
rect 16684 11815 16724 11824
rect 16780 14048 16820 14057
rect 16780 13964 16820 14008
rect 16300 11696 16340 11705
rect 16204 11108 16244 11117
rect 16204 10184 16244 11068
rect 16300 10436 16340 11656
rect 16780 11192 16820 13924
rect 16876 13712 16916 15940
rect 16876 13663 16916 13672
rect 16972 14636 17012 14645
rect 16876 13292 16916 13301
rect 16876 12704 16916 13252
rect 16876 12655 16916 12664
rect 16972 12536 17012 14596
rect 17068 13208 17108 18292
rect 17164 18080 17204 18089
rect 17164 16988 17204 18040
rect 17164 16939 17204 16948
rect 17260 16568 17300 18292
rect 17260 16519 17300 16528
rect 17260 16316 17300 16325
rect 17260 15728 17300 16276
rect 17260 15679 17300 15688
rect 17260 15560 17300 15569
rect 17068 13159 17108 13168
rect 17164 15392 17204 15401
rect 16972 12487 17012 12496
rect 17068 12788 17108 12797
rect 17068 12452 17108 12748
rect 17068 12200 17108 12412
rect 17068 12151 17108 12160
rect 16780 11143 16820 11152
rect 16972 12116 17012 12125
rect 16396 11024 16436 11033
rect 16396 10520 16436 10984
rect 16396 10471 16436 10480
rect 16780 11024 16820 11033
rect 16300 10387 16340 10396
rect 16204 10135 16244 10144
rect 16492 10184 16532 10193
rect 16108 9799 16148 9808
rect 16300 10016 16340 10025
rect 16012 9463 16052 9472
rect 16204 9596 16244 9605
rect 16204 9512 16244 9556
rect 16204 8672 16244 9472
rect 16204 8623 16244 8632
rect 16012 7160 16052 7169
rect 16012 6488 16052 7120
rect 16204 7160 16244 7169
rect 16204 6656 16244 7120
rect 16204 6607 16244 6616
rect 16012 6439 16052 6448
rect 15916 5599 15956 5608
rect 16300 5060 16340 9976
rect 16396 9512 16436 9521
rect 16396 8168 16436 9472
rect 16396 8119 16436 8128
rect 16492 8756 16532 10144
rect 16300 5011 16340 5020
rect 16492 5564 16532 8716
rect 16780 6656 16820 10984
rect 16972 11024 17012 12076
rect 17164 11780 17204 15352
rect 17260 14720 17300 15520
rect 17260 14671 17300 14680
rect 17164 11731 17204 11740
rect 17260 14552 17300 14561
rect 17260 12536 17300 14512
rect 17356 13124 17396 19132
rect 17452 16484 17492 20140
rect 17548 19844 17588 21484
rect 17548 19795 17588 19804
rect 17644 19760 17684 21559
rect 17740 21272 17780 22156
rect 17740 21223 17780 21232
rect 17836 21524 17876 21533
rect 17836 21020 17876 21484
rect 17836 20971 17876 20980
rect 17932 21440 17972 27196
rect 18028 26816 18068 27700
rect 23788 27740 23828 28120
rect 25420 27824 25460 28600
rect 25420 27775 25460 27784
rect 23788 27691 23828 27700
rect 24172 27740 24212 27749
rect 19660 27656 19700 27665
rect 19564 27488 19604 27497
rect 18316 27404 18356 27413
rect 18028 26767 18068 26776
rect 18220 26984 18260 26993
rect 18220 26900 18260 26944
rect 18028 26144 18068 26153
rect 18028 26060 18068 26104
rect 18028 25220 18068 26020
rect 18220 25556 18260 26860
rect 18316 26732 18356 27364
rect 18660 27236 19028 27245
rect 18660 27187 19028 27196
rect 19276 27152 19316 27161
rect 18316 26228 18356 26692
rect 18316 26179 18356 26188
rect 18412 27068 18452 27077
rect 18220 25507 18260 25516
rect 18316 26060 18356 26069
rect 18028 25085 18068 25180
rect 18220 25220 18260 25229
rect 18124 24800 18164 24809
rect 18124 24665 18164 24760
rect 18220 24632 18260 25180
rect 18316 24800 18356 26020
rect 18316 24751 18356 24760
rect 18220 24583 18260 24592
rect 18316 23960 18356 23969
rect 18124 23876 18164 23885
rect 18124 23288 18164 23836
rect 18316 23792 18356 23920
rect 18316 23456 18356 23752
rect 18316 23407 18356 23416
rect 18124 23239 18164 23248
rect 18316 23036 18356 23045
rect 18220 22868 18260 22877
rect 17836 20852 17876 20861
rect 17644 19711 17684 19720
rect 17740 20768 17780 20777
rect 17548 19508 17588 19517
rect 17548 18920 17588 19468
rect 17644 19256 17684 19265
rect 17740 19256 17780 20728
rect 17836 20264 17876 20812
rect 17932 20600 17972 21400
rect 18028 21524 18068 21533
rect 18028 21389 18068 21484
rect 18124 21356 18164 21365
rect 18124 21020 18164 21316
rect 18124 20971 18164 20980
rect 17932 20551 17972 20560
rect 18028 20768 18068 20777
rect 17836 20215 17876 20224
rect 18028 20516 18068 20728
rect 18124 20600 18164 20695
rect 18124 20551 18164 20560
rect 17932 20180 17972 20220
rect 17932 20096 17972 20140
rect 17932 20047 17972 20056
rect 18028 20012 18068 20476
rect 18220 20180 18260 22828
rect 18316 22616 18356 22996
rect 18316 22567 18356 22576
rect 18412 22280 18452 27028
rect 18796 26900 18836 26909
rect 18604 26732 18644 26741
rect 18604 26312 18644 26692
rect 18604 26263 18644 26272
rect 18796 26060 18836 26860
rect 18796 26011 18836 26020
rect 18892 26816 18932 26825
rect 18892 26648 18932 26776
rect 18892 25976 18932 26608
rect 19084 26564 19124 26575
rect 18988 26480 19028 26489
rect 18988 26144 19028 26440
rect 19084 26480 19124 26524
rect 19084 26431 19124 26440
rect 18988 26095 19028 26104
rect 19084 26312 19124 26321
rect 18892 25927 18932 25936
rect 18508 25892 18548 25901
rect 18508 25304 18548 25852
rect 18660 25724 19028 25733
rect 18660 25675 19028 25684
rect 18988 25472 19028 25481
rect 18508 25255 18548 25264
rect 18604 25388 18644 25397
rect 18508 24800 18548 24809
rect 18508 24632 18548 24760
rect 18508 24583 18548 24592
rect 18508 24464 18548 24473
rect 18604 24464 18644 25348
rect 18988 25337 19028 25432
rect 18796 25136 18836 25145
rect 18796 25001 18836 25096
rect 19084 25136 19124 26272
rect 19276 26144 19316 27112
rect 19180 25304 19220 25313
rect 19276 25304 19316 26104
rect 19372 26900 19412 26909
rect 19372 25388 19412 26860
rect 19564 26900 19604 27448
rect 19564 26816 19604 26860
rect 19564 26765 19604 26776
rect 19660 26900 19700 27616
rect 21868 27656 21908 27665
rect 21772 27572 21812 27581
rect 20428 27320 20468 27329
rect 19660 26816 19700 26860
rect 19660 26767 19700 26776
rect 19756 27152 19796 27161
rect 19756 26648 19796 27112
rect 20236 26816 20276 26911
rect 20236 26767 20276 26776
rect 20428 26732 20468 27280
rect 21388 27152 21428 27161
rect 19660 26608 19796 26648
rect 20236 26648 20276 26657
rect 20276 26608 20372 26648
rect 19372 25339 19412 25348
rect 19468 26480 19508 26489
rect 19220 25264 19316 25304
rect 19468 25304 19508 26440
rect 19660 25976 19700 26608
rect 20236 26599 20276 26608
rect 19900 26480 20268 26489
rect 19900 26431 20268 26440
rect 19948 26312 19988 26321
rect 19660 25927 19700 25936
rect 19756 26060 19796 26069
rect 19564 25724 19604 25733
rect 19564 25556 19604 25684
rect 19564 25507 19604 25516
rect 19660 25556 19700 25565
rect 19660 25388 19700 25516
rect 19660 25339 19700 25348
rect 19180 25255 19220 25264
rect 19468 25255 19508 25264
rect 19084 25087 19124 25096
rect 19564 25220 19604 25229
rect 19564 25085 19604 25180
rect 19276 25052 19316 25061
rect 19180 25012 19276 25052
rect 18796 24800 18836 24809
rect 18700 24632 18740 24643
rect 18700 24548 18740 24592
rect 18700 24499 18740 24508
rect 18548 24424 18644 24464
rect 18508 23960 18548 24424
rect 18796 24380 18836 24760
rect 18988 24632 19028 24641
rect 19180 24632 19220 25012
rect 19276 25003 19316 25012
rect 19028 24592 19220 24632
rect 19276 24884 19316 24893
rect 19276 24632 19316 24844
rect 19468 24800 19508 24809
rect 19468 24665 19508 24760
rect 19756 24716 19796 26020
rect 19852 25640 19892 25649
rect 19852 25388 19892 25600
rect 19948 25556 19988 26272
rect 20236 26144 20276 26153
rect 20332 26144 20372 26608
rect 20276 26104 20372 26144
rect 20236 26095 20276 26104
rect 19948 25507 19988 25516
rect 20044 25976 20084 25985
rect 19852 25339 19892 25348
rect 20044 25220 20084 25936
rect 20140 25892 20180 25901
rect 20140 25724 20180 25852
rect 20140 25675 20180 25684
rect 20140 25556 20180 25567
rect 20140 25472 20180 25516
rect 20140 25423 20180 25432
rect 20044 25171 20084 25180
rect 20140 25304 20180 25315
rect 20140 25220 20180 25264
rect 20140 25171 20180 25180
rect 19900 24968 20268 24977
rect 19900 24919 20268 24928
rect 18988 24583 19028 24592
rect 19276 24583 19316 24592
rect 18796 24331 18836 24340
rect 19564 24464 19604 24473
rect 18660 24212 19028 24221
rect 18660 24163 19028 24172
rect 18508 23911 18548 23920
rect 19084 23960 19124 23969
rect 18892 23792 18932 23801
rect 18412 22231 18452 22240
rect 18508 23624 18548 23633
rect 18412 22112 18452 22121
rect 18412 21608 18452 22072
rect 18412 20936 18452 21568
rect 18412 20887 18452 20896
rect 18412 20768 18452 20779
rect 18220 20131 18260 20140
rect 18316 20684 18356 20693
rect 18316 20096 18356 20644
rect 18412 20684 18452 20728
rect 18412 20635 18452 20644
rect 18316 20047 18356 20056
rect 18028 19963 18068 19972
rect 17932 19760 17972 19769
rect 17932 19340 17972 19720
rect 17932 19291 17972 19300
rect 17836 19256 17876 19265
rect 17740 19216 17836 19256
rect 17644 19172 17684 19216
rect 17644 19121 17684 19132
rect 17836 19004 17876 19216
rect 17836 18955 17876 18964
rect 18124 19256 18164 19265
rect 17548 18871 17588 18880
rect 17644 18500 17684 18509
rect 17452 16435 17492 16444
rect 17548 17996 17588 18005
rect 17548 16484 17588 17956
rect 17548 16435 17588 16444
rect 17644 17660 17684 18460
rect 17644 16316 17684 17620
rect 17452 16232 17492 16241
rect 17452 15392 17492 16192
rect 17548 16148 17588 16157
rect 17548 16013 17588 16108
rect 17644 15476 17684 16276
rect 17644 15427 17684 15436
rect 17740 18080 17780 18089
rect 17740 17072 17780 18040
rect 17836 17828 17876 17837
rect 17836 17156 17876 17788
rect 18028 17828 18068 17837
rect 17932 17744 17972 17753
rect 17932 17660 17972 17704
rect 18028 17693 18068 17788
rect 17932 17609 17972 17620
rect 17836 17107 17876 17116
rect 17740 16904 17780 17032
rect 17452 15343 17492 15352
rect 17452 15224 17492 15233
rect 17452 14720 17492 15184
rect 17452 14671 17492 14680
rect 17644 14552 17684 14561
rect 17644 14048 17684 14512
rect 17740 14216 17780 16864
rect 17932 16820 17972 16829
rect 17836 16232 17876 16241
rect 17836 15812 17876 16192
rect 17836 15763 17876 15772
rect 17932 15644 17972 16780
rect 17932 15595 17972 15604
rect 18028 15980 18068 15989
rect 17932 15476 17972 15485
rect 17932 14972 17972 15436
rect 17932 14923 17972 14932
rect 18028 15392 18068 15940
rect 18028 14384 18068 15352
rect 18124 14972 18164 19216
rect 18124 14923 18164 14932
rect 18220 19172 18260 19181
rect 18220 17156 18260 19132
rect 18220 15644 18260 17116
rect 18412 19004 18452 19013
rect 18412 15812 18452 18964
rect 18412 15763 18452 15772
rect 18508 16232 18548 23584
rect 18604 23372 18644 23381
rect 18604 23120 18644 23332
rect 18892 23204 18932 23752
rect 19084 23792 19124 23920
rect 19084 23743 19124 23752
rect 18892 23155 18932 23164
rect 19372 23540 19412 23549
rect 18604 22985 18644 23080
rect 19084 22868 19124 22877
rect 18660 22700 19028 22709
rect 18660 22651 19028 22660
rect 19084 22196 19124 22828
rect 19084 22147 19124 22156
rect 19180 22280 19220 22289
rect 18892 22028 18932 22037
rect 18892 21692 18932 21988
rect 18892 21643 18932 21652
rect 19084 22028 19124 22037
rect 19084 21524 19124 21988
rect 18660 21188 19028 21197
rect 18660 21139 19028 21148
rect 18604 20852 18644 20861
rect 18604 20264 18644 20812
rect 18988 20600 19028 20609
rect 18988 20432 19028 20560
rect 18988 20383 19028 20392
rect 18604 20215 18644 20224
rect 18700 20012 18740 20021
rect 18700 19877 18740 19972
rect 19084 20012 19124 21484
rect 19084 19963 19124 19972
rect 19084 19844 19124 19853
rect 18660 19676 19028 19685
rect 18660 19627 19028 19636
rect 18988 19424 19028 19433
rect 18988 19256 19028 19384
rect 18988 19207 19028 19216
rect 18700 19172 18740 19181
rect 18604 18920 18644 18929
rect 18604 18752 18644 18880
rect 18604 18703 18644 18712
rect 18700 18752 18740 19132
rect 18700 18332 18740 18712
rect 18988 18836 19028 18847
rect 18988 18752 19028 18796
rect 18988 18703 19028 18712
rect 18796 18668 18836 18677
rect 18796 18584 18836 18628
rect 18988 18584 19028 18593
rect 18796 18544 18988 18584
rect 18988 18535 19028 18544
rect 18700 18283 18740 18292
rect 18660 18164 19028 18173
rect 18660 18115 19028 18124
rect 18892 17828 18932 17837
rect 18700 17492 18740 17501
rect 18700 17072 18740 17452
rect 18700 17023 18740 17032
rect 18892 17072 18932 17788
rect 18892 17023 18932 17032
rect 18988 17744 19028 17753
rect 18988 16820 19028 17704
rect 18988 16771 19028 16780
rect 18660 16652 19028 16661
rect 18660 16603 19028 16612
rect 19084 16232 19124 19804
rect 19180 18668 19220 22240
rect 19276 21860 19316 21869
rect 19276 21440 19316 21820
rect 19276 21391 19316 21400
rect 19276 20600 19316 20609
rect 19276 20180 19316 20560
rect 19276 20131 19316 20140
rect 19180 18619 19220 18628
rect 19276 19928 19316 19937
rect 18220 14636 18260 15604
rect 18316 15728 18356 15737
rect 18316 14972 18356 15688
rect 18316 14923 18356 14932
rect 18412 15476 18452 15485
rect 18412 15308 18452 15436
rect 18220 14587 18260 14596
rect 18316 14804 18356 14813
rect 18028 14335 18068 14344
rect 17740 14176 18068 14216
rect 17644 13999 17684 14008
rect 17740 14048 17780 14057
rect 17740 13964 17780 14008
rect 17740 13913 17780 13924
rect 17644 13880 17684 13889
rect 17356 13075 17396 13084
rect 17548 13208 17588 13217
rect 17260 11444 17300 12496
rect 17452 12620 17492 12629
rect 17452 11864 17492 12580
rect 17548 11948 17588 13168
rect 17644 12704 17684 13840
rect 17644 12655 17684 12664
rect 17836 13124 17876 13133
rect 17836 12620 17876 13084
rect 17836 12571 17876 12580
rect 17548 11899 17588 11908
rect 17452 11815 17492 11824
rect 17740 11696 17780 11705
rect 17260 11395 17300 11404
rect 17452 11612 17492 11621
rect 17452 11192 17492 11572
rect 17740 11276 17780 11656
rect 17740 11227 17780 11236
rect 17932 11612 17972 11621
rect 17452 11143 17492 11152
rect 16972 10184 17012 10984
rect 17548 11024 17588 11033
rect 16972 10135 17012 10144
rect 17260 10184 17300 10193
rect 17260 9596 17300 10144
rect 17548 10184 17588 10984
rect 17548 10135 17588 10144
rect 17932 9680 17972 11572
rect 17932 9631 17972 9640
rect 17260 9547 17300 9556
rect 17836 9512 17876 9521
rect 17644 9472 17836 9512
rect 17356 9428 17396 9437
rect 17260 9260 17300 9269
rect 17260 8756 17300 9220
rect 17260 8707 17300 8716
rect 16780 6607 16820 6616
rect 17356 8000 17396 9388
rect 17644 9428 17684 9472
rect 17836 9463 17876 9472
rect 17644 9379 17684 9388
rect 17548 9344 17588 9353
rect 17548 8756 17588 9304
rect 17548 8707 17588 8716
rect 18028 8672 18068 14176
rect 18220 14048 18260 14057
rect 18124 12872 18164 12881
rect 18124 12368 18164 12832
rect 18124 12319 18164 12328
rect 18124 11024 18164 11033
rect 18124 10772 18164 10984
rect 18124 10723 18164 10732
rect 18220 10268 18260 14008
rect 18316 13376 18356 14764
rect 18412 14048 18452 15268
rect 18412 13913 18452 14008
rect 18412 13712 18452 13721
rect 18412 13577 18452 13672
rect 18316 13327 18356 13336
rect 18508 11696 18548 16192
rect 18892 16192 19124 16232
rect 19180 17576 19220 17585
rect 19180 17072 19220 17536
rect 18604 16064 18644 16073
rect 18604 15476 18644 16024
rect 18604 15427 18644 15436
rect 18700 15560 18740 15569
rect 18700 15425 18740 15520
rect 18892 15476 18932 16192
rect 19180 15644 19220 17032
rect 19276 15644 19316 19888
rect 19372 16484 19412 23500
rect 19468 23456 19508 23465
rect 19468 23288 19508 23416
rect 19468 23239 19508 23248
rect 19564 23204 19604 24424
rect 19756 24212 19796 24676
rect 20140 24716 20180 24725
rect 20140 24581 20180 24676
rect 19756 24163 19796 24172
rect 20332 24548 20372 24557
rect 20332 24380 20372 24508
rect 19852 24044 19892 24053
rect 19564 23155 19604 23164
rect 19660 23960 19700 23969
rect 19660 23120 19700 23920
rect 19852 23792 19892 24004
rect 19852 23743 19892 23752
rect 20236 23792 20276 23801
rect 19660 23071 19700 23080
rect 19756 23708 19796 23717
rect 19756 23060 19796 23668
rect 20236 23624 20276 23752
rect 20236 23575 20276 23584
rect 19900 23456 20268 23465
rect 19900 23407 20268 23416
rect 20236 23288 20276 23297
rect 19564 23036 19604 23045
rect 19756 23020 19892 23060
rect 19564 22901 19604 22996
rect 19852 22868 19892 23020
rect 19852 22819 19892 22828
rect 19468 22532 19508 22541
rect 19468 20180 19508 22492
rect 19564 22280 19604 22289
rect 19564 21692 19604 22240
rect 20236 22196 20276 23248
rect 20236 22147 20276 22156
rect 19900 21944 20268 21953
rect 19900 21895 20268 21904
rect 19564 21643 19604 21652
rect 19852 21776 19892 21785
rect 19852 21608 19892 21736
rect 20140 21776 20180 21785
rect 20140 21641 20180 21736
rect 19852 21104 19892 21568
rect 19852 21055 19892 21064
rect 20332 20936 20372 24340
rect 20428 21692 20468 26692
rect 20812 26816 20852 26825
rect 20428 21643 20468 21652
rect 20524 26480 20564 26489
rect 20524 23204 20564 26440
rect 20716 26060 20756 26069
rect 20620 25892 20660 25901
rect 20620 25220 20660 25852
rect 20716 25388 20756 26020
rect 20716 25339 20756 25348
rect 20620 25180 20756 25220
rect 19564 20684 19604 20693
rect 19564 20264 19604 20644
rect 19756 20684 19796 20693
rect 19564 20215 19604 20224
rect 19660 20432 19700 20441
rect 19468 20131 19508 20140
rect 19564 20012 19604 20021
rect 19468 19004 19508 19013
rect 19468 17744 19508 18964
rect 19468 17072 19508 17704
rect 19564 18836 19604 19972
rect 19564 17240 19604 18796
rect 19564 17191 19604 17200
rect 19468 16904 19508 17032
rect 19468 16855 19508 16864
rect 19564 16988 19604 16997
rect 19412 16444 19508 16484
rect 19372 16435 19412 16444
rect 19372 16316 19412 16325
rect 19372 16181 19412 16276
rect 19372 15644 19412 15653
rect 19276 15604 19372 15644
rect 19180 15595 19220 15604
rect 19372 15595 19412 15604
rect 18892 15427 18932 15436
rect 19084 15560 19124 15569
rect 18660 15140 19028 15149
rect 18660 15091 19028 15100
rect 18988 14972 19028 14981
rect 18796 14804 18836 14813
rect 18604 14720 18644 14729
rect 18604 14585 18644 14680
rect 18796 14552 18836 14764
rect 18796 14503 18836 14512
rect 18892 14636 18932 14647
rect 18892 14552 18932 14596
rect 18892 14503 18932 14512
rect 18892 14384 18932 14393
rect 18700 14132 18740 14141
rect 18700 13964 18740 14092
rect 18700 13915 18740 13924
rect 18796 14048 18836 14057
rect 18796 13796 18836 14008
rect 18892 13796 18932 14344
rect 18988 14132 19028 14932
rect 19084 14972 19124 15520
rect 19084 14923 19124 14932
rect 19180 15392 19220 15401
rect 19180 14720 19220 15352
rect 19180 14671 19220 14680
rect 19276 15308 19316 15317
rect 19084 14636 19124 14645
rect 19084 14216 19124 14596
rect 19180 14216 19220 14225
rect 19084 14176 19180 14216
rect 19180 14167 19220 14176
rect 18988 14092 19124 14132
rect 18988 13796 19028 13805
rect 18892 13756 18988 13796
rect 18796 13747 18836 13756
rect 18988 13747 19028 13756
rect 19084 13712 19124 14092
rect 19180 13712 19220 13721
rect 19084 13672 19180 13712
rect 18660 13628 19028 13637
rect 18660 13579 19028 13588
rect 18892 13460 18932 13469
rect 18700 13376 18740 13385
rect 18700 13241 18740 13336
rect 18796 13208 18836 13217
rect 18796 12956 18836 13168
rect 18796 12907 18836 12916
rect 18700 12536 18740 12545
rect 18700 12452 18740 12496
rect 18892 12536 18932 13420
rect 18892 12487 18932 12496
rect 18700 12401 18740 12412
rect 19084 12452 19124 13672
rect 19180 13663 19220 13672
rect 19276 13460 19316 15268
rect 19468 15056 19508 16444
rect 19564 15980 19604 16948
rect 19564 15308 19604 15940
rect 19564 15259 19604 15268
rect 19276 13411 19316 13420
rect 19372 15016 19508 15056
rect 19564 15056 19604 15065
rect 19372 13208 19412 15016
rect 19468 14888 19508 14897
rect 19468 14753 19508 14848
rect 19468 14636 19508 14645
rect 19468 14216 19508 14596
rect 19468 14167 19508 14176
rect 19468 14006 19508 14015
rect 19468 13628 19508 13966
rect 19468 13460 19508 13588
rect 19468 13411 19508 13420
rect 19276 13168 19412 13208
rect 19468 13292 19508 13301
rect 19276 13124 19316 13168
rect 19468 13124 19508 13252
rect 18660 12116 19028 12125
rect 18660 12067 19028 12076
rect 18892 11780 18932 11791
rect 18508 11647 18548 11656
rect 18700 11696 18740 11705
rect 18892 11696 18932 11740
rect 18700 11192 18740 11656
rect 18700 11143 18740 11152
rect 18796 11656 18892 11696
rect 18796 11108 18836 11656
rect 18892 11647 18932 11656
rect 18796 11059 18836 11068
rect 18660 10604 19028 10613
rect 18660 10555 19028 10564
rect 18316 10436 18356 10445
rect 18316 10301 18356 10396
rect 18988 10436 19028 10445
rect 18892 10268 18932 10277
rect 18220 9512 18260 10228
rect 18700 10228 18892 10268
rect 18028 8252 18068 8632
rect 18124 9472 18260 9512
rect 18412 9680 18452 9689
rect 18124 8504 18164 9472
rect 18412 8840 18452 9640
rect 18700 9428 18740 10228
rect 18892 10219 18932 10228
rect 18700 9379 18740 9388
rect 18892 10100 18932 10109
rect 18892 9344 18932 10060
rect 18988 9428 19028 10396
rect 19084 10184 19124 12412
rect 19180 13084 19316 13124
rect 19372 13084 19508 13124
rect 19180 11024 19220 13084
rect 19372 12704 19412 13084
rect 19372 12655 19412 12664
rect 19468 12956 19508 12965
rect 19372 12536 19412 12545
rect 19276 12032 19316 12041
rect 19276 11948 19316 11992
rect 19276 11897 19316 11908
rect 19180 10975 19220 10984
rect 19276 11696 19316 11705
rect 19084 10135 19124 10144
rect 19180 10856 19220 10865
rect 18988 9379 19028 9388
rect 18892 9295 18932 9304
rect 18412 8791 18452 8800
rect 18508 9260 18548 9269
rect 18508 8756 18548 9220
rect 18660 9092 19028 9101
rect 18660 9043 19028 9052
rect 18604 8756 18644 8765
rect 18508 8716 18604 8756
rect 18604 8707 18644 8716
rect 18124 8455 18164 8464
rect 18028 8084 18068 8212
rect 18028 8035 18068 8044
rect 19180 8084 19220 10816
rect 19276 9680 19316 11656
rect 19372 11444 19412 12496
rect 19468 11696 19508 12916
rect 19468 11647 19508 11656
rect 19372 11395 19412 11404
rect 19276 9631 19316 9640
rect 19372 11276 19412 11285
rect 19372 8084 19412 11236
rect 19564 11024 19604 15016
rect 19660 13292 19700 20392
rect 19756 20264 19796 20644
rect 20236 20600 20276 20695
rect 20236 20551 20276 20560
rect 19900 20432 20268 20441
rect 19900 20383 20268 20392
rect 19756 20215 19796 20224
rect 20332 20180 20372 20896
rect 20332 20131 20372 20140
rect 20428 20852 20468 20861
rect 20428 20096 20468 20812
rect 20428 20047 20468 20056
rect 20524 20600 20564 23164
rect 20620 23540 20660 23549
rect 20620 21524 20660 23500
rect 20716 23456 20756 25180
rect 20716 23407 20756 23416
rect 20812 23288 20852 26776
rect 21100 26648 21140 26657
rect 20908 25724 20948 25733
rect 20908 25472 20948 25684
rect 20908 25423 20948 25432
rect 21004 25556 21044 25565
rect 21004 25421 21044 25516
rect 20908 25304 20948 25313
rect 20908 24380 20948 25264
rect 21004 24884 21044 24893
rect 21004 24749 21044 24844
rect 20908 24331 20948 24340
rect 20812 23239 20852 23248
rect 20908 23960 20948 23969
rect 20908 23036 20948 23920
rect 20908 22987 20948 22996
rect 21004 23792 21044 23801
rect 20812 22952 20852 22961
rect 20812 22364 20852 22912
rect 21004 22532 21044 23752
rect 21100 23288 21140 26608
rect 21292 26144 21332 26153
rect 21292 26009 21332 26104
rect 21388 26060 21428 27112
rect 21388 26011 21428 26020
rect 21484 26732 21524 26741
rect 21484 25976 21524 26692
rect 21676 26480 21716 26489
rect 21676 26144 21716 26440
rect 21676 26095 21716 26104
rect 21484 25927 21524 25936
rect 21676 25976 21716 25985
rect 21292 25304 21332 25313
rect 21292 24800 21332 25264
rect 21580 25304 21620 25315
rect 21580 25220 21620 25264
rect 21388 25052 21428 25061
rect 21388 24917 21428 25012
rect 21292 24751 21332 24760
rect 21580 24716 21620 25180
rect 21580 24667 21620 24676
rect 21580 24548 21620 24557
rect 21580 24413 21620 24508
rect 21292 24128 21332 24137
rect 21292 23876 21332 24088
rect 21292 23827 21332 23836
rect 21388 23624 21428 23719
rect 21388 23575 21428 23584
rect 21100 23239 21140 23248
rect 21196 23456 21236 23465
rect 21004 22483 21044 22492
rect 21100 23120 21140 23129
rect 20812 22315 20852 22324
rect 20716 22112 20756 22121
rect 20716 21608 20756 22072
rect 20716 21559 20756 21568
rect 21100 21608 21140 23080
rect 21100 21559 21140 21568
rect 20620 21475 20660 21484
rect 20716 21440 20756 21449
rect 20524 20180 20564 20560
rect 20620 20768 20660 20777
rect 20620 20348 20660 20728
rect 20620 20299 20660 20308
rect 20332 19928 20372 19937
rect 19900 18920 20268 18929
rect 19900 18871 20268 18880
rect 20332 18500 20372 19888
rect 20524 19424 20564 20140
rect 20524 19375 20564 19384
rect 20716 19508 20756 21400
rect 21196 20180 21236 23416
rect 21580 23204 21620 23215
rect 21388 23120 21428 23129
rect 21388 21356 21428 23080
rect 21580 23120 21620 23164
rect 21580 23071 21620 23080
rect 21580 22868 21620 22877
rect 21484 22784 21524 22793
rect 21484 22364 21524 22744
rect 21484 22028 21524 22324
rect 21484 21979 21524 21988
rect 21580 21692 21620 22828
rect 21676 22532 21716 25936
rect 21772 25136 21812 27532
rect 21772 23792 21812 25096
rect 21772 23743 21812 23752
rect 21868 24632 21908 27616
rect 22252 27572 22292 27581
rect 22252 27068 22292 27532
rect 23692 27404 23732 27413
rect 23116 27320 23156 27329
rect 23156 27280 23444 27320
rect 23116 27271 23156 27280
rect 23404 27236 23444 27280
rect 23404 27187 23444 27196
rect 22252 27019 22292 27028
rect 22444 27068 22484 27077
rect 21676 22483 21716 22492
rect 21772 22532 21812 22541
rect 21772 22364 21812 22492
rect 21772 22315 21812 22324
rect 21676 22112 21716 22207
rect 21676 22063 21716 22072
rect 21580 21643 21620 21652
rect 21868 21608 21908 24592
rect 21868 21559 21908 21568
rect 21964 26732 22004 26741
rect 21388 21307 21428 21316
rect 21292 20768 21332 20777
rect 21292 20600 21332 20728
rect 21964 20768 22004 26692
rect 22444 26648 22484 27028
rect 23596 27068 23636 27077
rect 23020 26900 23060 26909
rect 23020 26816 23060 26860
rect 23020 26765 23060 26776
rect 22444 26599 22484 26608
rect 22636 26648 22676 26657
rect 22252 26480 22292 26489
rect 22156 26228 22196 26237
rect 22156 26060 22196 26188
rect 22156 26011 22196 26020
rect 22252 26144 22292 26440
rect 22636 26228 22676 26608
rect 22924 26396 22964 26405
rect 22636 26179 22676 26188
rect 22828 26228 22868 26237
rect 22156 25472 22196 25481
rect 22060 24296 22100 24305
rect 22060 23792 22100 24256
rect 22060 23743 22100 23752
rect 22060 22952 22100 22961
rect 22060 22364 22100 22912
rect 22060 22315 22100 22324
rect 22156 22280 22196 25432
rect 22156 22231 22196 22240
rect 21964 20719 22004 20728
rect 21292 20551 21332 20560
rect 21580 20684 21620 20693
rect 21388 20516 21428 20525
rect 21388 20381 21428 20476
rect 21580 20348 21620 20644
rect 21580 20299 21620 20308
rect 21676 20600 21716 20609
rect 20332 18451 20372 18460
rect 20428 19172 20468 19181
rect 20428 18416 20468 19132
rect 20716 18920 20756 19468
rect 20716 18871 20756 18880
rect 20908 20140 21236 20180
rect 21388 20264 21428 20273
rect 20908 19172 20948 20140
rect 20620 18752 20660 18761
rect 20620 18584 20660 18712
rect 20620 18535 20660 18544
rect 20812 18584 20852 18593
rect 20140 18332 20180 18341
rect 20140 17576 20180 18292
rect 20332 17912 20372 17921
rect 20428 17912 20468 18376
rect 20812 18416 20852 18544
rect 20716 18332 20756 18341
rect 20372 17872 20468 17912
rect 20524 18248 20564 18257
rect 20332 17863 20372 17872
rect 20140 17527 20180 17536
rect 20332 17744 20372 17753
rect 19900 17408 20268 17417
rect 19900 17359 20268 17368
rect 19852 17240 19892 17249
rect 19756 16904 19796 16913
rect 19756 16568 19796 16864
rect 19756 16519 19796 16528
rect 19852 16232 19892 17200
rect 20332 17240 20372 17704
rect 20524 17744 20564 18208
rect 20524 17695 20564 17704
rect 20332 17191 20372 17200
rect 20524 17576 20564 17585
rect 20428 17156 20468 17167
rect 19948 17072 19988 17081
rect 19948 16937 19988 17032
rect 20428 17072 20468 17116
rect 20428 17023 20468 17032
rect 20140 16988 20180 16997
rect 20140 16820 20180 16948
rect 20140 16771 20180 16780
rect 19852 16183 19892 16192
rect 19948 16736 19988 16745
rect 19948 16232 19988 16696
rect 20428 16400 20468 16409
rect 19948 16183 19988 16192
rect 20236 16316 20276 16325
rect 20236 16148 20276 16276
rect 20428 16265 20468 16360
rect 20236 16099 20276 16108
rect 20332 16148 20372 16159
rect 19756 16064 19796 16073
rect 19756 15476 19796 16024
rect 20332 16064 20372 16108
rect 20332 16015 20372 16024
rect 19900 15896 20268 15905
rect 20524 15896 20564 17536
rect 20620 17492 20660 17501
rect 20620 17072 20660 17452
rect 20620 16316 20660 17032
rect 20620 16267 20660 16276
rect 20716 16148 20756 18292
rect 20812 17828 20852 18376
rect 20908 17912 20948 19132
rect 21196 19760 21236 19769
rect 21196 19256 21236 19720
rect 21004 18500 21044 18509
rect 21004 18080 21044 18460
rect 21196 18332 21236 19216
rect 21196 18283 21236 18292
rect 21004 18031 21044 18040
rect 20908 17872 21044 17912
rect 20812 17779 20852 17788
rect 20908 17072 20948 17081
rect 20908 16820 20948 17032
rect 20908 16771 20948 16780
rect 20908 16316 20948 16325
rect 20908 16232 20948 16276
rect 20908 16181 20948 16192
rect 19900 15847 20268 15856
rect 20332 15856 20564 15896
rect 20620 16108 20756 16148
rect 21004 16148 21044 17872
rect 21388 17744 21428 20224
rect 19756 15427 19796 15436
rect 19852 15644 19892 15653
rect 19756 15308 19796 15317
rect 19756 14972 19796 15268
rect 19756 14923 19796 14932
rect 19756 14804 19796 14813
rect 19756 14669 19796 14764
rect 19852 14636 19892 15604
rect 19948 15560 19988 15569
rect 19948 14888 19988 15520
rect 20044 15392 20084 15487
rect 20044 15343 20084 15352
rect 19948 14839 19988 14848
rect 20044 15140 20084 15149
rect 20044 14804 20084 15100
rect 20044 14755 20084 14764
rect 19852 14552 19892 14596
rect 19756 14512 19892 14552
rect 20140 14552 20180 14647
rect 19756 14132 19796 14512
rect 20140 14503 20180 14512
rect 19900 14384 20268 14393
rect 19900 14335 20268 14344
rect 20140 14216 20180 14225
rect 19756 14092 19892 14132
rect 19756 13880 19796 13889
rect 19756 13745 19796 13840
rect 19660 13243 19700 13252
rect 19852 13292 19892 14092
rect 20140 14081 20180 14176
rect 20044 14048 20084 14057
rect 19948 13712 19988 13721
rect 19948 13460 19988 13672
rect 19948 13411 19988 13420
rect 20044 13376 20084 14008
rect 20044 13327 20084 13336
rect 20236 13964 20276 13973
rect 19756 13124 19796 13133
rect 19660 13040 19700 13049
rect 19660 12620 19700 13000
rect 19756 12956 19796 13084
rect 19852 13124 19892 13252
rect 19852 13075 19892 13084
rect 20236 13124 20276 13924
rect 20332 13544 20372 15856
rect 20428 15728 20468 15737
rect 20428 15560 20468 15688
rect 20428 15511 20468 15520
rect 20332 13292 20372 13504
rect 20332 13243 20372 13252
rect 20428 15392 20468 15401
rect 20428 13208 20468 15352
rect 20524 15308 20564 15317
rect 20524 14720 20564 15268
rect 20524 14671 20564 14680
rect 20620 14552 20660 16108
rect 20908 15560 20948 15569
rect 20812 15476 20852 15485
rect 20716 15392 20756 15401
rect 20716 14888 20756 15352
rect 20812 14972 20852 15436
rect 20908 15392 20948 15520
rect 20908 15343 20948 15352
rect 20812 14923 20852 14932
rect 20716 14839 20756 14848
rect 21004 14888 21044 16108
rect 21196 16904 21236 16913
rect 21196 16232 21236 16864
rect 21196 15560 21236 16192
rect 21292 16652 21332 16661
rect 21292 16148 21332 16612
rect 21292 16099 21332 16108
rect 21292 15560 21332 15569
rect 21196 15520 21292 15560
rect 21004 14839 21044 14848
rect 21100 15392 21140 15401
rect 21100 14804 21140 15352
rect 21100 14669 21140 14764
rect 20908 14636 20948 14645
rect 20524 14512 20660 14552
rect 20716 14552 20756 14561
rect 20524 14132 20564 14512
rect 20524 14083 20564 14092
rect 20620 14216 20660 14225
rect 20428 13159 20468 13168
rect 20524 13544 20564 13553
rect 20236 13075 20276 13084
rect 19756 12907 19796 12916
rect 19900 12872 20268 12881
rect 19900 12823 20268 12832
rect 19660 12571 19700 12580
rect 19948 12704 19988 12713
rect 19756 12536 19796 12545
rect 19756 12401 19796 12496
rect 19756 12284 19796 12293
rect 19756 12149 19796 12244
rect 19660 12116 19700 12125
rect 19660 11780 19700 12076
rect 19660 11731 19700 11740
rect 19948 11528 19988 12664
rect 20524 12704 20564 13504
rect 20620 13460 20660 14176
rect 20716 13628 20756 14512
rect 20812 14048 20852 14057
rect 20812 13913 20852 14008
rect 20716 13579 20756 13588
rect 20908 13628 20948 14596
rect 20908 13579 20948 13588
rect 21004 14636 21044 14645
rect 20620 13411 20660 13420
rect 20812 13460 20852 13555
rect 20812 13411 20852 13420
rect 20812 13292 20852 13301
rect 20524 12655 20564 12664
rect 20716 13124 20756 13133
rect 20524 12536 20564 12545
rect 20428 12452 20468 12461
rect 20236 12200 20276 12209
rect 20236 11780 20276 12160
rect 20236 11731 20276 11740
rect 19468 10016 19508 10025
rect 19468 9932 19508 9976
rect 19468 9881 19508 9892
rect 19564 8840 19604 10984
rect 19756 11488 19988 11528
rect 19756 9764 19796 11488
rect 19900 11360 20268 11369
rect 19900 11311 20268 11320
rect 20332 11024 20372 11033
rect 20140 10520 20180 10529
rect 20140 10436 20180 10480
rect 20140 10385 20180 10396
rect 20332 10016 20372 10984
rect 20332 9967 20372 9976
rect 19900 9848 20268 9857
rect 19900 9799 20268 9808
rect 19756 9715 19796 9724
rect 20428 9764 20468 12412
rect 20524 11192 20564 12496
rect 20716 12536 20756 13084
rect 20716 12487 20756 12496
rect 20812 12536 20852 13252
rect 20812 11696 20852 12496
rect 20812 11647 20852 11656
rect 21004 13124 21044 14596
rect 21196 14552 21236 14561
rect 21196 13964 21236 14512
rect 21196 13915 21236 13924
rect 21196 13796 21236 13807
rect 21196 13712 21236 13756
rect 21196 13663 21236 13672
rect 20524 11143 20564 11152
rect 20908 11528 20948 11537
rect 20908 11024 20948 11488
rect 20908 10975 20948 10984
rect 20524 9932 20564 9941
rect 20524 9797 20564 9892
rect 19564 8791 19604 8800
rect 19660 9512 19700 9521
rect 19660 8168 19700 9472
rect 20332 9512 20372 9521
rect 20140 9428 20180 9437
rect 20140 8924 20180 9388
rect 20140 8875 20180 8884
rect 19900 8336 20268 8345
rect 19900 8287 20268 8296
rect 19660 8119 19700 8128
rect 19372 8044 19508 8084
rect 19180 8035 19220 8044
rect 16492 4976 16532 5524
rect 16492 4927 16532 4936
rect 17356 5816 17396 7960
rect 17740 8000 17780 8009
rect 17356 4976 17396 5776
rect 17548 7160 17588 7169
rect 17548 6656 17588 7120
rect 17740 6992 17780 7960
rect 18124 8000 18164 8009
rect 18604 8000 18644 8009
rect 18124 7412 18164 7960
rect 18124 7363 18164 7372
rect 18508 7960 18604 8000
rect 17740 6943 17780 6952
rect 18124 7160 18164 7169
rect 17548 5732 17588 6616
rect 18124 6488 18164 7120
rect 18124 5900 18164 6448
rect 18316 7076 18356 7085
rect 18316 6488 18356 7036
rect 18508 6740 18548 7960
rect 18604 7951 18644 7960
rect 19180 7916 19220 7925
rect 18660 7580 19028 7589
rect 18660 7531 19028 7540
rect 18892 7412 18932 7421
rect 18700 7244 18740 7253
rect 18700 7160 18740 7204
rect 18700 7109 18740 7120
rect 18508 6691 18548 6700
rect 18604 7076 18644 7085
rect 18604 6656 18644 7036
rect 18604 6607 18644 6616
rect 18892 6656 18932 7372
rect 19180 7160 19220 7876
rect 19180 7076 19220 7120
rect 19372 7916 19412 7925
rect 19372 7244 19412 7876
rect 19372 7160 19412 7204
rect 19372 7080 19412 7120
rect 18892 6607 18932 6616
rect 18988 6992 19028 7001
rect 18316 6152 18356 6448
rect 18988 6488 19028 6952
rect 18988 6439 19028 6448
rect 19180 6488 19220 7036
rect 19468 6572 19508 8044
rect 20236 7748 20276 7757
rect 19564 7328 19604 7337
rect 19564 6824 19604 7288
rect 20236 7328 20276 7708
rect 20044 7244 20084 7253
rect 19564 6775 19604 6784
rect 19660 7076 19700 7085
rect 19660 6740 19700 7036
rect 20044 6992 20084 7204
rect 20236 7160 20276 7288
rect 20332 7244 20372 9472
rect 20428 8672 20468 9724
rect 20428 8623 20468 8632
rect 20812 8756 20852 8765
rect 20812 8504 20852 8716
rect 20620 8084 20660 8093
rect 20332 7195 20372 7204
rect 20524 7748 20564 7757
rect 20524 7244 20564 7708
rect 20524 7195 20564 7204
rect 20236 7111 20276 7120
rect 20044 6943 20084 6952
rect 20428 7076 20468 7085
rect 19900 6824 20268 6833
rect 19900 6775 20268 6784
rect 19660 6691 19700 6700
rect 19180 6439 19220 6448
rect 19372 6532 19508 6572
rect 18316 6103 18356 6112
rect 18660 6068 19028 6077
rect 18660 6019 19028 6028
rect 19372 5984 19412 6532
rect 20140 6488 20180 6497
rect 19372 5935 19412 5944
rect 19468 6404 19508 6413
rect 18124 5851 18164 5860
rect 17548 5683 17588 5692
rect 18220 5732 18260 5741
rect 17356 4927 17396 4936
rect 15052 4759 15092 4768
rect 18220 4808 18260 5692
rect 19468 5648 19508 6364
rect 20140 5900 20180 6448
rect 20428 5984 20468 7036
rect 20620 6656 20660 8044
rect 20812 7916 20852 8464
rect 20716 7328 20756 7337
rect 20716 7076 20756 7288
rect 20716 7027 20756 7036
rect 20620 6607 20660 6616
rect 20716 6488 20756 6497
rect 20428 5935 20468 5944
rect 20620 6236 20660 6245
rect 20140 5851 20180 5860
rect 20620 5900 20660 6196
rect 20620 5851 20660 5860
rect 20716 5732 20756 6448
rect 20716 5683 20756 5692
rect 20812 6236 20852 7876
rect 20908 8588 20948 8597
rect 20908 8000 20948 8548
rect 20908 7412 20948 7960
rect 20908 7363 20948 7372
rect 18220 4759 18260 4768
rect 19276 5564 19316 5573
rect 11980 4675 12020 4684
rect 10886 4556 11254 4565
rect 10886 4507 11254 4516
rect 18660 4556 19028 4565
rect 18660 4507 19028 4516
rect 19276 4388 19316 5524
rect 19468 5144 19508 5608
rect 20332 5648 20372 5657
rect 19900 5312 20268 5321
rect 19900 5263 20268 5272
rect 19468 5095 19508 5104
rect 19276 4339 19316 4348
rect 19852 4724 19892 4733
rect 9772 4087 9812 4096
rect 19852 4136 19892 4684
rect 20332 4388 20372 5608
rect 20332 4339 20372 4348
rect 20428 5480 20468 5489
rect 20428 4808 20468 5440
rect 20428 4220 20468 4768
rect 20524 4976 20564 4985
rect 20524 4388 20564 4936
rect 20524 4339 20564 4348
rect 20428 4171 20468 4180
rect 19852 4087 19892 4096
rect 20812 4136 20852 6196
rect 20908 5564 20948 5573
rect 20908 4976 20948 5524
rect 20908 4927 20948 4936
rect 21004 5396 21044 13084
rect 21196 13376 21236 13385
rect 21100 13040 21140 13049
rect 21100 12284 21140 13000
rect 21196 12788 21236 13336
rect 21196 12739 21236 12748
rect 21100 10940 21140 12244
rect 21292 11948 21332 15520
rect 21388 14636 21428 17704
rect 21484 20180 21524 20189
rect 21484 16484 21524 20140
rect 21676 20096 21716 20560
rect 21676 20047 21716 20056
rect 21772 19928 21812 19937
rect 21580 17744 21620 17753
rect 21580 16904 21620 17704
rect 21580 16855 21620 16864
rect 21484 16400 21524 16444
rect 21484 16320 21524 16360
rect 21676 15812 21716 15823
rect 21676 15728 21716 15772
rect 21676 15679 21716 15688
rect 21388 14587 21428 14596
rect 21484 15476 21524 15485
rect 21388 14468 21428 14477
rect 21388 14216 21428 14428
rect 21388 14167 21428 14176
rect 21388 14048 21428 14059
rect 21388 13964 21428 14008
rect 21388 13915 21428 13924
rect 21484 13880 21524 15436
rect 21580 15392 21620 15401
rect 21580 14804 21620 15352
rect 21580 14755 21620 14764
rect 21676 14888 21716 14897
rect 21676 14720 21716 14848
rect 21676 14671 21716 14680
rect 21580 14636 21620 14645
rect 21580 14132 21620 14596
rect 21580 14083 21620 14092
rect 21676 14552 21716 14561
rect 21388 12704 21428 12713
rect 21484 12704 21524 13840
rect 21676 13460 21716 14512
rect 21676 13411 21716 13420
rect 21580 13124 21620 13133
rect 21580 12956 21620 13084
rect 21772 12980 21812 19888
rect 22156 19424 22196 19433
rect 22156 19256 22196 19384
rect 22156 19207 22196 19216
rect 22156 19088 22196 19097
rect 22156 18584 22196 19048
rect 22252 18752 22292 26104
rect 22444 26144 22484 26153
rect 22444 25640 22484 26104
rect 22444 25591 22484 25600
rect 22828 25472 22868 26188
rect 22828 25423 22868 25432
rect 22924 25304 22964 26356
rect 23308 26228 23348 26237
rect 23020 26144 23060 26153
rect 23020 25472 23060 26104
rect 23116 25976 23156 25985
rect 23116 25556 23156 25936
rect 23116 25507 23156 25516
rect 23020 25423 23060 25432
rect 23212 25472 23252 25481
rect 22924 25220 22964 25264
rect 22924 25171 22964 25180
rect 23212 25304 23252 25432
rect 23308 25388 23348 26188
rect 23596 26144 23636 27028
rect 23692 26900 23732 27364
rect 23692 26851 23732 26860
rect 23596 26095 23636 26104
rect 23692 25976 23732 25985
rect 23692 25841 23732 25936
rect 24076 25892 24116 25901
rect 23308 25339 23348 25348
rect 23212 25136 23252 25264
rect 24076 25304 24116 25852
rect 24172 25556 24212 27700
rect 25804 27740 25844 27749
rect 24364 27656 24404 27665
rect 24172 25507 24212 25516
rect 24268 25808 24308 25817
rect 24076 25255 24116 25264
rect 22636 25052 22676 25061
rect 22636 24800 22676 25012
rect 22636 24751 22676 24760
rect 23020 24800 23060 24809
rect 22348 24716 22388 24725
rect 22348 24044 22388 24676
rect 22924 24716 22964 24725
rect 22924 24632 22964 24676
rect 22924 24581 22964 24592
rect 22348 23995 22388 24004
rect 22444 24464 22484 24473
rect 22348 23792 22388 23801
rect 22348 21440 22388 23752
rect 22444 23624 22484 24424
rect 22444 23575 22484 23584
rect 22540 24212 22580 24221
rect 22444 22280 22484 22289
rect 22444 21608 22484 22240
rect 22444 21559 22484 21568
rect 22348 21400 22484 21440
rect 22348 20768 22388 20777
rect 22348 19508 22388 20728
rect 22348 19172 22388 19468
rect 22348 19123 22388 19132
rect 22252 18703 22292 18712
rect 22156 18535 22196 18544
rect 22444 18500 22484 21400
rect 22540 19256 22580 24172
rect 22636 23876 22676 23885
rect 22636 23540 22676 23836
rect 22924 23792 22964 23801
rect 22924 23624 22964 23752
rect 22924 23575 22964 23584
rect 22636 23491 22676 23500
rect 22732 23540 22772 23549
rect 22732 23372 22772 23500
rect 22732 23323 22772 23332
rect 22732 23120 22772 23129
rect 22636 22196 22676 22205
rect 22636 21608 22676 22156
rect 22636 20768 22676 21568
rect 22732 21440 22772 23080
rect 23020 22028 23060 24760
rect 23212 24464 23252 25096
rect 23212 24415 23252 24424
rect 23308 25220 23348 25229
rect 23116 23792 23156 23887
rect 23116 23743 23156 23752
rect 23308 23624 23348 25180
rect 24268 25136 24308 25768
rect 24268 25087 24308 25096
rect 23308 23540 23348 23584
rect 23308 23489 23348 23500
rect 23596 24716 23636 24725
rect 23020 21979 23060 21988
rect 23500 21524 23540 21533
rect 22828 21440 22868 21449
rect 22732 21400 22828 21440
rect 22732 20852 22772 21400
rect 22828 21391 22868 21400
rect 23308 21188 23348 21197
rect 22732 20803 22772 20812
rect 22924 21104 22964 21113
rect 22924 20852 22964 21064
rect 22924 20803 22964 20812
rect 22636 20719 22676 20728
rect 23308 20768 23348 21148
rect 22732 20684 22772 20693
rect 22636 20600 22676 20609
rect 22636 20012 22676 20560
rect 22732 20549 22772 20644
rect 22636 19963 22676 19972
rect 22732 20180 22772 20189
rect 22540 19207 22580 19216
rect 22540 18752 22580 18761
rect 22540 18617 22580 18712
rect 22252 18460 22444 18500
rect 21868 17744 21908 17753
rect 21868 17324 21908 17704
rect 21868 16988 21908 17284
rect 21868 16939 21908 16948
rect 22060 17744 22100 17753
rect 21868 16820 21908 16829
rect 21868 16736 21908 16780
rect 21868 16685 21908 16696
rect 22060 16316 22100 17704
rect 22156 17576 22196 17585
rect 22156 17072 22196 17536
rect 22156 16484 22196 17032
rect 22156 16435 22196 16444
rect 22252 16400 22292 18460
rect 22444 18451 22484 18460
rect 22636 17660 22676 17669
rect 22444 17576 22484 17585
rect 22444 17156 22484 17536
rect 22444 17107 22484 17116
rect 22348 16484 22388 16579
rect 22348 16435 22388 16444
rect 22252 16351 22292 16360
rect 22060 16267 22100 16276
rect 22348 16316 22388 16325
rect 21964 16148 22004 16157
rect 21964 15980 22004 16108
rect 21964 15728 22004 15940
rect 21964 15679 22004 15688
rect 22060 16064 22100 16073
rect 21868 15560 21908 15569
rect 21868 14132 21908 15520
rect 21964 15476 22004 15485
rect 21964 14972 22004 15436
rect 21964 14923 22004 14932
rect 21868 14083 21908 14092
rect 21964 14636 22004 14645
rect 21964 13880 22004 14596
rect 22060 14552 22100 16024
rect 22348 15728 22388 16276
rect 22348 15679 22388 15688
rect 22156 15644 22196 15653
rect 22156 15392 22196 15604
rect 22444 15644 22484 15653
rect 22156 15343 22196 15352
rect 22252 15560 22292 15569
rect 22252 15140 22292 15520
rect 22444 15392 22484 15604
rect 22636 15644 22676 17620
rect 22636 15595 22676 15604
rect 22444 15343 22484 15352
rect 22540 15476 22580 15485
rect 22732 15476 22772 20140
rect 23116 20096 23156 20105
rect 22924 19844 22964 19853
rect 22924 19340 22964 19804
rect 23116 19592 23156 20056
rect 23116 19543 23156 19552
rect 23308 19424 23348 20728
rect 23308 19375 23348 19384
rect 23404 20516 23444 20525
rect 22924 19291 22964 19300
rect 23116 19256 23156 19265
rect 23116 19121 23156 19216
rect 23404 19172 23444 20476
rect 23500 20516 23540 21484
rect 23500 20467 23540 20476
rect 23596 20768 23636 24676
rect 24364 24632 24404 27616
rect 25228 27656 25268 27665
rect 24556 27572 24596 27583
rect 24556 27488 24596 27532
rect 24556 27439 24596 27448
rect 24748 27572 24788 27581
rect 24460 26312 24500 26321
rect 24460 26144 24500 26272
rect 24460 26095 24500 26104
rect 24748 25556 24788 27532
rect 24940 26900 24980 26909
rect 24844 26060 24884 26069
rect 24844 25925 24884 26020
rect 24748 25507 24788 25516
rect 24940 25472 24980 26860
rect 25132 26396 25172 26405
rect 25132 25892 25172 26356
rect 25132 25843 25172 25852
rect 25228 26060 25268 27616
rect 25804 27605 25844 27700
rect 26188 27740 26228 28600
rect 26764 28328 26804 28337
rect 26188 27691 26228 27700
rect 26380 27908 26420 27917
rect 26380 27656 26420 27868
rect 25900 27572 25940 27581
rect 24940 25423 24980 25432
rect 25228 25556 25268 26020
rect 23788 24548 23828 24557
rect 23788 23708 23828 24508
rect 24364 23960 24404 24592
rect 24940 25304 24980 25313
rect 24460 24380 24500 24389
rect 24460 24212 24500 24340
rect 24460 24163 24500 24172
rect 23788 23659 23828 23668
rect 24076 23876 24116 23885
rect 24076 23120 24116 23836
rect 24364 23792 24404 23920
rect 24364 23743 24404 23752
rect 24460 23792 24500 23801
rect 24076 23036 24116 23080
rect 24076 22364 24116 22996
rect 24076 21608 24116 22324
rect 23980 21568 24076 21608
rect 23884 21524 23924 21533
rect 23404 19123 23444 19132
rect 23020 19088 23060 19097
rect 22924 19048 23020 19088
rect 22924 18584 22964 19048
rect 23020 19020 23060 19048
rect 23500 19088 23540 19097
rect 22924 18535 22964 18544
rect 23212 18332 23252 18341
rect 23116 17744 23156 17753
rect 23116 17609 23156 17704
rect 23212 17576 23252 18292
rect 23500 17828 23540 19048
rect 23596 18332 23636 20728
rect 23788 21356 23828 21365
rect 23692 19340 23732 19435
rect 23692 19291 23732 19300
rect 23596 18283 23636 18292
rect 23692 19172 23732 19181
rect 23500 17779 23540 17788
rect 23020 17072 23060 17081
rect 23020 16568 23060 17032
rect 23020 16519 23060 16528
rect 22828 16316 22868 16325
rect 22828 16181 22868 16276
rect 23020 15728 23060 15737
rect 22252 15091 22292 15100
rect 22540 14804 22580 15436
rect 22060 14503 22100 14512
rect 22252 14720 22292 14729
rect 21964 13831 22004 13840
rect 22060 14048 22100 14057
rect 21868 13544 21908 13553
rect 21868 13208 21908 13504
rect 22060 13460 22100 14008
rect 22060 13411 22100 13420
rect 22156 13964 22196 13973
rect 22156 13712 22196 13924
rect 21868 13159 21908 13168
rect 22156 13208 22196 13672
rect 22156 13159 22196 13168
rect 22060 13124 22100 13135
rect 22060 13040 22100 13084
rect 22252 13124 22292 14680
rect 22444 14720 22484 14731
rect 22444 14636 22484 14680
rect 22444 14587 22484 14596
rect 22348 14552 22388 14561
rect 22348 13964 22388 14512
rect 22540 14468 22580 14764
rect 22540 14419 22580 14428
rect 22636 15436 22772 15476
rect 22924 15644 22964 15653
rect 22444 14048 22484 14143
rect 22444 13999 22484 14008
rect 22348 13915 22388 13924
rect 22636 13880 22676 15436
rect 22924 14888 22964 15604
rect 23020 15593 23060 15688
rect 22924 14839 22964 14848
rect 22924 14720 22964 14729
rect 22924 14048 22964 14680
rect 22924 13999 22964 14008
rect 23116 14552 23156 14561
rect 22444 13840 22676 13880
rect 22732 13964 22772 13973
rect 22348 13376 22388 13385
rect 22348 13241 22388 13336
rect 22252 13075 22292 13084
rect 22060 12991 22100 13000
rect 21580 12907 21620 12916
rect 21676 12940 21812 12980
rect 21428 12664 21524 12704
rect 21388 12655 21428 12664
rect 21292 11899 21332 11908
rect 21580 11612 21620 11621
rect 21100 10891 21140 10900
rect 21292 11360 21332 11369
rect 21292 10520 21332 11320
rect 21196 9428 21236 9437
rect 21100 8756 21140 8765
rect 21100 8084 21140 8716
rect 21196 8168 21236 9388
rect 21292 8756 21332 10480
rect 21484 11024 21524 11033
rect 21484 10520 21524 10984
rect 21484 10436 21524 10480
rect 21484 10385 21524 10396
rect 21484 10016 21524 10025
rect 21484 9596 21524 9976
rect 21484 9547 21524 9556
rect 21580 8924 21620 11572
rect 21676 10940 21716 12940
rect 21868 12536 21908 12545
rect 21772 12284 21812 12293
rect 21772 11612 21812 12244
rect 21772 11563 21812 11572
rect 21868 11696 21908 12496
rect 21676 10891 21716 10900
rect 21868 11108 21908 11656
rect 21580 8875 21620 8884
rect 21772 10772 21812 10781
rect 21292 8707 21332 8716
rect 21580 8756 21620 8765
rect 21196 8119 21236 8128
rect 21388 8672 21428 8681
rect 21388 8168 21428 8632
rect 21580 8672 21620 8716
rect 21580 8621 21620 8632
rect 21772 8672 21812 10732
rect 21868 10184 21908 11068
rect 21868 10135 21908 10144
rect 21964 11780 22004 11789
rect 21868 9932 21908 9941
rect 21868 9512 21908 9892
rect 21868 8756 21908 9472
rect 21868 8707 21908 8716
rect 21772 8623 21812 8632
rect 21388 8119 21428 8128
rect 21100 8035 21140 8044
rect 21292 6992 21332 7001
rect 20812 4087 20852 4096
rect 21004 4052 21044 5356
rect 21196 5984 21236 5993
rect 21196 5144 21236 5944
rect 21196 5095 21236 5104
rect 21292 5648 21332 6952
rect 21292 4220 21332 5608
rect 21388 6656 21428 6665
rect 21388 4976 21428 6616
rect 21388 4927 21428 4936
rect 21580 6404 21620 6413
rect 21580 4808 21620 6364
rect 21964 5816 22004 11740
rect 22444 11108 22484 13840
rect 22732 13829 22772 13924
rect 22828 13880 22868 13889
rect 22636 13712 22676 13721
rect 22540 13292 22580 13301
rect 22540 12788 22580 13252
rect 22636 13208 22676 13672
rect 22828 13460 22868 13840
rect 22828 13411 22868 13420
rect 22636 13159 22676 13168
rect 23116 13208 23156 14512
rect 23212 14468 23252 17536
rect 23308 17660 23348 17669
rect 23308 16064 23348 17620
rect 23500 17576 23540 17585
rect 23500 17072 23540 17536
rect 23500 17023 23540 17032
rect 23596 17492 23636 17501
rect 23692 17492 23732 19132
rect 23788 19004 23828 21316
rect 23884 20684 23924 21484
rect 23884 20635 23924 20644
rect 23884 20180 23924 20189
rect 23980 20180 24020 21568
rect 24076 21559 24116 21568
rect 24172 23456 24212 23465
rect 24172 21440 24212 23416
rect 24460 22532 24500 23752
rect 24940 23792 24980 25264
rect 25228 25304 25268 25516
rect 25804 27404 25844 27413
rect 25036 24800 25076 24809
rect 25036 24128 25076 24760
rect 25036 24079 25076 24088
rect 25132 24632 25172 24641
rect 24940 23743 24980 23752
rect 25132 23792 25172 24592
rect 25132 23743 25172 23752
rect 24460 22483 24500 22492
rect 24556 23708 24596 23717
rect 24460 22112 24500 22121
rect 24172 21391 24212 21400
rect 24268 21776 24308 21785
rect 24172 20768 24212 20777
rect 23924 20140 24020 20180
rect 24076 20516 24116 20525
rect 23884 20131 23924 20140
rect 24076 20096 24116 20476
rect 24076 20047 24116 20056
rect 24172 20012 24212 20728
rect 24268 20600 24308 21736
rect 24364 21524 24404 21533
rect 24364 20936 24404 21484
rect 24460 21524 24500 22072
rect 24460 21475 24500 21484
rect 24556 21692 24596 23668
rect 24748 23288 24788 23297
rect 24364 20684 24404 20896
rect 24364 20635 24404 20644
rect 24556 20852 24596 21652
rect 24268 20551 24308 20560
rect 24460 20600 24500 20609
rect 24364 20264 24404 20273
rect 24364 20096 24404 20224
rect 24364 20047 24404 20056
rect 24172 19963 24212 19972
rect 24460 19676 24500 20560
rect 24460 19627 24500 19636
rect 24076 19424 24116 19433
rect 24076 19256 24116 19384
rect 24076 19207 24116 19216
rect 24460 19256 24500 19265
rect 23788 18955 23828 18964
rect 24460 18752 24500 19216
rect 24556 19004 24596 20812
rect 24652 21860 24692 21869
rect 24652 21608 24692 21820
rect 24652 20768 24692 21568
rect 24652 20719 24692 20728
rect 24748 20096 24788 23248
rect 25228 23204 25268 25264
rect 25420 25388 25460 25399
rect 25420 25304 25460 25348
rect 25420 25255 25460 25264
rect 25324 24884 25364 24893
rect 25324 24548 25364 24844
rect 25708 24800 25748 24809
rect 25708 24548 25748 24760
rect 25804 24716 25844 27364
rect 25804 24667 25844 24676
rect 25708 24508 25844 24548
rect 25324 24499 25364 24508
rect 25708 24380 25748 24389
rect 25516 24296 25556 24305
rect 25516 24128 25556 24256
rect 25516 24079 25556 24088
rect 25708 23876 25748 24340
rect 25708 23827 25748 23836
rect 25804 23876 25844 24508
rect 25900 24044 25940 27532
rect 26188 27572 26228 27581
rect 25996 27236 26036 27245
rect 25996 26060 26036 27196
rect 25996 26011 26036 26020
rect 26188 25388 26228 27532
rect 26380 27404 26420 27616
rect 26764 27656 26804 28288
rect 26764 27607 26804 27616
rect 26476 27572 26516 27581
rect 26476 27437 26516 27532
rect 26860 27572 26900 27581
rect 26380 27355 26420 27364
rect 26434 27236 26802 27245
rect 26434 27187 26802 27196
rect 26380 27068 26420 27077
rect 26284 26900 26324 26909
rect 26284 25472 26324 26860
rect 26380 26732 26420 27028
rect 26764 26984 26804 26993
rect 26380 26683 26420 26692
rect 26476 26944 26764 26984
rect 26476 26228 26516 26944
rect 26764 26935 26804 26944
rect 26764 26648 26804 26657
rect 26476 26179 26516 26188
rect 26572 26228 26612 26237
rect 26668 26228 26708 26237
rect 26612 26188 26668 26228
rect 26572 26179 26612 26188
rect 26668 26179 26708 26188
rect 26764 26228 26804 26608
rect 26764 26144 26804 26188
rect 26764 26093 26804 26104
rect 26434 25724 26802 25733
rect 26434 25675 26802 25684
rect 26284 25432 26420 25472
rect 26188 25348 26324 25388
rect 25900 23995 25940 24004
rect 25996 25220 26036 25229
rect 25324 23624 25364 23633
rect 25324 23372 25364 23584
rect 25516 23624 25556 23633
rect 25516 23489 25556 23584
rect 25324 23323 25364 23332
rect 25804 23288 25844 23836
rect 25900 23876 25940 23885
rect 25900 23708 25940 23836
rect 25996 23792 26036 25180
rect 25996 23743 26036 23752
rect 26188 25220 26228 25229
rect 26188 24632 26228 25180
rect 26188 23792 26228 24592
rect 26188 23743 26228 23752
rect 26284 24716 26324 25348
rect 25900 23659 25940 23668
rect 26284 23708 26324 24676
rect 26380 24380 26420 25432
rect 26380 24331 26420 24340
rect 26860 24296 26900 27532
rect 26956 27404 26996 28600
rect 27244 28496 27284 28505
rect 26956 27355 26996 27364
rect 27052 27908 27092 27917
rect 26956 27236 26996 27245
rect 26956 26060 26996 27196
rect 26956 26011 26996 26020
rect 26860 24247 26900 24256
rect 26434 24212 26802 24221
rect 26434 24163 26802 24172
rect 26284 23659 26324 23668
rect 25804 23239 25844 23248
rect 25900 23540 25940 23549
rect 25228 23164 25364 23204
rect 24940 22868 24980 22877
rect 24940 22448 24980 22828
rect 24940 22280 24980 22408
rect 24940 21776 24980 22240
rect 24940 21727 24980 21736
rect 25228 21608 25268 21617
rect 25132 21440 25172 21449
rect 25132 20936 25172 21400
rect 25228 21020 25268 21568
rect 25228 20971 25268 20980
rect 25132 20887 25172 20896
rect 25036 20600 25076 20609
rect 25036 20465 25076 20560
rect 24748 20047 24788 20056
rect 25324 19592 25364 23164
rect 25900 22448 25940 23500
rect 26572 23372 26612 23381
rect 25804 22408 25940 22448
rect 26284 23120 26324 23129
rect 25804 22364 25844 22408
rect 25516 22112 25556 22121
rect 25516 21776 25556 22072
rect 25516 21727 25556 21736
rect 25804 21608 25844 22324
rect 25900 22280 25940 22289
rect 25900 22028 25940 22240
rect 25900 21979 25940 21988
rect 26092 22196 26132 22205
rect 26092 21692 26132 22156
rect 26188 22112 26228 22121
rect 26188 21860 26228 22072
rect 26188 21811 26228 21820
rect 26092 21643 26132 21652
rect 25804 21559 25844 21568
rect 25612 20936 25652 20945
rect 25420 20600 25460 20609
rect 25420 20180 25460 20560
rect 25420 20131 25460 20140
rect 25612 20180 25652 20896
rect 26092 20768 26132 20777
rect 25612 20131 25652 20140
rect 25900 20684 25940 20693
rect 25900 19928 25940 20644
rect 25900 19879 25940 19888
rect 26092 19844 26132 20728
rect 26092 19795 26132 19804
rect 26284 20096 26324 23080
rect 26572 23120 26612 23332
rect 27052 23204 27092 27868
rect 27244 27656 27284 28456
rect 27724 28160 27764 28600
rect 27724 28111 27764 28120
rect 27674 27992 28042 28001
rect 27674 27943 28042 27952
rect 27724 27824 27764 27833
rect 27244 27607 27284 27616
rect 27628 27740 27668 27749
rect 27436 27572 27476 27581
rect 27148 26984 27188 26993
rect 27148 26060 27188 26944
rect 27244 26984 27284 26993
rect 27244 26732 27284 26944
rect 27244 26683 27284 26692
rect 27436 26648 27476 27532
rect 27340 26608 27476 26648
rect 27532 27488 27572 27497
rect 27340 26396 27380 26608
rect 27148 26011 27188 26020
rect 27244 26356 27380 26396
rect 27436 26480 27476 26489
rect 27244 25808 27284 26356
rect 27436 26345 27476 26440
rect 27244 25759 27284 25768
rect 27340 26228 27380 26237
rect 27340 25304 27380 26188
rect 27532 26228 27572 27448
rect 27628 26732 27668 27700
rect 27724 27656 27764 27784
rect 28492 27740 28532 28600
rect 28972 28412 29012 28421
rect 28492 27691 28532 27700
rect 28684 28160 28724 28169
rect 27724 27607 27764 27616
rect 28684 27656 28724 28120
rect 28684 27607 28724 27616
rect 28876 28160 28916 28169
rect 28492 27572 28532 27581
rect 27916 27404 27956 27413
rect 27724 26984 27764 26993
rect 27724 26816 27764 26944
rect 27724 26767 27764 26776
rect 27916 26816 27956 27364
rect 27916 26767 27956 26776
rect 28108 27068 28148 27077
rect 27628 26683 27668 26692
rect 27674 26480 28042 26489
rect 27674 26431 28042 26440
rect 27532 26179 27572 26188
rect 27916 26228 27956 26323
rect 28108 26312 28148 27028
rect 28396 26900 28436 26909
rect 28300 26732 28340 26741
rect 28108 26263 28148 26272
rect 28204 26648 28244 26657
rect 27916 26179 27956 26188
rect 27628 26144 27668 26153
rect 28204 26144 28244 26608
rect 27628 26060 27668 26104
rect 28012 26104 28244 26144
rect 27532 26020 27668 26060
rect 27724 26060 27764 26069
rect 27532 25808 27572 26020
rect 27724 25892 27764 26020
rect 27916 26060 27956 26069
rect 27916 25976 27956 26020
rect 28012 26060 28052 26104
rect 28012 26011 28052 26020
rect 27916 25925 27956 25936
rect 27724 25843 27764 25852
rect 27532 25759 27572 25768
rect 27916 25808 27956 25817
rect 27340 25169 27380 25264
rect 27916 25136 27956 25768
rect 27916 25087 27956 25096
rect 28108 25220 28148 25229
rect 27674 24968 28042 24977
rect 27674 24919 28042 24928
rect 27436 24716 27476 24725
rect 27340 24632 27380 24641
rect 27052 23155 27092 23164
rect 27148 24380 27188 24389
rect 26572 23071 26612 23080
rect 26380 23036 26420 23045
rect 26380 22901 26420 22996
rect 26860 23036 26900 23045
rect 26434 22700 26802 22709
rect 26434 22651 26802 22660
rect 26380 22532 26420 22541
rect 26380 21692 26420 22492
rect 26860 22532 26900 22996
rect 26860 22483 26900 22492
rect 27052 22532 27092 22541
rect 27052 22397 27092 22492
rect 26764 22364 26804 22373
rect 27148 22364 27188 24340
rect 27244 23792 27284 23801
rect 27244 23288 27284 23752
rect 27244 23239 27284 23248
rect 27148 22324 27284 22364
rect 26764 22280 26804 22324
rect 26764 22229 26804 22240
rect 26956 22196 26996 22205
rect 26956 21860 26996 22156
rect 27148 22196 27188 22205
rect 27148 22028 27188 22156
rect 27148 21979 27188 21988
rect 26956 21811 26996 21820
rect 26380 21643 26420 21652
rect 26434 21188 26802 21197
rect 26434 21139 26802 21148
rect 27244 21188 27284 22324
rect 27340 22280 27380 24592
rect 27436 24044 27476 24676
rect 27436 23995 27476 24004
rect 28108 23624 28148 25180
rect 28204 24044 28244 24053
rect 28204 23792 28244 24004
rect 28204 23743 28244 23752
rect 28108 23575 28148 23584
rect 28204 23540 28244 23549
rect 27674 23456 28042 23465
rect 27674 23407 28042 23416
rect 28204 23204 28244 23500
rect 28204 23155 28244 23164
rect 27340 21608 27380 22240
rect 27532 22364 27572 22373
rect 27532 21776 27572 22324
rect 27674 21944 28042 21953
rect 27674 21895 28042 21904
rect 27532 21727 27572 21736
rect 27436 21608 27476 21617
rect 27340 21568 27436 21608
rect 27244 21139 27284 21148
rect 27244 20936 27284 20945
rect 27244 20264 27284 20896
rect 27244 20215 27284 20224
rect 25324 19543 25364 19552
rect 25516 19592 25556 19601
rect 25708 19592 25748 19601
rect 25556 19552 25708 19592
rect 25516 19543 25556 19552
rect 25708 19543 25748 19552
rect 25036 19340 25076 19349
rect 24556 18955 24596 18964
rect 24844 19172 24884 19181
rect 24172 17828 24212 17837
rect 23636 17452 23732 17492
rect 23788 17744 23828 17753
rect 23500 16484 23540 16493
rect 23500 16316 23540 16444
rect 23500 16232 23540 16276
rect 23500 16181 23540 16192
rect 23596 16316 23636 17452
rect 23308 16015 23348 16024
rect 23500 16064 23540 16073
rect 23308 15728 23348 15737
rect 23308 15056 23348 15688
rect 23308 14804 23348 15016
rect 23308 14755 23348 14764
rect 23404 15476 23444 15485
rect 23212 14419 23252 14428
rect 23308 14468 23348 14477
rect 23116 13159 23156 13168
rect 23212 14300 23252 14309
rect 22540 12739 22580 12748
rect 22732 13124 22772 13133
rect 22732 12956 22772 13084
rect 23212 13124 23252 14260
rect 23308 13964 23348 14428
rect 23308 13915 23348 13924
rect 23404 14216 23444 15436
rect 23404 14048 23444 14176
rect 23308 13460 23348 13469
rect 23308 13292 23348 13420
rect 23308 13243 23348 13252
rect 23212 13075 23252 13084
rect 23404 13040 23444 14008
rect 23404 12991 23444 13000
rect 23500 15476 23540 16024
rect 23500 13796 23540 15436
rect 23596 14552 23636 16276
rect 23692 16148 23732 16157
rect 23692 15812 23732 16108
rect 23788 15896 23828 17704
rect 23788 15847 23828 15856
rect 23692 15763 23732 15772
rect 23596 14503 23636 14512
rect 23692 15644 23732 15653
rect 23692 14804 23732 15604
rect 23788 15560 23828 15571
rect 23788 15476 23828 15520
rect 23788 15427 23828 15436
rect 23884 15392 23924 15401
rect 23596 14384 23636 14393
rect 23596 14132 23636 14344
rect 23596 14083 23636 14092
rect 22540 12620 22580 12629
rect 22540 11780 22580 12580
rect 22732 11864 22772 12916
rect 23500 12620 23540 13756
rect 23596 13964 23636 13973
rect 23596 13208 23636 13924
rect 23692 13964 23732 14764
rect 23788 15056 23828 15065
rect 23788 14048 23828 15016
rect 23884 14720 23924 15352
rect 23884 14671 23924 14680
rect 23980 15308 24020 15317
rect 23884 14552 23924 14561
rect 23884 14216 23924 14512
rect 23884 14167 23924 14176
rect 23788 13999 23828 14008
rect 23884 14048 23924 14057
rect 23692 13460 23732 13924
rect 23692 13411 23732 13420
rect 23596 13073 23636 13168
rect 23788 13124 23828 13133
rect 23884 13124 23924 14008
rect 23980 13544 24020 15268
rect 23980 13495 24020 13504
rect 24076 14972 24116 14981
rect 24076 14804 24116 14932
rect 23828 13084 23924 13124
rect 23980 13124 24020 13219
rect 23788 13075 23828 13084
rect 23980 13075 24020 13084
rect 23500 12571 23540 12580
rect 23116 12443 23156 12463
rect 23116 12368 23156 12403
rect 23116 12319 23156 12328
rect 23404 12452 23444 12461
rect 23404 12317 23444 12412
rect 23596 12284 23636 12293
rect 22732 11815 22772 11824
rect 22828 12116 22868 12125
rect 22540 11731 22580 11740
rect 22348 10940 22388 10949
rect 22348 8000 22388 10900
rect 22444 8252 22484 11068
rect 22732 10856 22772 10865
rect 22732 10100 22772 10816
rect 22732 10051 22772 10060
rect 22540 10016 22580 10025
rect 22540 9512 22580 9976
rect 22828 9680 22868 12076
rect 23596 11780 23636 12244
rect 23884 11780 23924 11789
rect 23596 11731 23636 11740
rect 23788 11740 23884 11780
rect 23308 11444 23348 11453
rect 23308 10184 23348 11404
rect 23788 11192 23828 11740
rect 23884 11731 23924 11740
rect 23788 11143 23828 11152
rect 23308 10135 23348 10144
rect 22828 9631 22868 9640
rect 23884 10016 23924 10025
rect 22540 9463 22580 9472
rect 23308 9512 23348 9521
rect 23116 8672 23156 8681
rect 22444 8084 22484 8212
rect 22444 8035 22484 8044
rect 22732 8504 22772 8513
rect 22348 7916 22388 7960
rect 22060 7160 22100 7169
rect 22060 6992 22100 7120
rect 22060 6943 22100 6952
rect 22252 7160 22292 7169
rect 22252 6656 22292 7120
rect 22252 6607 22292 6616
rect 21964 5767 22004 5776
rect 22348 5144 22388 7876
rect 22636 8000 22676 8009
rect 22636 7865 22676 7960
rect 22540 7832 22580 7841
rect 22540 7160 22580 7792
rect 22540 7111 22580 7120
rect 22732 6824 22772 8464
rect 22348 5095 22388 5104
rect 22636 5900 22676 5909
rect 22636 5060 22676 5860
rect 22732 5648 22772 6784
rect 22828 7916 22868 7925
rect 22828 7160 22868 7876
rect 23116 7832 23156 8632
rect 23020 7748 23060 7757
rect 23020 7244 23060 7708
rect 23116 7328 23156 7792
rect 23116 7279 23156 7288
rect 23212 8252 23252 8261
rect 23020 7195 23060 7204
rect 22828 6404 22868 7120
rect 22828 6355 22868 6364
rect 22732 5599 22772 5608
rect 22636 4976 22676 5020
rect 22636 4925 22676 4936
rect 22828 5228 22868 5237
rect 22828 4892 22868 5188
rect 23212 5060 23252 8212
rect 23308 8168 23348 9472
rect 23596 8756 23636 8765
rect 23596 8621 23636 8716
rect 23884 8756 23924 9976
rect 24076 9428 24116 14764
rect 24172 14216 24212 17788
rect 24460 17744 24500 18712
rect 24844 18332 24884 19132
rect 24940 19088 24980 19097
rect 24940 18668 24980 19048
rect 24940 18619 24980 18628
rect 24844 18283 24884 18292
rect 24460 17156 24500 17704
rect 24460 17107 24500 17116
rect 24940 17660 24980 17669
rect 24556 17072 24596 17081
rect 24364 16988 24404 16997
rect 24556 16988 24596 17032
rect 24404 16948 24596 16988
rect 24844 16988 24884 16997
rect 24364 16939 24404 16948
rect 24748 16820 24788 16829
rect 24556 16148 24596 16157
rect 24172 14167 24212 14176
rect 24268 16064 24308 16073
rect 24268 15812 24308 16024
rect 24172 13628 24212 13639
rect 24172 13544 24212 13588
rect 24172 13495 24212 13504
rect 24268 13124 24308 15772
rect 24364 15392 24404 15401
rect 24364 14048 24404 15352
rect 24364 13999 24404 14008
rect 24556 13292 24596 16108
rect 24748 15560 24788 16780
rect 24844 16316 24884 16948
rect 24844 16267 24884 16276
rect 24940 15728 24980 17620
rect 25036 16988 25076 19300
rect 25324 19256 25364 19265
rect 25324 18500 25364 19216
rect 25324 18451 25364 18460
rect 25708 19004 25748 19013
rect 25708 17744 25748 18964
rect 25996 18836 26036 18845
rect 25708 17240 25748 17704
rect 25036 16939 25076 16948
rect 25132 17072 25172 17081
rect 24940 15679 24980 15688
rect 24748 15511 24788 15520
rect 25132 14720 25172 17032
rect 25324 17072 25364 17081
rect 25324 16652 25364 17032
rect 25228 16232 25268 16241
rect 25228 15476 25268 16192
rect 25228 15427 25268 15436
rect 25132 14671 25172 14680
rect 24652 14636 24692 14645
rect 24652 13460 24692 14596
rect 25324 14132 25364 16612
rect 25420 16568 25460 16577
rect 25420 16400 25460 16528
rect 25420 15560 25460 16360
rect 25420 15511 25460 15520
rect 25612 16316 25652 16325
rect 25324 14083 25364 14092
rect 25516 14552 25556 14561
rect 24748 14048 24788 14057
rect 24748 13964 24788 14008
rect 24748 13924 24884 13964
rect 24844 13880 24884 13924
rect 24844 13831 24884 13840
rect 24652 13411 24692 13420
rect 24748 13796 24788 13805
rect 24556 13243 24596 13252
rect 24748 13208 24788 13756
rect 25324 13796 25364 13805
rect 24748 13159 24788 13168
rect 24940 13292 24980 13301
rect 24172 11696 24212 11705
rect 24172 11024 24212 11656
rect 24172 10975 24212 10984
rect 24172 10268 24212 10277
rect 24172 9680 24212 10228
rect 24268 9764 24308 13084
rect 24460 13124 24500 13133
rect 24460 12872 24500 13084
rect 24460 12823 24500 12832
rect 24652 13124 24692 13133
rect 24364 12788 24404 12797
rect 24364 11612 24404 12748
rect 24364 11192 24404 11572
rect 24652 12284 24692 13084
rect 24940 12704 24980 13252
rect 25324 13208 25364 13756
rect 25324 13159 25364 13168
rect 24940 12452 24980 12664
rect 24940 12403 24980 12412
rect 25036 13124 25076 13133
rect 25036 13040 25076 13084
rect 25036 12452 25076 13000
rect 25420 13124 25460 13133
rect 25420 12956 25460 13084
rect 25420 12907 25460 12916
rect 25516 12704 25556 14512
rect 25516 12569 25556 12664
rect 25036 12403 25076 12412
rect 25420 12536 25460 12545
rect 24364 11143 24404 11152
rect 24460 11444 24500 11453
rect 24460 11024 24500 11404
rect 24460 10975 24500 10984
rect 24268 9715 24308 9724
rect 24172 9631 24212 9640
rect 24652 9512 24692 12244
rect 25420 12284 25460 12496
rect 25420 12235 25460 12244
rect 24940 11528 24980 11537
rect 24940 10184 24980 11488
rect 25324 11192 25364 11201
rect 24940 10135 24980 10144
rect 25228 10772 25268 10781
rect 25228 10184 25268 10732
rect 24652 9463 24692 9472
rect 25228 9512 25268 10144
rect 25228 9463 25268 9472
rect 24076 9379 24116 9388
rect 24556 9428 24596 9437
rect 24460 9344 24500 9353
rect 24076 8924 24116 8933
rect 23884 8707 23924 8716
rect 23980 8884 24076 8924
rect 23980 8672 24020 8884
rect 24076 8875 24116 8884
rect 23980 8623 24020 8632
rect 24364 8756 24404 8765
rect 24076 8588 24116 8597
rect 23308 8119 23348 8128
rect 23404 8504 23444 8513
rect 23404 8000 23444 8464
rect 23404 7951 23444 7960
rect 23596 8168 23636 8177
rect 23596 8000 23636 8128
rect 23596 7951 23636 7960
rect 23788 8000 23828 8009
rect 23308 7832 23348 7841
rect 23308 6992 23348 7792
rect 23500 7664 23540 7673
rect 23500 7076 23540 7624
rect 23788 7412 23828 7960
rect 24076 8000 24116 8548
rect 24076 7951 24116 7960
rect 24172 8000 24212 8009
rect 23788 7363 23828 7372
rect 23500 7027 23540 7036
rect 23788 7076 23828 7085
rect 23308 6943 23348 6952
rect 23596 6656 23636 6665
rect 23308 6488 23348 6497
rect 23308 5228 23348 6448
rect 23308 5179 23348 5188
rect 23212 5011 23252 5020
rect 22828 4843 22868 4852
rect 23596 4892 23636 6616
rect 23788 6656 23828 7036
rect 23788 6607 23828 6616
rect 23596 4843 23636 4852
rect 23884 6488 23924 6497
rect 21580 4759 21620 4768
rect 23884 4808 23924 6448
rect 24172 5900 24212 7960
rect 24364 7412 24404 8716
rect 24460 7916 24500 9304
rect 24556 8672 24596 9388
rect 24556 8623 24596 8632
rect 24844 9428 24884 9437
rect 24844 8672 24884 9388
rect 24844 8623 24884 8632
rect 24556 8168 24596 8177
rect 24556 8000 24596 8128
rect 24556 7951 24596 7960
rect 24844 8000 24884 8009
rect 24460 7867 24500 7876
rect 24364 7363 24404 7372
rect 24172 5851 24212 5860
rect 24268 7076 24308 7085
rect 24268 6488 24308 7036
rect 24268 5060 24308 6448
rect 24652 6320 24692 6329
rect 24652 5648 24692 6280
rect 24844 6236 24884 7960
rect 25132 7748 25172 7757
rect 24844 6187 24884 6196
rect 24940 6488 24980 6497
rect 24940 5900 24980 6448
rect 24940 5851 24980 5860
rect 24652 5599 24692 5608
rect 25132 5648 25172 7708
rect 25324 6152 25364 11152
rect 25612 10940 25652 16276
rect 25708 16316 25748 17200
rect 25900 17828 25940 17837
rect 25900 17240 25940 17788
rect 25900 17191 25940 17200
rect 25708 16267 25748 16276
rect 25900 16232 25940 16241
rect 25708 16064 25748 16073
rect 25708 15560 25748 16024
rect 25708 15511 25748 15520
rect 25900 15728 25940 16192
rect 25900 14972 25940 15688
rect 25900 14923 25940 14932
rect 25996 14216 26036 18796
rect 26284 18584 26324 20056
rect 27340 20012 27380 20021
rect 26860 19844 26900 19853
rect 26434 19676 26802 19685
rect 26434 19627 26802 19636
rect 26380 19340 26420 19435
rect 26860 19424 26900 19804
rect 26860 19375 26900 19384
rect 27148 19844 27188 19853
rect 26380 19291 26420 19300
rect 26284 18535 26324 18544
rect 26668 19256 26708 19265
rect 26668 19004 26708 19216
rect 26668 18332 26708 18964
rect 26668 18283 26708 18292
rect 27148 19256 27188 19804
rect 26434 18164 26802 18173
rect 26434 18115 26802 18124
rect 26092 17996 26132 18005
rect 26092 15560 26132 17956
rect 27052 17660 27092 17669
rect 27052 17525 27092 17620
rect 26284 16988 26324 16997
rect 26188 16820 26228 16829
rect 26188 16400 26228 16780
rect 26188 16351 26228 16360
rect 26092 15511 26132 15520
rect 26284 16232 26324 16948
rect 26434 16652 26802 16661
rect 26434 16603 26802 16612
rect 26860 16316 26900 16325
rect 26476 16232 26516 16241
rect 26284 16192 26476 16232
rect 25996 14167 26036 14176
rect 26284 15224 26324 16192
rect 26476 16183 26516 16192
rect 26764 16232 26804 16241
rect 26764 15560 26804 16192
rect 26860 16181 26900 16276
rect 26764 15511 26804 15520
rect 26956 15728 26996 15737
rect 25900 14132 25940 14141
rect 25708 14048 25748 14057
rect 25708 12536 25748 14008
rect 25900 13292 25940 14092
rect 25900 13243 25940 13252
rect 25804 12956 25844 12965
rect 25804 12620 25844 12916
rect 25900 12872 25940 12881
rect 25900 12704 25940 12832
rect 25900 12655 25940 12664
rect 26188 12704 26228 12713
rect 25804 12571 25844 12580
rect 25708 12487 25748 12496
rect 26188 12536 26228 12664
rect 25804 12452 25844 12461
rect 25804 11276 25844 12412
rect 25804 11227 25844 11236
rect 25900 11864 25940 11873
rect 25612 10891 25652 10900
rect 25900 9596 25940 11824
rect 26188 11192 26228 12496
rect 26284 12032 26324 15184
rect 26434 15140 26802 15149
rect 26434 15091 26802 15100
rect 26860 13964 26900 13973
rect 26434 13628 26802 13637
rect 26434 13579 26802 13588
rect 26764 13460 26804 13469
rect 26764 12536 26804 13420
rect 26860 12704 26900 13924
rect 26860 12655 26900 12664
rect 26956 12620 26996 15688
rect 27148 15056 27188 19216
rect 27148 14804 27188 15016
rect 27148 14755 27188 14764
rect 27244 18752 27284 18761
rect 27052 14048 27092 14059
rect 27052 13964 27092 14008
rect 27052 13915 27092 13924
rect 26956 12571 26996 12580
rect 27148 13208 27188 13217
rect 26764 12487 26804 12496
rect 27052 12536 27092 12545
rect 26434 12116 26802 12125
rect 26434 12067 26802 12076
rect 26284 11983 26324 11992
rect 26188 11143 26228 11152
rect 26956 11696 26996 11705
rect 26956 11024 26996 11656
rect 26956 10975 26996 10984
rect 26434 10604 26802 10613
rect 26434 10555 26802 10564
rect 27052 10268 27092 12496
rect 27148 11696 27188 13168
rect 27244 12620 27284 18712
rect 27340 18416 27380 19972
rect 27436 19340 27476 21568
rect 28300 21188 28340 26692
rect 28396 26648 28436 26860
rect 28396 26599 28436 26608
rect 28396 26480 28436 26489
rect 28396 25136 28436 26440
rect 28396 25087 28436 25096
rect 28396 24380 28436 24389
rect 28396 23624 28436 24340
rect 28396 23575 28436 23584
rect 28492 21524 28532 27532
rect 28780 27572 28820 27581
rect 28780 27437 28820 27532
rect 28780 26984 28820 26993
rect 28876 26984 28916 28120
rect 28820 26944 28916 26984
rect 28780 26935 28820 26944
rect 28588 26816 28628 26825
rect 28588 25976 28628 26776
rect 28972 26816 29012 28372
rect 29260 27740 29300 28600
rect 30028 28580 30068 28600
rect 30028 28531 30068 28540
rect 30028 28244 30068 28253
rect 29260 27691 29300 27700
rect 29836 27740 29876 27749
rect 29260 27572 29300 27581
rect 29260 27437 29300 27532
rect 29644 27152 29684 27163
rect 29644 27068 29684 27112
rect 29644 27019 29684 27028
rect 29740 27068 29780 27077
rect 28972 26767 29012 26776
rect 29260 26984 29300 26993
rect 28780 26648 28820 26657
rect 28588 25927 28628 25936
rect 28684 26228 28724 26237
rect 28684 26060 28724 26188
rect 28780 26228 28820 26608
rect 29164 26480 29204 26489
rect 28780 26179 28820 26188
rect 28972 26228 29012 26237
rect 28972 26144 29012 26188
rect 28972 26093 29012 26104
rect 28588 25808 28628 25817
rect 28588 25388 28628 25768
rect 28684 25472 28724 26020
rect 28876 25892 28916 25901
rect 28876 25556 28916 25852
rect 29164 25808 29204 26440
rect 29164 25759 29204 25768
rect 28876 25507 28916 25516
rect 28684 25423 28724 25432
rect 28588 25339 28628 25348
rect 28876 25388 28916 25397
rect 28780 25304 28820 25313
rect 28780 24548 28820 25264
rect 28876 24800 28916 25348
rect 28972 25052 29012 25061
rect 28972 24917 29012 25012
rect 29164 25052 29204 25061
rect 29164 24884 29204 25012
rect 29164 24835 29204 24844
rect 28876 24751 28916 24760
rect 29260 24632 29300 26944
rect 29356 26900 29396 26909
rect 29356 26765 29396 26860
rect 29548 26900 29588 26909
rect 29356 26564 29396 26573
rect 29356 26060 29396 26524
rect 29356 25640 29396 26020
rect 29452 25976 29492 25985
rect 29452 25841 29492 25936
rect 29548 25892 29588 26860
rect 29356 25591 29396 25600
rect 29452 25556 29492 25565
rect 29260 24583 29300 24592
rect 29356 25472 29396 25481
rect 28684 24380 28724 24389
rect 28588 23456 28628 23465
rect 28588 23120 28628 23416
rect 28588 23071 28628 23080
rect 28492 21475 28532 21484
rect 27436 19291 27476 19300
rect 27532 20768 27572 20777
rect 27532 19172 27572 20728
rect 28108 20684 28148 20693
rect 27674 20432 28042 20441
rect 27674 20383 28042 20392
rect 28108 20012 28148 20644
rect 28300 20600 28340 21148
rect 28684 20684 28724 24340
rect 28780 22868 28820 24508
rect 29068 24548 29108 24557
rect 28972 24128 29012 24137
rect 28876 24044 28916 24053
rect 28876 23708 28916 24004
rect 28876 23659 28916 23668
rect 28972 23708 29012 24088
rect 28972 23659 29012 23668
rect 29068 23792 29108 24508
rect 29260 24464 29300 24473
rect 29164 24212 29204 24221
rect 29164 23876 29204 24172
rect 29164 23827 29204 23836
rect 28876 23540 28916 23549
rect 28876 23405 28916 23500
rect 28780 22819 28820 22828
rect 28972 23120 29012 23129
rect 28972 22532 29012 23080
rect 28972 22483 29012 22492
rect 28780 22280 28820 22289
rect 28780 21608 28820 22240
rect 28780 21559 28820 21568
rect 28972 21860 29012 21869
rect 28684 20635 28724 20644
rect 28972 20684 29012 21820
rect 28300 20551 28340 20560
rect 28108 19963 28148 19972
rect 28204 20096 28244 20105
rect 28204 19508 28244 20056
rect 27436 19132 27572 19172
rect 28108 19468 28244 19508
rect 28588 20096 28628 20105
rect 27436 18752 27476 19132
rect 27436 18703 27476 18712
rect 27532 19004 27572 19013
rect 27532 18584 27572 18964
rect 27674 18920 28042 18929
rect 27674 18871 28042 18880
rect 27532 18535 27572 18544
rect 28108 18500 28148 19468
rect 28588 18584 28628 20056
rect 28684 19424 28724 19433
rect 28684 18668 28724 19384
rect 28684 18619 28724 18628
rect 28588 18535 28628 18544
rect 28780 18584 28820 18593
rect 28108 18451 28148 18460
rect 28780 18449 28820 18544
rect 28972 18500 29012 20644
rect 29068 20096 29108 23752
rect 29164 23624 29204 23633
rect 29164 23489 29204 23584
rect 29164 23372 29204 23381
rect 29164 23204 29204 23332
rect 29164 23155 29204 23164
rect 29260 23036 29300 24424
rect 29260 22987 29300 22996
rect 29164 22952 29204 22961
rect 29164 22817 29204 22912
rect 29356 22364 29396 25432
rect 29452 25388 29492 25516
rect 29452 25339 29492 25348
rect 29452 24380 29492 24389
rect 29452 23120 29492 24340
rect 29548 24296 29588 25852
rect 29644 26900 29684 26909
rect 29644 26144 29684 26860
rect 29740 26312 29780 27028
rect 29740 26263 29780 26272
rect 29644 25556 29684 26104
rect 29644 25507 29684 25516
rect 29836 25472 29876 27700
rect 29932 27488 29972 27497
rect 29932 27353 29972 27448
rect 29932 26900 29972 26909
rect 29932 25640 29972 26860
rect 30028 26060 30068 28204
rect 30796 27656 30836 28600
rect 30796 27607 30836 27616
rect 30988 27572 31028 27581
rect 30220 27488 30260 27497
rect 30028 26011 30068 26020
rect 30124 26648 30164 26657
rect 30028 25892 30068 25901
rect 30028 25757 30068 25852
rect 29932 25591 29972 25600
rect 29836 25432 29972 25472
rect 29836 24716 29876 24725
rect 29548 24247 29588 24256
rect 29644 24632 29684 24641
rect 29644 24044 29684 24592
rect 29644 23995 29684 24004
rect 29740 24128 29780 24137
rect 29548 23876 29588 23885
rect 29548 23624 29588 23836
rect 29644 23792 29684 23887
rect 29644 23743 29684 23752
rect 29548 23575 29588 23584
rect 29644 23540 29684 23549
rect 29452 23071 29492 23080
rect 29548 23456 29588 23465
rect 29356 22315 29396 22324
rect 29548 22112 29588 23416
rect 29644 22952 29684 23500
rect 29740 23120 29780 24088
rect 29740 23071 29780 23080
rect 29836 23624 29876 24676
rect 29644 22903 29684 22912
rect 29548 22063 29588 22072
rect 29836 22196 29876 23584
rect 29260 21188 29300 21197
rect 29164 20768 29204 20777
rect 29164 20180 29204 20728
rect 29164 20131 29204 20140
rect 29068 20047 29108 20056
rect 29164 19172 29204 19183
rect 29164 19088 29204 19132
rect 29164 19039 29204 19048
rect 29260 18584 29300 21148
rect 29548 20852 29588 20861
rect 29548 19928 29588 20812
rect 29836 20096 29876 22156
rect 29932 20936 29972 25432
rect 30124 25220 30164 26608
rect 30220 25388 30260 27448
rect 30988 27320 31028 27532
rect 30988 27271 31028 27280
rect 30316 26900 30356 26909
rect 30316 26480 30356 26860
rect 30316 26431 30356 26440
rect 30412 26564 30452 26573
rect 30412 26144 30452 26524
rect 30988 26396 31028 26407
rect 30604 26312 30644 26321
rect 30604 26177 30644 26272
rect 30988 26312 31028 26356
rect 30988 26263 31028 26272
rect 30412 26095 30452 26104
rect 30220 25339 30260 25348
rect 30220 25220 30260 25229
rect 30124 25180 30220 25220
rect 30124 24632 30164 24641
rect 30028 24380 30068 24389
rect 30028 23036 30068 24340
rect 30028 22987 30068 22996
rect 30124 22784 30164 24592
rect 30220 23876 30260 25180
rect 30988 24464 31028 24473
rect 30988 24329 31028 24424
rect 30220 23827 30260 23836
rect 30508 23960 30548 23969
rect 30028 22280 30068 22375
rect 30124 22364 30164 22744
rect 30316 23708 30356 23717
rect 30316 22448 30356 23668
rect 30316 22399 30356 22408
rect 30412 22952 30452 22961
rect 30124 22315 30164 22324
rect 30028 22231 30068 22240
rect 30028 22112 30068 22121
rect 30028 21977 30068 22072
rect 30028 21776 30068 21785
rect 30028 21020 30068 21736
rect 30316 21440 30356 21449
rect 30316 21188 30356 21400
rect 30316 21139 30356 21148
rect 30028 20971 30068 20980
rect 29932 20887 29972 20896
rect 29932 20768 29972 20777
rect 29932 20264 29972 20728
rect 29932 20215 29972 20224
rect 30220 20684 30260 20693
rect 30220 20180 30260 20644
rect 30412 20516 30452 22912
rect 30508 22280 30548 23920
rect 30988 23624 31028 23633
rect 30508 22231 30548 22240
rect 30604 22448 30644 22457
rect 30604 21356 30644 22408
rect 30796 22448 30836 22457
rect 30604 21307 30644 21316
rect 30700 22280 30740 22289
rect 30508 21272 30548 21281
rect 30508 20768 30548 21232
rect 30604 21020 30644 21029
rect 30604 20885 30644 20980
rect 30508 20719 30548 20728
rect 30412 20467 30452 20476
rect 30700 20348 30740 22240
rect 30796 21524 30836 22408
rect 30988 21608 31028 23584
rect 30988 21559 31028 21568
rect 30796 21475 30836 21484
rect 30892 21440 30932 21449
rect 30892 21305 30932 21400
rect 30892 20936 30932 20945
rect 30892 20801 30932 20896
rect 30700 20299 30740 20308
rect 30220 20131 30260 20140
rect 29836 20047 29876 20056
rect 29548 19879 29588 19888
rect 29932 19928 29972 19937
rect 29932 19793 29972 19888
rect 29548 19088 29588 19097
rect 29548 18953 29588 19048
rect 29260 18535 29300 18544
rect 28972 18451 29012 18460
rect 27340 18367 27380 18376
rect 28684 18416 28724 18425
rect 27628 18332 27668 18341
rect 27628 18197 27668 18292
rect 28684 18281 28724 18376
rect 27436 17912 27476 17921
rect 27340 17576 27380 17585
rect 27340 17156 27380 17536
rect 27340 17107 27380 17116
rect 27436 16988 27476 17872
rect 28012 17912 28052 17921
rect 27532 17828 27572 17837
rect 27532 17240 27572 17788
rect 28012 17777 28052 17872
rect 27674 17408 28042 17417
rect 27674 17359 28042 17368
rect 28492 17240 28532 17249
rect 27532 17200 27668 17240
rect 27436 16939 27476 16948
rect 27532 17072 27572 17081
rect 27532 15644 27572 17032
rect 27628 16316 27668 17200
rect 27628 16267 27668 16276
rect 28108 16820 28148 16829
rect 28108 16064 28148 16780
rect 28300 16484 28340 16493
rect 28300 16232 28340 16444
rect 28300 16183 28340 16192
rect 28108 16015 28148 16024
rect 28492 16064 28532 17200
rect 28492 16015 28532 16024
rect 28780 16400 28820 16409
rect 27674 15896 28042 15905
rect 27674 15847 28042 15856
rect 27532 15595 27572 15604
rect 28300 15812 28340 15821
rect 27820 15560 27860 15569
rect 27820 14636 27860 15520
rect 28108 15560 28148 15569
rect 28108 15425 28148 15520
rect 28300 15476 28340 15772
rect 28780 15812 28820 16360
rect 28780 15763 28820 15772
rect 28300 15427 28340 15436
rect 28396 15560 28436 15569
rect 28396 14972 28436 15520
rect 28780 15560 28820 15569
rect 28396 14923 28436 14932
rect 28492 15476 28532 15485
rect 27820 14587 27860 14596
rect 27674 14384 28042 14393
rect 27674 14335 28042 14344
rect 27532 14048 27572 14057
rect 27532 13208 27572 14008
rect 27532 13159 27572 13168
rect 28396 13292 28436 13301
rect 28204 13124 28244 13133
rect 27340 13040 27380 13049
rect 27340 12704 27380 13000
rect 27674 12872 28042 12881
rect 27674 12823 28042 12832
rect 27340 12655 27380 12664
rect 28204 12704 28244 13084
rect 28204 12655 28244 12664
rect 27244 12571 27284 12580
rect 27436 12620 27476 12629
rect 27244 12452 27284 12461
rect 27244 12368 27284 12412
rect 27436 12452 27476 12580
rect 27436 12403 27476 12412
rect 27820 12536 27860 12545
rect 27820 12401 27860 12496
rect 27916 12452 27956 12461
rect 27244 12317 27284 12328
rect 27916 12317 27956 12412
rect 28108 12452 28148 12461
rect 27532 12284 27572 12293
rect 27148 11647 27188 11656
rect 27436 11696 27476 11705
rect 27436 11276 27476 11656
rect 27532 11528 27572 12244
rect 28108 12284 28148 12412
rect 28108 12235 28148 12244
rect 28204 12368 28244 12377
rect 27724 12200 27764 12209
rect 27628 11864 27668 11873
rect 27628 11729 27668 11824
rect 27724 11780 27764 12160
rect 27916 12032 27956 12041
rect 27916 11864 27956 11992
rect 27916 11815 27956 11824
rect 28204 11864 28244 12328
rect 28396 12368 28436 13252
rect 28396 12319 28436 12328
rect 28492 12956 28532 15436
rect 28684 14720 28724 14729
rect 28684 13376 28724 14680
rect 28780 13544 28820 15520
rect 28972 15308 29012 15317
rect 28876 14888 28916 14897
rect 28876 13880 28916 14848
rect 28876 13831 28916 13840
rect 28780 13495 28820 13504
rect 28684 13327 28724 13336
rect 28780 13292 28820 13301
rect 28780 13157 28820 13252
rect 28972 13208 29012 15268
rect 29836 14888 29876 14897
rect 29644 14720 29684 14729
rect 29644 14216 29684 14680
rect 29644 14167 29684 14176
rect 29836 13964 29876 14848
rect 29836 13915 29876 13924
rect 29068 13796 29108 13805
rect 29068 13661 29108 13756
rect 28972 13159 29012 13168
rect 28204 11815 28244 11824
rect 27724 11731 27764 11740
rect 27532 11479 27572 11488
rect 27674 11360 28042 11369
rect 27674 11311 28042 11320
rect 27436 11227 27476 11236
rect 28492 11024 28532 12916
rect 28876 12368 28916 12377
rect 28876 11948 28916 12328
rect 28876 11899 28916 11908
rect 28492 10975 28532 10984
rect 27148 10940 27188 10949
rect 27148 10352 27188 10900
rect 27148 10303 27188 10312
rect 27340 10940 27380 10949
rect 27052 10219 27092 10228
rect 25996 10184 26036 10193
rect 25996 9680 26036 10144
rect 25996 9631 26036 9640
rect 26092 10016 26132 10025
rect 25900 9547 25940 9556
rect 25996 9512 26036 9521
rect 25996 9377 26036 9472
rect 26092 9428 26132 9976
rect 26284 10016 26324 10025
rect 26284 9512 26324 9976
rect 27340 9680 27380 10900
rect 27674 9848 28042 9857
rect 27674 9799 28042 9808
rect 27340 9631 27380 9640
rect 26284 9463 26324 9472
rect 26092 9379 26132 9388
rect 25708 9344 25748 9353
rect 25708 8672 25748 9304
rect 26434 9092 26802 9101
rect 26434 9043 26802 9052
rect 26572 8756 26612 8765
rect 25900 8672 25940 8681
rect 25708 8623 25748 8632
rect 25804 8632 25900 8672
rect 25612 8084 25652 8124
rect 25612 8000 25652 8044
rect 25612 7496 25652 7960
rect 25612 7447 25652 7456
rect 25324 6103 25364 6112
rect 25804 6488 25844 8632
rect 25900 8537 25940 8632
rect 26476 8672 26516 8681
rect 26476 8504 26516 8632
rect 26572 8621 26612 8716
rect 27052 8672 27092 8681
rect 27052 8537 27092 8632
rect 26476 8455 26516 8464
rect 27674 8336 28042 8345
rect 27674 8287 28042 8296
rect 25900 8168 25940 8177
rect 25900 7832 25940 8128
rect 26284 8168 26324 8177
rect 25900 7783 25940 7792
rect 25996 8084 26036 8093
rect 25996 7664 26036 8044
rect 26284 8033 26324 8128
rect 26380 8084 26420 8093
rect 26380 7949 26420 8044
rect 26860 8000 26900 8009
rect 25996 7615 26036 7624
rect 26188 7916 26228 7925
rect 25804 5816 25844 6448
rect 25804 5767 25844 5776
rect 25132 5599 25172 5608
rect 24268 5011 24308 5020
rect 23884 4759 23924 4768
rect 26188 4724 26228 7876
rect 26764 7916 26804 7925
rect 26764 7781 26804 7876
rect 26860 7865 26900 7960
rect 26434 7580 26802 7589
rect 26434 7531 26802 7540
rect 27674 6824 28042 6833
rect 27674 6775 28042 6784
rect 26434 6068 26802 6077
rect 26434 6019 26802 6028
rect 27674 5312 28042 5321
rect 27674 5263 28042 5272
rect 26188 4675 26228 4684
rect 26434 4556 26802 4565
rect 26434 4507 26802 4516
rect 21292 4171 21332 4180
rect 21004 4003 21044 4012
rect 4352 3800 4720 3809
rect 4352 3751 4720 3760
rect 12126 3800 12494 3809
rect 12126 3751 12494 3760
rect 19900 3800 20268 3809
rect 19900 3751 20268 3760
rect 27674 3800 28042 3809
rect 27674 3751 28042 3760
rect 3112 3044 3480 3053
rect 3112 2995 3480 3004
rect 10886 3044 11254 3053
rect 10886 2995 11254 3004
rect 18660 3044 19028 3053
rect 18660 2995 19028 3004
rect 26434 3044 26802 3053
rect 26434 2995 26802 3004
rect 4352 2288 4720 2297
rect 4352 2239 4720 2248
rect 12126 2288 12494 2297
rect 12126 2239 12494 2248
rect 19900 2288 20268 2297
rect 19900 2239 20268 2248
rect 27674 2288 28042 2297
rect 27674 2239 28042 2248
rect 3112 1532 3480 1541
rect 3112 1483 3480 1492
rect 10886 1532 11254 1541
rect 10886 1483 11254 1492
rect 18660 1532 19028 1541
rect 18660 1483 19028 1492
rect 26434 1532 26802 1541
rect 26434 1483 26802 1492
rect 4352 776 4720 785
rect 4352 727 4720 736
rect 12126 776 12494 785
rect 12126 727 12494 736
rect 19900 776 20268 785
rect 19900 727 20268 736
rect 27674 776 28042 785
rect 27674 727 28042 736
<< via3 >>
rect 1132 26608 1172 26648
rect 1036 26356 1076 26396
rect 1228 26272 1268 26312
rect 844 26104 884 26144
rect 652 25600 692 25640
rect 76 20476 116 20516
rect 76 13840 116 13880
rect 1420 26020 1460 26060
rect 940 23836 980 23876
rect 1036 24592 1076 24632
rect 748 20812 788 20852
rect 556 20560 596 20600
rect 556 20308 596 20348
rect 652 18208 692 18248
rect 364 17956 404 17996
rect 460 18124 500 18164
rect 364 17284 404 17324
rect 652 17956 692 17996
rect 652 17368 692 17408
rect 556 13840 596 13880
rect 460 8044 500 8084
rect 268 7288 308 7328
rect 1036 21484 1076 21524
rect 1420 24088 1460 24128
rect 1804 26524 1844 26564
rect 1708 24508 1748 24548
rect 1804 24088 1844 24128
rect 2092 27700 2132 27740
rect 3148 28036 3188 28076
rect 2956 27784 2996 27824
rect 2572 27532 2612 27572
rect 2380 27364 2420 27404
rect 2284 27028 2324 27068
rect 2092 25852 2132 25892
rect 2476 26860 2516 26900
rect 3340 27448 3380 27488
rect 3112 27196 3480 27236
rect 3628 27196 3668 27236
rect 3724 27364 3764 27404
rect 2668 26188 2708 26228
rect 2668 25936 2708 25976
rect 2572 25180 2612 25220
rect 1900 23920 1940 23960
rect 1708 21484 1748 21524
rect 1132 20980 1172 21020
rect 1228 20224 1268 20264
rect 940 18460 980 18500
rect 940 17872 980 17912
rect 844 17368 884 17408
rect 1132 19552 1172 19592
rect 1132 17956 1172 17996
rect 1132 17200 1172 17240
rect 1228 16948 1268 16988
rect 940 12412 980 12452
rect 844 9724 884 9764
rect 1228 10144 1268 10184
rect 652 7624 692 7664
rect 940 8128 980 8168
rect 1036 7288 1076 7328
rect 748 6784 788 6824
rect 1228 7036 1268 7076
rect 1516 20812 1556 20852
rect 1516 20056 1556 20096
rect 1804 20896 1844 20936
rect 1900 20140 1940 20180
rect 1708 19972 1748 20012
rect 1708 18712 1748 18752
rect 1996 19804 2036 19844
rect 1900 19132 1940 19172
rect 1708 18292 1748 18332
rect 1804 18208 1844 18248
rect 1708 17788 1748 17828
rect 1804 17452 1844 17492
rect 2092 18292 2132 18332
rect 2188 17788 2228 17828
rect 2380 21064 2420 21104
rect 2668 23836 2708 23876
rect 3628 26944 3668 26984
rect 3148 26692 3188 26732
rect 3436 26020 3476 26060
rect 3112 25684 3480 25724
rect 3628 26020 3668 26060
rect 3148 25264 3188 25304
rect 3340 24508 3380 24548
rect 4684 28120 4724 28160
rect 4352 27952 4720 27992
rect 4396 27616 4436 27656
rect 3916 27364 3956 27404
rect 3820 26188 3860 26228
rect 3112 24172 3480 24212
rect 2764 23752 2804 23792
rect 2860 23164 2900 23204
rect 3724 24340 3764 24380
rect 3052 23164 3092 23204
rect 3340 22996 3380 23036
rect 3532 22912 3572 22952
rect 3112 22660 3480 22700
rect 2860 22072 2900 22112
rect 3436 21988 3476 22028
rect 2668 21568 2708 21608
rect 2572 21400 2612 21440
rect 2956 21484 2996 21524
rect 2860 21232 2900 21272
rect 3436 21316 3476 21356
rect 3112 21148 3480 21188
rect 2572 19300 2612 19340
rect 2476 18880 2516 18920
rect 2476 18376 2516 18416
rect 2380 17872 2420 17912
rect 2284 17704 2324 17744
rect 1420 16024 1460 16064
rect 1708 15688 1748 15728
rect 1420 15436 1460 15476
rect 1900 16948 1940 16988
rect 1996 17116 2036 17156
rect 1996 15604 2036 15644
rect 1612 14092 1652 14132
rect 1708 12412 1748 12452
rect 1612 10228 1652 10268
rect 2860 20728 2900 20768
rect 3148 20224 3188 20264
rect 2860 18964 2900 19004
rect 3244 20140 3284 20180
rect 3436 20392 3476 20432
rect 3112 19636 3480 19676
rect 3916 24424 3956 24464
rect 3820 23080 3860 23120
rect 3916 23164 3956 23204
rect 3724 21652 3764 21692
rect 3628 21484 3668 21524
rect 3148 19132 3188 19172
rect 2668 18700 2708 18740
rect 2860 18628 2900 18668
rect 3340 18880 3380 18920
rect 3052 18460 3092 18500
rect 2860 18376 2900 18416
rect 2764 18292 2804 18332
rect 2956 18292 2996 18332
rect 2668 17956 2708 17996
rect 2860 17704 2900 17744
rect 2668 17620 2708 17660
rect 3436 18292 3476 18332
rect 3532 19132 3572 19172
rect 3112 18124 3480 18164
rect 3244 17704 3284 17744
rect 2860 17452 2900 17492
rect 2476 17116 2516 17156
rect 2284 16948 2324 16988
rect 2572 16948 2612 16988
rect 2380 16780 2420 16820
rect 2380 16192 2420 16232
rect 2284 15604 2324 15644
rect 2764 16024 2804 16064
rect 3820 21232 3860 21272
rect 3724 20644 3764 20684
rect 3724 20140 3764 20180
rect 3724 19720 3764 19760
rect 3820 19216 3860 19256
rect 3724 18208 3764 18248
rect 3628 17704 3668 17744
rect 3724 17788 3764 17828
rect 3532 17620 3572 17660
rect 3112 16612 3480 16652
rect 3820 16360 3860 16400
rect 3820 16108 3860 16148
rect 3724 15772 3764 15812
rect 2476 15184 2516 15224
rect 2572 15016 2612 15056
rect 2668 15184 2708 15224
rect 3112 15100 3480 15140
rect 2380 14092 2420 14132
rect 1900 11656 1940 11696
rect 1804 7960 1844 8000
rect 1900 7120 1940 7160
rect 2092 10228 2132 10268
rect 2092 7876 2132 7916
rect 2380 11740 2420 11780
rect 2380 10984 2420 11024
rect 2476 10312 2516 10352
rect 2284 6616 2324 6656
rect 3436 13756 3476 13796
rect 3628 13756 3668 13796
rect 3112 13588 3480 13628
rect 3112 12076 3480 12116
rect 3340 11152 3380 11192
rect 3628 11068 3668 11108
rect 4972 27280 5012 27320
rect 4492 26776 4532 26816
rect 4352 26440 4720 26480
rect 4108 25180 4148 25220
rect 4352 24928 4720 24968
rect 4492 24760 4532 24800
rect 4204 24592 4244 24632
rect 4396 24592 4436 24632
rect 4972 24928 5012 24968
rect 5068 24844 5108 24884
rect 4300 23584 4340 23624
rect 4352 23416 4720 23456
rect 4108 23248 4148 23288
rect 4300 23080 4340 23120
rect 4108 22996 4148 23036
rect 4588 22660 4628 22700
rect 4108 22156 4148 22196
rect 4396 22240 4436 22280
rect 5068 22996 5108 23036
rect 4876 22660 4916 22700
rect 5260 26440 5300 26480
rect 5452 26272 5492 26312
rect 6220 27868 6260 27908
rect 5644 27616 5684 27656
rect 5356 26104 5396 26144
rect 5260 25768 5300 25808
rect 5260 24592 5300 24632
rect 5164 22576 5204 22616
rect 4588 22072 4628 22112
rect 4698 22072 4724 22112
rect 4724 22072 4738 22112
rect 4012 20140 4052 20180
rect 4352 21904 4720 21944
rect 4780 21820 4820 21860
rect 4492 21736 4532 21776
rect 4876 21568 4916 21608
rect 4588 21484 4628 21524
rect 4972 22240 5012 22280
rect 5068 21904 5108 21944
rect 5164 21736 5204 21776
rect 5164 21568 5204 21608
rect 4204 21232 4244 21272
rect 4300 21148 4340 21188
rect 4876 21148 4916 21188
rect 4204 21064 4244 21104
rect 4352 20392 4720 20432
rect 4492 20224 4532 20264
rect 4396 19972 4436 20012
rect 4492 19804 4532 19844
rect 4204 19720 4244 19760
rect 4876 19384 4916 19424
rect 4972 20560 5012 20600
rect 5164 21064 5204 21104
rect 5164 20560 5204 20600
rect 5068 20140 5108 20180
rect 4972 19468 5012 19508
rect 4396 19216 4436 19256
rect 4588 19132 4628 19172
rect 4352 18880 4720 18920
rect 4204 18796 4244 18836
rect 4972 18964 5012 19004
rect 4876 17872 4916 17912
rect 4204 17704 4244 17744
rect 4780 17452 4820 17492
rect 4876 17536 4916 17576
rect 4352 17368 4720 17408
rect 4780 17116 4820 17156
rect 4876 16528 4916 16568
rect 4012 15688 4052 15728
rect 4108 15604 4148 15644
rect 3112 10564 3480 10604
rect 3820 10732 3860 10772
rect 2956 10228 2996 10268
rect 2860 9976 2900 10016
rect 3628 10312 3668 10352
rect 3436 10144 3476 10184
rect 3820 10144 3860 10184
rect 3112 9052 3480 9092
rect 3052 7708 3092 7748
rect 3112 7540 3480 7580
rect 3052 7120 3092 7160
rect 3820 9472 3860 9512
rect 3820 8128 3860 8168
rect 3112 6028 3480 6068
rect 4492 16276 4532 16316
rect 4684 16276 4724 16316
rect 4684 16108 4724 16148
rect 4352 15856 4720 15896
rect 4396 15520 4436 15560
rect 4204 14932 4244 14972
rect 4204 14764 4244 14804
rect 4588 15100 4628 15140
rect 4108 14428 4148 14468
rect 4588 14512 4628 14552
rect 4108 14260 4148 14300
rect 4352 14344 4720 14384
rect 5164 19720 5204 19760
rect 5164 18712 5204 18752
rect 5068 17620 5108 17660
rect 5068 17284 5108 17324
rect 5068 16444 5108 16484
rect 4300 13840 4340 13880
rect 4684 13084 4724 13124
rect 4352 12832 4720 12872
rect 4396 12664 4436 12704
rect 4300 12496 4340 12536
rect 4108 11068 4148 11108
rect 4492 12580 4532 12620
rect 4352 11320 4720 11360
rect 4684 11152 4724 11192
rect 4588 11068 4628 11108
rect 4396 10984 4436 11024
rect 4492 10228 4532 10268
rect 4396 10144 4436 10184
rect 5164 15856 5204 15896
rect 5164 15268 5204 15308
rect 5452 26020 5492 26060
rect 6220 27616 6260 27656
rect 5932 27448 5972 27488
rect 5740 25600 5780 25640
rect 5548 22660 5588 22700
rect 5644 21400 5684 21440
rect 5836 23668 5876 23708
rect 5740 21148 5780 21188
rect 5740 20308 5780 20348
rect 5644 20140 5684 20180
rect 5836 20140 5876 20180
rect 5452 19972 5492 20012
rect 5452 19384 5492 19424
rect 5452 18712 5492 18752
rect 5740 19720 5780 19760
rect 5644 19300 5684 19340
rect 5740 18964 5780 19004
rect 5452 17452 5492 17492
rect 5548 17368 5588 17408
rect 5836 17284 5876 17324
rect 5740 17200 5780 17240
rect 5452 16948 5492 16988
rect 5548 16864 5588 16904
rect 5740 16864 5780 16904
rect 5836 16948 5876 16988
rect 5644 16444 5684 16484
rect 5548 15688 5588 15728
rect 5452 15352 5492 15392
rect 5452 14932 5492 14972
rect 5356 13840 5396 13880
rect 6700 27448 6740 27488
rect 6124 26608 6164 26648
rect 6028 26188 6068 26228
rect 6220 24508 6260 24548
rect 6220 23500 6260 23540
rect 6028 21820 6068 21860
rect 6028 21652 6068 21692
rect 6124 21568 6164 21608
rect 6028 21400 6068 21440
rect 6604 26104 6644 26144
rect 7756 27364 7796 27404
rect 8044 27616 8084 27656
rect 7180 27280 7220 27320
rect 7276 26356 7316 26396
rect 7084 26188 7124 26228
rect 6412 23584 6452 23624
rect 6412 22744 6452 22784
rect 6508 22408 6548 22448
rect 6604 22240 6644 22280
rect 6412 22072 6452 22112
rect 6604 21904 6644 21944
rect 6316 21736 6356 21776
rect 6028 19804 6068 19844
rect 6028 19636 6068 19676
rect 5836 15520 5876 15560
rect 5932 15688 5972 15728
rect 5836 15100 5876 15140
rect 5932 14596 5972 14636
rect 5836 14092 5876 14132
rect 5932 14428 5972 14468
rect 5644 13924 5684 13964
rect 5836 13420 5876 13460
rect 5548 13252 5588 13292
rect 5452 13168 5492 13208
rect 4972 11656 5012 11696
rect 5164 11656 5204 11696
rect 5068 10984 5108 11024
rect 5164 10564 5204 10604
rect 4684 9976 4724 10016
rect 4352 9808 4720 9848
rect 4684 8800 4724 8840
rect 4108 7876 4148 7916
rect 4684 8464 4724 8504
rect 4352 8296 4720 8336
rect 6220 20308 6260 20348
rect 6220 19468 6260 19508
rect 6508 21568 6548 21608
rect 6988 25348 7028 25388
rect 7372 26188 7412 26228
rect 7372 25264 7412 25304
rect 7852 25096 7892 25136
rect 7084 23836 7124 23876
rect 7468 23920 7508 23960
rect 6988 23332 7028 23372
rect 6796 22156 6836 22196
rect 6508 20896 6548 20936
rect 6892 21064 6932 21104
rect 6604 20812 6644 20852
rect 6412 20392 6452 20432
rect 6412 19972 6452 20012
rect 7276 23248 7316 23288
rect 7084 22492 7124 22532
rect 7564 22240 7604 22280
rect 7756 22408 7796 22448
rect 6700 19636 6740 19676
rect 6604 19300 6644 19340
rect 6316 19216 6356 19256
rect 6412 18880 6452 18920
rect 6604 18880 6644 18920
rect 6316 18628 6356 18668
rect 6604 18460 6644 18500
rect 6220 18040 6260 18080
rect 6796 18880 6836 18920
rect 6796 18460 6836 18500
rect 6700 17956 6740 17996
rect 6412 17452 6452 17492
rect 6508 17872 6548 17912
rect 6124 16528 6164 16568
rect 6316 17032 6356 17072
rect 6316 16444 6356 16484
rect 6412 16360 6452 16400
rect 6124 14092 6164 14132
rect 6316 15520 6356 15560
rect 6412 14764 6452 14804
rect 6412 14596 6452 14636
rect 6604 17536 6644 17576
rect 6700 17452 6740 17492
rect 6796 16276 6836 16316
rect 6604 15268 6644 15308
rect 6604 14596 6644 14636
rect 6220 13420 6260 13460
rect 6124 13336 6164 13376
rect 5644 12412 5684 12452
rect 5548 11656 5588 11696
rect 5548 10564 5588 10604
rect 5548 10312 5588 10352
rect 4780 8044 4820 8084
rect 4204 7960 4244 8000
rect 4108 7708 4148 7748
rect 4684 7876 4724 7916
rect 4352 6784 4720 6824
rect 4876 8380 4916 8420
rect 5068 8296 5108 8336
rect 5932 12328 5972 12368
rect 5740 11068 5780 11108
rect 5644 9892 5684 9932
rect 5644 8800 5684 8840
rect 6604 13336 6644 13376
rect 6316 13168 6356 13208
rect 6412 12412 6452 12452
rect 6028 10732 6068 10772
rect 5932 9724 5972 9764
rect 5836 9472 5876 9512
rect 6316 8044 6356 8084
rect 6796 11908 6836 11948
rect 6796 11740 6836 11780
rect 7084 20392 7124 20432
rect 7468 20728 7508 20768
rect 7468 20560 7508 20600
rect 7372 20140 7412 20180
rect 7852 21568 7892 21608
rect 8140 25012 8180 25052
rect 8620 27868 8660 27908
rect 8908 27448 8948 27488
rect 10060 28204 10100 28244
rect 9388 27784 9428 27824
rect 8524 26356 8564 26396
rect 8524 26104 8564 26144
rect 8332 24424 8372 24464
rect 8236 23920 8276 23960
rect 8332 23332 8372 23372
rect 8044 22744 8084 22784
rect 8236 22408 8276 22448
rect 7948 20812 7988 20852
rect 7756 20308 7796 20348
rect 7564 20140 7604 20180
rect 7084 19468 7124 19508
rect 7084 19300 7124 19340
rect 7372 19972 7412 20012
rect 7180 18880 7220 18920
rect 7276 19216 7316 19256
rect 7084 18208 7124 18248
rect 6988 17536 7028 17576
rect 7084 16444 7124 16484
rect 7372 18712 7412 18752
rect 7372 18040 7412 18080
rect 7276 17872 7316 17912
rect 7372 17704 7412 17744
rect 7372 17368 7412 17408
rect 7276 16528 7316 16568
rect 6988 16108 7028 16148
rect 7180 15520 7220 15560
rect 7276 15352 7316 15392
rect 7084 13084 7124 13124
rect 7372 15268 7412 15308
rect 8140 21820 8180 21860
rect 8140 21148 8180 21188
rect 8140 20812 8180 20852
rect 8140 20392 8180 20432
rect 7852 19720 7892 19760
rect 8044 19804 8084 19844
rect 8044 19384 8084 19424
rect 7660 18628 7700 18668
rect 7564 18460 7604 18500
rect 7564 18292 7604 18332
rect 7660 18208 7700 18248
rect 7564 17704 7604 17744
rect 7852 18880 7892 18920
rect 8140 18880 8180 18920
rect 8140 17956 8180 17996
rect 7948 17704 7988 17744
rect 7948 17200 7988 17240
rect 7660 17116 7700 17156
rect 7564 16108 7604 16148
rect 7660 15604 7700 15644
rect 7852 15352 7892 15392
rect 7468 13840 7508 13880
rect 7276 13168 7316 13208
rect 7180 12580 7220 12620
rect 7084 12412 7124 12452
rect 7276 12328 7316 12368
rect 7084 11656 7124 11696
rect 7468 12496 7508 12536
rect 7564 9976 7604 10016
rect 7756 13840 7796 13880
rect 8044 14008 8084 14048
rect 8044 12748 8084 12788
rect 8716 26440 8756 26480
rect 8812 26104 8852 26144
rect 8908 25264 8948 25304
rect 8908 25012 8948 25052
rect 8812 24676 8852 24716
rect 9100 26692 9140 26732
rect 9292 26440 9332 26480
rect 9196 25852 9236 25892
rect 9100 25264 9140 25304
rect 9100 24928 9140 24968
rect 9100 24760 9140 24800
rect 9292 24676 9332 24716
rect 8620 23500 8660 23540
rect 8812 23752 8852 23792
rect 8908 23668 8948 23708
rect 9004 23584 9044 23624
rect 8908 23332 8948 23372
rect 8812 22576 8852 22616
rect 8812 21904 8852 21944
rect 8620 21484 8660 21524
rect 9772 27700 9812 27740
rect 9292 22324 9332 22364
rect 9292 21988 9332 22028
rect 8812 21316 8852 21356
rect 9004 21148 9044 21188
rect 9100 21064 9140 21104
rect 8716 20476 8756 20516
rect 8812 20560 8852 20600
rect 8620 19216 8660 19256
rect 8524 18628 8564 18668
rect 8332 17956 8372 17996
rect 8332 17116 8372 17156
rect 8620 18460 8660 18500
rect 9004 20224 9044 20264
rect 8908 19720 8948 19760
rect 8812 18124 8852 18164
rect 8524 17704 8564 17744
rect 8524 17032 8564 17072
rect 8524 16528 8564 16568
rect 8236 16108 8276 16148
rect 8332 15604 8372 15644
rect 8908 17704 8948 17744
rect 8908 17284 8948 17324
rect 8524 15604 8564 15644
rect 8812 16780 8852 16820
rect 8044 11656 8084 11696
rect 7756 9892 7796 9932
rect 7084 9472 7124 9512
rect 8140 8884 8180 8924
rect 4352 5272 4720 5312
rect 8332 14008 8372 14048
rect 8524 13756 8564 13796
rect 9100 19216 9140 19256
rect 9100 18964 9140 19004
rect 9388 20812 9428 20852
rect 9676 26776 9716 26816
rect 10060 27196 10100 27236
rect 10156 26944 10196 26984
rect 9580 25600 9620 25640
rect 9580 25180 9620 25220
rect 9676 25096 9716 25136
rect 10060 24088 10100 24128
rect 10636 27028 10676 27068
rect 10828 27364 10868 27404
rect 10886 27196 11254 27236
rect 11308 26188 11348 26228
rect 11212 26104 11252 26144
rect 10886 25684 11254 25724
rect 11116 25516 11156 25556
rect 10828 25180 10868 25220
rect 10732 25012 10772 25052
rect 10636 24256 10676 24296
rect 10348 24088 10388 24128
rect 9868 22996 9908 23036
rect 10252 23248 10292 23288
rect 9580 21736 9620 21776
rect 9580 21064 9620 21104
rect 9676 20644 9716 20684
rect 10060 22324 10100 22364
rect 10060 21820 10100 21860
rect 9964 21148 10004 21188
rect 10060 21064 10100 21104
rect 9964 20812 10004 20852
rect 9196 18712 9236 18752
rect 9388 18880 9428 18920
rect 9580 19804 9620 19844
rect 10252 20476 10292 20516
rect 9772 19468 9812 19508
rect 9868 20308 9908 20348
rect 9580 19384 9620 19424
rect 9772 19216 9812 19256
rect 9196 18376 9236 18416
rect 8908 15184 8948 15224
rect 9004 16360 9044 16400
rect 9004 16108 9044 16148
rect 9196 17536 9236 17576
rect 9196 16780 9236 16820
rect 9292 16948 9332 16988
rect 9100 15688 9140 15728
rect 9484 17704 9524 17744
rect 9484 16780 9524 16820
rect 9484 15772 9524 15812
rect 9484 15604 9524 15644
rect 9388 15100 9428 15140
rect 9484 15016 9524 15056
rect 8908 14596 8948 14636
rect 8812 14092 8852 14132
rect 9388 14176 9428 14216
rect 8332 12580 8372 12620
rect 8716 12580 8756 12620
rect 8620 12412 8660 12452
rect 8524 9976 8564 10016
rect 9100 13672 9140 13712
rect 8908 13252 8948 13292
rect 9004 12580 9044 12620
rect 9004 11656 9044 11696
rect 9676 17956 9716 17996
rect 10060 19720 10100 19760
rect 9964 19552 10004 19592
rect 10156 19468 10196 19508
rect 9868 17704 9908 17744
rect 9868 17536 9908 17576
rect 9772 17368 9812 17408
rect 9772 17200 9812 17240
rect 9676 17032 9716 17072
rect 9676 16696 9716 16736
rect 9868 16780 9908 16820
rect 9772 14596 9812 14636
rect 9580 14092 9620 14132
rect 9580 13924 9620 13964
rect 9772 13924 9812 13964
rect 9964 15436 10004 15476
rect 9772 13168 9812 13208
rect 9868 13252 9908 13292
rect 11404 26020 11444 26060
rect 11404 25852 11444 25892
rect 10886 24172 11254 24212
rect 11404 25096 11444 25136
rect 11212 23836 11252 23876
rect 10886 22660 11254 22700
rect 10732 22492 10772 22532
rect 11116 22492 11156 22532
rect 10886 21148 11254 21188
rect 10732 20812 10772 20852
rect 11020 20728 11060 20768
rect 10252 18880 10292 18920
rect 10348 19468 10388 19508
rect 10924 20140 10964 20180
rect 11116 20140 11156 20180
rect 10636 19720 10676 19760
rect 11116 19972 11156 20012
rect 10886 19636 11254 19676
rect 10540 19216 10580 19256
rect 11500 23248 11540 23288
rect 12364 28288 12404 28328
rect 12126 27952 12494 27992
rect 11788 27532 11828 27572
rect 12364 27112 12404 27152
rect 11788 26776 11828 26816
rect 11692 26188 11732 26228
rect 12364 26860 12404 26900
rect 12556 26860 12596 26900
rect 12126 26440 12494 26480
rect 12076 25432 12116 25472
rect 11884 25180 11924 25220
rect 12126 24928 12494 24968
rect 11884 23248 11924 23288
rect 12364 24340 12404 24380
rect 13036 28288 13076 28328
rect 12844 26188 12884 26228
rect 12844 24256 12884 24296
rect 12652 23668 12692 23708
rect 12126 23416 12494 23456
rect 13132 28120 13172 28160
rect 13612 28120 13652 28160
rect 13516 26944 13556 26984
rect 13132 25936 13172 25976
rect 13516 26692 13556 26732
rect 13324 26020 13364 26060
rect 13228 24592 13268 24632
rect 13036 23920 13076 23960
rect 13228 24256 13268 24296
rect 12940 23332 12980 23372
rect 11980 23080 12020 23120
rect 11884 22828 11924 22868
rect 12126 21904 12494 21944
rect 11692 21316 11732 21356
rect 11596 21232 11636 21272
rect 11788 21064 11828 21104
rect 11404 19216 11444 19256
rect 10732 18880 10772 18920
rect 11020 18880 11060 18920
rect 10540 18292 10580 18332
rect 10348 16612 10388 16652
rect 10444 16444 10484 16484
rect 10252 15856 10292 15896
rect 10444 15856 10484 15896
rect 10444 15604 10484 15644
rect 10156 15520 10196 15560
rect 10156 14344 10196 14384
rect 10060 14008 10100 14048
rect 10348 15436 10388 15476
rect 10886 18124 11254 18164
rect 11596 19804 11636 19844
rect 11692 19468 11732 19508
rect 11500 18124 11540 18164
rect 10636 16528 10676 16568
rect 10732 17116 10772 17156
rect 11404 17536 11444 17576
rect 11692 18880 11732 18920
rect 11692 17704 11732 17744
rect 11500 17368 11540 17408
rect 10828 17032 10868 17072
rect 10886 16612 11254 16652
rect 11020 16360 11060 16400
rect 11212 16108 11252 16148
rect 11308 15772 11348 15812
rect 11404 15856 11444 15896
rect 10444 15100 10484 15140
rect 10348 14260 10388 14300
rect 10060 13252 10100 13292
rect 10060 11824 10100 11864
rect 10060 11656 10100 11696
rect 3112 4516 3480 4556
rect 10636 14428 10676 14468
rect 10636 13336 10676 13376
rect 11308 15352 11348 15392
rect 11212 15268 11252 15308
rect 10886 15100 11254 15140
rect 11116 14932 11156 14972
rect 10828 14764 10868 14804
rect 11308 14932 11348 14972
rect 11116 14512 11156 14552
rect 12126 20392 12494 20432
rect 12844 20308 12884 20348
rect 12364 19720 12404 19760
rect 12126 18880 12494 18920
rect 12652 20140 12692 20180
rect 13516 23836 13556 23876
rect 13420 23080 13460 23120
rect 13420 22324 13460 22364
rect 13900 26860 13940 26900
rect 13900 26356 13940 26396
rect 15340 27868 15380 27908
rect 14668 27028 14708 27068
rect 15244 26944 15284 26984
rect 15052 26776 15092 26816
rect 14572 26524 14612 26564
rect 13900 26020 13940 26060
rect 13996 26104 14036 26144
rect 13708 25180 13748 25220
rect 14188 25600 14228 25640
rect 14476 25852 14516 25892
rect 13900 24844 13940 24884
rect 14860 26692 14900 26732
rect 14956 26356 14996 26396
rect 14860 26104 14900 26144
rect 14668 25180 14708 25220
rect 14284 23920 14324 23960
rect 14764 25012 14804 25052
rect 14668 23584 14708 23624
rect 14476 23080 14516 23120
rect 13324 21568 13364 21608
rect 13324 21148 13364 21188
rect 13324 20560 13364 20600
rect 13516 20812 13556 20852
rect 13708 21316 13748 21356
rect 13708 20728 13748 20768
rect 13996 20560 14036 20600
rect 14572 20644 14612 20684
rect 14380 20308 14420 20348
rect 12652 19216 12692 19256
rect 11980 18292 12020 18332
rect 11788 17536 11828 17576
rect 12268 17956 12308 17996
rect 12556 17956 12596 17996
rect 12460 17872 12500 17912
rect 12268 17536 12308 17576
rect 12126 17368 12494 17408
rect 12652 17200 12692 17240
rect 11980 16780 12020 16820
rect 11884 16696 11924 16736
rect 11692 16612 11732 16652
rect 11788 16108 11828 16148
rect 12364 16780 12404 16820
rect 12460 16360 12500 16400
rect 12126 15856 12494 15896
rect 12460 15688 12500 15728
rect 11980 15436 12020 15476
rect 12172 15520 12212 15560
rect 11884 14932 11924 14972
rect 12172 15268 12212 15308
rect 11404 14176 11444 14216
rect 11500 14512 11540 14552
rect 11596 14344 11636 14384
rect 11500 14092 11540 14132
rect 10886 13588 11254 13628
rect 11404 13504 11444 13544
rect 11212 13252 11252 13292
rect 10828 12580 10868 12620
rect 10636 12244 10676 12284
rect 10540 11824 10580 11864
rect 10060 9892 10100 9932
rect 9772 8884 9812 8924
rect 10252 10564 10292 10604
rect 10886 12076 11254 12116
rect 10732 11992 10772 12032
rect 11404 13336 11444 13376
rect 11596 13084 11636 13124
rect 12364 15268 12404 15308
rect 11980 14596 12020 14636
rect 12126 14344 12494 14384
rect 11788 14260 11828 14300
rect 12268 14176 12308 14216
rect 12460 13924 12500 13964
rect 11788 13000 11828 13040
rect 10886 10564 11254 10604
rect 11020 10396 11060 10436
rect 11404 10984 11444 11024
rect 10886 9052 11254 9092
rect 10886 7540 11254 7580
rect 11500 9472 11540 9512
rect 11500 7960 11540 8000
rect 12652 15268 12692 15308
rect 13132 19720 13172 19760
rect 13324 19636 13364 19676
rect 12940 18964 12980 19004
rect 13132 18964 13172 19004
rect 13228 19384 13268 19424
rect 13132 17956 13172 17996
rect 12844 17536 12884 17576
rect 12940 17620 12980 17660
rect 13420 18040 13460 18080
rect 13804 18460 13844 18500
rect 12940 17032 12980 17072
rect 12844 16360 12884 16400
rect 13228 17032 13268 17072
rect 12844 15940 12884 15980
rect 12940 15856 12980 15896
rect 12844 15688 12884 15728
rect 12844 15436 12884 15476
rect 12940 15268 12980 15308
rect 12844 14932 12884 14972
rect 12940 14092 12980 14132
rect 12748 14008 12788 14048
rect 12748 13588 12788 13628
rect 12172 13168 12212 13208
rect 13132 16192 13172 16232
rect 13132 15268 13172 15308
rect 12126 12832 12494 12872
rect 13708 16444 13748 16484
rect 13228 14512 13268 14552
rect 13324 14344 13364 14384
rect 13324 13084 13364 13124
rect 12076 12580 12116 12620
rect 11980 11824 12020 11864
rect 12172 11656 12212 11696
rect 12126 11320 12494 11360
rect 12652 11068 12692 11108
rect 12268 10984 12308 11024
rect 13708 15772 13748 15812
rect 13516 13504 13556 13544
rect 13420 12664 13460 12704
rect 12940 11068 12980 11108
rect 12126 9808 12494 9848
rect 12460 9472 12500 9512
rect 11692 7960 11732 8000
rect 11980 9388 12020 9428
rect 12126 8296 12494 8336
rect 12126 6784 12494 6824
rect 10886 6028 11254 6068
rect 10252 5608 10292 5648
rect 12460 6448 12500 6488
rect 13132 9472 13172 9512
rect 12126 5272 12494 5312
rect 12940 5020 12980 5060
rect 13804 13084 13844 13124
rect 13804 12832 13844 12872
rect 13804 12328 13844 12368
rect 14284 18880 14324 18920
rect 14284 18628 14324 18668
rect 14092 17116 14132 17156
rect 14092 16444 14132 16484
rect 14476 16780 14516 16820
rect 14284 16024 14324 16064
rect 14476 15688 14516 15728
rect 14188 15268 14228 15308
rect 14284 15436 14324 15476
rect 14284 14932 14324 14972
rect 13996 14596 14036 14636
rect 14188 14512 14228 14552
rect 13996 14260 14036 14300
rect 13324 7204 13364 7244
rect 13708 7204 13748 7244
rect 15436 27196 15476 27236
rect 15436 26944 15476 26984
rect 15340 26104 15380 26144
rect 15244 25180 15284 25220
rect 14860 23752 14900 23792
rect 14860 20728 14900 20768
rect 15052 21484 15092 21524
rect 15244 21484 15284 21524
rect 15052 21316 15092 21356
rect 14956 19552 14996 19592
rect 15436 25180 15476 25220
rect 16204 26692 16244 26732
rect 16396 26524 16436 26564
rect 16204 26020 16244 26060
rect 15820 25852 15860 25892
rect 15628 24088 15668 24128
rect 15820 24088 15860 24128
rect 15628 23668 15668 23708
rect 15532 21820 15572 21860
rect 15340 21232 15380 21272
rect 15244 20560 15284 20600
rect 14956 19300 14996 19340
rect 14764 17788 14804 17828
rect 14668 16444 14708 16484
rect 15148 18964 15188 19004
rect 15340 19384 15380 19424
rect 15244 18880 15284 18920
rect 15340 18208 15380 18248
rect 15436 18460 15476 18500
rect 15244 18040 15284 18080
rect 15244 17536 15284 17576
rect 15148 16864 15188 16904
rect 15148 16528 15188 16568
rect 15244 16780 15284 16820
rect 15244 16108 15284 16148
rect 14668 14008 14708 14048
rect 14764 11824 14804 11864
rect 13996 6448 14036 6488
rect 13228 5608 13268 5648
rect 13804 5608 13844 5648
rect 13900 5020 13940 5060
rect 14956 14344 14996 14384
rect 14956 12076 14996 12116
rect 14956 11824 14996 11864
rect 15436 17032 15476 17072
rect 16396 25096 16436 25136
rect 16300 24004 16340 24044
rect 16300 23584 16340 23624
rect 16300 22240 16340 22280
rect 16396 22072 16436 22112
rect 16396 21568 16436 21608
rect 16012 20728 16052 20768
rect 15820 19972 15860 20012
rect 15820 19552 15860 19592
rect 15628 16528 15668 16568
rect 15436 15940 15476 15980
rect 15436 15772 15476 15812
rect 15340 14008 15380 14048
rect 15244 13252 15284 13292
rect 15148 13168 15188 13208
rect 15148 12412 15188 12452
rect 15148 11740 15188 11780
rect 15340 12664 15380 12704
rect 15148 10228 15188 10268
rect 15052 7960 15092 8000
rect 15148 7204 15188 7244
rect 15820 17956 15860 17996
rect 15916 18880 15956 18920
rect 15820 16780 15860 16820
rect 15820 14344 15860 14384
rect 15724 13252 15764 13292
rect 15628 13000 15668 13040
rect 15628 12664 15668 12704
rect 15820 12412 15860 12452
rect 15724 10144 15764 10184
rect 15628 6448 15668 6488
rect 16204 20140 16244 20180
rect 16300 19552 16340 19592
rect 16108 18628 16148 18668
rect 16204 19216 16244 19256
rect 16396 19300 16436 19340
rect 16108 18124 16148 18164
rect 16204 17704 16244 17744
rect 16012 17032 16052 17072
rect 16012 16696 16052 16736
rect 16108 16108 16148 16148
rect 16396 18964 16436 19004
rect 17164 28204 17204 28244
rect 16588 26608 16628 26648
rect 16588 26188 16628 26228
rect 16876 27532 16916 27572
rect 16876 27112 16916 27152
rect 16780 26860 16820 26900
rect 19900 27952 20268 27992
rect 17932 27196 17972 27236
rect 16780 25852 16820 25892
rect 16780 25432 16820 25472
rect 16972 25096 17012 25136
rect 16780 24844 16820 24884
rect 17260 26524 17300 26564
rect 17164 24844 17204 24884
rect 17164 24676 17204 24716
rect 17836 25516 17876 25556
rect 17356 24088 17396 24128
rect 16876 23836 16916 23876
rect 16972 23668 17012 23708
rect 17740 24508 17780 24548
rect 17356 23248 17396 23288
rect 17164 22240 17204 22280
rect 17068 21820 17108 21860
rect 16876 21736 16916 21776
rect 16972 21652 17012 21692
rect 16684 20812 16724 20852
rect 16588 19552 16628 19592
rect 16972 21148 17012 21188
rect 17836 23500 17876 23540
rect 17836 23080 17876 23120
rect 17260 21148 17300 21188
rect 17356 21652 17396 21692
rect 16876 19804 16916 19844
rect 16588 18460 16628 18500
rect 16684 18208 16724 18248
rect 16492 16864 16532 16904
rect 16300 15604 16340 15644
rect 16396 15184 16436 15224
rect 16108 14680 16148 14720
rect 16012 14092 16052 14132
rect 16012 13588 16052 13628
rect 17260 20476 17300 20516
rect 17452 20644 17492 20684
rect 17452 20140 17492 20180
rect 16972 18460 17012 18500
rect 16684 16444 16724 16484
rect 16876 16780 16916 16820
rect 16780 15520 16820 15560
rect 16876 15940 16916 15980
rect 16588 14596 16628 14636
rect 16300 13252 16340 13292
rect 16300 13084 16340 13124
rect 16396 13000 16436 13040
rect 16108 12328 16148 12368
rect 16780 14008 16820 14048
rect 16876 13672 16916 13712
rect 16972 14596 17012 14636
rect 17164 18040 17204 18080
rect 17260 16528 17300 16568
rect 17164 15352 17204 15392
rect 16972 12076 17012 12116
rect 16204 9472 16244 9512
rect 17260 14680 17300 14720
rect 17260 14512 17300 14552
rect 17548 19804 17588 19844
rect 18220 26944 18260 26984
rect 18028 26020 18068 26060
rect 18660 27196 19028 27236
rect 18220 25516 18260 25556
rect 18028 25180 18068 25220
rect 18124 24760 18164 24800
rect 18316 23416 18356 23456
rect 18124 23248 18164 23288
rect 18220 22828 18260 22868
rect 17836 20812 17876 20852
rect 17740 20728 17780 20768
rect 17548 19468 17588 19508
rect 17644 19216 17684 19256
rect 18028 21484 18068 21524
rect 18124 21316 18164 21356
rect 18124 20560 18164 20600
rect 18028 20476 18068 20516
rect 17932 20140 17972 20180
rect 18892 26776 18932 26816
rect 19084 26440 19124 26480
rect 18660 25684 19028 25724
rect 18988 25432 19028 25472
rect 18796 25096 18836 25136
rect 19564 26860 19604 26900
rect 21772 27532 21812 27572
rect 20428 27280 20468 27320
rect 19660 26776 19700 26816
rect 20236 26776 20276 26816
rect 21388 27112 21428 27152
rect 19468 26440 19508 26480
rect 19900 26440 20268 26480
rect 19756 26020 19796 26060
rect 19564 25684 19604 25724
rect 19660 25516 19700 25556
rect 19084 25096 19124 25136
rect 19564 25180 19604 25220
rect 18700 24508 18740 24548
rect 19468 24760 19508 24800
rect 19852 25600 19892 25640
rect 20140 25852 20180 25892
rect 20140 25516 20180 25556
rect 20140 25180 20180 25220
rect 19900 24928 20268 24968
rect 18796 24340 18836 24380
rect 18660 24172 19028 24212
rect 18508 23920 18548 23960
rect 19084 23920 19124 23960
rect 18412 21568 18452 21608
rect 18412 20644 18452 20684
rect 17836 18964 17876 19004
rect 18124 19216 18164 19256
rect 17548 16444 17588 16484
rect 17548 16108 17588 16148
rect 17644 15436 17684 15476
rect 17836 17788 17876 17828
rect 18028 17788 18068 17828
rect 17932 17704 17972 17744
rect 17452 15352 17492 15392
rect 18412 18964 18452 19004
rect 18604 23332 18644 23372
rect 18604 23080 18644 23120
rect 18660 22660 19028 22700
rect 19084 21988 19124 22028
rect 18660 21148 19028 21188
rect 18700 19972 18740 20012
rect 18660 19636 19028 19676
rect 18988 19384 19028 19424
rect 18604 18880 18644 18920
rect 18700 18712 18740 18752
rect 18988 18796 19028 18836
rect 18660 18124 19028 18164
rect 18892 17788 18932 17828
rect 18892 17032 18932 17072
rect 18988 16780 19028 16820
rect 18660 16612 19028 16652
rect 19276 21820 19316 21860
rect 18316 14932 18356 14972
rect 18412 15268 18452 15308
rect 18028 14344 18068 14384
rect 17740 14008 17780 14048
rect 17836 12580 17876 12620
rect 16972 10144 17012 10184
rect 18124 12832 18164 12872
rect 18412 14008 18452 14048
rect 18412 13672 18452 13712
rect 18700 15520 18740 15560
rect 19468 23416 19508 23456
rect 20140 24676 20180 24716
rect 19756 24172 19796 24212
rect 20332 24508 20372 24548
rect 20236 23584 20276 23624
rect 19900 23416 20268 23456
rect 19564 22996 19604 23036
rect 20236 22156 20276 22196
rect 19900 21904 20268 21944
rect 19564 21652 19604 21692
rect 19852 21736 19892 21776
rect 20140 21736 20180 21776
rect 19468 20140 19508 20180
rect 19468 16864 19508 16904
rect 19372 16276 19412 16316
rect 18660 15100 19028 15140
rect 18988 14932 19028 14972
rect 18796 14764 18836 14804
rect 18604 14680 18644 14720
rect 18892 14512 18932 14552
rect 18892 14344 18932 14384
rect 18700 13924 18740 13964
rect 19180 14680 19220 14720
rect 18660 13588 19028 13628
rect 18892 13420 18932 13460
rect 18700 13336 18740 13376
rect 18796 12916 18836 12956
rect 18700 12412 18740 12452
rect 19276 13420 19316 13460
rect 19468 14848 19508 14888
rect 19468 14176 19508 14216
rect 19468 13252 19508 13292
rect 18660 12076 19028 12116
rect 18892 11656 18932 11696
rect 18660 10564 19028 10604
rect 18316 10396 18356 10436
rect 18220 10228 18260 10268
rect 19372 12664 19412 12704
rect 19276 11992 19316 12032
rect 19276 11656 19316 11696
rect 19180 10816 19220 10856
rect 18660 9052 19028 9092
rect 19372 11236 19412 11276
rect 20236 20560 20276 20600
rect 19900 20392 20268 20432
rect 20620 23500 20660 23540
rect 20716 23416 20756 23456
rect 21004 25516 21044 25556
rect 21004 24844 21044 24884
rect 20908 23920 20948 23960
rect 20812 22912 20852 22952
rect 21292 26104 21332 26144
rect 21484 26692 21524 26732
rect 21580 25180 21620 25220
rect 21388 25012 21428 25052
rect 21580 24508 21620 24548
rect 21292 24088 21332 24128
rect 21388 23584 21428 23624
rect 21196 23416 21236 23456
rect 20716 22072 20756 22112
rect 20524 20560 20564 20600
rect 19900 18880 20268 18920
rect 21580 23080 21620 23120
rect 21772 25096 21812 25136
rect 21772 22492 21812 22532
rect 21676 22072 21716 22112
rect 23020 26776 23060 26816
rect 22252 26440 22292 26480
rect 22156 26020 22196 26060
rect 22828 26188 22868 26228
rect 22252 26104 22292 26144
rect 22156 25432 22196 25472
rect 21388 20476 21428 20516
rect 20620 18712 20660 18752
rect 19900 17368 20268 17408
rect 19948 17032 19988 17072
rect 20428 17032 20468 17072
rect 20140 16948 20180 16988
rect 20428 16360 20468 16400
rect 19948 16192 19988 16232
rect 20236 16108 20276 16148
rect 20332 16024 20372 16064
rect 20620 16276 20660 16316
rect 20908 17032 20948 17072
rect 20908 16780 20948 16820
rect 20908 16276 20948 16316
rect 19900 15856 20268 15896
rect 21388 17704 21428 17744
rect 21004 16108 21044 16148
rect 19756 14764 19796 14804
rect 20044 15352 20084 15392
rect 20044 14764 20084 14804
rect 20140 14512 20180 14552
rect 19900 14344 20268 14384
rect 20140 14176 20180 14216
rect 19756 13840 19796 13880
rect 19660 13252 19700 13292
rect 19948 13672 19988 13712
rect 19660 13000 19700 13040
rect 19852 13084 19892 13124
rect 20428 15352 20468 15392
rect 20908 15352 20948 15392
rect 20716 14848 20756 14888
rect 21196 16864 21236 16904
rect 21100 15352 21140 15392
rect 21100 14764 21140 14804
rect 20428 13168 20468 13208
rect 19900 12832 20268 12872
rect 19756 12496 19796 12536
rect 19756 12244 19796 12284
rect 19660 11740 19700 11780
rect 20812 14008 20852 14048
rect 21004 14596 21044 14636
rect 20812 13420 20852 13460
rect 20812 13252 20852 13292
rect 20428 12412 20468 12452
rect 19468 9892 19508 9932
rect 19900 11320 20268 11360
rect 20140 10396 20180 10436
rect 19900 9808 20268 9848
rect 20812 12496 20852 12536
rect 21196 13672 21236 13712
rect 20524 9892 20564 9932
rect 19900 8296 20268 8336
rect 17740 7960 17780 8000
rect 18124 7372 18164 7412
rect 18124 7120 18164 7160
rect 18660 7540 19028 7580
rect 18892 7372 18932 7412
rect 18700 7204 18740 7244
rect 19180 7120 19220 7160
rect 19372 7204 19412 7244
rect 19900 6784 20268 6824
rect 18660 6028 19028 6068
rect 10886 4516 11254 4556
rect 18660 4516 19028 4556
rect 19900 5272 20268 5312
rect 21484 20140 21524 20180
rect 21484 16444 21524 16484
rect 21676 15688 21716 15728
rect 21388 14596 21428 14636
rect 21388 14176 21428 14216
rect 21388 13924 21428 13964
rect 21580 15352 21620 15392
rect 21676 14848 21716 14888
rect 21484 13840 21524 13880
rect 22444 25600 22484 25640
rect 22828 25432 22868 25472
rect 23116 25516 23156 25556
rect 23212 25432 23252 25472
rect 22924 25180 22964 25220
rect 23692 25936 23732 25976
rect 24076 25852 24116 25892
rect 25804 27700 25844 27740
rect 22636 25012 22676 25052
rect 22924 24676 22964 24716
rect 22348 23752 22388 23792
rect 22540 24172 22580 24212
rect 22252 18712 22292 18752
rect 22924 23752 22964 23792
rect 22924 23584 22964 23624
rect 22636 23500 22676 23540
rect 22732 23332 22772 23372
rect 22636 22156 22676 22196
rect 23116 23752 23156 23792
rect 23308 23584 23348 23624
rect 23596 24676 23636 24716
rect 23020 21988 23060 22028
rect 22732 20644 22772 20684
rect 22540 18712 22580 18752
rect 21868 16696 21908 16736
rect 22348 16444 22388 16484
rect 22060 16276 22100 16316
rect 21964 14596 22004 14636
rect 22444 15604 22484 15644
rect 22156 15352 22196 15392
rect 23404 20476 23444 20516
rect 23116 19216 23156 19256
rect 24556 27448 24596 27488
rect 24460 26104 24500 26144
rect 24844 26020 24884 26060
rect 25228 26020 25268 26060
rect 25228 25516 25268 25556
rect 24940 25264 24980 25304
rect 24460 23752 24500 23792
rect 24076 22996 24116 23036
rect 24076 22324 24116 22364
rect 23116 17704 23156 17744
rect 23692 19300 23732 19340
rect 22828 16276 22868 16316
rect 23020 15688 23060 15728
rect 21964 13840 22004 13880
rect 21868 13504 21908 13544
rect 22060 13420 22100 13460
rect 22156 13672 22196 13712
rect 22444 14596 22484 14636
rect 22444 14008 22484 14048
rect 22348 13924 22388 13964
rect 22924 14848 22964 14888
rect 22924 14008 22964 14048
rect 22732 13924 22772 13964
rect 22348 13336 22388 13376
rect 22060 13000 22100 13040
rect 21580 12916 21620 12956
rect 21484 10480 21524 10520
rect 21580 8716 21620 8756
rect 21868 9472 21908 9512
rect 22540 13252 22580 13292
rect 22636 13168 22676 13208
rect 23308 17620 23348 17660
rect 23884 20644 23924 20684
rect 24172 23416 24212 23456
rect 25036 24088 25076 24128
rect 25132 24592 25172 24632
rect 24076 20476 24116 20516
rect 24364 21484 24404 21524
rect 24748 23248 24788 23288
rect 24268 20560 24308 20600
rect 24460 20560 24500 20600
rect 24652 21820 24692 21860
rect 25420 25264 25460 25304
rect 25708 24760 25748 24800
rect 25516 24088 25556 24128
rect 25708 23836 25748 23876
rect 25996 26020 26036 26060
rect 26476 27532 26516 27572
rect 26434 27196 26802 27236
rect 26380 27028 26420 27068
rect 26572 26188 26612 26228
rect 26764 26188 26804 26228
rect 26434 25684 26802 25724
rect 25516 23584 25556 23624
rect 25900 23836 25940 23876
rect 26188 25180 26228 25220
rect 26188 24592 26228 24632
rect 26284 24676 26324 24716
rect 26380 24340 26420 24380
rect 26956 27364 26996 27404
rect 26860 24256 26900 24296
rect 26434 24172 26802 24212
rect 25804 23248 25844 23288
rect 25900 23500 25940 23540
rect 24940 22408 24980 22448
rect 25036 20560 25076 20600
rect 26092 22156 26132 22196
rect 26188 22072 26228 22112
rect 27724 28120 27764 28160
rect 27674 27952 28042 27992
rect 27628 27700 27668 27740
rect 27244 26944 27284 26984
rect 27436 26440 27476 26480
rect 27244 25768 27284 25808
rect 27340 26188 27380 26228
rect 28684 28120 28724 28160
rect 27916 27364 27956 27404
rect 27724 26944 27764 26984
rect 27674 26440 28042 26480
rect 27916 26188 27956 26228
rect 27916 26020 27956 26060
rect 27724 25852 27764 25892
rect 27532 25768 27572 25808
rect 27340 25264 27380 25304
rect 27916 25096 27956 25136
rect 27674 24928 28042 24968
rect 27052 23164 27092 23204
rect 27148 24340 27188 24380
rect 26380 22996 26420 23036
rect 26434 22660 26802 22700
rect 27052 22492 27092 22532
rect 26764 22324 26804 22364
rect 27148 21988 27188 22028
rect 26956 21820 26996 21860
rect 26434 21148 26802 21188
rect 28108 23584 28148 23624
rect 27674 23416 28042 23456
rect 27674 21904 28042 21944
rect 25036 19300 25076 19340
rect 23500 16276 23540 16316
rect 23308 16024 23348 16064
rect 23404 15436 23444 15476
rect 23212 14428 23252 14468
rect 22540 12748 22580 12788
rect 23308 13924 23348 13964
rect 23404 14176 23444 14216
rect 23692 15772 23732 15812
rect 23596 14512 23636 14552
rect 23788 15436 23828 15476
rect 23884 15352 23924 15392
rect 23596 13924 23636 13964
rect 23884 14512 23924 14552
rect 23884 14008 23924 14048
rect 23596 13168 23636 13208
rect 23980 13504 24020 13544
rect 24076 14764 24116 14804
rect 23980 13084 24020 13124
rect 23500 12580 23540 12620
rect 23116 12328 23156 12368
rect 23404 12412 23444 12452
rect 22348 7876 22388 7916
rect 22636 7960 22676 8000
rect 23596 8716 23636 8756
rect 24172 13504 24212 13544
rect 24844 16276 24884 16316
rect 25708 18964 25748 19004
rect 25612 16276 25652 16316
rect 24844 13840 24884 13880
rect 24460 13084 24500 13124
rect 24460 12832 24500 12872
rect 24364 12748 24404 12788
rect 24940 12412 24980 12452
rect 25036 13000 25076 13040
rect 25420 12916 25460 12956
rect 25516 12664 25556 12704
rect 25420 12496 25460 12536
rect 24652 12244 24692 12284
rect 24652 9472 24692 9512
rect 24076 9388 24116 9428
rect 24556 9388 24596 9428
rect 24172 7960 24212 8000
rect 24556 8128 24596 8168
rect 26434 19636 26802 19676
rect 26380 19300 26420 19340
rect 26668 18964 26708 19004
rect 26668 18292 26708 18332
rect 26434 18124 26802 18164
rect 27052 17620 27092 17660
rect 26092 15520 26132 15560
rect 26434 16612 26802 16652
rect 26860 16276 26900 16316
rect 25804 12916 25844 12956
rect 25900 12832 25940 12872
rect 26188 12664 26228 12704
rect 25708 12496 25748 12536
rect 25900 11824 25940 11864
rect 26434 15100 26802 15140
rect 26434 13588 26802 13628
rect 26764 13420 26804 13460
rect 27244 18712 27284 18752
rect 27052 13924 27092 13964
rect 27052 12496 27092 12536
rect 26434 12076 26802 12116
rect 26434 10564 26802 10604
rect 28396 26608 28436 26648
rect 28396 23584 28436 23624
rect 28780 27532 28820 27572
rect 28588 26776 28628 26816
rect 29260 27700 29300 27740
rect 29836 27700 29876 27740
rect 29260 27532 29300 27572
rect 29644 27112 29684 27152
rect 29740 27028 29780 27068
rect 28780 26608 28820 26648
rect 28684 26188 28724 26228
rect 28972 26104 29012 26144
rect 29164 25768 29204 25808
rect 28780 25264 28820 25304
rect 28972 25012 29012 25052
rect 29164 24844 29204 24884
rect 28876 24760 28916 24800
rect 29356 26860 29396 26900
rect 29452 25936 29492 25976
rect 29356 25600 29396 25640
rect 29452 25516 29492 25556
rect 29260 24592 29300 24632
rect 28492 21484 28532 21524
rect 28300 21148 28340 21188
rect 27674 20392 28042 20432
rect 28972 24088 29012 24128
rect 28876 23668 28916 23708
rect 29164 24172 29204 24212
rect 28876 23500 28916 23540
rect 28972 21820 29012 21860
rect 28684 20644 28724 20684
rect 28300 20560 28340 20600
rect 28588 20056 28628 20096
rect 27674 18880 28042 18920
rect 28780 18544 28820 18584
rect 29164 23584 29204 23624
rect 29164 23332 29204 23372
rect 29260 22996 29300 23036
rect 29164 22912 29204 22952
rect 29644 26860 29684 26900
rect 29932 27448 29972 27488
rect 30028 25852 30068 25892
rect 29932 25600 29972 25640
rect 29548 24256 29588 24296
rect 29548 23836 29588 23876
rect 29644 23752 29684 23792
rect 29644 23500 29684 23540
rect 29548 22072 29588 22112
rect 29836 22156 29876 22196
rect 29260 21148 29300 21188
rect 29164 19132 29204 19172
rect 30988 27280 31028 27320
rect 30412 26524 30452 26564
rect 30988 26356 31028 26396
rect 30604 26272 30644 26312
rect 30220 25348 30260 25388
rect 30988 24424 31028 24464
rect 30028 22240 30068 22280
rect 30028 22072 30068 22112
rect 30028 21736 30068 21776
rect 30604 20980 30644 21020
rect 30892 21400 30932 21440
rect 30892 20896 30932 20936
rect 29932 19888 29972 19928
rect 29548 19048 29588 19088
rect 28684 18376 28724 18416
rect 27628 18292 27668 18332
rect 28012 17872 28052 17912
rect 27674 17368 28042 17408
rect 27674 15856 28042 15896
rect 28108 15520 28148 15560
rect 27674 14344 28042 14384
rect 27674 12832 28042 12872
rect 27244 12412 27284 12452
rect 27820 12496 27860 12536
rect 27916 12412 27956 12452
rect 28108 12244 28148 12284
rect 28204 12328 28244 12368
rect 27628 11824 27668 11864
rect 28780 13504 28820 13544
rect 28780 13252 28820 13292
rect 29068 13756 29108 13796
rect 27674 11320 28042 11360
rect 25996 9472 26036 9512
rect 27674 9808 28042 9848
rect 26434 9052 26802 9092
rect 26572 8716 26612 8756
rect 25900 8632 25940 8672
rect 25612 8044 25652 8084
rect 27052 8632 27092 8672
rect 27674 8296 28042 8336
rect 26284 8128 26324 8168
rect 26380 8044 26420 8084
rect 26860 7960 26900 8000
rect 26764 7876 26804 7916
rect 26434 7540 26802 7580
rect 27674 6784 28042 6824
rect 26434 6028 26802 6068
rect 27674 5272 28042 5312
rect 26434 4516 26802 4556
rect 4352 3760 4720 3800
rect 12126 3760 12494 3800
rect 19900 3760 20268 3800
rect 27674 3760 28042 3800
rect 3112 3004 3480 3044
rect 10886 3004 11254 3044
rect 18660 3004 19028 3044
rect 26434 3004 26802 3044
rect 4352 2248 4720 2288
rect 12126 2248 12494 2288
rect 19900 2248 20268 2288
rect 27674 2248 28042 2288
rect 3112 1492 3480 1532
rect 10886 1492 11254 1532
rect 18660 1492 19028 1532
rect 26434 1492 26802 1532
rect 4352 736 4720 776
rect 12126 736 12494 776
rect 19900 736 20268 776
rect 27674 736 28042 776
<< metal4 >>
rect 12355 28288 12364 28328
rect 12404 28288 13036 28328
rect 13076 28288 13085 28328
rect 10051 28204 10060 28244
rect 10100 28204 17164 28244
rect 17204 28204 17213 28244
rect 4675 28120 4684 28160
rect 4724 28120 4876 28160
rect 4916 28120 4925 28160
rect 13123 28120 13132 28160
rect 13172 28120 13612 28160
rect 13652 28120 13661 28160
rect 27715 28120 27724 28160
rect 27764 28120 28684 28160
rect 28724 28120 28733 28160
rect 3139 28036 3148 28076
rect 3188 28036 6700 28076
rect 6740 28036 6749 28076
rect 4343 27952 4352 27992
rect 4720 27952 4729 27992
rect 12117 27952 12126 27992
rect 12494 27952 12503 27992
rect 19891 27952 19900 27992
rect 20268 27952 20277 27992
rect 27665 27952 27674 27992
rect 28042 27952 28051 27992
rect 6125 27868 6220 27908
rect 6260 27868 6269 27908
rect 8611 27868 8620 27908
rect 8660 27868 15340 27908
rect 15380 27868 15389 27908
rect 2947 27784 2956 27824
rect 2996 27784 9388 27824
rect 9428 27784 9437 27824
rect 2083 27700 2092 27740
rect 2132 27700 9772 27740
rect 9812 27700 9821 27740
rect 25795 27700 25804 27740
rect 25844 27700 27628 27740
rect 27668 27700 27677 27740
rect 29251 27700 29260 27740
rect 29300 27700 29836 27740
rect 29876 27700 29885 27740
rect 4387 27616 4396 27656
rect 4436 27616 5644 27656
rect 5684 27616 5693 27656
rect 6211 27616 6220 27656
rect 6260 27616 8044 27656
rect 8084 27616 8093 27656
rect 2563 27532 2572 27572
rect 2612 27532 11788 27572
rect 11828 27532 11837 27572
rect 16867 27532 16876 27572
rect 16916 27532 16972 27572
rect 17012 27532 17021 27572
rect 21763 27532 21772 27572
rect 21812 27532 26476 27572
rect 26516 27532 27532 27572
rect 27572 27532 27581 27572
rect 28685 27532 28780 27572
rect 28820 27532 28829 27572
rect 29165 27532 29260 27572
rect 29300 27532 29309 27572
rect 3331 27448 3340 27488
rect 3380 27448 5932 27488
rect 5972 27448 5981 27488
rect 6691 27448 6700 27488
rect 6740 27448 8908 27488
rect 8948 27448 8957 27488
rect 24547 27448 24556 27488
rect 24596 27448 29932 27488
rect 29972 27448 29981 27488
rect 2371 27364 2380 27404
rect 2420 27364 3724 27404
rect 3764 27364 3773 27404
rect 3821 27364 3916 27404
rect 3956 27364 3965 27404
rect 7661 27364 7756 27404
rect 7796 27364 7805 27404
rect 10243 27364 10252 27404
rect 10292 27364 10828 27404
rect 10868 27364 10877 27404
rect 26947 27364 26956 27404
rect 26996 27364 27916 27404
rect 27956 27364 27965 27404
rect 4963 27280 4972 27320
rect 5012 27280 7180 27320
rect 7220 27280 7229 27320
rect 20419 27280 20428 27320
rect 20468 27280 30988 27320
rect 31028 27280 31037 27320
rect 3103 27196 3112 27236
rect 3480 27196 3489 27236
rect 3619 27196 3628 27236
rect 3668 27196 10060 27236
rect 10100 27196 10109 27236
rect 10877 27196 10886 27236
rect 11254 27196 11263 27236
rect 15427 27196 15436 27236
rect 15476 27196 17932 27236
rect 17972 27196 17981 27236
rect 18651 27196 18660 27236
rect 19028 27196 19037 27236
rect 26425 27196 26434 27236
rect 26802 27196 26811 27236
rect 12355 27112 12364 27152
rect 12404 27112 16876 27152
rect 16916 27112 16925 27152
rect 21379 27112 21388 27152
rect 21428 27112 29644 27152
rect 29684 27112 29693 27152
rect 2275 27028 2284 27068
rect 2324 27028 10636 27068
rect 10676 27028 10685 27068
rect 14659 27028 14668 27068
rect 14708 27028 18124 27068
rect 18164 27028 18173 27068
rect 26371 27028 26380 27068
rect 26420 27028 29740 27068
rect 29780 27028 29789 27068
rect 3619 26944 3628 26984
rect 3668 26944 10156 26984
rect 10196 26944 10205 26984
rect 13507 26944 13516 26984
rect 13556 26944 15244 26984
rect 15284 26944 15293 26984
rect 15427 26944 15436 26984
rect 15476 26944 18220 26984
rect 18260 26944 18269 26984
rect 27149 26944 27244 26984
rect 27284 26944 27293 26984
rect 27715 26944 27724 26984
rect 27764 26944 29684 26984
rect 29644 26900 29684 26944
rect 2467 26860 2476 26900
rect 2516 26860 12364 26900
rect 12404 26860 12413 26900
rect 12547 26860 12556 26900
rect 12596 26860 13900 26900
rect 13940 26860 16780 26900
rect 16820 26860 16829 26900
rect 19555 26860 19564 26900
rect 19604 26860 29356 26900
rect 29396 26860 29405 26900
rect 29635 26860 29644 26900
rect 29684 26860 29693 26900
rect 4483 26776 4492 26816
rect 4532 26776 9676 26816
rect 9716 26776 9725 26816
rect 11779 26776 11788 26816
rect 11828 26776 15052 26816
rect 15092 26776 15101 26816
rect 18883 26776 18892 26816
rect 18932 26776 19660 26816
rect 19700 26776 19709 26816
rect 20227 26776 20236 26816
rect 20276 26776 20428 26816
rect 20468 26776 20477 26816
rect 23011 26776 23020 26816
rect 23060 26776 28588 26816
rect 28628 26776 28637 26816
rect 3139 26692 3148 26732
rect 3188 26692 9100 26732
rect 9140 26692 9149 26732
rect 13507 26692 13516 26732
rect 13556 26692 14860 26732
rect 14900 26692 14909 26732
rect 16195 26692 16204 26732
rect 16244 26692 19564 26732
rect 19604 26692 19613 26732
rect 21475 26692 21484 26732
rect 21524 26692 28820 26732
rect 28780 26648 28820 26692
rect 1123 26608 1132 26648
rect 1172 26608 6124 26648
rect 6164 26608 6173 26648
rect 12940 26608 16532 26648
rect 16579 26608 16588 26648
rect 16628 26608 28396 26648
rect 28436 26608 28445 26648
rect 28771 26608 28780 26648
rect 28820 26608 28829 26648
rect 12940 26564 12980 26608
rect 16492 26564 16532 26608
rect 1795 26524 1804 26564
rect 1844 26524 12980 26564
rect 14563 26524 14572 26564
rect 14612 26524 16396 26564
rect 16436 26524 16445 26564
rect 16492 26524 17260 26564
rect 17300 26524 30412 26564
rect 30452 26524 30461 26564
rect 4343 26440 4352 26480
rect 4720 26440 4729 26480
rect 5251 26440 5260 26480
rect 5300 26440 8716 26480
rect 8756 26440 9292 26480
rect 9332 26440 9341 26480
rect 12117 26440 12126 26480
rect 12494 26440 12503 26480
rect 12556 26440 17972 26480
rect 19075 26440 19084 26480
rect 19124 26440 19468 26480
rect 19508 26440 19517 26480
rect 19891 26440 19900 26480
rect 20268 26440 20277 26480
rect 22243 26440 22252 26480
rect 22292 26440 27436 26480
rect 27476 26440 27485 26480
rect 27665 26440 27674 26480
rect 28042 26440 28051 26480
rect 12556 26396 12596 26440
rect 17932 26396 17972 26440
rect 1027 26356 1036 26396
rect 1076 26356 7276 26396
rect 7316 26356 7325 26396
rect 8515 26356 8524 26396
rect 8564 26356 12596 26396
rect 13891 26356 13900 26396
rect 13940 26356 14956 26396
rect 14996 26356 15005 26396
rect 17932 26356 30988 26396
rect 31028 26356 31037 26396
rect 1219 26272 1228 26312
rect 1268 26272 4148 26312
rect 5443 26272 5452 26312
rect 5492 26272 30604 26312
rect 30644 26272 30653 26312
rect 4108 26228 4148 26272
rect 2659 26188 2668 26228
rect 2708 26188 3820 26228
rect 3860 26188 3869 26228
rect 4108 26188 5492 26228
rect 5933 26188 6028 26228
rect 6068 26188 6077 26228
rect 7075 26188 7084 26228
rect 7124 26188 7372 26228
rect 7412 26188 7421 26228
rect 11299 26188 11308 26228
rect 11348 26188 11692 26228
rect 11732 26188 11741 26228
rect 12835 26188 12844 26228
rect 12884 26188 16588 26228
rect 16628 26188 16637 26228
rect 22819 26188 22828 26228
rect 22868 26188 26572 26228
rect 26612 26188 26621 26228
rect 26755 26188 26764 26228
rect 26804 26188 27340 26228
rect 27380 26188 27389 26228
rect 27523 26188 27532 26228
rect 27572 26188 27916 26228
rect 27956 26188 28684 26228
rect 28724 26188 28733 26228
rect 835 26104 844 26144
rect 884 26104 5356 26144
rect 5396 26104 5405 26144
rect 5452 26060 5492 26188
rect 12844 26144 12884 26188
rect 6595 26104 6604 26144
rect 6644 26104 8524 26144
rect 8564 26104 8812 26144
rect 8852 26104 8861 26144
rect 11203 26104 11212 26144
rect 11252 26104 12884 26144
rect 13987 26104 13996 26144
rect 14036 26104 14860 26144
rect 14900 26104 14909 26144
rect 15245 26104 15340 26144
rect 15380 26104 15389 26144
rect 21283 26104 21292 26144
rect 21332 26104 22252 26144
rect 22292 26104 22301 26144
rect 24451 26104 24460 26144
rect 24500 26104 28972 26144
rect 29012 26104 29021 26144
rect 1411 26020 1420 26060
rect 1460 26020 3436 26060
rect 3476 26020 3485 26060
rect 3533 26020 3628 26060
rect 3668 26020 3677 26060
rect 5443 26020 5452 26060
rect 5492 26020 5501 26060
rect 11395 26020 11404 26060
rect 11444 26020 13324 26060
rect 13364 26020 13373 26060
rect 13891 26020 13900 26060
rect 13940 26020 16204 26060
rect 16244 26020 16253 26060
rect 18019 26020 18028 26060
rect 18068 26020 19756 26060
rect 19796 26020 19805 26060
rect 22147 26020 22156 26060
rect 22196 26020 24844 26060
rect 24884 26020 25228 26060
rect 25268 26020 25277 26060
rect 25987 26020 25996 26060
rect 26036 26020 27916 26060
rect 27956 26020 27965 26060
rect 2659 25936 2668 25976
rect 2708 25936 13132 25976
rect 13172 25936 13181 25976
rect 13900 25892 13940 26020
rect 23683 25936 23692 25976
rect 23732 25936 29300 25976
rect 29357 25936 29452 25976
rect 29492 25936 29501 25976
rect 29260 25892 29300 25936
rect 2083 25852 2092 25892
rect 2132 25852 9196 25892
rect 9236 25852 9245 25892
rect 11395 25852 11404 25892
rect 11444 25852 13940 25892
rect 14467 25852 14476 25892
rect 14516 25852 15820 25892
rect 15860 25852 15869 25892
rect 16771 25852 16780 25892
rect 16820 25852 20140 25892
rect 20180 25852 20189 25892
rect 24067 25852 24076 25892
rect 24116 25852 27724 25892
rect 27764 25852 27773 25892
rect 29260 25852 30028 25892
rect 30068 25852 30077 25892
rect 5251 25768 5260 25808
rect 5300 25768 27244 25808
rect 27284 25768 27293 25808
rect 27523 25768 27532 25808
rect 27572 25768 29164 25808
rect 29204 25768 29213 25808
rect 3103 25684 3112 25724
rect 3480 25684 3489 25724
rect 10877 25684 10886 25724
rect 11254 25684 11263 25724
rect 18651 25684 18660 25724
rect 19028 25684 19037 25724
rect 19555 25684 19564 25724
rect 19604 25684 20180 25724
rect 26425 25684 26434 25724
rect 26802 25684 26811 25724
rect 643 25600 652 25640
rect 692 25600 5740 25640
rect 5780 25600 5789 25640
rect 9571 25600 9580 25640
rect 9620 25600 14188 25640
rect 14228 25600 14237 25640
rect 17836 25600 19852 25640
rect 19892 25600 19901 25640
rect 17836 25556 17876 25600
rect 20140 25556 20180 25684
rect 22435 25600 22444 25640
rect 22484 25600 29356 25640
rect 29396 25600 29405 25640
rect 29923 25600 29932 25640
rect 29972 25600 29981 25640
rect 11107 25516 11116 25556
rect 11156 25516 17836 25556
rect 17876 25516 17885 25556
rect 18211 25516 18220 25556
rect 18260 25516 19660 25556
rect 19700 25516 19709 25556
rect 20131 25516 20140 25556
rect 20180 25516 20189 25556
rect 20995 25516 21004 25556
rect 21044 25516 23116 25556
rect 23156 25516 23165 25556
rect 25219 25516 25228 25556
rect 25268 25516 29452 25556
rect 29492 25516 29501 25556
rect 29932 25472 29972 25600
rect 12067 25432 12076 25472
rect 12116 25432 16780 25472
rect 16820 25432 16829 25472
rect 18979 25432 18988 25472
rect 19028 25432 22156 25472
rect 22196 25432 22828 25472
rect 22868 25432 22877 25472
rect 23203 25432 23212 25472
rect 23252 25432 29972 25472
rect 6979 25348 6988 25388
rect 7028 25348 30220 25388
rect 30260 25348 30269 25388
rect 2947 25264 2956 25304
rect 2996 25264 3148 25304
rect 3188 25264 3197 25304
rect 7363 25264 7372 25304
rect 7412 25264 8332 25304
rect 8372 25264 8908 25304
rect 8948 25264 8957 25304
rect 9091 25264 9100 25304
rect 9140 25264 24940 25304
rect 24980 25264 25420 25304
rect 25460 25264 25469 25304
rect 27331 25264 27340 25304
rect 27380 25264 28780 25304
rect 28820 25264 28829 25304
rect 2563 25180 2572 25220
rect 2612 25180 4108 25220
rect 4148 25180 7276 25220
rect 7316 25180 7325 25220
rect 9571 25180 9580 25220
rect 9620 25180 10828 25220
rect 10868 25180 10877 25220
rect 11875 25180 11884 25220
rect 11924 25180 13708 25220
rect 13748 25180 14668 25220
rect 14708 25180 15244 25220
rect 15284 25180 15436 25220
rect 15476 25180 15485 25220
rect 16300 25180 18028 25220
rect 18068 25180 18077 25220
rect 19555 25180 19564 25220
rect 19604 25180 20140 25220
rect 20180 25180 20189 25220
rect 21475 25180 21484 25220
rect 21524 25180 21580 25220
rect 21620 25180 21629 25220
rect 22915 25180 22924 25220
rect 22964 25180 26188 25220
rect 26228 25180 26237 25220
rect 16300 25136 16340 25180
rect 7843 25096 7852 25136
rect 7892 25096 9676 25136
rect 9716 25096 9725 25136
rect 11395 25096 11404 25136
rect 11444 25096 16340 25136
rect 16387 25096 16396 25136
rect 16436 25096 16972 25136
rect 17012 25096 17021 25136
rect 18787 25096 18796 25136
rect 18836 25096 19084 25136
rect 19124 25096 21772 25136
rect 21812 25096 21821 25136
rect 22540 25096 27916 25136
rect 27956 25096 27965 25136
rect 22540 25052 22580 25096
rect 8131 25012 8140 25052
rect 8180 25012 8908 25052
rect 8948 25012 8957 25052
rect 10723 25012 10732 25052
rect 10772 25012 14764 25052
rect 14804 25012 14813 25052
rect 21379 25012 21388 25052
rect 21428 25012 22580 25052
rect 22627 25012 22636 25052
rect 22676 25012 28972 25052
rect 29012 25012 29021 25052
rect 4343 24928 4352 24968
rect 4720 24928 4729 24968
rect 4963 24928 4972 24968
rect 5012 24928 9100 24968
rect 9140 24928 9149 24968
rect 12117 24928 12126 24968
rect 12494 24928 12503 24968
rect 19891 24928 19900 24968
rect 20268 24928 20277 24968
rect 27665 24928 27674 24968
rect 28042 24928 28051 24968
rect 5059 24844 5068 24884
rect 5108 24844 13900 24884
rect 13940 24844 13949 24884
rect 16771 24844 16780 24884
rect 16820 24844 17164 24884
rect 17204 24844 17213 24884
rect 20995 24844 21004 24884
rect 21044 24844 29164 24884
rect 29204 24844 29213 24884
rect 4483 24760 4492 24800
rect 4532 24760 9100 24800
rect 9140 24760 9149 24800
rect 18115 24760 18124 24800
rect 18164 24760 19468 24800
rect 19508 24760 19517 24800
rect 25699 24760 25708 24800
rect 25748 24760 28876 24800
rect 28916 24760 28925 24800
rect 8803 24676 8812 24716
rect 8852 24676 9292 24716
rect 9332 24676 9341 24716
rect 17155 24676 17164 24716
rect 17204 24676 20140 24716
rect 20180 24676 20189 24716
rect 22915 24676 22924 24716
rect 22964 24676 23596 24716
rect 23636 24676 26284 24716
rect 26324 24676 26333 24716
rect 1027 24592 1036 24632
rect 1076 24592 4204 24632
rect 4244 24592 4253 24632
rect 4387 24592 4396 24632
rect 4436 24592 5260 24632
rect 5300 24592 5309 24632
rect 13219 24592 13228 24632
rect 13268 24592 25132 24632
rect 25172 24592 25181 24632
rect 26179 24592 26188 24632
rect 26228 24592 29260 24632
rect 29300 24592 29309 24632
rect 1613 24508 1708 24548
rect 1748 24508 1757 24548
rect 3331 24508 3340 24548
rect 3380 24508 6220 24548
rect 6260 24508 6269 24548
rect 17731 24508 17740 24548
rect 17780 24508 18700 24548
rect 18740 24508 20332 24548
rect 20372 24508 20381 24548
rect 21571 24508 21580 24548
rect 21620 24508 29644 24548
rect 29684 24508 29693 24548
rect 3907 24424 3916 24464
rect 3956 24424 3965 24464
rect 8323 24424 8332 24464
rect 8372 24424 30988 24464
rect 31028 24424 31037 24464
rect 3916 24380 3956 24424
rect 3715 24340 3724 24380
rect 3764 24340 3956 24380
rect 12355 24340 12364 24380
rect 12404 24340 18796 24380
rect 18836 24340 18845 24380
rect 26371 24340 26380 24380
rect 26420 24340 27148 24380
rect 27188 24340 27197 24380
rect 10627 24256 10636 24296
rect 10676 24256 12844 24296
rect 12884 24256 12893 24296
rect 13219 24256 13228 24296
rect 13268 24256 26860 24296
rect 26900 24256 26909 24296
rect 29539 24256 29548 24296
rect 29588 24256 29597 24296
rect 3103 24172 3112 24212
rect 3480 24172 3489 24212
rect 10877 24172 10886 24212
rect 11254 24172 11263 24212
rect 18651 24172 18660 24212
rect 19028 24172 19037 24212
rect 19747 24172 19756 24212
rect 19796 24172 22540 24212
rect 22580 24172 22589 24212
rect 26425 24172 26434 24212
rect 26802 24172 26811 24212
rect 27235 24172 27244 24212
rect 27284 24172 29164 24212
rect 29204 24172 29213 24212
rect 1411 24088 1420 24128
rect 1460 24088 1804 24128
rect 1844 24088 10060 24128
rect 10100 24088 10109 24128
rect 10339 24088 10348 24128
rect 10388 24088 10732 24128
rect 10772 24088 15628 24128
rect 15668 24088 15677 24128
rect 15811 24088 15820 24128
rect 15860 24088 17356 24128
rect 17396 24088 17405 24128
rect 21283 24088 21292 24128
rect 21332 24088 25036 24128
rect 25076 24088 25085 24128
rect 25507 24088 25516 24128
rect 25556 24088 28972 24128
rect 29012 24088 29021 24128
rect 12940 24004 16300 24044
rect 16340 24004 29260 24044
rect 29300 24004 29309 24044
rect 12940 23960 12980 24004
rect 29548 23960 29588 24256
rect 1891 23920 1900 23960
rect 1940 23920 7468 23960
rect 7508 23920 8236 23960
rect 8276 23920 12980 23960
rect 13027 23920 13036 23960
rect 13076 23920 14284 23960
rect 14324 23920 14333 23960
rect 18499 23920 18508 23960
rect 18548 23920 19084 23960
rect 19124 23920 19133 23960
rect 20899 23920 20908 23960
rect 20948 23920 29588 23960
rect 931 23836 940 23876
rect 980 23836 2668 23876
rect 2708 23836 2956 23876
rect 2996 23836 7084 23876
rect 7124 23836 7133 23876
rect 11203 23836 11212 23876
rect 11252 23836 13516 23876
rect 13556 23836 13565 23876
rect 16867 23836 16876 23876
rect 16916 23836 25708 23876
rect 25748 23836 25757 23876
rect 25891 23836 25900 23876
rect 25940 23836 29548 23876
rect 29588 23836 29597 23876
rect 2755 23752 2764 23792
rect 2804 23752 8812 23792
rect 8852 23752 8861 23792
rect 14851 23752 14860 23792
rect 14900 23752 22348 23792
rect 22388 23752 22924 23792
rect 22964 23752 22973 23792
rect 23107 23752 23116 23792
rect 23156 23752 24460 23792
rect 24500 23752 29644 23792
rect 29684 23752 29693 23792
rect 5827 23668 5836 23708
rect 5876 23668 8908 23708
rect 8948 23668 8957 23708
rect 12643 23668 12652 23708
rect 12692 23668 15628 23708
rect 15668 23668 15677 23708
rect 16963 23668 16972 23708
rect 17012 23668 28876 23708
rect 28916 23668 28925 23708
rect 4291 23584 4300 23624
rect 4340 23584 4349 23624
rect 6403 23584 6412 23624
rect 6452 23584 9004 23624
rect 9044 23584 9053 23624
rect 14659 23584 14668 23624
rect 14708 23584 16300 23624
rect 16340 23584 19756 23624
rect 19796 23584 19805 23624
rect 20227 23584 20236 23624
rect 20276 23584 21388 23624
rect 21428 23584 21437 23624
rect 22915 23584 22924 23624
rect 22964 23584 23308 23624
rect 23348 23584 23357 23624
rect 25507 23584 25516 23624
rect 25556 23584 28108 23624
rect 28148 23584 28157 23624
rect 28387 23584 28396 23624
rect 28436 23584 29164 23624
rect 29204 23584 29213 23624
rect 4300 23540 4340 23584
rect 4204 23500 4340 23540
rect 6211 23500 6220 23540
rect 6260 23500 8620 23540
rect 8660 23500 8669 23540
rect 17827 23500 17836 23540
rect 17876 23500 20620 23540
rect 20660 23500 22580 23540
rect 22627 23500 22636 23540
rect 22676 23500 22685 23540
rect 25891 23500 25900 23540
rect 25940 23500 28876 23540
rect 28916 23500 28925 23540
rect 29549 23500 29644 23540
rect 29684 23500 29693 23540
rect 4204 23288 4244 23500
rect 4343 23416 4352 23456
rect 4720 23416 4729 23456
rect 12117 23416 12126 23456
rect 12494 23416 12503 23456
rect 18307 23416 18316 23456
rect 18356 23416 19468 23456
rect 19508 23416 19517 23456
rect 19891 23416 19900 23456
rect 20268 23416 20277 23456
rect 20707 23416 20716 23456
rect 20756 23416 21196 23456
rect 21236 23416 21245 23456
rect 22540 23372 22580 23500
rect 22636 23456 22676 23500
rect 22636 23416 24172 23456
rect 24212 23416 24221 23456
rect 27665 23416 27674 23456
rect 28042 23416 28051 23456
rect 6979 23332 6988 23372
rect 7028 23332 8332 23372
rect 8372 23332 8908 23372
rect 8948 23332 8957 23372
rect 12931 23332 12940 23372
rect 12980 23332 18604 23372
rect 18644 23332 18653 23372
rect 22540 23332 22732 23372
rect 22772 23332 29164 23372
rect 29204 23332 29213 23372
rect 4099 23248 4108 23288
rect 4148 23248 4244 23288
rect 7267 23248 7276 23288
rect 7316 23248 10252 23288
rect 10292 23248 11500 23288
rect 11540 23248 11549 23288
rect 11875 23248 11884 23288
rect 11924 23248 17356 23288
rect 17396 23248 17405 23288
rect 18115 23248 18124 23288
rect 18164 23248 24748 23288
rect 24788 23248 25804 23288
rect 25844 23248 25853 23288
rect 2851 23164 2860 23204
rect 2900 23164 3052 23204
rect 3092 23164 3916 23204
rect 3956 23164 27052 23204
rect 27092 23164 27101 23204
rect 3725 23080 3820 23120
rect 3860 23080 3869 23120
rect 4012 23080 4244 23120
rect 4291 23080 4300 23120
rect 4340 23080 6164 23120
rect 4012 23036 4052 23080
rect 4204 23036 4244 23080
rect 6124 23036 6164 23080
rect 7180 23080 11980 23120
rect 12020 23080 13420 23120
rect 13460 23080 13469 23120
rect 14467 23080 14476 23120
rect 14516 23080 17836 23120
rect 17876 23080 17885 23120
rect 18595 23080 18604 23120
rect 18644 23080 21580 23120
rect 21620 23080 21629 23120
rect 7180 23036 7220 23080
rect 3331 22996 3340 23036
rect 3380 22996 4052 23036
rect 4099 22996 4108 23036
rect 4148 22996 4157 23036
rect 4204 22996 5068 23036
rect 5108 22996 5117 23036
rect 6124 22996 7220 23036
rect 9773 22996 9868 23036
rect 9908 22996 9917 23036
rect 19469 22996 19564 23036
rect 19604 22996 19613 23036
rect 19747 22996 19756 23036
rect 19796 22996 24076 23036
rect 24116 22996 24125 23036
rect 26371 22996 26380 23036
rect 26420 22996 29260 23036
rect 29300 22996 29309 23036
rect 4108 22952 4148 22996
rect 3523 22912 3532 22952
rect 3572 22912 4148 22952
rect 6019 22912 6028 22952
rect 6068 22912 7412 22952
rect 7372 22868 7412 22912
rect 19564 22868 19604 22996
rect 20803 22912 20812 22952
rect 20852 22912 29164 22952
rect 29204 22912 29213 22952
rect 7372 22828 11884 22868
rect 11924 22828 11933 22868
rect 18211 22828 18220 22868
rect 18260 22828 19604 22868
rect 6403 22744 6412 22784
rect 6452 22744 8044 22784
rect 8084 22744 8093 22784
rect 3103 22660 3112 22700
rect 3480 22660 3489 22700
rect 4579 22660 4588 22700
rect 4628 22660 4876 22700
rect 4916 22660 5548 22700
rect 5588 22660 5597 22700
rect 10877 22660 10886 22700
rect 11254 22660 11263 22700
rect 18651 22660 18660 22700
rect 19028 22660 19037 22700
rect 26425 22660 26434 22700
rect 26802 22660 26811 22700
rect 5155 22576 5164 22616
rect 5204 22576 8812 22616
rect 8852 22576 8861 22616
rect 7075 22492 7084 22532
rect 7124 22492 9772 22532
rect 9812 22492 9821 22532
rect 10723 22492 10732 22532
rect 10772 22492 11116 22532
rect 11156 22492 15340 22532
rect 15380 22492 15389 22532
rect 21763 22492 21772 22532
rect 21812 22492 27052 22532
rect 27092 22492 27101 22532
rect 6499 22408 6508 22448
rect 6548 22408 7756 22448
rect 7796 22408 7805 22448
rect 8141 22408 8236 22448
rect 8276 22408 8285 22448
rect 24931 22408 24940 22448
rect 24980 22408 27244 22448
rect 27284 22408 27293 22448
rect 1219 22324 1228 22364
rect 1268 22324 9292 22364
rect 9332 22324 9341 22364
rect 10051 22324 10060 22364
rect 10100 22324 13420 22364
rect 13460 22324 13469 22364
rect 24067 22324 24076 22364
rect 24116 22324 26764 22364
rect 26804 22324 26813 22364
rect 4195 22240 4204 22280
rect 4244 22240 4396 22280
rect 4436 22240 4445 22280
rect 4963 22240 4972 22280
rect 5012 22240 6604 22280
rect 6644 22240 7564 22280
rect 7604 22240 7613 22280
rect 16291 22240 16300 22280
rect 16340 22240 17164 22280
rect 17204 22240 28780 22280
rect 28820 22240 28829 22280
rect 30019 22240 30028 22280
rect 30068 22240 30077 22280
rect 30028 22196 30068 22240
rect 4099 22156 4108 22196
rect 4148 22156 6604 22196
rect 6644 22156 6796 22196
rect 6836 22156 6845 22196
rect 20227 22156 20236 22196
rect 20276 22156 22636 22196
rect 22676 22156 22685 22196
rect 26083 22156 26092 22196
rect 26132 22156 29836 22196
rect 29876 22156 30068 22196
rect 2851 22072 2860 22112
rect 2900 22072 4588 22112
rect 4628 22072 4637 22112
rect 4689 22072 4698 22112
rect 4738 22072 4972 22112
rect 5012 22072 5021 22112
rect 5251 22072 5260 22112
rect 5300 22072 6412 22112
rect 6452 22072 6461 22112
rect 16387 22072 16396 22112
rect 16436 22072 19124 22112
rect 20707 22072 20716 22112
rect 20756 22072 21676 22112
rect 21716 22072 21725 22112
rect 26179 22072 26188 22112
rect 26228 22072 29548 22112
rect 29588 22072 30028 22112
rect 30068 22072 30077 22112
rect 19084 22028 19124 22072
rect 3427 21988 3436 22028
rect 3476 21988 9292 22028
rect 9332 21988 9341 22028
rect 19075 21988 19084 22028
rect 19124 21988 19133 22028
rect 23011 21988 23020 22028
rect 23060 21988 27148 22028
rect 27188 21988 27197 22028
rect 4343 21904 4352 21944
rect 4720 21904 4729 21944
rect 5059 21904 5068 21944
rect 5108 21904 6604 21944
rect 6644 21904 8812 21944
rect 8852 21904 8861 21944
rect 12117 21904 12126 21944
rect 12494 21904 12503 21944
rect 19891 21904 19900 21944
rect 20268 21904 20277 21944
rect 27665 21904 27674 21944
rect 28042 21904 28051 21944
rect 4195 21820 4204 21860
rect 4244 21820 4780 21860
rect 4820 21820 4829 21860
rect 6019 21820 6028 21860
rect 6068 21820 6164 21860
rect 8131 21820 8140 21860
rect 8180 21820 10060 21860
rect 10100 21820 10109 21860
rect 15523 21820 15532 21860
rect 15572 21820 17068 21860
rect 17108 21820 19276 21860
rect 19316 21820 19325 21860
rect 24643 21820 24652 21860
rect 24692 21820 26956 21860
rect 26996 21820 28972 21860
rect 29012 21820 29021 21860
rect 4483 21736 4492 21776
rect 4532 21736 5164 21776
rect 5204 21736 5213 21776
rect 3715 21652 3724 21692
rect 3764 21652 6028 21692
rect 6068 21652 6077 21692
rect 6124 21608 6164 21820
rect 6307 21736 6316 21776
rect 6356 21736 6365 21776
rect 9571 21736 9580 21776
rect 9620 21736 12652 21776
rect 12692 21736 12701 21776
rect 16867 21736 16876 21776
rect 16916 21736 19852 21776
rect 19892 21736 19901 21776
rect 20131 21736 20140 21776
rect 20180 21736 20428 21776
rect 20468 21736 30028 21776
rect 30068 21736 30077 21776
rect 6316 21608 6356 21736
rect 16877 21652 16972 21692
rect 17012 21652 17021 21692
rect 17347 21652 17356 21692
rect 17396 21652 19564 21692
rect 19604 21652 19613 21692
rect 2659 21568 2668 21608
rect 2708 21568 4628 21608
rect 4867 21568 4876 21608
rect 4916 21568 5164 21608
rect 5204 21568 5213 21608
rect 6115 21568 6124 21608
rect 6164 21568 6173 21608
rect 6316 21568 6508 21608
rect 6548 21568 6557 21608
rect 7843 21568 7852 21608
rect 7892 21568 13324 21608
rect 13364 21568 13373 21608
rect 16387 21568 16396 21608
rect 16436 21568 18412 21608
rect 18452 21568 18461 21608
rect 4588 21524 4628 21568
rect 7852 21524 7892 21568
rect 1027 21484 1036 21524
rect 1076 21484 1708 21524
rect 1748 21484 1757 21524
rect 2947 21484 2956 21524
rect 2996 21484 3628 21524
rect 3668 21484 3677 21524
rect 4579 21484 4588 21524
rect 4628 21484 7892 21524
rect 8611 21484 8620 21524
rect 8660 21484 15052 21524
rect 15092 21484 15101 21524
rect 15235 21484 15244 21524
rect 15284 21484 18028 21524
rect 18068 21484 18077 21524
rect 24355 21484 24364 21524
rect 24404 21484 28492 21524
rect 28532 21484 28541 21524
rect 2477 21400 2572 21440
rect 2612 21400 2621 21440
rect 5635 21400 5644 21440
rect 5684 21400 6028 21440
rect 6068 21400 6077 21440
rect 6691 21400 6700 21440
rect 6740 21400 30892 21440
rect 30932 21400 30941 21440
rect 3427 21316 3436 21356
rect 3476 21316 8812 21356
rect 8852 21316 8861 21356
rect 11683 21316 11692 21356
rect 11732 21316 13708 21356
rect 13748 21316 13757 21356
rect 15043 21316 15052 21356
rect 15092 21316 18124 21356
rect 18164 21316 18173 21356
rect 2736 21232 2764 21272
rect 2804 21232 2860 21272
rect 2900 21232 3572 21272
rect 3725 21232 3820 21272
rect 3860 21232 3869 21272
rect 4195 21232 4204 21272
rect 4244 21232 8908 21272
rect 8948 21232 8957 21272
rect 11587 21232 11596 21272
rect 11636 21232 15340 21272
rect 15380 21232 15389 21272
rect 3532 21188 3572 21232
rect 3103 21148 3112 21188
rect 3480 21148 3489 21188
rect 3532 21148 4300 21188
rect 4340 21148 4349 21188
rect 4867 21148 4876 21188
rect 4916 21148 4972 21188
rect 5012 21148 5021 21188
rect 5731 21148 5740 21188
rect 5780 21148 8140 21188
rect 8180 21148 8189 21188
rect 8995 21148 9004 21188
rect 9044 21148 9964 21188
rect 10004 21148 10013 21188
rect 10877 21148 10886 21188
rect 11254 21148 11263 21188
rect 13315 21148 13324 21188
rect 13364 21148 16972 21188
rect 17012 21148 17260 21188
rect 17300 21148 17309 21188
rect 18651 21148 18660 21188
rect 19028 21148 19037 21188
rect 26425 21148 26434 21188
rect 26802 21148 26811 21188
rect 28291 21148 28300 21188
rect 28340 21148 29260 21188
rect 29300 21148 29309 21188
rect 2371 21064 2380 21104
rect 2420 21064 4204 21104
rect 4244 21064 4253 21104
rect 5155 21064 5164 21104
rect 5204 21064 6892 21104
rect 6932 21064 6941 21104
rect 9091 21064 9100 21104
rect 9140 21064 9580 21104
rect 9620 21064 9629 21104
rect 10051 21064 10060 21104
rect 10100 21064 11788 21104
rect 11828 21064 11837 21104
rect 1123 20980 1132 21020
rect 1172 20980 30604 21020
rect 30644 20980 30653 21020
rect 1507 20896 1516 20936
rect 1556 20896 1804 20936
rect 1844 20896 1853 20936
rect 6499 20896 6508 20936
rect 6548 20896 30892 20936
rect 30932 20896 30941 20936
rect 739 20812 748 20852
rect 788 20812 1516 20852
rect 1556 20812 1565 20852
rect 6509 20812 6604 20852
rect 6644 20812 6653 20852
rect 7939 20812 7948 20852
rect 7988 20812 8140 20852
rect 8180 20812 8189 20852
rect 9379 20812 9388 20852
rect 9428 20812 9964 20852
rect 10004 20812 10013 20852
rect 10060 20812 10732 20852
rect 10772 20812 11636 20852
rect 13507 20812 13516 20852
rect 13556 20812 16052 20852
rect 16675 20812 16684 20852
rect 16724 20812 17836 20852
rect 17876 20812 29452 20852
rect 29492 20812 29501 20852
rect 2851 20728 2860 20768
rect 2900 20728 7468 20768
rect 7508 20728 8948 20768
rect 3715 20644 3724 20684
rect 3764 20644 8524 20684
rect 8564 20644 8573 20684
rect 8908 20600 8948 20728
rect 10060 20684 10100 20812
rect 10723 20728 10732 20768
rect 10772 20728 11020 20768
rect 11060 20728 11069 20768
rect 9667 20644 9676 20684
rect 9716 20644 10100 20684
rect 11596 20684 11636 20812
rect 16012 20768 16052 20812
rect 13699 20728 13708 20768
rect 13748 20728 14860 20768
rect 14900 20728 14909 20768
rect 16003 20728 16012 20768
rect 16052 20728 17740 20768
rect 17780 20728 17789 20768
rect 11596 20644 14572 20684
rect 14612 20644 14621 20684
rect 17443 20644 17452 20684
rect 17492 20644 17932 20684
rect 17972 20644 18412 20684
rect 18452 20644 18461 20684
rect 22723 20644 22732 20684
rect 22772 20644 23884 20684
rect 23924 20644 28684 20684
rect 28724 20644 28733 20684
rect 547 20560 556 20600
rect 596 20560 4972 20600
rect 5012 20560 5021 20600
rect 5155 20560 5164 20600
rect 5204 20560 7468 20600
rect 7508 20560 7517 20600
rect 8707 20560 8716 20600
rect 8756 20560 8812 20600
rect 8852 20560 8861 20600
rect 8908 20560 13324 20600
rect 13364 20560 13373 20600
rect 13987 20560 13996 20600
rect 14036 20560 15244 20600
rect 15284 20560 15293 20600
rect 18029 20560 18124 20600
rect 18164 20560 18173 20600
rect 20227 20560 20236 20600
rect 20276 20560 20524 20600
rect 20564 20560 20573 20600
rect 24259 20560 24268 20600
rect 24308 20560 24460 20600
rect 24500 20560 25036 20600
rect 25076 20560 28300 20600
rect 28340 20560 28349 20600
rect 13324 20516 13364 20560
rect 67 20476 76 20516
rect 116 20476 8716 20516
rect 8756 20476 8765 20516
rect 9772 20476 10252 20516
rect 10292 20476 10301 20516
rect 13324 20476 17068 20516
rect 17108 20476 17117 20516
rect 17251 20476 17260 20516
rect 17300 20476 18028 20516
rect 18068 20476 18077 20516
rect 21379 20476 21388 20516
rect 21428 20476 23404 20516
rect 23444 20476 24076 20516
rect 24116 20476 24125 20516
rect 9772 20432 9812 20476
rect 2563 20392 2572 20432
rect 2612 20392 3436 20432
rect 3476 20392 3485 20432
rect 4343 20392 4352 20432
rect 4720 20392 4729 20432
rect 6403 20392 6412 20432
rect 6452 20392 7084 20432
rect 7124 20392 7133 20432
rect 8131 20392 8140 20432
rect 8180 20392 9812 20432
rect 9859 20392 9868 20432
rect 9908 20392 9919 20432
rect 12117 20392 12126 20432
rect 12494 20392 12503 20432
rect 19891 20392 19900 20432
rect 20268 20392 20277 20432
rect 27665 20392 27674 20432
rect 28042 20392 28051 20432
rect 9868 20348 9908 20392
rect 547 20308 556 20348
rect 596 20308 5740 20348
rect 5780 20308 5789 20348
rect 6211 20308 6220 20348
rect 6260 20308 7756 20348
rect 7796 20308 7805 20348
rect 9859 20308 9868 20348
rect 9908 20308 9917 20348
rect 12835 20308 12844 20348
rect 12884 20308 14380 20348
rect 14420 20308 14429 20348
rect 1219 20224 1228 20264
rect 1268 20224 3148 20264
rect 3188 20224 3197 20264
rect 4483 20224 4492 20264
rect 4532 20224 9004 20264
rect 9044 20224 9053 20264
rect 1805 20140 1900 20180
rect 1940 20140 1949 20180
rect 3235 20140 3244 20180
rect 3284 20140 3724 20180
rect 3764 20140 3773 20180
rect 3917 20140 4012 20180
rect 4052 20140 4061 20180
rect 4973 20140 5068 20180
rect 5108 20140 5117 20180
rect 5549 20140 5644 20180
rect 5684 20140 5693 20180
rect 5827 20140 5836 20180
rect 5876 20140 5971 20180
rect 7277 20140 7372 20180
rect 7412 20140 7421 20180
rect 7555 20140 7564 20180
rect 7604 20140 7699 20180
rect 9868 20140 10196 20180
rect 10723 20140 10732 20180
rect 10772 20140 10924 20180
rect 10964 20140 10973 20180
rect 11107 20140 11116 20180
rect 11156 20140 12652 20180
rect 12692 20140 12701 20180
rect 16195 20140 16204 20180
rect 16244 20140 17452 20180
rect 17492 20140 17501 20180
rect 17837 20140 17932 20180
rect 17972 20140 17981 20180
rect 19373 20140 19468 20180
rect 19508 20140 19517 20180
rect 21389 20140 21484 20180
rect 21524 20140 21533 20180
rect 9868 20096 9908 20140
rect 1507 20056 1516 20096
rect 1556 20056 9908 20096
rect 10156 20096 10196 20140
rect 10156 20056 28588 20096
rect 28628 20056 28637 20096
rect 1699 19972 1708 20012
rect 1748 19972 1757 20012
rect 4387 19972 4396 20012
rect 4436 19972 5452 20012
rect 5492 19972 5501 20012
rect 6403 19972 6412 20012
rect 6452 19972 7372 20012
rect 7412 19972 7421 20012
rect 11107 19972 11116 20012
rect 11156 19972 12652 20012
rect 12692 19972 12701 20012
rect 15811 19972 15820 20012
rect 15860 19972 18700 20012
rect 18740 19972 18749 20012
rect 1708 19760 1748 19972
rect 2860 19888 29932 19928
rect 29972 19888 29981 19928
rect 2860 19844 2900 19888
rect 1987 19804 1996 19844
rect 2036 19804 2900 19844
rect 4195 19804 4204 19844
rect 4244 19804 4492 19844
rect 4532 19804 4541 19844
rect 5059 19804 5068 19844
rect 5108 19804 6028 19844
rect 6068 19804 6077 19844
rect 8035 19804 8044 19844
rect 8084 19804 9580 19844
rect 9620 19804 9629 19844
rect 9763 19804 9772 19844
rect 9812 19804 11596 19844
rect 11636 19804 11645 19844
rect 16867 19804 16876 19844
rect 16916 19804 17548 19844
rect 17588 19804 17597 19844
rect 1708 19720 3724 19760
rect 3764 19720 3773 19760
rect 4195 19720 4204 19760
rect 4244 19720 5164 19760
rect 5204 19720 5213 19760
rect 5731 19720 5740 19760
rect 5780 19720 7852 19760
rect 7892 19720 7901 19760
rect 8899 19720 8908 19760
rect 8948 19720 10060 19760
rect 10100 19720 10636 19760
rect 10676 19720 10685 19760
rect 12355 19720 12364 19760
rect 12404 19720 13132 19760
rect 13172 19720 13181 19760
rect 5164 19676 5204 19720
rect 3103 19636 3112 19676
rect 3480 19636 3489 19676
rect 5164 19636 6028 19676
rect 6068 19636 6700 19676
rect 6740 19636 6749 19676
rect 10877 19636 10886 19676
rect 11254 19636 11263 19676
rect 13315 19636 13324 19676
rect 13364 19636 16340 19676
rect 18651 19636 18660 19676
rect 19028 19636 19037 19676
rect 26425 19636 26434 19676
rect 26802 19636 26811 19676
rect 16300 19592 16340 19636
rect 1123 19552 1132 19592
rect 1172 19552 9964 19592
rect 10004 19552 10013 19592
rect 14947 19552 14956 19592
rect 14996 19552 15820 19592
rect 15860 19552 15869 19592
rect 16291 19552 16300 19592
rect 16340 19552 16588 19592
rect 16628 19552 16637 19592
rect 4963 19468 4972 19508
rect 5012 19468 5021 19508
rect 6211 19468 6220 19508
rect 6260 19468 7084 19508
rect 7124 19468 7133 19508
rect 9763 19468 9772 19508
rect 9812 19468 10156 19508
rect 10196 19468 10205 19508
rect 10339 19468 10348 19508
rect 10388 19468 10636 19508
rect 10676 19468 10685 19508
rect 11683 19468 11692 19508
rect 11732 19468 17548 19508
rect 17588 19468 17597 19508
rect 4972 19424 5012 19468
rect 2467 19384 2476 19424
rect 2516 19384 4876 19424
rect 4916 19384 4925 19424
rect 4972 19384 5452 19424
rect 5492 19384 8044 19424
rect 8084 19384 8093 19424
rect 9571 19384 9580 19424
rect 9620 19384 13228 19424
rect 13268 19384 13277 19424
rect 15331 19384 15340 19424
rect 15380 19384 18988 19424
rect 19028 19384 19037 19424
rect 2563 19300 2572 19340
rect 2612 19300 2956 19340
rect 2996 19300 3005 19340
rect 5347 19300 5356 19340
rect 5396 19300 5644 19340
rect 5684 19300 5693 19340
rect 6595 19300 6604 19340
rect 6644 19300 7084 19340
rect 7124 19300 7852 19340
rect 7892 19300 7901 19340
rect 14947 19300 14956 19340
rect 14996 19300 16396 19340
rect 16436 19300 16445 19340
rect 23683 19300 23692 19340
rect 23732 19300 25036 19340
rect 25076 19300 25085 19340
rect 26371 19300 26380 19340
rect 26420 19300 26429 19340
rect 26380 19256 26420 19300
rect 3725 19216 3820 19256
rect 3860 19216 3869 19256
rect 4387 19216 4396 19256
rect 4436 19216 6316 19256
rect 6356 19216 6365 19256
rect 7181 19216 7276 19256
rect 7316 19216 7325 19256
rect 8611 19216 8620 19256
rect 8660 19216 9100 19256
rect 9140 19216 9772 19256
rect 9812 19216 9821 19256
rect 10531 19216 10540 19256
rect 10580 19216 11404 19256
rect 11444 19216 11453 19256
rect 12643 19216 12652 19256
rect 12692 19216 16204 19256
rect 16244 19216 16253 19256
rect 17059 19216 17068 19256
rect 17108 19216 17644 19256
rect 17684 19216 18124 19256
rect 18164 19216 18173 19256
rect 23107 19216 23116 19256
rect 23156 19216 26420 19256
rect 1603 19132 1612 19172
rect 1652 19132 1900 19172
rect 1940 19132 1949 19172
rect 3139 19132 3148 19172
rect 3188 19132 3532 19172
rect 3572 19132 3581 19172
rect 4579 19132 4588 19172
rect 4628 19132 4637 19172
rect 6211 19132 6220 19172
rect 6260 19132 29164 19172
rect 29204 19132 29213 19172
rect 4588 19004 4628 19132
rect 4867 19048 4876 19088
rect 4916 19048 29548 19088
rect 29588 19048 29597 19088
rect 2659 18964 2668 19004
rect 2708 18964 2860 19004
rect 2900 18964 2909 19004
rect 4588 18964 4972 19004
rect 5012 18964 5021 19004
rect 5731 18964 5740 19004
rect 5780 18964 9100 19004
rect 9140 18964 9149 19004
rect 9196 18964 12940 19004
rect 12980 18964 12989 19004
rect 13123 18964 13132 19004
rect 13172 18964 15148 19004
rect 15188 18964 15197 19004
rect 15244 18964 16396 19004
rect 16436 18964 16445 19004
rect 17827 18964 17836 19004
rect 17876 18964 18412 19004
rect 18452 18964 18461 19004
rect 25699 18964 25708 19004
rect 25748 18964 26668 19004
rect 26708 18964 26717 19004
rect 9196 18920 9236 18964
rect 15244 18920 15284 18964
rect 2467 18880 2476 18920
rect 2516 18880 2572 18920
rect 2612 18880 3340 18920
rect 3380 18880 3389 18920
rect 4343 18880 4352 18920
rect 4720 18880 4729 18920
rect 5827 18880 5836 18920
rect 5876 18880 6412 18920
rect 6452 18880 6461 18920
rect 6595 18880 6604 18920
rect 6644 18880 6796 18920
rect 6836 18880 6845 18920
rect 7171 18880 7180 18920
rect 7220 18880 7852 18920
rect 7892 18880 7901 18920
rect 8045 18880 8140 18920
rect 8180 18880 8189 18920
rect 8236 18880 9236 18920
rect 9379 18880 9388 18920
rect 9428 18880 9523 18920
rect 10243 18880 10252 18920
rect 10292 18880 10732 18920
rect 10772 18880 10781 18920
rect 11011 18880 11020 18920
rect 11060 18880 11692 18920
rect 11732 18880 11741 18920
rect 12117 18880 12126 18920
rect 12494 18880 12503 18920
rect 12643 18880 12652 18920
rect 12692 18880 14284 18920
rect 14324 18880 14333 18920
rect 15235 18880 15244 18920
rect 15284 18880 15293 18920
rect 15907 18880 15916 18920
rect 15956 18880 18604 18920
rect 18644 18880 18653 18920
rect 19891 18880 19900 18920
rect 20268 18880 20277 18920
rect 27665 18880 27674 18920
rect 28042 18880 28051 18920
rect 8236 18836 8276 18880
rect 4195 18796 4204 18836
rect 4244 18796 8276 18836
rect 8707 18796 8716 18836
rect 8756 18796 18412 18836
rect 18452 18796 18988 18836
rect 19028 18796 19037 18836
rect 1699 18712 1708 18752
rect 1748 18712 2380 18752
rect 2420 18712 2429 18752
rect 2659 18700 2668 18740
rect 2708 18700 2804 18740
rect 5069 18712 5164 18752
rect 5204 18712 5213 18752
rect 5357 18712 5452 18752
rect 5492 18712 5501 18752
rect 7363 18712 7372 18752
rect 7412 18712 9196 18752
rect 9236 18712 9245 18752
rect 12940 18712 18700 18752
rect 18740 18712 18749 18752
rect 20611 18712 20620 18752
rect 20660 18712 22252 18752
rect 22292 18712 22540 18752
rect 22580 18712 27244 18752
rect 27284 18712 27293 18752
rect 2764 18668 2804 18700
rect 12940 18668 12980 18712
rect 2764 18628 2860 18668
rect 2900 18628 2909 18668
rect 6307 18628 6316 18668
rect 6356 18628 7372 18668
rect 7412 18628 7421 18668
rect 7565 18628 7660 18668
rect 7700 18628 7709 18668
rect 8515 18628 8524 18668
rect 8564 18628 12980 18668
rect 14275 18628 14284 18668
rect 14324 18628 16108 18668
rect 16148 18628 16157 18668
rect 2860 18544 28780 18584
rect 28820 18544 28829 18584
rect 2860 18500 2900 18544
rect 931 18460 940 18500
rect 980 18460 2900 18500
rect 2947 18460 2956 18500
rect 2996 18460 3052 18500
rect 3092 18460 3101 18500
rect 6509 18460 6604 18500
rect 6644 18460 6653 18500
rect 6787 18460 6796 18500
rect 6836 18460 7564 18500
rect 7604 18460 7988 18500
rect 8419 18460 8428 18500
rect 8468 18460 8620 18500
rect 8660 18460 8669 18500
rect 13795 18460 13804 18500
rect 13844 18460 15436 18500
rect 15476 18460 15485 18500
rect 16579 18460 16588 18500
rect 16628 18460 16972 18500
rect 17012 18460 17021 18500
rect 7948 18416 7988 18460
rect 2467 18376 2476 18416
rect 2516 18376 2668 18416
rect 2708 18376 2717 18416
rect 2851 18376 2860 18416
rect 2900 18376 7700 18416
rect 7948 18376 9196 18416
rect 9236 18376 9245 18416
rect 9388 18376 28684 18416
rect 28724 18376 28733 18416
rect 7660 18332 7700 18376
rect 1699 18292 1708 18332
rect 1748 18292 2092 18332
rect 2132 18292 2764 18332
rect 2804 18292 2813 18332
rect 2947 18292 2956 18332
rect 2996 18292 3436 18332
rect 3476 18292 3485 18332
rect 5827 18292 5836 18332
rect 5876 18292 7564 18332
rect 7604 18292 7613 18332
rect 7660 18292 8660 18332
rect 8620 18248 8660 18292
rect 9388 18248 9428 18376
rect 10445 18292 10540 18332
rect 10580 18292 10589 18332
rect 11885 18292 11980 18332
rect 12020 18292 12029 18332
rect 26659 18292 26668 18332
rect 26708 18292 27628 18332
rect 27668 18292 27677 18332
rect 460 18208 652 18248
rect 692 18208 701 18248
rect 1795 18208 1804 18248
rect 1844 18208 3724 18248
rect 3764 18208 3773 18248
rect 7075 18208 7084 18248
rect 7124 18208 7660 18248
rect 7700 18208 7709 18248
rect 8620 18208 9428 18248
rect 10435 18208 10444 18248
rect 10484 18208 15340 18248
rect 15380 18208 16684 18248
rect 16724 18208 16733 18248
rect 460 18164 500 18208
rect 451 18124 460 18164
rect 500 18124 509 18164
rect 3103 18124 3112 18164
rect 3480 18124 3489 18164
rect 7468 18124 8812 18164
rect 8852 18124 8861 18164
rect 10877 18124 10886 18164
rect 11254 18124 11263 18164
rect 11491 18124 11500 18164
rect 11540 18124 16108 18164
rect 16148 18124 16157 18164
rect 18651 18124 18660 18164
rect 19028 18124 19037 18164
rect 26425 18124 26434 18164
rect 26802 18124 26811 18164
rect 6211 18040 6220 18080
rect 6260 18040 7276 18080
rect 7316 18040 7372 18080
rect 7412 18040 7421 18080
rect 7468 17996 7508 18124
rect 7555 18040 7564 18080
rect 7604 18040 13420 18080
rect 13460 18040 13469 18080
rect 15235 18040 15244 18080
rect 15284 18040 17164 18080
rect 17204 18040 17213 18080
rect 355 17956 364 17996
rect 404 17956 652 17996
rect 692 17956 701 17996
rect 1123 17956 1132 17996
rect 1172 17956 2668 17996
rect 2708 17956 2717 17996
rect 6691 17956 6700 17996
rect 6740 17956 7508 17996
rect 8131 17956 8140 17996
rect 8180 17956 8332 17996
rect 8372 17956 8381 17996
rect 9667 17956 9676 17996
rect 9716 17956 9772 17996
rect 9812 17956 9821 17996
rect 12259 17956 12268 17996
rect 12308 17956 12556 17996
rect 12596 17956 13132 17996
rect 13172 17956 13181 17996
rect 15811 17956 15820 17996
rect 15860 17956 16876 17996
rect 16916 17956 16925 17996
rect 931 17872 940 17912
rect 980 17872 1804 17912
rect 1844 17872 2380 17912
rect 2420 17872 2572 17912
rect 2612 17872 2621 17912
rect 3907 17872 3916 17912
rect 3956 17872 4532 17912
rect 4867 17872 4876 17912
rect 4916 17872 6508 17912
rect 6548 17872 6557 17912
rect 7267 17872 7276 17912
rect 7316 17872 12460 17912
rect 12500 17872 12509 17912
rect 12940 17872 28012 17912
rect 28052 17872 28061 17912
rect 4492 17828 4532 17872
rect 12940 17828 12980 17872
rect 1699 17788 1708 17828
rect 1748 17788 2188 17828
rect 2228 17788 2237 17828
rect 3715 17788 3724 17828
rect 3764 17788 4436 17828
rect 4492 17788 12980 17828
rect 14755 17788 14764 17828
rect 14804 17788 16780 17828
rect 16820 17788 17836 17828
rect 17876 17788 18028 17828
rect 18068 17788 18077 17828
rect 18499 17788 18508 17828
rect 18548 17788 18892 17828
rect 18932 17788 18941 17828
rect 4396 17744 4436 17788
rect 2275 17704 2284 17744
rect 2324 17704 2860 17744
rect 2900 17704 2909 17744
rect 3235 17704 3244 17744
rect 3284 17704 3628 17744
rect 3668 17704 3677 17744
rect 4195 17704 4204 17744
rect 4244 17704 4253 17744
rect 4396 17704 7372 17744
rect 7412 17704 7421 17744
rect 7555 17704 7564 17744
rect 7604 17704 7660 17744
rect 7700 17704 7709 17744
rect 7939 17704 7948 17744
rect 7988 17704 8524 17744
rect 8564 17704 8573 17744
rect 8899 17704 8908 17744
rect 8948 17704 9484 17744
rect 9524 17704 9533 17744
rect 9773 17704 9868 17744
rect 9908 17704 9917 17744
rect 11683 17704 11692 17744
rect 11732 17704 16204 17744
rect 16244 17704 17932 17744
rect 17972 17704 17981 17744
rect 21379 17704 21388 17744
rect 21428 17704 23116 17744
rect 23156 17704 23165 17744
rect 3244 17660 3284 17704
rect 4204 17660 4244 17704
rect 2659 17620 2668 17660
rect 2708 17620 3284 17660
rect 3523 17620 3532 17660
rect 3572 17620 4244 17660
rect 4973 17620 5068 17660
rect 5108 17620 5117 17660
rect 7363 17620 7372 17660
rect 7412 17620 8044 17660
rect 8084 17620 12940 17660
rect 12980 17620 12989 17660
rect 23299 17620 23308 17660
rect 23348 17620 27052 17660
rect 27092 17620 27101 17660
rect 4867 17536 4876 17576
rect 4916 17536 6604 17576
rect 6644 17536 6653 17576
rect 6979 17536 6988 17576
rect 7028 17536 8524 17576
rect 8564 17536 8573 17576
rect 9187 17536 9196 17576
rect 9236 17536 9868 17576
rect 9908 17536 9917 17576
rect 11395 17536 11404 17576
rect 11444 17536 11788 17576
rect 11828 17536 11837 17576
rect 11884 17536 12268 17576
rect 12308 17536 12317 17576
rect 12835 17536 12844 17576
rect 12884 17536 15244 17576
rect 15284 17536 15436 17576
rect 15476 17536 15485 17576
rect 1795 17452 1804 17492
rect 1844 17452 2860 17492
rect 2900 17452 2909 17492
rect 4771 17452 4780 17492
rect 4820 17452 5452 17492
rect 5492 17452 5501 17492
rect 6403 17452 6412 17492
rect 6452 17452 6700 17492
rect 6740 17452 6749 17492
rect 6988 17408 7028 17536
rect 11884 17492 11924 17536
rect 8995 17452 9004 17492
rect 9044 17452 9388 17492
rect 9428 17452 11924 17492
rect 643 17368 652 17408
rect 692 17368 844 17408
rect 884 17368 893 17408
rect 4343 17368 4352 17408
rect 4720 17368 4729 17408
rect 4780 17368 5260 17408
rect 5300 17368 5309 17408
rect 5539 17368 5548 17408
rect 5588 17368 7028 17408
rect 7363 17368 7372 17408
rect 7412 17368 9772 17408
rect 9812 17368 9821 17408
rect 11405 17368 11500 17408
rect 11540 17368 11549 17408
rect 12117 17368 12126 17408
rect 12494 17368 12503 17408
rect 19891 17368 19900 17408
rect 20268 17368 20277 17408
rect 27665 17368 27674 17408
rect 28042 17368 28051 17408
rect 4780 17324 4820 17368
rect 355 17284 364 17324
rect 404 17284 4820 17324
rect 5059 17284 5068 17324
rect 5108 17284 5836 17324
rect 5876 17284 5885 17324
rect 8899 17284 8908 17324
rect 8948 17284 9868 17324
rect 9908 17284 9917 17324
rect 1123 17200 1132 17240
rect 1172 17200 1228 17240
rect 1268 17200 1277 17240
rect 5731 17200 5740 17240
rect 5780 17200 7948 17240
rect 7988 17200 7997 17240
rect 9763 17200 9772 17240
rect 9812 17200 12652 17240
rect 12692 17200 12701 17240
rect 1987 17116 1996 17156
rect 2036 17116 2476 17156
rect 2516 17116 2525 17156
rect 4771 17116 4780 17156
rect 4820 17116 7660 17156
rect 7700 17116 7709 17156
rect 8323 17116 8332 17156
rect 8372 17116 8428 17156
rect 8468 17116 8477 17156
rect 10723 17116 10732 17156
rect 10772 17116 14092 17156
rect 14132 17116 14141 17156
rect 5059 17032 5068 17072
rect 5108 17032 6316 17072
rect 6356 17032 6365 17072
rect 8515 17032 8524 17072
rect 8564 17032 9676 17072
rect 9716 17032 9725 17072
rect 10819 17032 10828 17072
rect 10868 17032 12940 17072
rect 12980 17032 13228 17072
rect 13268 17032 13277 17072
rect 15427 17032 15436 17072
rect 15476 17032 16012 17072
rect 16052 17032 16061 17072
rect 18883 17032 18892 17072
rect 18932 17032 19948 17072
rect 19988 17032 20428 17072
rect 20468 17032 20477 17072
rect 20899 17032 20908 17072
rect 20948 17032 23116 17072
rect 23156 17032 23165 17072
rect 1219 16948 1228 16988
rect 1268 16948 1900 16988
rect 1940 16948 2284 16988
rect 2324 16948 2572 16988
rect 2612 16948 2621 16988
rect 5443 16948 5452 16988
rect 5492 16948 5836 16988
rect 5876 16948 5885 16988
rect 6316 16904 6356 17032
rect 9283 16948 9292 16988
rect 9332 16948 20140 16988
rect 20180 16948 20189 16988
rect 5539 16864 5548 16904
rect 5588 16864 5740 16904
rect 5780 16864 5789 16904
rect 6316 16864 10444 16904
rect 10484 16864 10493 16904
rect 15139 16864 15148 16904
rect 15188 16864 16492 16904
rect 16532 16864 16541 16904
rect 19459 16864 19468 16904
rect 19508 16864 21196 16904
rect 21236 16864 21245 16904
rect 2371 16780 2380 16820
rect 2420 16780 2668 16820
rect 2708 16780 2717 16820
rect 8803 16780 8812 16820
rect 8852 16780 9196 16820
rect 9236 16780 9484 16820
rect 9524 16780 9533 16820
rect 9859 16780 9868 16820
rect 9908 16780 11980 16820
rect 12020 16780 12029 16820
rect 12355 16780 12364 16820
rect 12404 16780 13420 16820
rect 13460 16780 13469 16820
rect 14467 16780 14476 16820
rect 14516 16780 15244 16820
rect 15284 16780 15293 16820
rect 15811 16780 15820 16820
rect 15860 16780 16876 16820
rect 16916 16780 16925 16820
rect 18979 16780 18988 16820
rect 19028 16780 19180 16820
rect 19220 16780 20908 16820
rect 20948 16780 20957 16820
rect 9667 16696 9676 16736
rect 9716 16696 11884 16736
rect 11924 16696 11933 16736
rect 15820 16652 15860 16780
rect 15917 16696 16012 16736
rect 16052 16696 21868 16736
rect 21908 16696 21917 16736
rect 3103 16612 3112 16652
rect 3480 16612 3489 16652
rect 10339 16612 10348 16652
rect 10388 16612 10772 16652
rect 10877 16612 10886 16652
rect 11254 16612 11263 16652
rect 11683 16612 11692 16652
rect 11732 16612 15860 16652
rect 18651 16612 18660 16652
rect 19028 16612 19037 16652
rect 26425 16612 26434 16652
rect 26802 16612 26811 16652
rect 10732 16568 10772 16612
rect 11692 16568 11732 16612
rect 4867 16528 4876 16568
rect 4916 16528 6124 16568
rect 6164 16528 6173 16568
rect 7267 16528 7276 16568
rect 7316 16528 8524 16568
rect 8564 16528 8573 16568
rect 10541 16528 10636 16568
rect 10676 16528 10685 16568
rect 10732 16528 11732 16568
rect 12940 16528 15148 16568
rect 15188 16528 15197 16568
rect 15619 16528 15628 16568
rect 15668 16528 17260 16568
rect 17300 16528 17309 16568
rect 12940 16484 12980 16528
rect 5059 16444 5068 16484
rect 5108 16444 5644 16484
rect 5684 16444 5693 16484
rect 6307 16444 6316 16484
rect 6356 16444 7084 16484
rect 7124 16444 7133 16484
rect 10435 16444 10444 16484
rect 10484 16444 12980 16484
rect 13699 16444 13708 16484
rect 13748 16444 14092 16484
rect 14132 16444 14141 16484
rect 14659 16444 14668 16484
rect 14708 16444 16684 16484
rect 16724 16444 17548 16484
rect 17588 16444 17597 16484
rect 21475 16444 21484 16484
rect 21524 16444 22348 16484
rect 22388 16444 22397 16484
rect 3811 16360 3820 16400
rect 3860 16360 6412 16400
rect 6452 16360 6461 16400
rect 8995 16360 9004 16400
rect 9044 16360 9196 16400
rect 9236 16360 11020 16400
rect 11060 16360 11069 16400
rect 12451 16360 12460 16400
rect 12500 16360 12652 16400
rect 12692 16360 12701 16400
rect 12835 16360 12844 16400
rect 12884 16360 20428 16400
rect 20468 16360 20477 16400
rect 3811 16276 3820 16316
rect 3860 16276 4492 16316
rect 4532 16276 4541 16316
rect 4675 16276 4684 16316
rect 4724 16276 6796 16316
rect 6836 16276 6845 16316
rect 8131 16276 8140 16316
rect 8180 16276 19372 16316
rect 19412 16276 19421 16316
rect 20611 16276 20620 16316
rect 20660 16276 20908 16316
rect 20948 16276 22060 16316
rect 22100 16276 22828 16316
rect 22868 16276 22877 16316
rect 23491 16276 23500 16316
rect 23540 16276 24844 16316
rect 24884 16276 25612 16316
rect 25652 16276 26860 16316
rect 26900 16276 26909 16316
rect 2371 16192 2380 16232
rect 2420 16192 13132 16232
rect 13172 16192 13181 16232
rect 13900 16192 19948 16232
rect 19988 16192 19997 16232
rect 13900 16148 13940 16192
rect 3811 16108 3820 16148
rect 3860 16108 4684 16148
rect 4724 16108 4733 16148
rect 6979 16108 6988 16148
rect 7028 16108 7564 16148
rect 7604 16108 7613 16148
rect 8227 16108 8236 16148
rect 8276 16108 9004 16148
rect 9044 16108 9053 16148
rect 11203 16108 11212 16148
rect 11252 16108 11788 16148
rect 11828 16108 13940 16148
rect 15235 16108 15244 16148
rect 15284 16108 16108 16148
rect 16148 16108 16157 16148
rect 16387 16108 16396 16148
rect 16436 16108 17548 16148
rect 17588 16108 17597 16148
rect 20227 16108 20236 16148
rect 20276 16108 21004 16148
rect 21044 16108 21053 16148
rect 16396 16064 16436 16108
rect 1325 16024 1420 16064
rect 1460 16024 1469 16064
rect 2755 16024 2764 16064
rect 2804 16024 13324 16064
rect 13364 16024 13373 16064
rect 14275 16024 14284 16064
rect 14324 16024 16436 16064
rect 20323 16024 20332 16064
rect 20372 16024 20524 16064
rect 20564 16024 23308 16064
rect 23348 16024 23357 16064
rect 3619 15940 3628 15980
rect 3668 15940 12844 15980
rect 12884 15940 12893 15980
rect 12940 15940 15436 15980
rect 15476 15940 15485 15980
rect 16781 15940 16876 15980
rect 16916 15940 16925 15980
rect 12940 15896 12980 15940
rect 4343 15856 4352 15896
rect 4720 15856 4729 15896
rect 5155 15856 5164 15896
rect 5204 15856 5356 15896
rect 5396 15856 10252 15896
rect 10292 15856 10301 15896
rect 10435 15856 10444 15896
rect 10484 15856 11404 15896
rect 11444 15856 11453 15896
rect 12117 15856 12126 15896
rect 12494 15856 12503 15896
rect 12931 15856 12940 15896
rect 12980 15856 12989 15896
rect 19891 15856 19900 15896
rect 20268 15856 20277 15896
rect 27665 15856 27674 15896
rect 28042 15856 28051 15896
rect 3715 15772 3724 15812
rect 3764 15772 6028 15812
rect 6068 15772 6077 15812
rect 6124 15772 9484 15812
rect 9524 15772 9533 15812
rect 6124 15728 6164 15772
rect 10252 15728 10292 15856
rect 11299 15772 11308 15812
rect 11348 15772 13708 15812
rect 13748 15772 13757 15812
rect 15341 15772 15436 15812
rect 15476 15772 15485 15812
rect 23683 15772 23692 15812
rect 23732 15772 23741 15812
rect 1699 15688 1708 15728
rect 1748 15688 1804 15728
rect 1844 15688 1853 15728
rect 4003 15688 4012 15728
rect 4052 15688 5068 15728
rect 5108 15688 5548 15728
rect 5588 15688 5597 15728
rect 5923 15688 5932 15728
rect 5972 15688 6164 15728
rect 7564 15688 9100 15728
rect 9140 15688 9149 15728
rect 10252 15688 12460 15728
rect 12500 15688 12509 15728
rect 12835 15688 12844 15728
rect 12884 15688 14476 15728
rect 14516 15688 14525 15728
rect 21667 15688 21676 15728
rect 21716 15688 23020 15728
rect 23060 15688 23069 15728
rect 7564 15644 7604 15688
rect 23692 15644 23732 15772
rect 1987 15604 1996 15644
rect 2036 15604 2284 15644
rect 2324 15604 2333 15644
rect 4099 15604 4108 15644
rect 4148 15604 7604 15644
rect 7651 15604 7660 15644
rect 7700 15604 8332 15644
rect 8372 15604 8381 15644
rect 8515 15604 8524 15644
rect 8564 15604 9484 15644
rect 9524 15604 9533 15644
rect 10435 15604 10444 15644
rect 10484 15604 16300 15644
rect 16340 15604 16349 15644
rect 22435 15604 22444 15644
rect 22484 15604 23732 15644
rect 4387 15520 4396 15560
rect 4436 15520 5836 15560
rect 5876 15520 5885 15560
rect 6307 15520 6316 15560
rect 6356 15520 7180 15560
rect 7220 15520 7229 15560
rect 10147 15520 10156 15560
rect 10196 15520 12172 15560
rect 12212 15520 16780 15560
rect 16820 15520 16829 15560
rect 18403 15520 18412 15560
rect 18452 15520 18700 15560
rect 18740 15520 18749 15560
rect 26083 15520 26092 15560
rect 26132 15520 28108 15560
rect 28148 15520 28157 15560
rect 1411 15436 1420 15476
rect 1460 15436 8236 15476
rect 8276 15436 8285 15476
rect 9955 15436 9964 15476
rect 10004 15436 10348 15476
rect 10388 15436 10397 15476
rect 11971 15436 11980 15476
rect 12020 15436 12844 15476
rect 12884 15436 12893 15476
rect 14275 15436 14284 15476
rect 14324 15436 17644 15476
rect 17684 15436 17693 15476
rect 23395 15436 23404 15476
rect 23444 15436 23788 15476
rect 23828 15436 23837 15476
rect 5443 15352 5452 15392
rect 5492 15352 7276 15392
rect 7316 15352 7325 15392
rect 7757 15352 7852 15392
rect 7892 15352 7901 15392
rect 11299 15352 11308 15392
rect 11348 15352 12308 15392
rect 17155 15352 17164 15392
rect 17204 15352 17452 15392
rect 17492 15352 17501 15392
rect 19459 15352 19468 15392
rect 19508 15352 20044 15392
rect 20084 15352 20093 15392
rect 20419 15352 20428 15392
rect 20468 15352 20908 15392
rect 20948 15352 21100 15392
rect 21140 15352 21149 15392
rect 21571 15352 21580 15392
rect 21620 15352 22156 15392
rect 22196 15352 23884 15392
rect 23924 15352 23933 15392
rect 5155 15268 5164 15308
rect 5204 15268 6604 15308
rect 6644 15268 7372 15308
rect 7412 15268 7421 15308
rect 11203 15268 11212 15308
rect 11252 15268 12172 15308
rect 12212 15268 12221 15308
rect 12268 15224 12308 15352
rect 12355 15268 12364 15308
rect 12404 15268 12652 15308
rect 12692 15268 12701 15308
rect 12931 15268 12940 15308
rect 12980 15268 13132 15308
rect 13172 15268 13181 15308
rect 14179 15268 14188 15308
rect 14228 15268 18412 15308
rect 18452 15268 18461 15308
rect 2381 15184 2476 15224
rect 2516 15184 2525 15224
rect 2659 15184 2668 15224
rect 2708 15184 8908 15224
rect 8948 15184 8957 15224
rect 12268 15184 16396 15224
rect 16436 15184 16445 15224
rect 3103 15100 3112 15140
rect 3480 15100 3489 15140
rect 4579 15100 4588 15140
rect 4628 15100 5644 15140
rect 5684 15100 5693 15140
rect 5827 15100 5836 15140
rect 5876 15100 9388 15140
rect 9428 15100 9437 15140
rect 10435 15100 10444 15140
rect 10484 15100 10732 15140
rect 10772 15100 10781 15140
rect 10877 15100 10886 15140
rect 11254 15100 11263 15140
rect 18651 15100 18660 15140
rect 19028 15100 19037 15140
rect 26425 15100 26434 15140
rect 26802 15100 26811 15140
rect 10732 15056 10772 15100
rect 2563 15016 2572 15056
rect 2612 15016 9484 15056
rect 9524 15016 9533 15056
rect 10732 15016 11348 15056
rect 11308 14972 11348 15016
rect 4195 14932 4204 14972
rect 4244 14932 5452 14972
rect 5492 14932 5501 14972
rect 10435 14932 10444 14972
rect 10484 14932 11116 14972
rect 11156 14932 11165 14972
rect 11299 14932 11308 14972
rect 11348 14932 11357 14972
rect 11875 14932 11884 14972
rect 11924 14932 12844 14972
rect 12884 14932 14284 14972
rect 14324 14932 14333 14972
rect 18307 14932 18316 14972
rect 18356 14932 18988 14972
rect 19028 14932 19037 14972
rect 1699 14848 1708 14888
rect 1748 14848 19468 14888
rect 19508 14848 19517 14888
rect 20707 14848 20716 14888
rect 20756 14848 21676 14888
rect 21716 14848 22924 14888
rect 22964 14848 22973 14888
rect 4195 14764 4204 14804
rect 4244 14764 6412 14804
rect 6452 14764 6461 14804
rect 7747 14764 7756 14804
rect 7796 14764 8948 14804
rect 10627 14764 10636 14804
rect 10676 14764 10828 14804
rect 10868 14764 10877 14804
rect 12940 14764 18796 14804
rect 18836 14764 18845 14804
rect 19267 14764 19276 14804
rect 19316 14764 19756 14804
rect 19796 14764 20044 14804
rect 20084 14764 20093 14804
rect 21091 14764 21100 14804
rect 21140 14764 24076 14804
rect 24116 14764 24125 14804
rect 8908 14720 8948 14764
rect 12940 14720 12980 14764
rect 8908 14680 12980 14720
rect 16099 14680 16108 14720
rect 16148 14680 17260 14720
rect 17300 14680 17309 14720
rect 18595 14680 18604 14720
rect 18644 14680 19180 14720
rect 19220 14680 19229 14720
rect 5923 14596 5932 14636
rect 5972 14596 6412 14636
rect 6452 14596 6461 14636
rect 6595 14596 6604 14636
rect 6644 14596 8908 14636
rect 8948 14596 8957 14636
rect 9763 14596 9772 14636
rect 9812 14596 11980 14636
rect 12020 14596 12404 14636
rect 13987 14596 13996 14636
rect 14036 14596 16588 14636
rect 16628 14596 16972 14636
rect 17012 14596 17021 14636
rect 20995 14596 21004 14636
rect 21044 14596 21388 14636
rect 21428 14596 21437 14636
rect 21955 14596 21964 14636
rect 22004 14596 22444 14636
rect 22484 14596 22493 14636
rect 4012 14512 4588 14552
rect 4628 14512 4637 14552
rect 11107 14512 11116 14552
rect 11156 14512 11500 14552
rect 11540 14512 11549 14552
rect 4012 14300 4052 14512
rect 12364 14468 12404 14596
rect 13219 14512 13228 14552
rect 13268 14512 14188 14552
rect 14228 14512 17260 14552
rect 17300 14512 17309 14552
rect 18883 14512 18892 14552
rect 18932 14512 19660 14552
rect 19700 14512 20140 14552
rect 20180 14512 20189 14552
rect 23587 14512 23596 14552
rect 23636 14512 23884 14552
rect 23924 14512 23933 14552
rect 4099 14428 4108 14468
rect 4148 14428 4204 14468
rect 4244 14428 5932 14468
rect 5972 14428 10636 14468
rect 10676 14428 10685 14468
rect 12364 14428 13076 14468
rect 23203 14428 23212 14468
rect 23252 14428 23924 14468
rect 13036 14384 13076 14428
rect 4343 14344 4352 14384
rect 4720 14344 4729 14384
rect 10147 14344 10156 14384
rect 10196 14344 11596 14384
rect 11636 14344 11645 14384
rect 12117 14344 12126 14384
rect 12494 14344 12503 14384
rect 13036 14344 13324 14384
rect 13364 14344 13373 14384
rect 14947 14344 14956 14384
rect 14996 14344 15820 14384
rect 15860 14344 15869 14384
rect 18019 14344 18028 14384
rect 18068 14344 18892 14384
rect 18932 14344 18941 14384
rect 19891 14344 19900 14384
rect 20268 14344 20277 14384
rect 4012 14260 4108 14300
rect 4148 14260 4157 14300
rect 10339 14260 10348 14300
rect 10388 14260 11788 14300
rect 11828 14260 11980 14300
rect 12020 14260 13996 14300
rect 14036 14260 14045 14300
rect 18028 14216 18068 14344
rect 9379 14176 9388 14216
rect 9428 14176 10100 14216
rect 11395 14176 11404 14216
rect 11444 14176 12268 14216
rect 12308 14176 18068 14216
rect 18604 14176 19180 14216
rect 19220 14176 19468 14216
rect 19508 14176 19517 14216
rect 20131 14176 20140 14216
rect 20180 14176 20189 14216
rect 21379 14176 21388 14216
rect 21428 14176 23404 14216
rect 23444 14176 23453 14216
rect 1603 14092 1612 14132
rect 1652 14092 1900 14132
rect 1940 14092 1949 14132
rect 2371 14092 2380 14132
rect 2420 14092 5836 14132
rect 5876 14092 5885 14132
rect 6115 14092 6124 14132
rect 6164 14092 6604 14132
rect 6644 14092 6653 14132
rect 8803 14092 8812 14132
rect 8852 14092 9580 14132
rect 9620 14092 9629 14132
rect 10060 14048 10100 14176
rect 11491 14092 11500 14132
rect 11540 14092 12940 14132
rect 12980 14092 12989 14132
rect 15917 14092 16012 14132
rect 16052 14092 16061 14132
rect 7949 14008 8044 14048
rect 8084 14008 8093 14048
rect 8323 14008 8332 14048
rect 8372 14008 8716 14048
rect 8756 14008 8765 14048
rect 10051 14008 10060 14048
rect 10100 14008 10540 14048
rect 10580 14008 12748 14048
rect 12788 14008 12797 14048
rect 14659 14008 14668 14048
rect 14708 14008 15340 14048
rect 15380 14008 15389 14048
rect 16685 14008 16780 14048
rect 16820 14008 16829 14048
rect 17731 14008 17740 14048
rect 17780 14008 18412 14048
rect 18452 14008 18461 14048
rect 5635 13924 5644 13964
rect 5684 13924 9580 13964
rect 9620 13924 9772 13964
rect 9812 13924 9821 13964
rect 12451 13924 12460 13964
rect 12500 13924 18508 13964
rect 18548 13924 18557 13964
rect 18604 13880 18644 14176
rect 20140 14048 20180 14176
rect 23884 14048 23924 14428
rect 27665 14344 27674 14384
rect 28042 14344 28051 14384
rect 20140 14008 20812 14048
rect 20852 14008 22444 14048
rect 22484 14008 22924 14048
rect 22964 14008 22973 14048
rect 23875 14008 23884 14048
rect 23924 14008 23933 14048
rect 18691 13924 18700 13964
rect 18740 13924 21388 13964
rect 21428 13924 22348 13964
rect 22388 13924 22397 13964
rect 22723 13924 22732 13964
rect 22772 13924 23308 13964
rect 23348 13924 23357 13964
rect 23587 13924 23596 13964
rect 23636 13924 27052 13964
rect 27092 13924 27101 13964
rect 67 13840 76 13880
rect 116 13840 556 13880
rect 596 13840 605 13880
rect 4291 13840 4300 13880
rect 4340 13840 5356 13880
rect 5396 13840 7276 13880
rect 7316 13840 7468 13880
rect 7508 13840 7517 13880
rect 7747 13840 7756 13880
rect 7796 13840 18644 13880
rect 19747 13840 19756 13880
rect 19796 13840 21484 13880
rect 21524 13840 21533 13880
rect 21955 13840 21964 13880
rect 22004 13840 24844 13880
rect 24884 13840 24893 13880
rect 3427 13756 3436 13796
rect 3476 13756 3628 13796
rect 3668 13756 3677 13796
rect 8429 13756 8524 13796
rect 8564 13756 8573 13796
rect 10243 13756 10252 13796
rect 10292 13756 29068 13796
rect 29108 13756 29117 13796
rect 9091 13672 9100 13712
rect 9140 13672 16876 13712
rect 16916 13672 16925 13712
rect 18403 13672 18412 13712
rect 18452 13672 19948 13712
rect 19988 13672 19997 13712
rect 21187 13672 21196 13712
rect 21236 13672 22156 13712
rect 22196 13672 22205 13712
rect 3103 13588 3112 13628
rect 3480 13588 3489 13628
rect 10877 13588 10886 13628
rect 11254 13588 11263 13628
rect 12739 13588 12748 13628
rect 12788 13588 16012 13628
rect 16052 13588 16061 13628
rect 18651 13588 18660 13628
rect 19028 13588 19037 13628
rect 26425 13588 26434 13628
rect 26802 13588 26811 13628
rect 11395 13504 11404 13544
rect 11444 13504 13516 13544
rect 13556 13504 13565 13544
rect 21859 13504 21868 13544
rect 21908 13504 23980 13544
rect 24020 13504 24029 13544
rect 24163 13504 24172 13544
rect 24212 13504 28780 13544
rect 28820 13504 28829 13544
rect 26764 13460 26804 13504
rect 5827 13420 5836 13460
rect 5876 13420 6220 13460
rect 6260 13420 6269 13460
rect 18883 13420 18892 13460
rect 18932 13420 19276 13460
rect 19316 13420 19325 13460
rect 20803 13420 20812 13460
rect 20852 13420 22060 13460
rect 22100 13420 22109 13460
rect 26755 13420 26764 13460
rect 26804 13420 26813 13460
rect 6115 13336 6124 13376
rect 6164 13336 6604 13376
rect 6644 13336 6653 13376
rect 8611 13336 8620 13376
rect 8660 13336 8908 13376
rect 8948 13336 8957 13376
rect 10627 13336 10636 13376
rect 10676 13336 11404 13376
rect 11444 13336 11453 13376
rect 18403 13336 18412 13376
rect 18452 13336 18700 13376
rect 18740 13336 18749 13376
rect 22339 13336 22348 13376
rect 22388 13336 28820 13376
rect 28780 13292 28820 13336
rect 5539 13252 5548 13292
rect 5588 13252 8908 13292
rect 8948 13252 9868 13292
rect 9908 13252 9917 13292
rect 10051 13252 10060 13292
rect 10100 13252 11212 13292
rect 11252 13252 11261 13292
rect 15235 13252 15244 13292
rect 15284 13252 15724 13292
rect 15764 13252 16300 13292
rect 16340 13252 16349 13292
rect 19459 13252 19468 13292
rect 19508 13252 19660 13292
rect 19700 13252 19709 13292
rect 20803 13252 20812 13292
rect 20852 13252 22540 13292
rect 22580 13252 22589 13292
rect 28771 13252 28780 13292
rect 28820 13252 28829 13292
rect 5443 13168 5452 13208
rect 5492 13168 6316 13208
rect 6356 13168 6365 13208
rect 7267 13168 7276 13208
rect 7316 13168 7564 13208
rect 7604 13168 7613 13208
rect 9763 13168 9772 13208
rect 9812 13168 12172 13208
rect 12212 13168 12980 13208
rect 12940 13124 12980 13168
rect 13036 13168 15148 13208
rect 15188 13168 15197 13208
rect 20332 13168 20428 13208
rect 20468 13168 20477 13208
rect 22627 13168 22636 13208
rect 22676 13168 23596 13208
rect 23636 13168 23645 13208
rect 13036 13124 13076 13168
rect 4675 13084 4684 13124
rect 4724 13084 5452 13124
rect 5492 13084 7084 13124
rect 7124 13084 11500 13124
rect 11540 13084 11596 13124
rect 11636 13084 11645 13124
rect 12940 13084 13076 13124
rect 13229 13084 13324 13124
rect 13364 13084 13373 13124
rect 13795 13084 13804 13124
rect 13844 13084 16300 13124
rect 16340 13084 16349 13124
rect 19747 13084 19756 13124
rect 19796 13084 19852 13124
rect 19892 13084 19901 13124
rect 20332 13040 20372 13168
rect 23971 13084 23980 13124
rect 24020 13084 24460 13124
rect 24500 13084 24509 13124
rect 11779 13000 11788 13040
rect 11828 13000 15628 13040
rect 15668 13000 16396 13040
rect 16436 13000 16445 13040
rect 19651 13000 19660 13040
rect 19700 13000 20372 13040
rect 22051 13000 22060 13040
rect 22100 13000 25036 13040
rect 25076 13000 25085 13040
rect 18787 12916 18796 12956
rect 18836 12916 21580 12956
rect 21620 12916 25420 12956
rect 25460 12916 25804 12956
rect 25844 12916 25853 12956
rect 4343 12832 4352 12872
rect 4720 12832 4729 12872
rect 12117 12832 12126 12872
rect 12494 12832 12503 12872
rect 13795 12832 13804 12872
rect 13844 12832 18124 12872
rect 18164 12832 18173 12872
rect 19891 12832 19900 12872
rect 20268 12832 20277 12872
rect 24451 12832 24460 12872
rect 24500 12832 25900 12872
rect 25940 12832 25949 12872
rect 27665 12832 27674 12872
rect 28042 12832 28051 12872
rect 4396 12748 8044 12788
rect 8084 12748 8093 12788
rect 22531 12748 22540 12788
rect 22580 12748 24364 12788
rect 24404 12748 24413 12788
rect 4396 12704 4436 12748
rect 4387 12664 4396 12704
rect 4436 12664 4445 12704
rect 13325 12664 13420 12704
rect 13460 12664 13469 12704
rect 15331 12664 15340 12704
rect 15380 12664 15628 12704
rect 15668 12664 15677 12704
rect 19277 12664 19372 12704
rect 19412 12664 19421 12704
rect 25507 12664 25516 12704
rect 25556 12664 26188 12704
rect 26228 12664 26237 12704
rect 4483 12580 4492 12620
rect 4532 12580 4876 12620
rect 4916 12580 7180 12620
rect 7220 12580 7229 12620
rect 8237 12580 8332 12620
rect 8372 12580 8381 12620
rect 8621 12580 8716 12620
rect 8756 12580 8765 12620
rect 8909 12580 9004 12620
rect 9044 12580 9053 12620
rect 10243 12580 10252 12620
rect 10292 12580 10828 12620
rect 10868 12580 12076 12620
rect 12116 12580 17836 12620
rect 17876 12580 17885 12620
rect 23491 12580 23500 12620
rect 23540 12580 27092 12620
rect 27052 12536 27092 12580
rect 4195 12496 4204 12536
rect 4244 12496 4300 12536
rect 4340 12496 7468 12536
rect 7508 12496 7517 12536
rect 19747 12496 19756 12536
rect 19796 12496 20812 12536
rect 20852 12496 20861 12536
rect 25411 12496 25420 12536
rect 25460 12496 25708 12536
rect 25748 12496 25757 12536
rect 27043 12496 27052 12536
rect 27092 12496 27820 12536
rect 27860 12496 27869 12536
rect 931 12412 940 12452
rect 980 12412 1708 12452
rect 1748 12412 5644 12452
rect 5684 12412 5693 12452
rect 6403 12412 6412 12452
rect 6452 12412 7084 12452
rect 7124 12412 7133 12452
rect 8525 12412 8620 12452
rect 8660 12412 8669 12452
rect 15139 12412 15148 12452
rect 15188 12412 15820 12452
rect 15860 12412 15869 12452
rect 18691 12412 18700 12452
rect 18740 12412 20428 12452
rect 20468 12412 20477 12452
rect 23107 12412 23116 12452
rect 23156 12412 23404 12452
rect 23444 12412 23453 12452
rect 24931 12412 24940 12452
rect 24980 12412 27244 12452
rect 27284 12412 27916 12452
rect 27956 12412 27965 12452
rect 5923 12328 5932 12368
rect 5972 12328 7276 12368
rect 7316 12328 7325 12368
rect 13795 12328 13804 12368
rect 13844 12328 16108 12368
rect 16148 12328 16157 12368
rect 23107 12328 23116 12368
rect 23156 12328 28204 12368
rect 28244 12328 28253 12368
rect 10627 12244 10636 12284
rect 10676 12244 19756 12284
rect 19796 12244 19805 12284
rect 24643 12244 24652 12284
rect 24692 12244 28108 12284
rect 28148 12244 28157 12284
rect 3103 12076 3112 12116
rect 3480 12076 3489 12116
rect 10877 12076 10886 12116
rect 11254 12076 11263 12116
rect 14947 12076 14956 12116
rect 14996 12076 16972 12116
rect 17012 12076 17021 12116
rect 18651 12076 18660 12116
rect 19028 12076 19037 12116
rect 26425 12076 26434 12116
rect 26802 12076 26811 12116
rect 10723 11992 10732 12032
rect 10772 11992 19276 12032
rect 19316 11992 19325 12032
rect 6787 11908 6796 11948
rect 6836 11908 10732 11948
rect 10772 11908 14804 11948
rect 14764 11864 14804 11908
rect 10051 11824 10060 11864
rect 10100 11824 10540 11864
rect 10580 11824 11980 11864
rect 12020 11824 12029 11864
rect 14755 11824 14764 11864
rect 14804 11824 14956 11864
rect 14996 11824 15005 11864
rect 25891 11824 25900 11864
rect 25940 11824 27628 11864
rect 27668 11824 27677 11864
rect 2371 11740 2380 11780
rect 2420 11740 6796 11780
rect 6836 11740 6845 11780
rect 15139 11740 15148 11780
rect 15188 11740 19660 11780
rect 19700 11740 19709 11780
rect 1891 11656 1900 11696
rect 1940 11656 4972 11696
rect 5012 11656 5021 11696
rect 5155 11656 5164 11696
rect 5204 11656 5548 11696
rect 5588 11656 5597 11696
rect 7075 11656 7084 11696
rect 7124 11656 8044 11696
rect 8084 11656 9004 11696
rect 9044 11656 9053 11696
rect 10051 11656 10060 11696
rect 10100 11656 12172 11696
rect 12212 11656 12221 11696
rect 18883 11656 18892 11696
rect 18932 11656 19276 11696
rect 19316 11656 19325 11696
rect 4343 11320 4352 11360
rect 4720 11320 4729 11360
rect 12117 11320 12126 11360
rect 12494 11320 12503 11360
rect 19891 11320 19900 11360
rect 20268 11320 20277 11360
rect 27665 11320 27674 11360
rect 28042 11320 28051 11360
rect 19277 11236 19372 11276
rect 19412 11236 19421 11276
rect 3331 11152 3340 11192
rect 3380 11152 4684 11192
rect 4724 11152 4733 11192
rect 3619 11068 3628 11108
rect 3668 11068 4108 11108
rect 4148 11068 4157 11108
rect 4579 11068 4588 11108
rect 4628 11068 5740 11108
rect 5780 11068 5789 11108
rect 12643 11068 12652 11108
rect 12692 11068 12940 11108
rect 12980 11068 12989 11108
rect 2371 10984 2380 11024
rect 2420 10984 4396 11024
rect 4436 10984 5068 11024
rect 5108 10984 5117 11024
rect 11395 10984 11404 11024
rect 11444 10984 12268 11024
rect 12308 10984 12317 11024
rect 19171 10816 19180 10856
rect 19220 10816 19660 10856
rect 19700 10816 19709 10856
rect 3811 10732 3820 10772
rect 3860 10732 6028 10772
rect 6068 10732 6077 10772
rect 3103 10564 3112 10604
rect 3480 10564 3489 10604
rect 5155 10564 5164 10604
rect 5204 10564 5548 10604
rect 5588 10564 5597 10604
rect 10157 10564 10252 10604
rect 10292 10564 10301 10604
rect 10877 10564 10886 10604
rect 11254 10564 11263 10604
rect 18651 10564 18660 10604
rect 19028 10564 19037 10604
rect 26425 10564 26434 10604
rect 26802 10564 26811 10604
rect 18499 10480 18508 10520
rect 18548 10480 21484 10520
rect 21524 10480 21533 10520
rect 10723 10396 10732 10436
rect 10772 10396 11020 10436
rect 11060 10396 11069 10436
rect 18307 10396 18316 10436
rect 18356 10396 20140 10436
rect 20180 10396 20189 10436
rect 2467 10312 2476 10352
rect 2516 10312 3628 10352
rect 3668 10312 3677 10352
rect 3724 10312 5548 10352
rect 5588 10312 5597 10352
rect 3724 10268 3764 10312
rect 1603 10228 1612 10268
rect 1652 10228 2092 10268
rect 2132 10228 2141 10268
rect 2947 10228 2956 10268
rect 2996 10228 3764 10268
rect 4195 10228 4204 10268
rect 4244 10228 4492 10268
rect 4532 10228 4541 10268
rect 15139 10228 15148 10268
rect 15188 10228 18220 10268
rect 18260 10228 18269 10268
rect 1219 10144 1228 10184
rect 1268 10144 3436 10184
rect 3476 10144 3820 10184
rect 3860 10144 3869 10184
rect 4003 10144 4012 10184
rect 4052 10144 4244 10184
rect 4387 10144 4396 10184
rect 4436 10144 4876 10184
rect 4916 10144 4925 10184
rect 15715 10144 15724 10184
rect 15764 10144 16972 10184
rect 17012 10144 17021 10184
rect 4204 10016 4244 10144
rect 2851 9976 2860 10016
rect 2900 9976 4244 10016
rect 4675 9976 4684 10016
rect 4724 9976 5068 10016
rect 5108 9976 5117 10016
rect 7555 9976 7564 10016
rect 7604 9976 8524 10016
rect 8564 9976 8573 10016
rect 5635 9892 5644 9932
rect 5684 9892 7756 9932
rect 7796 9892 7805 9932
rect 10051 9892 10060 9932
rect 10100 9892 19468 9932
rect 19508 9892 19517 9932
rect 20429 9892 20524 9932
rect 20564 9892 20573 9932
rect 4343 9808 4352 9848
rect 4720 9808 4729 9848
rect 12117 9808 12126 9848
rect 12494 9808 12503 9848
rect 19891 9808 19900 9848
rect 20268 9808 20277 9848
rect 27665 9808 27674 9848
rect 28042 9808 28051 9848
rect 835 9724 844 9764
rect 884 9724 5932 9764
rect 5972 9724 5981 9764
rect 3811 9472 3820 9512
rect 3860 9472 5836 9512
rect 5876 9472 7084 9512
rect 7124 9472 7133 9512
rect 11491 9472 11500 9512
rect 11540 9472 12460 9512
rect 12500 9472 13132 9512
rect 13172 9472 16204 9512
rect 16244 9472 16253 9512
rect 21859 9472 21868 9512
rect 21908 9472 24652 9512
rect 24692 9472 25996 9512
rect 26036 9472 26045 9512
rect 11980 9428 12020 9472
rect 11971 9388 11980 9428
rect 12020 9388 12060 9428
rect 24067 9388 24076 9428
rect 24116 9388 24556 9428
rect 24596 9388 24605 9428
rect 3103 9052 3112 9092
rect 3480 9052 3489 9092
rect 10877 9052 10886 9092
rect 11254 9052 11263 9092
rect 18651 9052 18660 9092
rect 19028 9052 19037 9092
rect 26425 9052 26434 9092
rect 26802 9052 26811 9092
rect 8131 8884 8140 8924
rect 8180 8884 9772 8924
rect 9812 8884 9821 8924
rect 4675 8800 4684 8840
rect 4724 8800 5644 8840
rect 5684 8800 5693 8840
rect 21571 8716 21580 8756
rect 21620 8716 23596 8756
rect 23636 8716 26572 8756
rect 26612 8716 26621 8756
rect 25891 8632 25900 8672
rect 25940 8632 27052 8672
rect 27092 8632 27101 8672
rect 4675 8464 4684 8504
rect 4724 8464 4916 8504
rect 4876 8420 4916 8464
rect 4867 8380 4876 8420
rect 4916 8380 4925 8420
rect 4343 8296 4352 8336
rect 4720 8296 4729 8336
rect 4973 8296 5068 8336
rect 5108 8296 5117 8336
rect 12117 8296 12126 8336
rect 12494 8296 12503 8336
rect 19891 8296 19900 8336
rect 20268 8296 20277 8336
rect 27665 8296 27674 8336
rect 28042 8296 28051 8336
rect 931 8128 940 8168
rect 980 8128 3820 8168
rect 3860 8128 3869 8168
rect 24547 8128 24556 8168
rect 24596 8128 26284 8168
rect 26324 8128 26333 8168
rect 451 8044 460 8084
rect 500 8044 1612 8084
rect 1652 8044 1661 8084
rect 4771 8044 4780 8084
rect 4820 8044 6316 8084
rect 6356 8044 6365 8084
rect 25603 8044 25612 8084
rect 25652 8044 26380 8084
rect 26420 8044 26429 8084
rect 1795 7960 1804 8000
rect 1844 7960 4204 8000
rect 4244 7960 4253 8000
rect 11491 7960 11500 8000
rect 11540 7960 11692 8000
rect 11732 7960 11741 8000
rect 15043 7960 15052 8000
rect 15092 7960 17740 8000
rect 17780 7960 17789 8000
rect 22627 7960 22636 8000
rect 22676 7960 24172 8000
rect 24212 7960 26860 8000
rect 26900 7960 26909 8000
rect 2083 7876 2092 7916
rect 2132 7876 4108 7916
rect 4148 7876 4684 7916
rect 4724 7876 4733 7916
rect 22339 7876 22348 7916
rect 22388 7876 26764 7916
rect 26804 7876 26813 7916
rect 3043 7708 3052 7748
rect 3092 7708 4108 7748
rect 4148 7708 4157 7748
rect 643 7624 652 7664
rect 692 7624 1516 7664
rect 1556 7624 1565 7664
rect 3103 7540 3112 7580
rect 3480 7540 3489 7580
rect 10877 7540 10886 7580
rect 11254 7540 11263 7580
rect 18651 7540 18660 7580
rect 19028 7540 19037 7580
rect 26425 7540 26434 7580
rect 26802 7540 26811 7580
rect 18115 7372 18124 7412
rect 18164 7372 18892 7412
rect 18932 7372 18941 7412
rect 259 7288 268 7328
rect 308 7288 1036 7328
rect 1076 7288 1085 7328
rect 13315 7204 13324 7244
rect 13364 7204 13708 7244
rect 13748 7204 15148 7244
rect 15188 7204 15197 7244
rect 18691 7204 18700 7244
rect 18740 7204 19372 7244
rect 19412 7204 19421 7244
rect 1891 7120 1900 7160
rect 1940 7120 3052 7160
rect 3092 7120 3101 7160
rect 18115 7120 18124 7160
rect 18164 7120 19180 7160
rect 19220 7120 19229 7160
rect 1219 7036 1228 7076
rect 1268 7036 2764 7076
rect 2804 7036 2813 7076
rect 739 6784 748 6824
rect 788 6784 1420 6824
rect 1460 6784 1469 6824
rect 4343 6784 4352 6824
rect 4720 6784 4729 6824
rect 12117 6784 12126 6824
rect 12494 6784 12503 6824
rect 19891 6784 19900 6824
rect 20268 6784 20277 6824
rect 27665 6784 27674 6824
rect 28042 6784 28051 6824
rect 2275 6616 2284 6656
rect 2324 6616 2380 6656
rect 2420 6616 2429 6656
rect 12451 6448 12460 6488
rect 12500 6448 13996 6488
rect 14036 6448 15628 6488
rect 15668 6448 15677 6488
rect 3103 6028 3112 6068
rect 3480 6028 3489 6068
rect 10877 6028 10886 6068
rect 11254 6028 11263 6068
rect 18651 6028 18660 6068
rect 19028 6028 19037 6068
rect 26425 6028 26434 6068
rect 26802 6028 26811 6068
rect 10243 5608 10252 5648
rect 10292 5608 13228 5648
rect 13268 5608 13804 5648
rect 13844 5608 13853 5648
rect 4343 5272 4352 5312
rect 4720 5272 4729 5312
rect 12117 5272 12126 5312
rect 12494 5272 12503 5312
rect 19891 5272 19900 5312
rect 20268 5272 20277 5312
rect 27665 5272 27674 5312
rect 28042 5272 28051 5312
rect 12931 5020 12940 5060
rect 12980 5020 13900 5060
rect 13940 5020 13949 5060
rect 3103 4516 3112 4556
rect 3480 4516 3489 4556
rect 10877 4516 10886 4556
rect 11254 4516 11263 4556
rect 18651 4516 18660 4556
rect 19028 4516 19037 4556
rect 26425 4516 26434 4556
rect 26802 4516 26811 4556
rect 4343 3760 4352 3800
rect 4720 3760 4729 3800
rect 12117 3760 12126 3800
rect 12494 3760 12503 3800
rect 19891 3760 19900 3800
rect 20268 3760 20277 3800
rect 27665 3760 27674 3800
rect 28042 3760 28051 3800
rect 3103 3004 3112 3044
rect 3480 3004 3489 3044
rect 10877 3004 10886 3044
rect 11254 3004 11263 3044
rect 18651 3004 18660 3044
rect 19028 3004 19037 3044
rect 26425 3004 26434 3044
rect 26802 3004 26811 3044
rect 4343 2248 4352 2288
rect 4720 2248 4729 2288
rect 12117 2248 12126 2288
rect 12494 2248 12503 2288
rect 19891 2248 19900 2288
rect 20268 2248 20277 2288
rect 27665 2248 27674 2288
rect 28042 2248 28051 2288
rect 3103 1492 3112 1532
rect 3480 1492 3489 1532
rect 10877 1492 10886 1532
rect 11254 1492 11263 1532
rect 18651 1492 18660 1532
rect 19028 1492 19037 1532
rect 26425 1492 26434 1532
rect 26802 1492 26811 1532
rect 4343 736 4352 776
rect 4720 736 4729 776
rect 12117 736 12126 776
rect 12494 736 12503 776
rect 19891 736 19900 776
rect 20268 736 20277 776
rect 27665 736 27674 776
rect 28042 736 28051 776
<< via4 >>
rect 4876 28120 4916 28160
rect 6700 28036 6740 28076
rect 4352 27952 4720 27992
rect 12126 27952 12494 27992
rect 19900 27952 20268 27992
rect 27674 27952 28042 27992
rect 6220 27868 6260 27908
rect 16972 27532 17012 27572
rect 27532 27532 27572 27572
rect 28780 27532 28820 27572
rect 29260 27532 29300 27572
rect 3916 27364 3956 27404
rect 7756 27364 7796 27404
rect 10252 27364 10292 27404
rect 3112 27196 3480 27236
rect 10886 27196 11254 27236
rect 18660 27196 19028 27236
rect 26434 27196 26802 27236
rect 18124 27028 18164 27068
rect 27244 26944 27284 26984
rect 20428 26776 20468 26816
rect 19564 26692 19604 26732
rect 4352 26440 4720 26480
rect 12126 26440 12494 26480
rect 19900 26440 20268 26480
rect 27674 26440 28042 26480
rect 6028 26188 6068 26228
rect 27532 26188 27572 26228
rect 15340 26104 15380 26144
rect 3628 26020 3668 26060
rect 29452 25936 29492 25976
rect 3112 25684 3480 25724
rect 10886 25684 11254 25724
rect 18660 25684 19028 25724
rect 26434 25684 26802 25724
rect 2956 25264 2996 25304
rect 8332 25264 8372 25304
rect 7276 25180 7316 25220
rect 21484 25180 21524 25220
rect 4352 24928 4720 24968
rect 12126 24928 12494 24968
rect 19900 24928 20268 24968
rect 27674 24928 28042 24968
rect 1708 24508 1748 24548
rect 29644 24508 29684 24548
rect 3112 24172 3480 24212
rect 10886 24172 11254 24212
rect 18660 24172 19028 24212
rect 26434 24172 26802 24212
rect 27244 24172 27284 24212
rect 10732 24088 10772 24128
rect 29260 24004 29300 24044
rect 2956 23836 2996 23876
rect 19756 23584 19796 23624
rect 29644 23500 29684 23540
rect 4352 23416 4720 23456
rect 12126 23416 12494 23456
rect 19900 23416 20268 23456
rect 27674 23416 28042 23456
rect 3820 23080 3860 23120
rect 9868 22996 9908 23036
rect 19564 22996 19604 23036
rect 19756 22996 19796 23036
rect 6028 22912 6068 22952
rect 3112 22660 3480 22700
rect 10886 22660 11254 22700
rect 18660 22660 19028 22700
rect 26434 22660 26802 22700
rect 9772 22492 9812 22532
rect 15340 22492 15380 22532
rect 8236 22408 8276 22448
rect 27244 22408 27284 22448
rect 1228 22324 1268 22364
rect 4204 22240 4244 22280
rect 28780 22240 28820 22280
rect 6604 22156 6644 22196
rect 4972 22072 5012 22112
rect 5260 22072 5300 22112
rect 4352 21904 4720 21944
rect 12126 21904 12494 21944
rect 19900 21904 20268 21944
rect 27674 21904 28042 21944
rect 4204 21820 4244 21860
rect 12652 21736 12692 21776
rect 20428 21736 20468 21776
rect 16972 21652 17012 21692
rect 2572 21400 2612 21440
rect 6700 21400 6740 21440
rect 2764 21232 2804 21272
rect 3820 21232 3860 21272
rect 8908 21232 8948 21272
rect 3112 21148 3480 21188
rect 4972 21148 5012 21188
rect 10886 21148 11254 21188
rect 18660 21148 19028 21188
rect 26434 21148 26802 21188
rect 1516 20896 1556 20936
rect 6604 20812 6644 20852
rect 29452 20812 29492 20852
rect 8524 20644 8564 20684
rect 10732 20728 10772 20768
rect 17932 20644 17972 20684
rect 8716 20560 8756 20600
rect 18124 20560 18164 20600
rect 17068 20476 17108 20516
rect 2572 20392 2612 20432
rect 4352 20392 4720 20432
rect 9868 20392 9908 20432
rect 12126 20392 12494 20432
rect 19900 20392 20268 20432
rect 27674 20392 28042 20432
rect 1900 20140 1940 20180
rect 4012 20140 4052 20180
rect 5068 20140 5108 20180
rect 5644 20140 5684 20180
rect 5836 20140 5876 20180
rect 7372 20140 7412 20180
rect 7564 20140 7604 20180
rect 10732 20140 10772 20180
rect 17932 20140 17972 20180
rect 19468 20140 19508 20180
rect 21484 20140 21524 20180
rect 12652 19972 12692 20012
rect 4204 19804 4244 19844
rect 5068 19804 5108 19844
rect 9772 19804 9812 19844
rect 3112 19636 3480 19676
rect 10886 19636 11254 19676
rect 18660 19636 19028 19676
rect 26434 19636 26802 19676
rect 10636 19468 10676 19508
rect 2476 19384 2516 19424
rect 2956 19300 2996 19340
rect 5356 19300 5396 19340
rect 7852 19300 7892 19340
rect 3820 19216 3860 19256
rect 7276 19216 7316 19256
rect 17068 19216 17108 19256
rect 1612 19132 1652 19172
rect 6220 19132 6260 19172
rect 4876 19048 4916 19088
rect 2668 18964 2708 19004
rect 16396 18964 16436 19004
rect 2572 18880 2612 18920
rect 4352 18880 4720 18920
rect 5836 18880 5876 18920
rect 8140 18880 8180 18920
rect 9388 18880 9428 18920
rect 12126 18880 12494 18920
rect 12652 18880 12692 18920
rect 19900 18880 20268 18920
rect 27674 18880 28042 18920
rect 8716 18796 8756 18836
rect 18412 18796 18452 18836
rect 2380 18712 2420 18752
rect 5164 18712 5204 18752
rect 5452 18712 5492 18752
rect 7372 18628 7412 18668
rect 7660 18628 7700 18668
rect 2956 18460 2996 18500
rect 6604 18460 6644 18500
rect 8428 18460 8468 18500
rect 2668 18376 2708 18416
rect 9196 18376 9236 18416
rect 5836 18292 5876 18332
rect 10540 18292 10580 18332
rect 11980 18292 12020 18332
rect 10444 18208 10484 18248
rect 3112 18124 3480 18164
rect 10886 18124 11254 18164
rect 18660 18124 19028 18164
rect 26434 18124 26802 18164
rect 7276 18040 7316 18080
rect 7564 18040 7604 18080
rect 9772 17956 9812 17996
rect 16876 17956 16916 17996
rect 1804 17872 1844 17912
rect 2572 17872 2612 17912
rect 3916 17872 3956 17912
rect 16780 17788 16820 17828
rect 18508 17788 18548 17828
rect 7660 17704 7700 17744
rect 9868 17704 9908 17744
rect 5068 17620 5108 17660
rect 7372 17620 7412 17660
rect 8044 17620 8084 17660
rect 8524 17536 8564 17576
rect 15436 17536 15476 17576
rect 9004 17452 9044 17492
rect 9388 17452 9428 17492
rect 4352 17368 4720 17408
rect 5260 17368 5300 17408
rect 11500 17368 11540 17408
rect 12126 17368 12494 17408
rect 19900 17368 20268 17408
rect 27674 17368 28042 17408
rect 9868 17284 9908 17324
rect 1228 17200 1268 17240
rect 8428 17116 8468 17156
rect 5068 17032 5108 17072
rect 23116 17032 23156 17072
rect 10444 16864 10484 16904
rect 2668 16780 2708 16820
rect 13420 16780 13460 16820
rect 19180 16780 19220 16820
rect 16012 16696 16052 16736
rect 3112 16612 3480 16652
rect 10886 16612 11254 16652
rect 18660 16612 19028 16652
rect 26434 16612 26802 16652
rect 10636 16528 10676 16568
rect 9196 16360 9236 16400
rect 12652 16360 12692 16400
rect 3820 16276 3860 16316
rect 8140 16276 8180 16316
rect 16396 16108 16436 16148
rect 1420 16024 1460 16064
rect 13324 16024 13364 16064
rect 20524 16024 20564 16064
rect 3628 15940 3668 15980
rect 16876 15940 16916 15980
rect 4352 15856 4720 15896
rect 5356 15856 5396 15896
rect 12126 15856 12494 15896
rect 19900 15856 20268 15896
rect 27674 15856 28042 15896
rect 6028 15772 6068 15812
rect 15436 15772 15476 15812
rect 1804 15688 1844 15728
rect 5068 15688 5108 15728
rect 18412 15520 18452 15560
rect 8236 15436 8276 15476
rect 7852 15352 7892 15392
rect 19468 15352 19508 15392
rect 2476 15184 2516 15224
rect 3112 15100 3480 15140
rect 5644 15100 5684 15140
rect 10732 15100 10772 15140
rect 10886 15100 11254 15140
rect 18660 15100 19028 15140
rect 26434 15100 26802 15140
rect 10444 14932 10484 14972
rect 1708 14848 1748 14888
rect 7756 14764 7796 14804
rect 10636 14764 10676 14804
rect 19276 14764 19316 14804
rect 19660 14512 19700 14552
rect 4204 14428 4244 14468
rect 4352 14344 4720 14384
rect 12126 14344 12494 14384
rect 19900 14344 20268 14384
rect 11980 14260 12020 14300
rect 19180 14176 19220 14216
rect 1900 14092 1940 14132
rect 6604 14092 6644 14132
rect 16012 14092 16052 14132
rect 8044 14008 8084 14048
rect 8716 14008 8756 14048
rect 10540 14008 10580 14048
rect 16780 14008 16820 14048
rect 18508 13924 18548 13964
rect 27674 14344 28042 14384
rect 7276 13840 7316 13880
rect 8524 13756 8564 13796
rect 10252 13756 10292 13796
rect 3112 13588 3480 13628
rect 10886 13588 11254 13628
rect 18660 13588 19028 13628
rect 26434 13588 26802 13628
rect 8620 13336 8660 13376
rect 8908 13336 8948 13376
rect 18412 13336 18452 13376
rect 7564 13168 7604 13208
rect 5452 13084 5492 13124
rect 11500 13084 11540 13124
rect 13324 13084 13364 13124
rect 19756 13084 19796 13124
rect 4352 12832 4720 12872
rect 12126 12832 12494 12872
rect 19900 12832 20268 12872
rect 27674 12832 28042 12872
rect 13420 12664 13460 12704
rect 19372 12664 19412 12704
rect 4876 12580 4916 12620
rect 8332 12580 8372 12620
rect 8716 12580 8756 12620
rect 9004 12580 9044 12620
rect 10252 12580 10292 12620
rect 4204 12496 4244 12536
rect 8620 12412 8660 12452
rect 23116 12412 23156 12452
rect 19756 12244 19796 12284
rect 3112 12076 3480 12116
rect 10886 12076 11254 12116
rect 18660 12076 19028 12116
rect 26434 12076 26802 12116
rect 19276 11992 19316 12032
rect 10732 11908 10772 11948
rect 4352 11320 4720 11360
rect 12126 11320 12494 11360
rect 19900 11320 20268 11360
rect 27674 11320 28042 11360
rect 19372 11236 19412 11276
rect 19660 10816 19700 10856
rect 3112 10564 3480 10604
rect 10252 10564 10292 10604
rect 10886 10564 11254 10604
rect 18660 10564 19028 10604
rect 26434 10564 26802 10604
rect 18508 10480 18548 10520
rect 10732 10396 10772 10436
rect 4204 10228 4244 10268
rect 4012 10144 4052 10184
rect 4876 10144 4916 10184
rect 5068 9976 5108 10016
rect 20524 9892 20564 9932
rect 4352 9808 4720 9848
rect 12126 9808 12494 9848
rect 19900 9808 20268 9848
rect 27674 9808 28042 9848
rect 3112 9052 3480 9092
rect 10886 9052 11254 9092
rect 18660 9052 19028 9092
rect 26434 9052 26802 9092
rect 4352 8296 4720 8336
rect 5068 8296 5108 8336
rect 12126 8296 12494 8336
rect 19900 8296 20268 8336
rect 27674 8296 28042 8336
rect 1612 8044 1652 8084
rect 1516 7624 1556 7664
rect 3112 7540 3480 7580
rect 10886 7540 11254 7580
rect 18660 7540 19028 7580
rect 26434 7540 26802 7580
rect 2764 7036 2804 7076
rect 1420 6784 1460 6824
rect 4352 6784 4720 6824
rect 12126 6784 12494 6824
rect 19900 6784 20268 6824
rect 27674 6784 28042 6824
rect 2380 6616 2420 6656
rect 3112 6028 3480 6068
rect 10886 6028 11254 6068
rect 18660 6028 19028 6068
rect 26434 6028 26802 6068
rect 4352 5272 4720 5312
rect 12126 5272 12494 5312
rect 19900 5272 20268 5312
rect 27674 5272 28042 5312
rect 3112 4516 3480 4556
rect 10886 4516 11254 4556
rect 18660 4516 19028 4556
rect 26434 4516 26802 4556
rect 4352 3760 4720 3800
rect 12126 3760 12494 3800
rect 19900 3760 20268 3800
rect 27674 3760 28042 3800
rect 3112 3004 3480 3044
rect 10886 3004 11254 3044
rect 18660 3004 19028 3044
rect 26434 3004 26802 3044
rect 4352 2248 4720 2288
rect 12126 2248 12494 2288
rect 19900 2248 20268 2288
rect 27674 2248 28042 2288
rect 3112 1492 3480 1532
rect 10886 1492 11254 1532
rect 18660 1492 19028 1532
rect 26434 1492 26802 1532
rect 4352 736 4720 776
rect 12126 736 12494 776
rect 19900 736 20268 776
rect 27674 736 28042 776
<< metal5 >>
rect 4876 28160 4916 28169
rect 3076 27236 3516 28016
rect 4316 27992 4756 28016
rect 4316 27952 4352 27992
rect 4720 27952 4756 27992
rect 3076 27196 3112 27236
rect 3480 27196 3516 27236
rect 3076 25724 3516 27196
rect 3916 27404 3956 27413
rect 3076 25684 3112 25724
rect 3480 25684 3516 25724
rect 2956 25304 2996 25313
rect 1708 24548 1748 24557
rect 1228 22364 1268 22373
rect 1228 17240 1268 22324
rect 1228 17191 1268 17200
rect 1516 20936 1556 20945
rect 1420 16064 1460 16073
rect 1420 6824 1460 16024
rect 1516 7664 1556 20896
rect 1612 19172 1652 19181
rect 1612 8084 1652 19132
rect 1708 14888 1748 24508
rect 2956 23876 2996 25264
rect 2956 23827 2996 23836
rect 3076 24212 3516 25684
rect 3076 24172 3112 24212
rect 3480 24172 3516 24212
rect 3076 22700 3516 24172
rect 3076 22660 3112 22700
rect 3480 22660 3516 22700
rect 2572 21440 2612 21449
rect 2572 20432 2612 21400
rect 1900 20180 1940 20189
rect 1804 17912 1844 17921
rect 1804 15728 1844 17872
rect 1804 15679 1844 15688
rect 1708 14839 1748 14848
rect 1900 14132 1940 20140
rect 2476 19424 2516 19433
rect 1900 14083 1940 14092
rect 2380 18752 2420 18761
rect 1612 8035 1652 8044
rect 1516 7615 1556 7624
rect 1420 6775 1460 6784
rect 2380 6656 2420 18712
rect 2476 15224 2516 19384
rect 2572 18920 2612 20392
rect 2764 21272 2804 21281
rect 2572 17912 2612 18880
rect 2572 17863 2612 17872
rect 2668 19004 2708 19013
rect 2668 18416 2708 18964
rect 2668 16820 2708 18376
rect 2668 16771 2708 16780
rect 2476 15175 2516 15184
rect 2764 7076 2804 21232
rect 3076 21188 3516 22660
rect 3076 21148 3112 21188
rect 3480 21148 3516 21188
rect 3076 19676 3516 21148
rect 3076 19636 3112 19676
rect 3480 19636 3516 19676
rect 2956 19340 2996 19349
rect 2956 18500 2996 19300
rect 2956 18451 2996 18460
rect 2764 7027 2804 7036
rect 3076 18164 3516 19636
rect 3076 18124 3112 18164
rect 3480 18124 3516 18164
rect 3076 16652 3516 18124
rect 3076 16612 3112 16652
rect 3480 16612 3516 16652
rect 3076 15140 3516 16612
rect 3628 26060 3668 26069
rect 3628 15980 3668 26020
rect 3820 23120 3860 23129
rect 3820 21272 3860 23080
rect 3820 21223 3860 21232
rect 3820 19256 3860 19265
rect 3820 16316 3860 19216
rect 3916 17912 3956 27364
rect 4316 26480 4756 27952
rect 4316 26440 4352 26480
rect 4720 26440 4756 26480
rect 4316 24968 4756 26440
rect 4316 24928 4352 24968
rect 4720 24928 4756 24968
rect 4316 23456 4756 24928
rect 4316 23416 4352 23456
rect 4720 23416 4756 23456
rect 4204 22280 4244 22289
rect 4204 21860 4244 22240
rect 4204 21811 4244 21820
rect 4316 21944 4756 23416
rect 4316 21904 4352 21944
rect 4720 21904 4756 21944
rect 4316 20432 4756 21904
rect 4316 20392 4352 20432
rect 4720 20392 4756 20432
rect 3916 17863 3956 17872
rect 4012 20180 4052 20189
rect 3820 16267 3860 16276
rect 3628 15931 3668 15940
rect 3076 15100 3112 15140
rect 3480 15100 3516 15140
rect 3076 13628 3516 15100
rect 3076 13588 3112 13628
rect 3480 13588 3516 13628
rect 3076 12116 3516 13588
rect 3076 12076 3112 12116
rect 3480 12076 3516 12116
rect 3076 10604 3516 12076
rect 3076 10564 3112 10604
rect 3480 10564 3516 10604
rect 3076 9092 3516 10564
rect 4012 10184 4052 20140
rect 4204 19844 4244 19853
rect 4204 14468 4244 19804
rect 4204 14419 4244 14428
rect 4316 18920 4756 20392
rect 4876 19088 4916 28120
rect 6700 28076 6740 28085
rect 6220 27908 6260 27917
rect 6028 26228 6068 26237
rect 6028 22952 6068 26188
rect 4972 22112 5012 22121
rect 4972 21188 5012 22072
rect 4972 21139 5012 21148
rect 5260 22112 5300 22121
rect 5068 20180 5108 20189
rect 5068 19844 5108 20140
rect 5068 19795 5108 19804
rect 4876 19039 4916 19048
rect 4316 18880 4352 18920
rect 4720 18880 4756 18920
rect 4316 17408 4756 18880
rect 5164 18752 5204 18761
rect 4316 17368 4352 17408
rect 4720 17368 4756 17408
rect 4316 15896 4756 17368
rect 4316 15856 4352 15896
rect 4720 15856 4756 15896
rect 4316 14384 4756 15856
rect 5068 18712 5164 18740
rect 5068 18700 5204 18712
rect 5068 17660 5108 18700
rect 5068 17072 5108 17620
rect 5260 17408 5300 22072
rect 5644 20180 5684 20189
rect 5260 17359 5300 17368
rect 5356 19340 5396 19349
rect 5068 15728 5108 17032
rect 5356 15896 5396 19300
rect 5356 15847 5396 15856
rect 5452 18752 5492 18761
rect 5068 15679 5108 15688
rect 4316 14344 4352 14384
rect 4720 14344 4756 14384
rect 4316 12872 4756 14344
rect 5452 13124 5492 18712
rect 5644 15140 5684 20140
rect 5836 20180 5876 20189
rect 5836 18920 5876 20140
rect 5836 18332 5876 18880
rect 5836 18283 5876 18292
rect 6028 15812 6068 22912
rect 6220 19172 6260 27868
rect 6604 22196 6644 22205
rect 6604 20852 6644 22156
rect 6700 21440 6740 28036
rect 7756 27404 7796 27413
rect 6700 21391 6740 21400
rect 7276 25220 7316 25229
rect 6604 20803 6644 20812
rect 7276 19256 7316 25180
rect 7276 19207 7316 19216
rect 7372 20180 7412 20189
rect 6220 19123 6260 19132
rect 7372 18668 7412 20140
rect 6028 15763 6068 15772
rect 6604 18500 6644 18509
rect 5644 15091 5684 15100
rect 6604 14132 6644 18460
rect 6604 14083 6644 14092
rect 7276 18080 7316 18089
rect 7276 13880 7316 18040
rect 7372 17660 7412 18628
rect 7372 17611 7412 17620
rect 7564 20180 7604 20189
rect 7564 18080 7604 20140
rect 7276 13831 7316 13840
rect 7564 13208 7604 18040
rect 7660 18668 7700 18677
rect 7660 17744 7700 18628
rect 7660 17695 7700 17704
rect 7756 14804 7796 27364
rect 10252 27404 10292 27413
rect 8332 25304 8372 25313
rect 8236 22448 8276 22457
rect 7852 19340 7892 19349
rect 7852 15392 7892 19300
rect 8140 18920 8180 18929
rect 7852 15343 7892 15352
rect 8044 17660 8084 17669
rect 7756 14755 7796 14764
rect 8044 14048 8084 17620
rect 8140 16316 8180 18880
rect 8140 16267 8180 16276
rect 8236 15476 8276 22408
rect 8236 15427 8276 15436
rect 8044 13999 8084 14008
rect 7564 13159 7604 13168
rect 5452 13075 5492 13084
rect 4316 12832 4352 12872
rect 4720 12832 4756 12872
rect 4204 12536 4244 12545
rect 4204 10268 4244 12496
rect 4204 10219 4244 10228
rect 4316 11360 4756 12832
rect 4316 11320 4352 11360
rect 4720 11320 4756 11360
rect 4012 10135 4052 10144
rect 3076 9052 3112 9092
rect 3480 9052 3516 9092
rect 3076 7580 3516 9052
rect 3076 7540 3112 7580
rect 3480 7540 3516 7580
rect 2380 6607 2420 6616
rect 3076 6068 3516 7540
rect 3076 6028 3112 6068
rect 3480 6028 3516 6068
rect 3076 4556 3516 6028
rect 3076 4516 3112 4556
rect 3480 4516 3516 4556
rect 3076 3044 3516 4516
rect 3076 3004 3112 3044
rect 3480 3004 3516 3044
rect 3076 1532 3516 3004
rect 3076 1492 3112 1532
rect 3480 1492 3516 1532
rect 3076 712 3516 1492
rect 4316 9848 4756 11320
rect 4876 12620 4916 12629
rect 4876 10184 4916 12580
rect 8332 12620 8372 25264
rect 9868 23036 9908 23045
rect 9772 22532 9812 22541
rect 8908 21272 8948 21281
rect 8524 20684 8564 20693
rect 8524 20180 8564 20644
rect 8716 20600 8756 20609
rect 8524 20140 8660 20180
rect 8428 18500 8468 18509
rect 8428 17156 8468 18460
rect 8428 17107 8468 17116
rect 8524 17576 8564 17585
rect 8524 13796 8564 17536
rect 8524 13747 8564 13756
rect 8620 13536 8660 20140
rect 8716 18836 8756 20560
rect 8716 14048 8756 18796
rect 8716 13999 8756 14008
rect 8620 13496 8756 13536
rect 8332 12571 8372 12580
rect 8620 13376 8660 13385
rect 8620 12452 8660 13336
rect 8716 12620 8756 13496
rect 8908 13376 8948 21232
rect 9772 19844 9812 22492
rect 9868 20432 9908 22996
rect 9868 20383 9908 20392
rect 9388 18920 9428 18929
rect 9196 18416 9236 18425
rect 8908 13327 8948 13336
rect 9004 17492 9044 17501
rect 8716 12571 8756 12580
rect 9004 12620 9044 17452
rect 9196 16400 9236 18376
rect 9388 17492 9428 18880
rect 9772 17996 9812 19804
rect 9772 17947 9812 17956
rect 9388 17443 9428 17452
rect 9868 17744 9908 17753
rect 9868 17324 9908 17704
rect 9868 17275 9908 17284
rect 9196 16351 9236 16360
rect 10252 13796 10292 27364
rect 10850 27236 11290 28016
rect 10850 27196 10886 27236
rect 11254 27196 11290 27236
rect 10850 25724 11290 27196
rect 10850 25684 10886 25724
rect 11254 25684 11290 25724
rect 10850 24212 11290 25684
rect 10850 24172 10886 24212
rect 11254 24172 11290 24212
rect 10732 24128 10772 24137
rect 10732 20768 10772 24088
rect 10636 20728 10732 20768
rect 10636 19508 10676 20728
rect 10732 20719 10772 20728
rect 10850 22700 11290 24172
rect 10850 22660 10886 22700
rect 11254 22660 11290 22700
rect 10850 21188 11290 22660
rect 10850 21148 10886 21188
rect 11254 21148 11290 21188
rect 10636 19459 10676 19468
rect 10732 20180 10772 20189
rect 10540 18332 10580 18341
rect 10444 18248 10484 18257
rect 10444 16904 10484 18208
rect 10444 14972 10484 16864
rect 10444 14923 10484 14932
rect 10540 14048 10580 18292
rect 10636 16568 10676 16577
rect 10636 14804 10676 16528
rect 10732 15140 10772 20140
rect 10732 15091 10772 15100
rect 10850 19676 11290 21148
rect 10850 19636 10886 19676
rect 11254 19636 11290 19676
rect 10850 18164 11290 19636
rect 12090 27992 12530 28016
rect 12090 27952 12126 27992
rect 12494 27952 12530 27992
rect 12090 26480 12530 27952
rect 12090 26440 12126 26480
rect 12494 26440 12530 26480
rect 12090 24968 12530 26440
rect 16972 27572 17012 27581
rect 12090 24928 12126 24968
rect 12494 24928 12530 24968
rect 12090 23456 12530 24928
rect 12090 23416 12126 23456
rect 12494 23416 12530 23456
rect 12090 21944 12530 23416
rect 15340 26144 15380 26153
rect 15340 22532 15380 26104
rect 15340 22483 15380 22492
rect 12090 21904 12126 21944
rect 12494 21904 12530 21944
rect 12090 20432 12530 21904
rect 12090 20392 12126 20432
rect 12494 20392 12530 20432
rect 12090 18920 12530 20392
rect 12090 18880 12126 18920
rect 12494 18880 12530 18920
rect 10850 18124 10886 18164
rect 11254 18124 11290 18164
rect 10850 16652 11290 18124
rect 11980 18332 12020 18341
rect 10850 16612 10886 16652
rect 11254 16612 11290 16652
rect 10850 15140 11290 16612
rect 10850 15100 10886 15140
rect 11254 15100 11290 15140
rect 10636 14755 10676 14764
rect 10540 13999 10580 14008
rect 10252 13747 10292 13756
rect 10850 13628 11290 15100
rect 10850 13588 10886 13628
rect 11254 13588 11290 13628
rect 9004 12571 9044 12580
rect 10252 12620 10292 12629
rect 8620 12403 8660 12412
rect 10252 10604 10292 12580
rect 10850 12116 11290 13588
rect 11500 17408 11540 17417
rect 11500 13124 11540 17368
rect 11980 14300 12020 18292
rect 11980 14251 12020 14260
rect 12090 17408 12530 18880
rect 12090 17368 12126 17408
rect 12494 17368 12530 17408
rect 12090 15896 12530 17368
rect 12652 21776 12692 21785
rect 12652 20012 12692 21736
rect 16972 21692 17012 27532
rect 18624 27236 19064 28016
rect 18624 27196 18660 27236
rect 19028 27196 19064 27236
rect 16972 21643 17012 21652
rect 18124 27068 18164 27077
rect 17932 20684 17972 20693
rect 12652 18920 12692 19972
rect 17068 20516 17108 20525
rect 17068 19256 17108 20476
rect 17932 20180 17972 20644
rect 18124 20600 18164 27028
rect 18124 20551 18164 20560
rect 18624 25724 19064 27196
rect 19864 27992 20304 28016
rect 19864 27952 19900 27992
rect 20268 27952 20304 27992
rect 18624 25684 18660 25724
rect 19028 25684 19064 25724
rect 18624 24212 19064 25684
rect 18624 24172 18660 24212
rect 19028 24172 19064 24212
rect 18624 22700 19064 24172
rect 19564 26732 19604 26741
rect 19564 23036 19604 26692
rect 19864 26480 20304 27952
rect 26398 27236 26838 28016
rect 27638 27992 28078 28016
rect 27638 27952 27674 27992
rect 28042 27952 28078 27992
rect 26398 27196 26434 27236
rect 26802 27196 26838 27236
rect 19864 26440 19900 26480
rect 20268 26440 20304 26480
rect 19864 24968 20304 26440
rect 19864 24928 19900 24968
rect 20268 24928 20304 24968
rect 19564 22987 19604 22996
rect 19756 23624 19796 23633
rect 19756 23036 19796 23584
rect 19756 22987 19796 22996
rect 19864 23456 20304 24928
rect 19864 23416 19900 23456
rect 20268 23416 20304 23456
rect 18624 22660 18660 22700
rect 19028 22660 19064 22700
rect 18624 21188 19064 22660
rect 18624 21148 18660 21188
rect 19028 21148 19064 21188
rect 17932 20131 17972 20140
rect 17068 19207 17108 19216
rect 18624 19676 19064 21148
rect 19864 21944 20304 23416
rect 19864 21904 19900 21944
rect 20268 21904 20304 21944
rect 19864 20432 20304 21904
rect 20428 26816 20468 26825
rect 20428 21776 20468 26776
rect 26398 25724 26838 27196
rect 27532 27572 27572 27581
rect 26398 25684 26434 25724
rect 26802 25684 26838 25724
rect 20428 21727 20468 21736
rect 21484 25220 21524 25229
rect 19864 20392 19900 20432
rect 20268 20392 20304 20432
rect 18624 19636 18660 19676
rect 19028 19636 19064 19676
rect 12652 16400 12692 18880
rect 16396 19004 16436 19013
rect 15436 17576 15476 17585
rect 12652 16351 12692 16360
rect 13420 16820 13460 16829
rect 12090 15856 12126 15896
rect 12494 15856 12530 15896
rect 12090 14384 12530 15856
rect 12090 14344 12126 14384
rect 12494 14344 12530 14384
rect 11500 13075 11540 13084
rect 10850 12076 10886 12116
rect 11254 12076 11290 12116
rect 10252 10555 10292 10564
rect 10732 11948 10772 11957
rect 10732 10436 10772 11908
rect 10732 10387 10772 10396
rect 10850 10604 11290 12076
rect 10850 10564 10886 10604
rect 11254 10564 11290 10604
rect 4876 10135 4916 10144
rect 4316 9808 4352 9848
rect 4720 9808 4756 9848
rect 4316 8336 4756 9808
rect 4316 8296 4352 8336
rect 4720 8296 4756 8336
rect 4316 6824 4756 8296
rect 5068 10016 5108 10025
rect 5068 8336 5108 9976
rect 5068 8287 5108 8296
rect 10850 9092 11290 10564
rect 10850 9052 10886 9092
rect 11254 9052 11290 9092
rect 4316 6784 4352 6824
rect 4720 6784 4756 6824
rect 4316 5312 4756 6784
rect 4316 5272 4352 5312
rect 4720 5272 4756 5312
rect 4316 3800 4756 5272
rect 4316 3760 4352 3800
rect 4720 3760 4756 3800
rect 4316 2288 4756 3760
rect 4316 2248 4352 2288
rect 4720 2248 4756 2288
rect 4316 776 4756 2248
rect 4316 736 4352 776
rect 4720 736 4756 776
rect 4316 712 4756 736
rect 10850 7580 11290 9052
rect 10850 7540 10886 7580
rect 11254 7540 11290 7580
rect 10850 6068 11290 7540
rect 10850 6028 10886 6068
rect 11254 6028 11290 6068
rect 10850 4556 11290 6028
rect 10850 4516 10886 4556
rect 11254 4516 11290 4556
rect 10850 3044 11290 4516
rect 10850 3004 10886 3044
rect 11254 3004 11290 3044
rect 10850 1532 11290 3004
rect 10850 1492 10886 1532
rect 11254 1492 11290 1532
rect 10850 712 11290 1492
rect 12090 12872 12530 14344
rect 13324 16064 13364 16073
rect 13324 13124 13364 16024
rect 13324 13075 13364 13084
rect 12090 12832 12126 12872
rect 12494 12832 12530 12872
rect 12090 11360 12530 12832
rect 13420 12704 13460 16780
rect 15436 15812 15476 17536
rect 15436 15763 15476 15772
rect 16012 16736 16052 16745
rect 16012 14132 16052 16696
rect 16396 16148 16436 18964
rect 18412 18836 18452 18845
rect 16876 17996 16916 18005
rect 16396 16099 16436 16108
rect 16780 17828 16820 17837
rect 16012 14083 16052 14092
rect 16780 14048 16820 17788
rect 16876 15980 16916 17956
rect 16876 15931 16916 15940
rect 16780 13999 16820 14008
rect 18412 15560 18452 18796
rect 18624 18164 19064 19636
rect 18624 18124 18660 18164
rect 19028 18124 19064 18164
rect 18412 13376 18452 15520
rect 18412 13327 18452 13336
rect 18508 17828 18548 17837
rect 18508 13964 18548 17788
rect 13420 12655 13460 12664
rect 12090 11320 12126 11360
rect 12494 11320 12530 11360
rect 12090 9848 12530 11320
rect 18508 10520 18548 13924
rect 18508 10471 18548 10480
rect 18624 16652 19064 18124
rect 19468 20180 19508 20189
rect 18624 16612 18660 16652
rect 19028 16612 19064 16652
rect 18624 15140 19064 16612
rect 18624 15100 18660 15140
rect 19028 15100 19064 15140
rect 18624 13628 19064 15100
rect 19180 16820 19220 16829
rect 19180 14216 19220 16780
rect 19468 15392 19508 20140
rect 19468 15343 19508 15352
rect 19864 18920 20304 20392
rect 21484 20180 21524 25180
rect 21484 20131 21524 20140
rect 26398 24212 26838 25684
rect 26398 24172 26434 24212
rect 26802 24172 26838 24212
rect 26398 22700 26838 24172
rect 26398 22660 26434 22700
rect 26802 22660 26838 22700
rect 26398 21188 26838 22660
rect 27244 26984 27284 26993
rect 27244 24212 27284 26944
rect 27532 26228 27572 27532
rect 27532 26179 27572 26188
rect 27638 26480 28078 27952
rect 27638 26440 27674 26480
rect 28042 26440 28078 26480
rect 27244 22448 27284 24172
rect 27244 22399 27284 22408
rect 27638 24968 28078 26440
rect 27638 24928 27674 24968
rect 28042 24928 28078 24968
rect 27638 23456 28078 24928
rect 27638 23416 27674 23456
rect 28042 23416 28078 23456
rect 26398 21148 26434 21188
rect 26802 21148 26838 21188
rect 19864 18880 19900 18920
rect 20268 18880 20304 18920
rect 19864 17408 20304 18880
rect 19864 17368 19900 17408
rect 20268 17368 20304 17408
rect 19864 15896 20304 17368
rect 26398 19676 26838 21148
rect 26398 19636 26434 19676
rect 26802 19636 26838 19676
rect 26398 18164 26838 19636
rect 26398 18124 26434 18164
rect 26802 18124 26838 18164
rect 23116 17072 23156 17081
rect 19864 15856 19900 15896
rect 20268 15856 20304 15896
rect 19180 14167 19220 14176
rect 19276 14804 19316 14813
rect 18624 13588 18660 13628
rect 19028 13588 19064 13628
rect 18624 12116 19064 13588
rect 18624 12076 18660 12116
rect 19028 12076 19064 12116
rect 18624 10604 19064 12076
rect 19276 12032 19316 14764
rect 19660 14552 19700 14561
rect 19276 11983 19316 11992
rect 19372 12704 19412 12713
rect 19372 11276 19412 12664
rect 19372 11227 19412 11236
rect 19660 10856 19700 14512
rect 19864 14384 20304 15856
rect 19864 14344 19900 14384
rect 20268 14344 20304 14384
rect 19756 13124 19796 13133
rect 19756 12284 19796 13084
rect 19756 12235 19796 12244
rect 19864 12872 20304 14344
rect 19864 12832 19900 12872
rect 20268 12832 20304 12872
rect 19660 10807 19700 10816
rect 19864 11360 20304 12832
rect 19864 11320 19900 11360
rect 20268 11320 20304 11360
rect 18624 10564 18660 10604
rect 19028 10564 19064 10604
rect 12090 9808 12126 9848
rect 12494 9808 12530 9848
rect 12090 8336 12530 9808
rect 12090 8296 12126 8336
rect 12494 8296 12530 8336
rect 12090 6824 12530 8296
rect 12090 6784 12126 6824
rect 12494 6784 12530 6824
rect 12090 5312 12530 6784
rect 12090 5272 12126 5312
rect 12494 5272 12530 5312
rect 12090 3800 12530 5272
rect 12090 3760 12126 3800
rect 12494 3760 12530 3800
rect 12090 2288 12530 3760
rect 12090 2248 12126 2288
rect 12494 2248 12530 2288
rect 12090 776 12530 2248
rect 12090 736 12126 776
rect 12494 736 12530 776
rect 12090 712 12530 736
rect 18624 9092 19064 10564
rect 18624 9052 18660 9092
rect 19028 9052 19064 9092
rect 18624 7580 19064 9052
rect 18624 7540 18660 7580
rect 19028 7540 19064 7580
rect 18624 6068 19064 7540
rect 18624 6028 18660 6068
rect 19028 6028 19064 6068
rect 18624 4556 19064 6028
rect 18624 4516 18660 4556
rect 19028 4516 19064 4556
rect 18624 3044 19064 4516
rect 18624 3004 18660 3044
rect 19028 3004 19064 3044
rect 18624 1532 19064 3004
rect 18624 1492 18660 1532
rect 19028 1492 19064 1532
rect 18624 712 19064 1492
rect 19864 9848 20304 11320
rect 20524 16064 20564 16073
rect 20524 9932 20564 16024
rect 23116 12452 23156 17032
rect 23116 12403 23156 12412
rect 26398 16652 26838 18124
rect 26398 16612 26434 16652
rect 26802 16612 26838 16652
rect 26398 15140 26838 16612
rect 26398 15100 26434 15140
rect 26802 15100 26838 15140
rect 26398 13628 26838 15100
rect 26398 13588 26434 13628
rect 26802 13588 26838 13628
rect 20524 9883 20564 9892
rect 26398 12116 26838 13588
rect 26398 12076 26434 12116
rect 26802 12076 26838 12116
rect 26398 10604 26838 12076
rect 26398 10564 26434 10604
rect 26802 10564 26838 10604
rect 19864 9808 19900 9848
rect 20268 9808 20304 9848
rect 19864 8336 20304 9808
rect 19864 8296 19900 8336
rect 20268 8296 20304 8336
rect 19864 6824 20304 8296
rect 19864 6784 19900 6824
rect 20268 6784 20304 6824
rect 19864 5312 20304 6784
rect 19864 5272 19900 5312
rect 20268 5272 20304 5312
rect 19864 3800 20304 5272
rect 19864 3760 19900 3800
rect 20268 3760 20304 3800
rect 19864 2288 20304 3760
rect 19864 2248 19900 2288
rect 20268 2248 20304 2288
rect 19864 776 20304 2248
rect 19864 736 19900 776
rect 20268 736 20304 776
rect 19864 712 20304 736
rect 26398 9092 26838 10564
rect 26398 9052 26434 9092
rect 26802 9052 26838 9092
rect 26398 7580 26838 9052
rect 26398 7540 26434 7580
rect 26802 7540 26838 7580
rect 26398 6068 26838 7540
rect 26398 6028 26434 6068
rect 26802 6028 26838 6068
rect 26398 4556 26838 6028
rect 26398 4516 26434 4556
rect 26802 4516 26838 4556
rect 26398 3044 26838 4516
rect 26398 3004 26434 3044
rect 26802 3004 26838 3044
rect 26398 1532 26838 3004
rect 26398 1492 26434 1532
rect 26802 1492 26838 1532
rect 26398 712 26838 1492
rect 27638 21944 28078 23416
rect 28780 27572 28820 27581
rect 28780 22280 28820 27532
rect 29260 27572 29300 27581
rect 29260 24044 29300 27532
rect 29260 23995 29300 24004
rect 29452 25976 29492 25985
rect 28780 22231 28820 22240
rect 27638 21904 27674 21944
rect 28042 21904 28078 21944
rect 27638 20432 28078 21904
rect 29452 20852 29492 25936
rect 29644 24548 29684 24557
rect 29644 23540 29684 24508
rect 29644 23491 29684 23500
rect 29452 20803 29492 20812
rect 27638 20392 27674 20432
rect 28042 20392 28078 20432
rect 27638 18920 28078 20392
rect 27638 18880 27674 18920
rect 28042 18880 28078 18920
rect 27638 17408 28078 18880
rect 27638 17368 27674 17408
rect 28042 17368 28078 17408
rect 27638 15896 28078 17368
rect 27638 15856 27674 15896
rect 28042 15856 28078 15896
rect 27638 14384 28078 15856
rect 27638 14344 27674 14384
rect 28042 14344 28078 14384
rect 27638 12872 28078 14344
rect 27638 12832 27674 12872
rect 28042 12832 28078 12872
rect 27638 11360 28078 12832
rect 27638 11320 27674 11360
rect 28042 11320 28078 11360
rect 27638 9848 28078 11320
rect 27638 9808 27674 9848
rect 28042 9808 28078 9848
rect 27638 8336 28078 9808
rect 27638 8296 27674 8336
rect 28042 8296 28078 8336
rect 27638 6824 28078 8296
rect 27638 6784 27674 6824
rect 28042 6784 28078 6824
rect 27638 5312 28078 6784
rect 27638 5272 27674 5312
rect 28042 5272 28078 5312
rect 27638 3800 28078 5272
rect 27638 3760 27674 3800
rect 28042 3760 28078 3800
rect 27638 2288 28078 3760
rect 27638 2248 27674 2288
rect 28042 2248 28078 2288
rect 27638 776 28078 2248
rect 27638 736 27674 776
rect 28042 736 28078 776
rect 27638 712 28078 736
use sg13g2_inv_2  _1056_
timestamp 1747056038
transform -1 0 5088 0 -1 24948
box -48 -56 432 834
use sg13g2_inv_1  _1057_
timestamp 1747056038
transform -1 0 20928 0 1 3780
box -48 -56 336 834
use sg13g2_inv_1  _1058_
timestamp 1747056038
transform -1 0 21120 0 -1 5292
box -48 -56 336 834
use sg13g2_inv_1  _1059_
timestamp 1747056038
transform 1 0 8928 0 -1 12852
box -48 -56 336 834
use sg13g2_inv_1  _1060_
timestamp 1747056038
transform -1 0 29184 0 -1 18900
box -48 -56 336 834
use sg13g2_inv_1  _1061_
timestamp 1747056038
transform -1 0 20736 0 1 20412
box -48 -56 336 834
use sg13g2_inv_2  _1062_
timestamp 1747056038
transform 1 0 20928 0 1 18900
box -48 -56 432 834
use sg13g2_inv_2  _1063_
timestamp 1747056038
transform 1 0 19680 0 -1 12852
box -48 -56 432 834
use sg13g2_inv_2  _1064_
timestamp 1747056038
transform -1 0 19584 0 1 11340
box -48 -56 432 834
use sg13g2_inv_1  _1065_
timestamp 1747056038
transform 1 0 19488 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _1066_
timestamp 1747056038
transform -1 0 18528 0 1 14364
box -48 -56 336 834
use sg13g2_inv_1  _1067_
timestamp 1747056038
transform 1 0 22560 0 1 14364
box -48 -56 336 834
use sg13g2_inv_1  _1068_
timestamp 1747056038
transform -1 0 24288 0 1 12852
box -48 -56 336 834
use sg13g2_inv_1  _1069_
timestamp 1747056038
transform 1 0 20256 0 1 17388
box -48 -56 336 834
use sg13g2_inv_2  _1070_
timestamp 1747056038
transform -1 0 7008 0 -1 23436
box -48 -56 432 834
use sg13g2_inv_1  _1071_
timestamp 1747056038
transform -1 0 8160 0 -1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1072_
timestamp 1747056038
transform -1 0 17568 0 -1 20412
box -48 -56 336 834
use sg13g2_inv_1  _1073_
timestamp 1747056038
transform 1 0 15648 0 -1 26460
box -48 -56 336 834
use sg13g2_inv_1  _1074_
timestamp 1747056038
transform 1 0 12480 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _1075_
timestamp 1747056038
transform 1 0 22368 0 -1 24948
box -48 -56 336 834
use sg13g2_inv_1  _1076_
timestamp 1747056038
transform 1 0 2112 0 1 24948
box -48 -56 336 834
use sg13g2_inv_1  _1077_
timestamp 1747056038
transform -1 0 8928 0 -1 6804
box -48 -56 336 834
use sg13g2_inv_2  _1078_
timestamp 1747056038
transform -1 0 10656 0 -1 5292
box -48 -56 432 834
use sg13g2_o21ai_1  _1079_
timestamp 1747056038
transform -1 0 20736 0 -1 15876
box -48 -56 538 834
use sg13g2_nand3_1  _1080_
timestamp 1747056038
transform -1 0 24192 0 -1 15876
box -48 -56 528 834
use sg13g2_nor2_1  _1081_
timestamp 1747056038
transform 1 0 21504 0 1 12852
box -48 -56 432 834
use sg13g2_a21oi_1  _1082_
timestamp 1747056038
transform -1 0 22944 0 -1 15876
box -48 -56 528 834
use sg13g2_a21oi_1  _1083_
timestamp 1747056038
transform -1 0 20640 0 1 14364
box -48 -56 528 834
use sg13g2_nor2_1  _1084_
timestamp 1747056038
transform -1 0 20160 0 1 12852
box -48 -56 432 834
use sg13g2_nand2b_1  _1085_
timestamp 1747056038
transform -1 0 21600 0 1 14364
box -48 -56 528 834
use sg13g2_nor3_1  _1086_
timestamp 1747056038
transform 1 0 20256 0 -1 14364
box -48 -56 528 834
use sg13g2_nor2_1  _1087_
timestamp 1747056038
transform -1 0 19776 0 1 12852
box -48 -56 432 834
use sg13g2_nand3_1  _1088_
timestamp 1747056038
transform 1 0 20640 0 1 14364
box -48 -56 528 834
use sg13g2_a21oi_1  _1089_
timestamp 1747056038
transform -1 0 21216 0 -1 15876
box -48 -56 528 834
use sg13g2_a22oi_1  _1090_
timestamp 1747056038
transform 1 0 19680 0 -1 15876
box -48 -56 624 834
use sg13g2_inv_1  _1091_
timestamp 1747056038
transform 1 0 15168 0 1 21924
box -48 -56 336 834
use sg13g2_and2_2  _1092_
timestamp 1747056038
transform -1 0 19872 0 -1 27972
box -48 -56 624 834
use sg13g2_nand2_1  _1093_
timestamp 1747056038
transform -1 0 11136 0 1 24948
box -48 -56 432 834
use sg13g2_nor2_1  _1094_
timestamp 1747056038
transform 1 0 4992 0 -1 27972
box -48 -56 432 834
use sg13g2_or2_1  _1095_
timestamp 1747056038
transform -1 0 18624 0 -1 24948
box -48 -56 528 834
use sg13g2_nor2_1  _1096_
timestamp 1747056038
transform -1 0 28608 0 -1 26460
box -48 -56 432 834
use sg13g2_a21o_1  _1097_
timestamp 1747056038
transform -1 0 16608 0 -1 26460
box -48 -56 720 834
use sg13g2_nand2_1  _1098_
timestamp 1747056038
transform -1 0 29952 0 1 24948
box -48 -56 432 834
use sg13g2_nand3_1  _1099_
timestamp 1747056038
transform 1 0 18336 0 -1 26460
box -48 -56 528 834
use sg13g2_nor3_2  _1100_
timestamp 1747056038
transform 1 0 17856 0 1 24948
box -48 -56 912 834
use sg13g2_inv_1  _1101_
timestamp 1747056038
transform -1 0 15840 0 1 26460
box -48 -56 336 834
use sg13g2_nor2_1  _1102_
timestamp 1747056038
transform 1 0 2304 0 -1 27972
box -48 -56 432 834
use sg13g2_and2_1  _1103_
timestamp 1747056038
transform 1 0 16704 0 1 26460
box -48 -56 528 834
use sg13g2_nor2b_1  _1104_
timestamp 1747056038
transform -1 0 25344 0 1 24948
box -54 -56 528 834
use sg13g2_a221oi_1  _1105_
timestamp 1747056038
transform -1 0 18144 0 -1 26460
box -48 -56 816 834
use sg13g2_a21oi_2  _1106_
timestamp 1747056038
transform 1 0 16608 0 -1 26460
box -48 -56 816 834
use sg13g2_and2_1  _1107_
timestamp 1747056038
transform 1 0 18720 0 -1 21924
box -48 -56 528 834
use sg13g2_nand2_1  _1108_
timestamp 1747056038
transform -1 0 20736 0 1 26460
box -48 -56 432 834
use sg13g2_nor2_1  _1109_
timestamp 1747056038
transform -1 0 30048 0 1 20412
box -48 -56 432 834
use sg13g2_a21oi_1  _1110_
timestamp 1747056038
transform -1 0 25344 0 1 20412
box -48 -56 528 834
use sg13g2_nand2_1  _1111_
timestamp 1747056038
transform 1 0 2688 0 -1 27972
box -48 -56 432 834
use sg13g2_nor2_1  _1112_
timestamp 1747056038
transform 1 0 17376 0 -1 23436
box -48 -56 432 834
use sg13g2_a21oi_2  _1113_
timestamp 1747056038
transform 1 0 16896 0 1 21924
box -48 -56 816 834
use sg13g2_o21ai_1  _1114_
timestamp 1747056038
transform -1 0 17376 0 -1 23436
box -48 -56 538 834
use sg13g2_nor2_1  _1115_
timestamp 1747056038
transform 1 0 27744 0 -1 18900
box -48 -56 432 834
use sg13g2_a21oi_1  _1116_
timestamp 1747056038
transform -1 0 24672 0 1 20412
box -48 -56 528 834
use sg13g2_nor2_1  _1117_
timestamp 1747056038
transform 1 0 30144 0 1 21924
box -48 -56 432 834
use sg13g2_or2_1  _1118_
timestamp 1747056038
transform 1 0 24960 0 -1 21924
box -48 -56 528 834
use sg13g2_inv_1  _1119_
timestamp 1747056038
transform -1 0 30528 0 -1 20412
box -48 -56 336 834
use sg13g2_nor2_1  _1120_
timestamp 1747056038
transform -1 0 30144 0 -1 24948
box -48 -56 432 834
use sg13g2_nor2_1  _1121_
timestamp 1747056038
transform -1 0 30816 0 1 23436
box -48 -56 432 834
use sg13g2_a21oi_1  _1122_
timestamp 1747056038
transform 1 0 29664 0 1 21924
box -48 -56 528 834
use sg13g2_nor2_1  _1123_
timestamp 1747056038
transform 1 0 30048 0 1 23436
box -48 -56 432 834
use sg13g2_xnor2_1  _1124_
timestamp 1747056038
transform 1 0 12384 0 -1 27972
box -48 -56 816 834
use sg13g2_nor2_2  _1125_
timestamp 1747056038
transform -1 0 9408 0 1 23436
box -48 -56 624 834
use sg13g2_and2_1  _1126_
timestamp 1747056038
transform -1 0 10080 0 1 21924
box -48 -56 528 834
use sg13g2_nand2_1  _1127_
timestamp 1747056038
transform 1 0 6144 0 1 20412
box -48 -56 432 834
use sg13g2_nand2_1  _1128_
timestamp 1747056038
transform 1 0 2496 0 1 26460
box -48 -56 432 834
use sg13g2_o21ai_1  _1129_
timestamp 1747056038
transform 1 0 16416 0 1 21924
box -48 -56 538 834
use sg13g2_and2_2  _1130_
timestamp 1747056038
transform -1 0 18240 0 1 21924
box -48 -56 624 834
use sg13g2_o21ai_1  _1131_
timestamp 1747056038
transform 1 0 7392 0 -1 23436
box -48 -56 538 834
use sg13g2_nand3b_1  _1132_
timestamp 1747056038
transform -1 0 24576 0 1 14364
box -48 -56 720 834
use sg13g2_nor2_2  _1133_
timestamp 1747056038
transform -1 0 23712 0 -1 15876
box -48 -56 624 834
use sg13g2_nor2_1  _1134_
timestamp 1747056038
transform -1 0 1920 0 -1 27972
box -48 -56 432 834
use sg13g2_xnor2_1  _1135_
timestamp 1747056038
transform -1 0 22176 0 1 20412
box -48 -56 816 834
use sg13g2_nand2_1  _1136_
timestamp 1747056038
transform 1 0 27936 0 1 18900
box -48 -56 432 834
use sg13g2_xnor2_1  _1137_
timestamp 1747056038
transform -1 0 23520 0 -1 20412
box -48 -56 816 834
use sg13g2_inv_1  _1138_
timestamp 1747056038
transform -1 0 22944 0 1 18900
box -48 -56 336 834
use sg13g2_nand2_1  _1139_
timestamp 1747056038
transform 1 0 2880 0 1 26460
box -48 -56 432 834
use sg13g2_nand2_1  _1140_
timestamp 1747056038
transform 1 0 8160 0 -1 12852
box -48 -56 432 834
use sg13g2_xnor2_1  _1141_
timestamp 1747056038
transform -1 0 9696 0 1 24948
box -48 -56 816 834
use sg13g2_o21ai_1  _1142_
timestamp 1747056038
transform 1 0 9696 0 1 24948
box -48 -56 538 834
use sg13g2_and2_1  _1143_
timestamp 1747056038
transform 1 0 12096 0 -1 26460
box -48 -56 528 834
use sg13g2_xor2_1  _1144_
timestamp 1747056038
transform -1 0 11904 0 1 24948
box -48 -56 816 834
use sg13g2_nand2_1  _1145_
timestamp 1747056038
transform 1 0 4224 0 -1 27972
box -48 -56 432 834
use sg13g2_a21oi_1  _1146_
timestamp 1747056038
transform -1 0 15168 0 1 24948
box -48 -56 528 834
use sg13g2_a22oi_1  _1147_
timestamp 1747056038
transform 1 0 15360 0 1 23436
box -48 -56 624 834
use sg13g2_and2_1  _1148_
timestamp 1747056038
transform -1 0 21216 0 1 23436
box -48 -56 528 834
use sg13g2_or2_1  _1149_
timestamp 1747056038
transform -1 0 20736 0 1 23436
box -48 -56 528 834
use sg13g2_xnor2_1  _1150_
timestamp 1747056038
transform 1 0 18720 0 1 23436
box -48 -56 816 834
use sg13g2_nand2_1  _1151_
timestamp 1747056038
transform 1 0 29664 0 1 23436
box -48 -56 432 834
use sg13g2_xnor2_1  _1152_
timestamp 1747056038
transform -1 0 22464 0 1 23436
box -48 -56 816 834
use sg13g2_nor2_1  _1153_
timestamp 1747056038
transform -1 0 26016 0 -1 24948
box -48 -56 432 834
use sg13g2_inv_1  _1154_
timestamp 1747056038
transform -1 0 16992 0 1 23436
box -48 -56 336 834
use sg13g2_a221oi_1  _1155_
timestamp 1747056038
transform -1 0 16224 0 -1 23436
box -48 -56 816 834
use sg13g2_o21ai_1  _1156_
timestamp 1747056038
transform -1 0 21696 0 1 23436
box -48 -56 538 834
use sg13g2_nand2_1  _1157_
timestamp 1747056038
transform 1 0 28992 0 -1 24948
box -48 -56 432 834
use sg13g2_nor2_1  _1158_
timestamp 1747056038
transform 1 0 23520 0 -1 21924
box -48 -56 432 834
use sg13g2_o21ai_1  _1159_
timestamp 1747056038
transform -1 0 22656 0 1 20412
box -48 -56 538 834
use sg13g2_a21oi_2  _1160_
timestamp 1747056038
transform -1 0 22752 0 -1 20412
box -48 -56 816 834
use sg13g2_a21o_1  _1161_
timestamp 1747056038
transform 1 0 20736 0 1 20412
box -48 -56 720 834
use sg13g2_a21oi_1  _1162_
timestamp 1747056038
transform 1 0 19968 0 1 20412
box -48 -56 528 834
use sg13g2_and3_1  _1163_
timestamp 1747056038
transform -1 0 20160 0 -1 20412
box -48 -56 720 834
use sg13g2_nor3_1  _1164_
timestamp 1747056038
transform 1 0 19008 0 -1 20412
box -48 -56 528 834
use sg13g2_xor2_1  _1165_
timestamp 1747056038
transform -1 0 20928 0 -1 20412
box -48 -56 816 834
use sg13g2_nor2_1  _1166_
timestamp 1747056038
transform -1 0 19392 0 1 14364
box -48 -56 432 834
use sg13g2_o21ai_1  _1167_
timestamp 1747056038
transform 1 0 18720 0 -1 15876
box -48 -56 538 834
use sg13g2_o21ai_1  _1168_
timestamp 1747056038
transform 1 0 19200 0 -1 15876
box -48 -56 538 834
use sg13g2_xor2_1  _1169_
timestamp 1747056038
transform -1 0 14016 0 -1 24948
box -48 -56 816 834
use sg13g2_a21oi_1  _1170_
timestamp 1747056038
transform -1 0 12096 0 -1 26460
box -48 -56 528 834
use sg13g2_xnor2_1  _1171_
timestamp 1747056038
transform 1 0 11904 0 1 24948
box -48 -56 816 834
use sg13g2_nor2_1  _1172_
timestamp 1747056038
transform -1 0 19392 0 1 12852
box -48 -56 432 834
use sg13g2_xnor2_1  _1173_
timestamp 1747056038
transform -1 0 11712 0 1 23436
box -48 -56 816 834
use sg13g2_inv_1  _1174_
timestamp 1747056038
transform 1 0 7104 0 -1 11340
box -48 -56 336 834
use sg13g2_nor2b_1  _1175_
timestamp 1747056038
transform -1 0 20640 0 1 12852
box -54 -56 528 834
use sg13g2_xor2_1  _1176_
timestamp 1747056038
transform 1 0 7296 0 1 24948
box -48 -56 816 834
use sg13g2_xor2_1  _1177_
timestamp 1747056038
transform 1 0 7584 0 -1 24948
box -48 -56 816 834
use sg13g2_xnor2_1  _1178_
timestamp 1747056038
transform -1 0 8832 0 -1 26460
box -48 -56 816 834
use sg13g2_and2_1  _1179_
timestamp 1747056038
transform 1 0 20544 0 -1 12852
box -48 -56 528 834
use sg13g2_nand2_1  _1180_
timestamp 1747056038
transform -1 0 21408 0 -1 12852
box -48 -56 432 834
use sg13g2_mux4_1  _1181_
timestamp 1747056038
transform 1 0 7200 0 1 12852
box -48 -56 2064 834
use sg13g2_nand3_1  _1182_
timestamp 1747056038
transform 1 0 23712 0 1 11340
box -48 -56 528 834
use sg13g2_inv_1  _1183_
timestamp 1747056038
transform 1 0 21888 0 1 12852
box -48 -56 336 834
use sg13g2_nand3b_1  _1184_
timestamp 1747056038
transform 1 0 17568 0 1 12852
box -48 -56 720 834
use sg13g2_and3_2  _1185_
timestamp 1747056038
transform 1 0 21312 0 -1 20412
box -48 -56 720 834
use sg13g2_nor2_2  _1186_
timestamp 1747056038
transform -1 0 23136 0 -1 11340
box -48 -56 624 834
use sg13g2_nor2b_1  _1187_
timestamp 1747056038
transform -1 0 20256 0 -1 14364
box -54 -56 528 834
use sg13g2_xnor2_1  _1188_
timestamp 1747056038
transform 1 0 21504 0 1 18900
box -48 -56 816 834
use sg13g2_inv_1  _1189_
timestamp 1747056038
transform -1 0 18048 0 1 8316
box -48 -56 336 834
use sg13g2_a21oi_1  _1190_
timestamp 1747056038
transform -1 0 20064 0 -1 23436
box -48 -56 528 834
use sg13g2_xnor2_1  _1191_
timestamp 1747056038
transform -1 0 20256 0 1 23436
box -48 -56 816 834
use sg13g2_xnor2_1  _1192_
timestamp 1747056038
transform 1 0 17952 0 1 23436
box -48 -56 816 834
use sg13g2_a22oi_1  _1193_
timestamp 1747056038
transform -1 0 18816 0 -1 14364
box -48 -56 624 834
use sg13g2_o21ai_1  _1194_
timestamp 1747056038
transform -1 0 19296 0 -1 14364
box -48 -56 538 834
use sg13g2_o21ai_1  _1195_
timestamp 1747056038
transform -1 0 19776 0 -1 14364
box -48 -56 538 834
use sg13g2_nand3_1  _1196_
timestamp 1747056038
transform -1 0 19008 0 1 14364
box -48 -56 528 834
use sg13g2_o21ai_1  _1197_
timestamp 1747056038
transform -1 0 7392 0 -1 21924
box -48 -56 538 834
use sg13g2_mux4_1  _1198_
timestamp 1747056038
transform 1 0 18240 0 1 17388
box -48 -56 2064 834
use sg13g2_nor2b_1  _1199_
timestamp 1747056038
transform 1 0 9888 0 1 17388
box -54 -56 528 834
use sg13g2_nand2_2  _1200_
timestamp 1747056038
transform 1 0 7680 0 -1 17388
box -48 -56 624 834
use sg13g2_nor2_2  _1201_
timestamp 1747056038
transform 1 0 9504 0 -1 17388
box -48 -56 624 834
use sg13g2_or2_2  _1202_
timestamp 1747056038
transform 1 0 9600 0 1 18900
box -48 -56 624 834
use sg13g2_nor2_1  _1203_
timestamp 1747056038
transform 1 0 5760 0 1 20412
box -48 -56 432 834
use sg13g2_a221oi_1  _1204_
timestamp 1747056038
transform 1 0 7680 0 1 18900
box -48 -56 816 834
use sg13g2_nor2b_2  _1205_
timestamp 1747056038
transform 1 0 9408 0 1 23436
box -54 -56 720 834
use sg13g2_and2_1  _1206_
timestamp 1747056038
transform 1 0 10656 0 1 18900
box -48 -56 528 834
use sg13g2_nand2_2  _1207_
timestamp 1747056038
transform 1 0 11616 0 -1 18900
box -48 -56 624 834
use sg13g2_nor2_1  _1208_
timestamp 1747056038
transform -1 0 22656 0 1 18900
box -48 -56 432 834
use sg13g2_mux2_2  _1209_
timestamp 1747056038
transform -1 0 19488 0 1 18900
box -48 -56 1104 834
use sg13g2_and2_2  _1210_
timestamp 1747056038
transform 1 0 13344 0 1 18900
box -48 -56 624 834
use sg13g2_nand2_2  _1211_
timestamp 1747056038
transform -1 0 15648 0 -1 18900
box -48 -56 624 834
use sg13g2_nand2_1  _1212_
timestamp 1747056038
transform -1 0 8256 0 -1 20412
box -48 -56 432 834
use sg13g2_nor2_1  _1213_
timestamp 1747056038
transform 1 0 16512 0 1 17388
box -48 -56 432 834
use sg13g2_nand2b_2  _1214_
timestamp 1747056038
transform -1 0 14016 0 -1 18900
box -48 -56 816 834
use sg13g2_o21ai_1  _1215_
timestamp 1747056038
transform 1 0 8256 0 -1 20412
box -48 -56 538 834
use sg13g2_inv_1  _1216_
timestamp 1747056038
transform -1 0 9408 0 -1 20412
box -48 -56 336 834
use sg13g2_nor2b_2  _1217_
timestamp 1747056038
transform 1 0 10080 0 1 23436
box -54 -56 720 834
use sg13g2_and2_1  _1218_
timestamp 1747056038
transform 1 0 10848 0 1 20412
box -48 -56 528 834
use sg13g2_nand2_1  _1219_
timestamp 1747056038
transform -1 0 15648 0 -1 26460
box -48 -56 432 834
use sg13g2_xnor2_1  _1220_
timestamp 1747056038
transform -1 0 8736 0 1 23436
box -48 -56 816 834
use sg13g2_nand2b_1  _1221_
timestamp 1747056038
transform -1 0 7872 0 1 20412
box -48 -56 528 834
use sg13g2_and2_2  _1222_
timestamp 1747056038
transform 1 0 9984 0 1 20412
box -48 -56 624 834
use sg13g2_nand2_1  _1223_
timestamp 1747056038
transform 1 0 7008 0 -1 23436
box -48 -56 432 834
use sg13g2_a21oi_1  _1224_
timestamp 1747056038
transform -1 0 9120 0 1 20412
box -48 -56 528 834
use sg13g2_a221oi_1  _1225_
timestamp 1747056038
transform 1 0 7872 0 1 20412
box -48 -56 816 834
use sg13g2_a21oi_1  _1226_
timestamp 1747056038
transform 1 0 7392 0 -1 21924
box -48 -56 528 834
use sg13g2_o21ai_1  _1227_
timestamp 1747056038
transform 1 0 6816 0 1 21924
box -48 -56 538 834
use sg13g2_a21oi_2  _1228_
timestamp 1747056038
transform 1 0 7296 0 1 21924
box -48 -56 816 834
use sg13g2_o21ai_1  _1229_
timestamp 1747056038
transform 1 0 4320 0 -1 21924
box -48 -56 538 834
use sg13g2_nor2_1  _1230_
timestamp 1747056038
transform -1 0 1152 0 -1 27972
box -48 -56 432 834
use sg13g2_o21ai_1  _1231_
timestamp 1747056038
transform 1 0 5760 0 -1 21924
box -48 -56 538 834
use sg13g2_nand2_1  _1232_
timestamp 1747056038
transform -1 0 3072 0 -1 11340
box -48 -56 432 834
use sg13g2_nor2_1  _1233_
timestamp 1747056038
transform 1 0 672 0 1 9828
box -48 -56 432 834
use sg13g2_xor2_1  _1234_
timestamp 1747056038
transform 1 0 2496 0 1 21924
box -48 -56 816 834
use sg13g2_xnor2_1  _1235_
timestamp 1747056038
transform 1 0 3264 0 1 21924
box -48 -56 816 834
use sg13g2_nand2_1  _1236_
timestamp 1747056038
transform -1 0 12864 0 1 17388
box -48 -56 432 834
use sg13g2_nand2_1  _1237_
timestamp 1747056038
transform -1 0 8928 0 -1 12852
box -48 -56 432 834
use sg13g2_xnor2_1  _1238_
timestamp 1747056038
transform 1 0 3264 0 -1 21924
box -48 -56 816 834
use sg13g2_xnor2_1  _1239_
timestamp 1747056038
transform 1 0 3840 0 1 20412
box -48 -56 816 834
use sg13g2_xnor2_1  _1240_
timestamp 1747056038
transform 1 0 4128 0 1 14364
box -48 -56 816 834
use sg13g2_xnor2_1  _1241_
timestamp 1747056038
transform -1 0 8736 0 -1 14364
box -48 -56 816 834
use sg13g2_and2_1  _1242_
timestamp 1747056038
transform -1 0 12864 0 1 18900
box -48 -56 528 834
use sg13g2_nand2_1  _1243_
timestamp 1747056038
transform -1 0 10176 0 -1 18900
box -48 -56 432 834
use sg13g2_a21oi_1  _1244_
timestamp 1747056038
transform -1 0 6624 0 -1 15876
box -48 -56 528 834
use sg13g2_o21ai_1  _1245_
timestamp 1747056038
transform 1 0 5472 0 -1 14364
box -48 -56 538 834
use sg13g2_nor2b_2  _1246_
timestamp 1747056038
transform -1 0 10848 0 -1 18900
box -54 -56 720 834
use sg13g2_nand2b_2  _1247_
timestamp 1747056038
transform -1 0 11616 0 -1 18900
box -48 -56 816 834
use sg13g2_a21o_1  _1248_
timestamp 1747056038
transform 1 0 8736 0 -1 14364
box -48 -56 720 834
use sg13g2_nor2_1  _1249_
timestamp 1747056038
transform -1 0 8352 0 -1 15876
box -48 -56 432 834
use sg13g2_mux2_1  _1250_
timestamp 1747056038
transform 1 0 20736 0 1 15876
box -48 -56 1008 834
use sg13g2_mux2_1  _1251_
timestamp 1747056038
transform 1 0 20448 0 -1 17388
box -48 -56 1008 834
use sg13g2_mux2_2  _1252_
timestamp 1747056038
transform -1 0 22080 0 1 17388
box -48 -56 1104 834
use sg13g2_a221oi_1  _1253_
timestamp 1747056038
transform -1 0 7968 0 1 17388
box -48 -56 816 834
use sg13g2_inv_1  _1254_
timestamp 1747056038
transform -1 0 5472 0 -1 18900
box -48 -56 336 834
use sg13g2_a22oi_1  _1255_
timestamp 1747056038
transform 1 0 4800 0 1 17388
box -48 -56 624 834
use sg13g2_o21ai_1  _1256_
timestamp 1747056038
transform 1 0 4512 0 -1 20412
box -48 -56 538 834
use sg13g2_nor2_2  _1257_
timestamp 1747056038
transform 1 0 9024 0 1 18900
box -48 -56 624 834
use sg13g2_nand2_2  _1258_
timestamp 1747056038
transform 1 0 5088 0 1 18900
box -48 -56 624 834
use sg13g2_a221oi_1  _1259_
timestamp 1747056038
transform -1 0 5760 0 -1 20412
box -48 -56 816 834
use sg13g2_nor2_1  _1260_
timestamp 1747056038
transform 1 0 960 0 1 26460
box -48 -56 432 834
use sg13g2_o21ai_1  _1261_
timestamp 1747056038
transform -1 0 6240 0 1 21924
box -48 -56 538 834
use sg13g2_a21oi_2  _1262_
timestamp 1747056038
transform -1 0 6048 0 -1 23436
box -48 -56 816 834
use sg13g2_o21ai_1  _1263_
timestamp 1747056038
transform -1 0 2592 0 1 18900
box -48 -56 538 834
use sg13g2_nor2_1  _1264_
timestamp 1747056038
transform -1 0 3744 0 -1 17388
box -48 -56 432 834
use sg13g2_o21ai_1  _1265_
timestamp 1747056038
transform -1 0 3072 0 1 18900
box -48 -56 538 834
use sg13g2_mux4_1  _1266_
timestamp 1747056038
transform -1 0 20256 0 -1 17388
box -48 -56 2064 834
use sg13g2_inv_1  _1267_
timestamp 1747056038
transform -1 0 12288 0 -1 15876
box -48 -56 336 834
use sg13g2_nor2_1  _1268_
timestamp 1747056038
transform 1 0 7584 0 -1 15876
box -48 -56 432 834
use sg13g2_a221oi_1  _1269_
timestamp 1747056038
transform -1 0 7872 0 1 15876
box -48 -56 816 834
use sg13g2_and2_1  _1270_
timestamp 1747056038
transform -1 0 4128 0 -1 15876
box -48 -56 528 834
use sg13g2_o21ai_1  _1271_
timestamp 1747056038
transform -1 0 3840 0 1 20412
box -48 -56 538 834
use sg13g2_and2_1  _1272_
timestamp 1747056038
transform 1 0 768 0 -1 12852
box -48 -56 528 834
use sg13g2_xor2_1  _1273_
timestamp 1747056038
transform 1 0 1248 0 -1 12852
box -48 -56 816 834
use sg13g2_xnor2_1  _1274_
timestamp 1747056038
transform 1 0 2016 0 1 12852
box -48 -56 816 834
use sg13g2_o21ai_1  _1275_
timestamp 1747056038
transform 1 0 2688 0 -1 12852
box -48 -56 538 834
use sg13g2_nor2b_1  _1276_
timestamp 1747056038
transform 1 0 2880 0 1 12852
box -54 -56 528 834
use sg13g2_xnor2_1  _1277_
timestamp 1747056038
transform 1 0 2400 0 -1 14364
box -48 -56 816 834
use sg13g2_xor2_1  _1278_
timestamp 1747056038
transform 1 0 3168 0 -1 14364
box -48 -56 816 834
use sg13g2_xnor2_1  _1279_
timestamp 1747056038
transform 1 0 5376 0 -1 12852
box -48 -56 816 834
use sg13g2_o21ai_1  _1280_
timestamp 1747056038
transform 1 0 6144 0 1 12852
box -48 -56 538 834
use sg13g2_nand2_1  _1281_
timestamp 1747056038
transform 1 0 864 0 -1 9828
box -48 -56 432 834
use sg13g2_nand2_1  _1282_
timestamp 1747056038
transform 1 0 960 0 -1 8316
box -48 -56 432 834
use sg13g2_xnor2_1  _1283_
timestamp 1747056038
transform 1 0 960 0 -1 11340
box -48 -56 816 834
use sg13g2_xnor2_1  _1284_
timestamp 1747056038
transform 1 0 1248 0 1 11340
box -48 -56 816 834
use sg13g2_nand2_1  _1285_
timestamp 1747056038
transform 1 0 576 0 -1 8316
box -48 -56 432 834
use sg13g2_xnor2_1  _1286_
timestamp 1747056038
transform 1 0 2592 0 1 9828
box -48 -56 816 834
use sg13g2_nand2_1  _1287_
timestamp 1747056038
transform -1 0 3744 0 1 9828
box -48 -56 432 834
use sg13g2_xor2_1  _1288_
timestamp 1747056038
transform -1 0 3840 0 -1 11340
box -48 -56 816 834
use sg13g2_a21oi_1  _1289_
timestamp 1747056038
transform -1 0 3456 0 1 11340
box -48 -56 528 834
use sg13g2_o21ai_1  _1290_
timestamp 1747056038
transform 1 0 3456 0 1 11340
box -48 -56 538 834
use sg13g2_a221oi_1  _1291_
timestamp 1747056038
transform -1 0 4704 0 -1 14364
box -48 -56 816 834
use sg13g2_o21ai_1  _1292_
timestamp 1747056038
transform 1 0 4128 0 -1 15876
box -48 -56 538 834
use sg13g2_o21ai_1  _1293_
timestamp 1747056038
transform -1 0 4896 0 1 15876
box -48 -56 538 834
use sg13g2_a21oi_1  _1294_
timestamp 1747056038
transform 1 0 3072 0 1 18900
box -48 -56 528 834
use sg13g2_o21ai_1  _1295_
timestamp 1747056038
transform 1 0 864 0 1 18900
box -48 -56 538 834
use sg13g2_a21oi_2  _1296_
timestamp 1747056038
transform 1 0 1344 0 1 18900
box -48 -56 816 834
use sg13g2_o21ai_1  _1297_
timestamp 1747056038
transform -1 0 2880 0 -1 21924
box -48 -56 538 834
use sg13g2_nor2_1  _1298_
timestamp 1747056038
transform -1 0 1344 0 1 6804
box -48 -56 432 834
use sg13g2_nand2_1  _1299_
timestamp 1747056038
transform 1 0 9600 0 1 20412
box -48 -56 432 834
use sg13g2_o21ai_1  _1300_
timestamp 1747056038
transform -1 0 1248 0 1 20412
box -48 -56 538 834
use sg13g2_nand2_1  _1301_
timestamp 1747056038
transform -1 0 23808 0 1 18900
box -48 -56 432 834
use sg13g2_o21ai_1  _1302_
timestamp 1747056038
transform 1 0 22080 0 1 17388
box -48 -56 538 834
use sg13g2_mux2_2  _1303_
timestamp 1747056038
transform -1 0 22560 0 -1 17388
box -48 -56 1104 834
use sg13g2_a22oi_1  _1304_
timestamp 1747056038
transform -1 0 8928 0 -1 17388
box -48 -56 624 834
use sg13g2_o21ai_1  _1305_
timestamp 1747056038
transform -1 0 8736 0 -1 18900
box -48 -56 538 834
use sg13g2_a21oi_1  _1306_
timestamp 1747056038
transform -1 0 3936 0 1 12852
box -48 -56 528 834
use sg13g2_xor2_1  _1307_
timestamp 1747056038
transform 1 0 8928 0 1 11340
box -48 -56 816 834
use sg13g2_nand2b_1  _1308_
timestamp 1747056038
transform 1 0 8736 0 -1 11340
box -48 -56 528 834
use sg13g2_xnor2_1  _1309_
timestamp 1747056038
transform -1 0 8928 0 1 11340
box -48 -56 816 834
use sg13g2_a21o_1  _1310_
timestamp 1747056038
transform -1 0 2688 0 -1 12852
box -48 -56 720 834
use sg13g2_nand2_1  _1311_
timestamp 1747056038
transform 1 0 7104 0 -1 12852
box -48 -56 432 834
use sg13g2_nor2_1  _1312_
timestamp 1747056038
transform 1 0 4224 0 1 9828
box -48 -56 432 834
use sg13g2_xnor2_1  _1313_
timestamp 1747056038
transform 1 0 3936 0 -1 12852
box -48 -56 816 834
use sg13g2_xnor2_1  _1314_
timestamp 1747056038
transform 1 0 4224 0 1 12852
box -48 -56 816 834
use sg13g2_xnor2_1  _1315_
timestamp 1747056038
transform -1 0 7488 0 1 14364
box -48 -56 816 834
use sg13g2_o21ai_1  _1316_
timestamp 1747056038
transform 1 0 6240 0 1 14364
box -48 -56 538 834
use sg13g2_o21ai_1  _1317_
timestamp 1747056038
transform 1 0 3840 0 -1 11340
box -48 -56 538 834
use sg13g2_xnor2_1  _1318_
timestamp 1747056038
transform 1 0 6048 0 1 9828
box -48 -56 816 834
use sg13g2_xor2_1  _1319_
timestamp 1747056038
transform -1 0 7104 0 -1 11340
box -48 -56 816 834
use sg13g2_nor2_1  _1320_
timestamp 1747056038
transform -1 0 8160 0 -1 12852
box -48 -56 432 834
use sg13g2_xor2_1  _1321_
timestamp 1747056038
transform -1 0 8160 0 1 11340
box -48 -56 816 834
use sg13g2_o21ai_1  _1322_
timestamp 1747056038
transform 1 0 2016 0 1 11340
box -48 -56 538 834
use sg13g2_xnor2_1  _1323_
timestamp 1747056038
transform -1 0 7392 0 1 11340
box -48 -56 816 834
use sg13g2_a21oi_1  _1324_
timestamp 1747056038
transform 1 0 6624 0 -1 12852
box -48 -56 528 834
use sg13g2_o21ai_1  _1325_
timestamp 1747056038
transform -1 0 6624 0 1 11340
box -48 -56 538 834
use sg13g2_a21oi_1  _1326_
timestamp 1747056038
transform -1 0 7104 0 1 12852
box -48 -56 528 834
use sg13g2_o21ai_1  _1327_
timestamp 1747056038
transform 1 0 5184 0 1 12852
box -48 -56 538 834
use sg13g2_o21ai_1  _1328_
timestamp 1747056038
transform -1 0 5376 0 1 15876
box -48 -56 538 834
use sg13g2_a22oi_1  _1329_
timestamp 1747056038
transform -1 0 6240 0 -1 17388
box -48 -56 624 834
use sg13g2_nor2_1  _1330_
timestamp 1747056038
transform 1 0 3072 0 -1 27972
box -48 -56 432 834
use sg13g2_nor2_1  _1331_
timestamp 1747056038
transform 1 0 1440 0 -1 6804
box -48 -56 432 834
use sg13g2_o21ai_1  _1332_
timestamp 1747056038
transform 1 0 1152 0 -1 21924
box -48 -56 538 834
use sg13g2_a21oi_2  _1333_
timestamp 1747056038
transform 1 0 1248 0 1 20412
box -48 -56 816 834
use sg13g2_o21ai_1  _1334_
timestamp 1747056038
transform -1 0 3264 0 1 17388
box -48 -56 538 834
use sg13g2_nor2_1  _1335_
timestamp 1747056038
transform -1 0 2304 0 1 17388
box -48 -56 432 834
use sg13g2_o21ai_1  _1336_
timestamp 1747056038
transform -1 0 2592 0 -1 18900
box -48 -56 538 834
use sg13g2_mux4_1  _1337_
timestamp 1747056038
transform -1 0 25728 0 -1 17388
box -48 -56 2064 834
use sg13g2_a22oi_1  _1338_
timestamp 1747056038
transform 1 0 11520 0 1 15876
box -48 -56 624 834
use sg13g2_o21ai_1  _1339_
timestamp 1747056038
transform -1 0 10464 0 1 15876
box -48 -56 538 834
use sg13g2_o21ai_1  _1340_
timestamp 1747056038
transform 1 0 4704 0 -1 12852
box -48 -56 538 834
use sg13g2_nand2_1  _1341_
timestamp 1747056038
transform 1 0 10848 0 1 8316
box -48 -56 432 834
use sg13g2_nor2_1  _1342_
timestamp 1747056038
transform 1 0 9696 0 1 11340
box -48 -56 432 834
use sg13g2_xor2_1  _1343_
timestamp 1747056038
transform -1 0 12480 0 1 11340
box -48 -56 816 834
use sg13g2_xnor2_1  _1344_
timestamp 1747056038
transform -1 0 11712 0 1 11340
box -48 -56 816 834
use sg13g2_o21ai_1  _1345_
timestamp 1747056038
transform 1 0 9216 0 -1 11340
box -48 -56 538 834
use sg13g2_and2_1  _1346_
timestamp 1747056038
transform -1 0 10272 0 -1 11340
box -48 -56 528 834
use sg13g2_or2_1  _1347_
timestamp 1747056038
transform -1 0 10752 0 -1 11340
box -48 -56 528 834
use sg13g2_nand2b_1  _1348_
timestamp 1747056038
transform -1 0 9696 0 -1 12852
box -48 -56 528 834
use sg13g2_xnor2_1  _1349_
timestamp 1747056038
transform -1 0 10464 0 -1 12852
box -48 -56 816 834
use sg13g2_xnor2_1  _1350_
timestamp 1747056038
transform -1 0 10752 0 1 12852
box -48 -56 816 834
use sg13g2_inv_1  _1351_
timestamp 1747056038
transform 1 0 8352 0 -1 15876
box -48 -56 336 834
use sg13g2_a21oi_1  _1352_
timestamp 1747056038
transform -1 0 10368 0 -1 14364
box -48 -56 528 834
use sg13g2_a22oi_1  _1353_
timestamp 1747056038
transform 1 0 6912 0 1 9828
box -48 -56 624 834
use sg13g2_nand2b_1  _1354_
timestamp 1747056038
transform 1 0 10560 0 1 9828
box -48 -56 528 834
use sg13g2_nor2b_1  _1355_
timestamp 1747056038
transform 1 0 10368 0 -1 9828
box -54 -56 528 834
use sg13g2_xnor2_1  _1356_
timestamp 1747056038
transform 1 0 7488 0 1 9828
box -48 -56 816 834
use sg13g2_xnor2_1  _1357_
timestamp 1747056038
transform 1 0 8256 0 1 9828
box -48 -56 816 834
use sg13g2_nand2_1  _1358_
timestamp 1747056038
transform 1 0 7872 0 -1 11340
box -48 -56 432 834
use sg13g2_xnor2_1  _1359_
timestamp 1747056038
transform -1 0 10560 0 1 9828
box -48 -56 816 834
use sg13g2_a21oi_1  _1360_
timestamp 1747056038
transform -1 0 7872 0 -1 11340
box -48 -56 528 834
use sg13g2_xnor2_1  _1361_
timestamp 1747056038
transform -1 0 9792 0 1 9828
box -48 -56 816 834
use sg13g2_o21ai_1  _1362_
timestamp 1747056038
transform 1 0 9120 0 -1 9828
box -48 -56 538 834
use sg13g2_a21oi_1  _1363_
timestamp 1747056038
transform -1 0 8736 0 -1 11340
box -48 -56 528 834
use sg13g2_o21ai_1  _1364_
timestamp 1747056038
transform 1 0 10752 0 1 12852
box -48 -56 538 834
use sg13g2_a21o_1  _1365_
timestamp 1747056038
transform 1 0 9312 0 1 12852
box -48 -56 720 834
use sg13g2_o21ai_1  _1366_
timestamp 1747056038
transform -1 0 6144 0 -1 15876
box -48 -56 538 834
use sg13g2_a22oi_1  _1367_
timestamp 1747056038
transform 1 0 5088 0 -1 17388
box -48 -56 624 834
use sg13g2_nor2_1  _1368_
timestamp 1747056038
transform 1 0 4032 0 -1 17388
box -48 -56 432 834
use sg13g2_nor2_1  _1369_
timestamp 1747056038
transform 1 0 2976 0 -1 17388
box -48 -56 432 834
use sg13g2_o21ai_1  _1370_
timestamp 1747056038
transform 1 0 1056 0 -1 18900
box -48 -56 538 834
use sg13g2_a21oi_2  _1371_
timestamp 1747056038
transform 1 0 1152 0 1 17388
box -48 -56 816 834
use sg13g2_o21ai_1  _1372_
timestamp 1747056038
transform -1 0 2784 0 1 17388
box -48 -56 538 834
use sg13g2_nor2_1  _1373_
timestamp 1747056038
transform -1 0 3168 0 -1 15876
box -48 -56 432 834
use sg13g2_o21ai_1  _1374_
timestamp 1747056038
transform -1 0 2304 0 -1 17388
box -48 -56 538 834
use sg13g2_nand2_1  _1375_
timestamp 1747056038
transform 1 0 13344 0 1 15876
box -48 -56 432 834
use sg13g2_mux2_1  _1376_
timestamp 1747056038
transform 1 0 23040 0 1 15876
box -48 -56 1008 834
use sg13g2_mux2_2  _1377_
timestamp 1747056038
transform -1 0 23616 0 -1 17388
box -48 -56 1104 834
use sg13g2_a22oi_1  _1378_
timestamp 1747056038
transform -1 0 13344 0 -1 15876
box -48 -56 624 834
use sg13g2_a21oi_1  _1379_
timestamp 1747056038
transform -1 0 13728 0 1 14364
box -48 -56 528 834
use sg13g2_nand3_1  _1380_
timestamp 1747056038
transform -1 0 13248 0 1 14364
box -48 -56 528 834
use sg13g2_a21oi_1  _1381_
timestamp 1747056038
transform -1 0 10560 0 1 11340
box -48 -56 528 834
use sg13g2_and2_1  _1382_
timestamp 1747056038
transform 1 0 12288 0 1 8316
box -48 -56 528 834
use sg13g2_xor2_1  _1383_
timestamp 1747056038
transform 1 0 13056 0 -1 8316
box -48 -56 816 834
use sg13g2_xor2_1  _1384_
timestamp 1747056038
transform -1 0 13824 0 -1 11340
box -48 -56 816 834
use sg13g2_o21ai_1  _1385_
timestamp 1747056038
transform 1 0 12000 0 -1 11340
box -48 -56 538 834
use sg13g2_nand2_1  _1386_
timestamp 1747056038
transform 1 0 10560 0 1 11340
box -48 -56 432 834
use sg13g2_xnor2_1  _1387_
timestamp 1747056038
transform -1 0 13344 0 1 11340
box -48 -56 816 834
use sg13g2_xnor2_1  _1388_
timestamp 1747056038
transform 1 0 12480 0 -1 12852
box -48 -56 816 834
use sg13g2_xor2_1  _1389_
timestamp 1747056038
transform 1 0 11808 0 -1 14364
box -48 -56 816 834
use sg13g2_a21o_1  _1390_
timestamp 1747056038
transform -1 0 13248 0 -1 14364
box -48 -56 720 834
use sg13g2_o21ai_1  _1391_
timestamp 1747056038
transform 1 0 11520 0 1 9828
box -48 -56 538 834
use sg13g2_xor2_1  _1392_
timestamp 1747056038
transform 1 0 10944 0 -1 9828
box -48 -56 816 834
use sg13g2_xnor2_1  _1393_
timestamp 1747056038
transform 1 0 11712 0 -1 9828
box -48 -56 816 834
use sg13g2_and2_1  _1394_
timestamp 1747056038
transform 1 0 10272 0 1 6804
box -48 -56 528 834
use sg13g2_xor2_1  _1395_
timestamp 1747056038
transform 1 0 11424 0 -1 6804
box -48 -56 816 834
use sg13g2_o21ai_1  _1396_
timestamp 1747056038
transform 1 0 9696 0 -1 9828
box -48 -56 538 834
use sg13g2_xor2_1  _1397_
timestamp 1747056038
transform 1 0 12000 0 1 6804
box -48 -56 816 834
use sg13g2_a21oi_1  _1398_
timestamp 1747056038
transform 1 0 12000 0 1 9828
box -48 -56 528 834
use sg13g2_o21ai_1  _1399_
timestamp 1747056038
transform 1 0 12480 0 1 9828
box -48 -56 538 834
use sg13g2_a21oi_1  _1400_
timestamp 1747056038
transform 1 0 11136 0 -1 12852
box -48 -56 528 834
use sg13g2_o21ai_1  _1401_
timestamp 1747056038
transform -1 0 13824 0 1 11340
box -48 -56 538 834
use sg13g2_a21oi_1  _1402_
timestamp 1747056038
transform 1 0 12288 0 -1 15876
box -48 -56 528 834
use sg13g2_o21ai_1  _1403_
timestamp 1747056038
transform -1 0 12768 0 1 15876
box -48 -56 538 834
use sg13g2_nor2b_1  _1404_
timestamp 1747056038
transform -1 0 2304 0 -1 15876
box -54 -56 528 834
use sg13g2_o21ai_1  _1405_
timestamp 1747056038
transform 1 0 2304 0 -1 17388
box -48 -56 538 834
use sg13g2_a21oi_2  _1406_
timestamp 1747056038
transform -1 0 2016 0 1 15876
box -48 -56 816 834
use sg13g2_o21ai_1  _1407_
timestamp 1747056038
transform 1 0 12768 0 1 20412
box -48 -56 538 834
use sg13g2_nor2_1  _1408_
timestamp 1747056038
transform 1 0 8160 0 -1 23436
box -48 -56 432 834
use sg13g2_o21ai_1  _1409_
timestamp 1747056038
transform 1 0 13248 0 1 20412
box -48 -56 538 834
use sg13g2_o21ai_1  _1410_
timestamp 1747056038
transform 1 0 12576 0 -1 11340
box -48 -56 538 834
use sg13g2_and2_1  _1411_
timestamp 1747056038
transform -1 0 18144 0 1 9828
box -48 -56 528 834
use sg13g2_xor2_1  _1412_
timestamp 1747056038
transform 1 0 15648 0 1 6804
box -48 -56 816 834
use sg13g2_xor2_1  _1413_
timestamp 1747056038
transform -1 0 15360 0 -1 11340
box -48 -56 816 834
use sg13g2_a21oi_1  _1414_
timestamp 1747056038
transform 1 0 13632 0 1 9828
box -48 -56 528 834
use sg13g2_nor2_1  _1415_
timestamp 1747056038
transform 1 0 11616 0 -1 11340
box -48 -56 432 834
use sg13g2_xor2_1  _1416_
timestamp 1747056038
transform -1 0 14592 0 -1 11340
box -48 -56 816 834
use sg13g2_nor2_1  _1417_
timestamp 1747056038
transform -1 0 14496 0 1 9828
box -48 -56 432 834
use sg13g2_nand2_1  _1418_
timestamp 1747056038
transform 1 0 13824 0 1 11340
box -48 -56 432 834
use sg13g2_nor2_1  _1419_
timestamp 1747056038
transform -1 0 15072 0 1 11340
box -48 -56 432 834
use sg13g2_xnor2_1  _1420_
timestamp 1747056038
transform -1 0 18048 0 -1 14364
box -48 -56 816 834
use sg13g2_o21ai_1  _1421_
timestamp 1747056038
transform -1 0 14496 0 1 12852
box -48 -56 538 834
use sg13g2_a22oi_1  _1422_
timestamp 1747056038
transform -1 0 13056 0 -1 9828
box -48 -56 624 834
use sg13g2_xor2_1  _1423_
timestamp 1747056038
transform -1 0 15648 0 -1 9828
box -48 -56 816 834
use sg13g2_nand2b_1  _1424_
timestamp 1747056038
transform 1 0 14496 0 1 9828
box -48 -56 528 834
use sg13g2_xor2_1  _1425_
timestamp 1747056038
transform -1 0 14880 0 -1 9828
box -48 -56 816 834
use sg13g2_xnor2_1  _1426_
timestamp 1747056038
transform 1 0 12960 0 1 6804
box -48 -56 816 834
use sg13g2_a21o_1  _1427_
timestamp 1747056038
transform -1 0 12768 0 -1 8316
box -48 -56 720 834
use sg13g2_nor2b_1  _1428_
timestamp 1747056038
transform 1 0 14880 0 -1 6804
box -54 -56 528 834
use sg13g2_xnor2_1  _1429_
timestamp 1747056038
transform -1 0 14496 0 1 6804
box -48 -56 816 834
use sg13g2_a21oi_1  _1430_
timestamp 1747056038
transform 1 0 13632 0 -1 9828
box -48 -56 528 834
use sg13g2_o21ai_1  _1431_
timestamp 1747056038
transform -1 0 13632 0 1 9828
box -48 -56 538 834
use sg13g2_a221oi_1  _1432_
timestamp 1747056038
transform 1 0 13824 0 -1 12852
box -48 -56 816 834
use sg13g2_nor2_1  _1433_
timestamp 1747056038
transform -1 0 16896 0 -1 17388
box -48 -56 432 834
use sg13g2_mux4_1  _1434_
timestamp 1747056038
transform 1 0 26208 0 1 15876
box -48 -56 2064 834
use sg13g2_a221oi_1  _1435_
timestamp 1747056038
transform -1 0 16032 0 -1 17388
box -48 -56 816 834
use sg13g2_nor2_1  _1436_
timestamp 1747056038
transform -1 0 13344 0 1 18900
box -48 -56 432 834
use sg13g2_a21oi_1  _1437_
timestamp 1747056038
transform -1 0 12768 0 -1 20412
box -48 -56 528 834
use sg13g2_or3_1  _1438_
timestamp 1747056038
transform 1 0 13248 0 -1 20412
box -48 -56 720 834
use sg13g2_a21oi_1  _1439_
timestamp 1747056038
transform 1 0 14400 0 -1 20412
box -48 -56 528 834
use sg13g2_a21oi_1  _1440_
timestamp 1747056038
transform 1 0 13920 0 -1 20412
box -48 -56 528 834
use sg13g2_o21ai_1  _1441_
timestamp 1747056038
transform 1 0 13632 0 -1 21924
box -48 -56 538 834
use sg13g2_a21oi_2  _1442_
timestamp 1747056038
transform 1 0 14112 0 -1 21924
box -48 -56 816 834
use sg13g2_o21ai_1  _1443_
timestamp 1747056038
transform 1 0 16704 0 1 20412
box -48 -56 538 834
use sg13g2_nor2_1  _1444_
timestamp 1747056038
transform -1 0 16896 0 -1 21924
box -48 -56 432 834
use sg13g2_o21ai_1  _1445_
timestamp 1747056038
transform 1 0 17568 0 1 18900
box -48 -56 538 834
use sg13g2_xnor2_1  _1446_
timestamp 1747056038
transform -1 0 17280 0 -1 14364
box -48 -56 816 834
use sg13g2_a21oi_1  _1447_
timestamp 1747056038
transform 1 0 15840 0 -1 14364
box -48 -56 528 834
use sg13g2_o21ai_1  _1448_
timestamp 1747056038
transform 1 0 15744 0 -1 9828
box -48 -56 538 834
use sg13g2_xor2_1  _1449_
timestamp 1747056038
transform -1 0 17280 0 -1 8316
box -48 -56 816 834
use sg13g2_a21oi_1  _1450_
timestamp 1747056038
transform 1 0 15168 0 1 6804
box -48 -56 528 834
use sg13g2_xor2_1  _1451_
timestamp 1747056038
transform 1 0 15552 0 -1 6804
box -48 -56 816 834
use sg13g2_xnor2_1  _1452_
timestamp 1747056038
transform -1 0 17184 0 1 6804
box -48 -56 816 834
use sg13g2_xnor2_1  _1453_
timestamp 1747056038
transform 1 0 15744 0 -1 8316
box -48 -56 816 834
use sg13g2_xnor2_1  _1454_
timestamp 1747056038
transform -1 0 16992 0 -1 9828
box -48 -56 816 834
use sg13g2_a21oi_1  _1455_
timestamp 1747056038
transform -1 0 15648 0 1 12852
box -48 -56 528 834
use sg13g2_a21oi_1  _1456_
timestamp 1747056038
transform -1 0 14688 0 1 11340
box -48 -56 528 834
use sg13g2_a21o_1  _1457_
timestamp 1747056038
transform -1 0 15648 0 1 9828
box -48 -56 720 834
use sg13g2_xnor2_1  _1458_
timestamp 1747056038
transform -1 0 17184 0 1 9828
box -48 -56 816 834
use sg13g2_xnor2_1  _1459_
timestamp 1747056038
transform -1 0 18912 0 -1 12852
box -48 -56 816 834
use sg13g2_xnor2_1  _1460_
timestamp 1747056038
transform -1 0 16320 0 1 11340
box -48 -56 816 834
use sg13g2_xnor2_1  _1461_
timestamp 1747056038
transform 1 0 15360 0 -1 12852
box -48 -56 816 834
use sg13g2_mux2_1  _1462_
timestamp 1747056038
transform -1 0 16608 0 1 12852
box -48 -56 1008 834
use sg13g2_nor2_1  _1463_
timestamp 1747056038
transform -1 0 15840 0 -1 15876
box -48 -56 432 834
use sg13g2_nor2b_1  _1464_
timestamp 1747056038
transform -1 0 24480 0 -1 14364
box -54 -56 528 834
use sg13g2_nor2_1  _1465_
timestamp 1747056038
transform -1 0 28608 0 1 15876
box -48 -56 432 834
use sg13g2_a21oi_2  _1466_
timestamp 1747056038
transform 1 0 23712 0 1 17388
box -48 -56 816 834
use sg13g2_a221oi_1  _1467_
timestamp 1747056038
transform 1 0 15552 0 1 15876
box -48 -56 816 834
use sg13g2_nor2_1  _1468_
timestamp 1747056038
transform 1 0 16224 0 1 20412
box -48 -56 432 834
use sg13g2_a221oi_1  _1469_
timestamp 1747056038
transform -1 0 17760 0 -1 18900
box -48 -56 816 834
use sg13g2_o21ai_1  _1470_
timestamp 1747056038
transform 1 0 15744 0 -1 18900
box -48 -56 538 834
use sg13g2_a21oi_1  _1471_
timestamp 1747056038
transform 1 0 16608 0 1 18900
box -48 -56 528 834
use sg13g2_a21oi_1  _1472_
timestamp 1747056038
transform -1 0 17280 0 -1 20412
box -48 -56 528 834
use sg13g2_o21ai_1  _1473_
timestamp 1747056038
transform 1 0 18336 0 -1 20412
box -48 -56 538 834
use sg13g2_a21oi_2  _1474_
timestamp 1747056038
transform -1 0 18720 0 1 20412
box -48 -56 816 834
use sg13g2_nor2_1  _1475_
timestamp 1747056038
transform 1 0 8544 0 1 15876
box -48 -56 432 834
use sg13g2_nand2b_2  _1476_
timestamp 1747056038
transform 1 0 9120 0 1 17388
box -48 -56 816 834
use sg13g2_nor2_1  _1477_
timestamp 1747056038
transform 1 0 5952 0 -1 18900
box -48 -56 432 834
use sg13g2_a221oi_1  _1478_
timestamp 1747056038
transform 1 0 6912 0 -1 18900
box -48 -56 816 834
use sg13g2_nand2b_1  _1479_
timestamp 1747056038
transform -1 0 6720 0 -1 17388
box -48 -56 528 834
use sg13g2_nor2_1  _1480_
timestamp 1747056038
transform -1 0 9120 0 -1 20412
box -48 -56 432 834
use sg13g2_nand2_2  _1481_
timestamp 1747056038
transform -1 0 14688 0 -1 14364
box -48 -56 624 834
use sg13g2_nor2_1  _1482_
timestamp 1747056038
transform 1 0 4704 0 -1 17388
box -48 -56 432 834
use sg13g2_or2_1  _1483_
timestamp 1747056038
transform -1 0 7200 0 1 17388
box -48 -56 528 834
use sg13g2_a22oi_1  _1484_
timestamp 1747056038
transform 1 0 6144 0 1 17388
box -48 -56 624 834
use sg13g2_o21ai_1  _1485_
timestamp 1747056038
transform -1 0 5952 0 -1 18900
box -48 -56 538 834
use sg13g2_a221oi_1  _1486_
timestamp 1747056038
transform 1 0 5376 0 1 17388
box -48 -56 816 834
use sg13g2_nor2_1  _1487_
timestamp 1747056038
transform 1 0 2880 0 -1 21924
box -48 -56 432 834
use sg13g2_o21ai_1  _1488_
timestamp 1747056038
transform 1 0 7872 0 -1 21924
box -48 -56 538 834
use sg13g2_a21oi_2  _1489_
timestamp 1747056038
transform -1 0 8832 0 1 21924
box -48 -56 816 834
use sg13g2_a22oi_1  _1490_
timestamp 1747056038
transform -1 0 8256 0 -1 18900
box -48 -56 624 834
use sg13g2_o21ai_1  _1491_
timestamp 1747056038
transform 1 0 6912 0 -1 20412
box -48 -56 538 834
use sg13g2_nor2_1  _1492_
timestamp 1747056038
transform -1 0 6336 0 -1 14364
box -48 -56 432 834
use sg13g2_and2_1  _1493_
timestamp 1747056038
transform 1 0 4128 0 1 11340
box -48 -56 528 834
use sg13g2_xnor2_1  _1494_
timestamp 1747056038
transform 1 0 4608 0 1 11340
box -48 -56 816 834
use sg13g2_xnor2_1  _1495_
timestamp 1747056038
transform 1 0 4800 0 -1 11340
box -48 -56 816 834
use sg13g2_nand2_1  _1496_
timestamp 1747056038
transform -1 0 960 0 1 6804
box -48 -56 432 834
use sg13g2_nand2_1  _1497_
timestamp 1747056038
transform 1 0 1344 0 1 6804
box -48 -56 432 834
use sg13g2_nor2_1  _1498_
timestamp 1747056038
transform 1 0 1056 0 -1 6804
box -48 -56 432 834
use sg13g2_xor2_1  _1499_
timestamp 1747056038
transform 1 0 1056 0 1 9828
box -48 -56 816 834
use sg13g2_xnor2_1  _1500_
timestamp 1747056038
transform 1 0 1728 0 -1 11340
box -48 -56 816 834
use sg13g2_a21oi_1  _1501_
timestamp 1747056038
transform -1 0 4800 0 -1 11340
box -48 -56 528 834
use sg13g2_o21ai_1  _1502_
timestamp 1747056038
transform 1 0 5472 0 1 11340
box -48 -56 538 834
use sg13g2_o21ai_1  _1503_
timestamp 1747056038
transform 1 0 6336 0 -1 14364
box -48 -56 538 834
use sg13g2_nand3b_1  _1504_
timestamp 1747056038
transform -1 0 7968 0 -1 14364
box -48 -56 720 834
use sg13g2_nand3_1  _1505_
timestamp 1747056038
transform 1 0 6816 0 -1 14364
box -48 -56 528 834
use sg13g2_o21ai_1  _1506_
timestamp 1747056038
transform -1 0 7872 0 -1 20412
box -48 -56 538 834
use sg13g2_a22oi_1  _1507_
timestamp 1747056038
transform 1 0 6336 0 -1 20412
box -48 -56 624 834
use sg13g2_nor2_1  _1508_
timestamp 1747056038
transform 1 0 4128 0 -1 20412
box -48 -56 432 834
use sg13g2_nor2_1  _1509_
timestamp 1747056038
transform 1 0 576 0 -1 26460
box -48 -56 432 834
use sg13g2_o21ai_1  _1510_
timestamp 1747056038
transform -1 0 5760 0 1 21924
box -48 -56 538 834
use sg13g2_a21oi_2  _1511_
timestamp 1747056038
transform -1 0 5280 0 1 21924
box -48 -56 816 834
use sg13g2_a22oi_1  _1512_
timestamp 1747056038
transform 1 0 6528 0 1 15876
box -48 -56 624 834
use sg13g2_o21ai_1  _1513_
timestamp 1747056038
transform -1 0 7488 0 -1 17388
box -48 -56 538 834
use sg13g2_nor2_1  _1514_
timestamp 1747056038
transform -1 0 10272 0 1 14364
box -48 -56 432 834
use sg13g2_nor2_1  _1515_
timestamp 1747056038
transform 1 0 6720 0 -1 15876
box -48 -56 432 834
use sg13g2_a22oi_1  _1516_
timestamp 1747056038
transform -1 0 6144 0 -1 11340
box -48 -56 624 834
use sg13g2_xor2_1  _1517_
timestamp 1747056038
transform 1 0 5760 0 -1 9828
box -48 -56 816 834
use sg13g2_xnor2_1  _1518_
timestamp 1747056038
transform 1 0 6528 0 -1 9828
box -48 -56 816 834
use sg13g2_and2_1  _1519_
timestamp 1747056038
transform 1 0 1728 0 1 6804
box -48 -56 528 834
use sg13g2_or2_1  _1520_
timestamp 1747056038
transform -1 0 4320 0 1 5292
box -48 -56 528 834
use sg13g2_nand2b_1  _1521_
timestamp 1747056038
transform 1 0 2208 0 1 6804
box -48 -56 528 834
use sg13g2_o21ai_1  _1522_
timestamp 1747056038
transform 1 0 1824 0 1 9828
box -48 -56 538 834
use sg13g2_xnor2_1  _1523_
timestamp 1747056038
transform 1 0 2880 0 -1 8316
box -48 -56 816 834
use sg13g2_o21ai_1  _1524_
timestamp 1747056038
transform 1 0 7104 0 1 8316
box -48 -56 538 834
use sg13g2_a21oi_1  _1525_
timestamp 1747056038
transform -1 0 7776 0 -1 9828
box -48 -56 528 834
use sg13g2_nor3_1  _1526_
timestamp 1747056038
transform -1 0 11808 0 -1 14364
box -48 -56 528 834
use sg13g2_nor2_1  _1527_
timestamp 1747056038
transform -1 0 10752 0 -1 14364
box -48 -56 432 834
use sg13g2_o21ai_1  _1528_
timestamp 1747056038
transform 1 0 7488 0 1 14364
box -48 -56 538 834
use sg13g2_o21ai_1  _1529_
timestamp 1747056038
transform -1 0 6528 0 1 15876
box -48 -56 538 834
use sg13g2_a22oi_1  _1530_
timestamp 1747056038
transform 1 0 5376 0 1 15876
box -48 -56 624 834
use sg13g2_nor2_1  _1531_
timestamp 1747056038
transform 1 0 4032 0 -1 18900
box -48 -56 432 834
use sg13g2_nor2_1  _1532_
timestamp 1747056038
transform 1 0 3552 0 -1 18900
box -48 -56 432 834
use sg13g2_o21ai_1  _1533_
timestamp 1747056038
transform 1 0 1728 0 -1 20412
box -48 -56 538 834
use sg13g2_a21oi_1  _1534_
timestamp 1747056038
transform -1 0 2688 0 -1 20412
box -48 -56 528 834
use sg13g2_a22oi_1  _1535_
timestamp 1747056038
transform -1 0 9504 0 -1 17388
box -48 -56 624 834
use sg13g2_o21ai_1  _1536_
timestamp 1747056038
transform 1 0 8544 0 1 18900
box -48 -56 538 834
use sg13g2_o21ai_1  _1537_
timestamp 1747056038
transform 1 0 9408 0 -1 14364
box -48 -56 538 834
use sg13g2_and2_1  _1538_
timestamp 1747056038
transform 1 0 6816 0 -1 6804
box -48 -56 528 834
use sg13g2_xor2_1  _1539_
timestamp 1747056038
transform 1 0 7296 0 -1 6804
box -48 -56 816 834
use sg13g2_a21o_1  _1540_
timestamp 1747056038
transform -1 0 3360 0 1 6804
box -48 -56 720 834
use sg13g2_xor2_1  _1541_
timestamp 1747056038
transform 1 0 8064 0 1 6804
box -48 -56 816 834
use sg13g2_or2_1  _1542_
timestamp 1747056038
transform 1 0 6144 0 1 8316
box -48 -56 528 834
use sg13g2_o21ai_1  _1543_
timestamp 1747056038
transform 1 0 6624 0 1 8316
box -48 -56 538 834
use sg13g2_and2_1  _1544_
timestamp 1747056038
transform -1 0 8448 0 -1 9828
box -48 -56 528 834
use sg13g2_xnor2_1  _1545_
timestamp 1747056038
transform -1 0 8832 0 1 8316
box -48 -56 816 834
use sg13g2_xnor2_1  _1546_
timestamp 1747056038
transform 1 0 8064 0 -1 8316
box -48 -56 816 834
use sg13g2_xnor2_1  _1547_
timestamp 1747056038
transform 1 0 8832 0 -1 8316
box -48 -56 816 834
use sg13g2_o21ai_1  _1548_
timestamp 1747056038
transform 1 0 9408 0 1 14364
box -48 -56 538 834
use sg13g2_nor2_1  _1549_
timestamp 1747056038
transform -1 0 18432 0 1 18900
box -48 -56 432 834
use sg13g2_a21oi_1  _1550_
timestamp 1747056038
transform 1 0 11136 0 1 18900
box -48 -56 528 834
use sg13g2_a21oi_1  _1551_
timestamp 1747056038
transform -1 0 9888 0 -1 20412
box -48 -56 528 834
use sg13g2_o21ai_1  _1552_
timestamp 1747056038
transform 1 0 9888 0 -1 20412
box -48 -56 538 834
use sg13g2_a21oi_1  _1553_
timestamp 1747056038
transform 1 0 10176 0 1 18900
box -48 -56 528 834
use sg13g2_o21ai_1  _1554_
timestamp 1747056038
transform -1 0 11328 0 -1 20412
box -48 -56 538 834
use sg13g2_o21ai_1  _1555_
timestamp 1747056038
transform -1 0 10848 0 -1 20412
box -48 -56 538 834
use sg13g2_nand2b_1  _1556_
timestamp 1747056038
transform 1 0 768 0 -1 20412
box -48 -56 528 834
use sg13g2_nand2_1  _1557_
timestamp 1747056038
transform -1 0 28896 0 -1 18900
box -48 -56 432 834
use sg13g2_a21oi_2  _1558_
timestamp 1747056038
transform -1 0 2784 0 1 20412
box -48 -56 816 834
use sg13g2_nor2_1  _1559_
timestamp 1747056038
transform -1 0 10848 0 1 17388
box -48 -56 432 834
use sg13g2_a221oi_1  _1560_
timestamp 1747056038
transform 1 0 10464 0 -1 15876
box -48 -56 816 834
use sg13g2_or2_1  _1561_
timestamp 1747056038
transform 1 0 10464 0 1 15876
box -48 -56 528 834
use sg13g2_nor2_1  _1562_
timestamp 1747056038
transform -1 0 12288 0 1 14364
box -48 -56 432 834
use sg13g2_a21oi_1  _1563_
timestamp 1747056038
transform -1 0 8064 0 1 8316
box -48 -56 528 834
use sg13g2_xnor2_1  _1564_
timestamp 1747056038
transform -1 0 12096 0 -1 8316
box -48 -56 816 834
use sg13g2_xor2_1  _1565_
timestamp 1747056038
transform 1 0 11232 0 1 8316
box -48 -56 816 834
use sg13g2_nand2_1  _1566_
timestamp 1747056038
transform -1 0 12288 0 -1 5292
box -48 -56 432 834
use sg13g2_xnor2_1  _1567_
timestamp 1747056038
transform 1 0 10752 0 1 6804
box -48 -56 816 834
use sg13g2_a21oi_1  _1568_
timestamp 1747056038
transform -1 0 8640 0 -1 6804
box -48 -56 528 834
use sg13g2_xnor2_1  _1569_
timestamp 1747056038
transform -1 0 11424 0 -1 6804
box -48 -56 816 834
use sg13g2_a21oi_1  _1570_
timestamp 1747056038
transform 1 0 10368 0 -1 8316
box -48 -56 528 834
use sg13g2_o21ai_1  _1571_
timestamp 1747056038
transform -1 0 12000 0 1 6804
box -48 -56 538 834
use sg13g2_o21ai_1  _1572_
timestamp 1747056038
transform 1 0 11424 0 1 14364
box -48 -56 538 834
use sg13g2_nor2_1  _1573_
timestamp 1747056038
transform -1 0 18240 0 1 14364
box -48 -56 432 834
use sg13g2_a21oi_1  _1574_
timestamp 1747056038
transform 1 0 17184 0 -1 15876
box -48 -56 528 834
use sg13g2_a22oi_1  _1575_
timestamp 1747056038
transform -1 0 12000 0 -1 15876
box -48 -56 624 834
use sg13g2_o21ai_1  _1576_
timestamp 1747056038
transform -1 0 11328 0 -1 17388
box -48 -56 538 834
use sg13g2_a21oi_1  _1577_
timestamp 1747056038
transform 1 0 3744 0 1 17388
box -48 -56 528 834
use sg13g2_o21ai_1  _1578_
timestamp 1747056038
transform -1 0 2016 0 -1 18900
box -48 -56 538 834
use sg13g2_a21oi_1  _1579_
timestamp 1747056038
transform 1 0 864 0 -1 17388
box -48 -56 528 834
use sg13g2_and2_1  _1580_
timestamp 1747056038
transform -1 0 14208 0 -1 17388
box -48 -56 528 834
use sg13g2_a221oi_1  _1581_
timestamp 1747056038
transform 1 0 13728 0 1 15876
box -48 -56 816 834
use sg13g2_or2_1  _1582_
timestamp 1747056038
transform -1 0 15264 0 -1 15876
box -48 -56 528 834
use sg13g2_nor2_1  _1583_
timestamp 1747056038
transform 1 0 13248 0 -1 14364
box -48 -56 432 834
use sg13g2_nand2b_1  _1584_
timestamp 1747056038
transform -1 0 13536 0 -1 9828
box -48 -56 528 834
use sg13g2_o21ai_1  _1585_
timestamp 1747056038
transform 1 0 10848 0 -1 8316
box -48 -56 538 834
use sg13g2_nor2_1  _1586_
timestamp 1747056038
transform 1 0 17280 0 1 8316
box -48 -56 432 834
use sg13g2_xnor2_1  _1587_
timestamp 1747056038
transform 1 0 12768 0 1 8316
box -48 -56 816 834
use sg13g2_xnor2_1  _1588_
timestamp 1747056038
transform -1 0 15072 0 1 8316
box -48 -56 816 834
use sg13g2_and2_1  _1589_
timestamp 1747056038
transform 1 0 12384 0 -1 6804
box -48 -56 528 834
use sg13g2_xor2_1  _1590_
timestamp 1747056038
transform -1 0 14112 0 -1 6804
box -48 -56 816 834
use sg13g2_o21ai_1  _1591_
timestamp 1747056038
transform 1 0 11424 0 -1 5292
box -48 -56 538 834
use sg13g2_xor2_1  _1592_
timestamp 1747056038
transform 1 0 14112 0 -1 6804
box -48 -56 816 834
use sg13g2_a21oi_1  _1593_
timestamp 1747056038
transform 1 0 14496 0 1 6804
box -48 -56 528 834
use sg13g2_o21ai_1  _1594_
timestamp 1747056038
transform -1 0 14592 0 -1 8316
box -48 -56 538 834
use sg13g2_o21ai_1  _1595_
timestamp 1747056038
transform 1 0 13632 0 -1 14364
box -48 -56 538 834
use sg13g2_nor3_1  _1596_
timestamp 1747056038
transform -1 0 18624 0 -1 15876
box -48 -56 528 834
use sg13g2_nor2_1  _1597_
timestamp 1747056038
transform 1 0 17184 0 1 14364
box -48 -56 432 834
use sg13g2_a22oi_1  _1598_
timestamp 1747056038
transform 1 0 14208 0 -1 15876
box -48 -56 624 834
use sg13g2_o21ai_1  _1599_
timestamp 1747056038
transform -1 0 14208 0 -1 15876
box -48 -56 538 834
use sg13g2_a21oi_1  _1600_
timestamp 1747056038
transform 1 0 2016 0 1 15876
box -48 -56 528 834
use sg13g2_o21ai_1  _1601_
timestamp 1747056038
transform 1 0 768 0 1 15876
box -48 -56 538 834
use sg13g2_a21oi_1  _1602_
timestamp 1747056038
transform -1 0 1824 0 -1 17388
box -48 -56 528 834
use sg13g2_o21ai_1  _1603_
timestamp 1747056038
transform -1 0 15840 0 -1 14364
box -48 -56 538 834
use sg13g2_nand2_1  _1604_
timestamp 1747056038
transform -1 0 21504 0 -1 5292
box -48 -56 432 834
use sg13g2_nor2_1  _1605_
timestamp 1747056038
transform 1 0 19200 0 -1 6804
box -48 -56 432 834
use sg13g2_xnor2_1  _1606_
timestamp 1747056038
transform -1 0 18144 0 -1 6804
box -48 -56 816 834
use sg13g2_a21oi_1  _1607_
timestamp 1747056038
transform 1 0 12864 0 -1 6804
box -48 -56 528 834
use sg13g2_xnor2_1  _1608_
timestamp 1747056038
transform -1 0 17376 0 -1 6804
box -48 -56 816 834
use sg13g2_a21oi_2  _1609_
timestamp 1747056038
transform 1 0 13536 0 1 8316
box -48 -56 816 834
use sg13g2_nand2b_1  _1610_
timestamp 1747056038
transform 1 0 17184 0 1 9828
box -48 -56 528 834
use sg13g2_nor2b_1  _1611_
timestamp 1747056038
transform 1 0 17184 0 -1 11340
box -54 -56 528 834
use sg13g2_xnor2_1  _1612_
timestamp 1747056038
transform 1 0 15648 0 1 9828
box -48 -56 816 834
use sg13g2_xnor2_1  _1613_
timestamp 1747056038
transform 1 0 15648 0 -1 11340
box -48 -56 816 834
use sg13g2_xnor2_1  _1614_
timestamp 1747056038
transform -1 0 17184 0 -1 11340
box -48 -56 816 834
use sg13g2_o21ai_1  _1615_
timestamp 1747056038
transform 1 0 14880 0 -1 14364
box -48 -56 538 834
use sg13g2_nor2_1  _1616_
timestamp 1747056038
transform -1 0 15264 0 1 14364
box -48 -56 432 834
use sg13g2_a21oi_1  _1617_
timestamp 1747056038
transform 1 0 14496 0 -1 18900
box -48 -56 528 834
use sg13g2_a22oi_1  _1618_
timestamp 1747056038
transform 1 0 14688 0 -1 17388
box -48 -56 624 834
use sg13g2_o21ai_1  _1619_
timestamp 1747056038
transform -1 0 15072 0 1 17388
box -48 -56 538 834
use sg13g2_o21ai_1  _1620_
timestamp 1747056038
transform 1 0 13344 0 1 17388
box -48 -56 538 834
use sg13g2_a221oi_1  _1621_
timestamp 1747056038
transform 1 0 13824 0 1 17388
box -48 -56 816 834
use sg13g2_o21ai_1  _1622_
timestamp 1747056038
transform 1 0 14016 0 -1 18900
box -48 -56 538 834
use sg13g2_nor2_1  _1623_
timestamp 1747056038
transform 1 0 14208 0 -1 17388
box -48 -56 432 834
use sg13g2_nor2_1  _1624_
timestamp 1747056038
transform -1 0 16032 0 -1 21924
box -48 -56 432 834
use sg13g2_o21ai_1  _1625_
timestamp 1747056038
transform 1 0 13728 0 1 20412
box -48 -56 538 834
use sg13g2_a21oi_2  _1626_
timestamp 1747056038
transform 1 0 14208 0 1 20412
box -48 -56 816 834
use sg13g2_nor2_1  _1627_
timestamp 1747056038
transform -1 0 16224 0 -1 15876
box -48 -56 432 834
use sg13g2_a221oi_1  _1628_
timestamp 1747056038
transform -1 0 15552 0 1 15876
box -48 -56 816 834
use sg13g2_or2_1  _1629_
timestamp 1747056038
transform 1 0 16512 0 -1 15876
box -48 -56 528 834
use sg13g2_o21ai_1  _1630_
timestamp 1747056038
transform 1 0 14688 0 1 12852
box -48 -56 538 834
use sg13g2_nor2_1  _1631_
timestamp 1747056038
transform -1 0 16896 0 1 14364
box -48 -56 432 834
use sg13g2_or2_1  _1632_
timestamp 1747056038
transform 1 0 16320 0 1 11340
box -48 -56 528 834
use sg13g2_o21ai_1  _1633_
timestamp 1747056038
transform 1 0 18144 0 -1 11340
box -48 -56 538 834
use sg13g2_xnor2_1  _1634_
timestamp 1747056038
transform 1 0 18528 0 1 9828
box -48 -56 816 834
use sg13g2_o21ai_1  _1635_
timestamp 1747056038
transform 1 0 19584 0 1 6804
box -48 -56 538 834
use sg13g2_xnor2_1  _1636_
timestamp 1747056038
transform 1 0 19584 0 1 8316
box -48 -56 816 834
use sg13g2_xnor2_1  _1637_
timestamp 1747056038
transform -1 0 21024 0 -1 9828
box -48 -56 816 834
use sg13g2_xnor2_1  _1638_
timestamp 1747056038
transform -1 0 19488 0 -1 9828
box -48 -56 816 834
use sg13g2_and2_1  _1639_
timestamp 1747056038
transform -1 0 18144 0 -1 11340
box -48 -56 528 834
use sg13g2_o21ai_1  _1640_
timestamp 1747056038
transform 1 0 18720 0 1 11340
box -48 -56 538 834
use sg13g2_o21ai_1  _1641_
timestamp 1747056038
transform -1 0 17376 0 1 11340
box -48 -56 538 834
use sg13g2_nor2_1  _1642_
timestamp 1747056038
transform -1 0 18240 0 -1 17388
box -48 -56 432 834
use sg13g2_a21oi_1  _1643_
timestamp 1747056038
transform 1 0 17664 0 -1 15876
box -48 -56 528 834
use sg13g2_a22oi_1  _1644_
timestamp 1747056038
transform -1 0 17664 0 1 15876
box -48 -56 624 834
use sg13g2_o21ai_1  _1645_
timestamp 1747056038
transform 1 0 17664 0 1 15876
box -48 -56 538 834
use sg13g2_a21oi_1  _1646_
timestamp 1747056038
transform -1 0 16800 0 -1 20412
box -48 -56 528 834
use sg13g2_o21ai_1  _1647_
timestamp 1747056038
transform 1 0 17376 0 -1 21924
box -48 -56 538 834
use sg13g2_a21oi_2  _1648_
timestamp 1747056038
transform -1 0 17952 0 1 20412
box -48 -56 816 834
use sg13g2_nor2_2  _1649_
timestamp 1747056038
transform 1 0 8736 0 -1 18900
box -48 -56 624 834
use sg13g2_nor2_1  _1650_
timestamp 1747056038
transform 1 0 6528 0 1 20412
box -48 -56 432 834
use sg13g2_a221oi_1  _1651_
timestamp 1747056038
transform 1 0 6912 0 1 18900
box -48 -56 816 834
use sg13g2_and2_1  _1652_
timestamp 1747056038
transform -1 0 5184 0 -1 18900
box -48 -56 528 834
use sg13g2_nand2_1  _1653_
timestamp 1747056038
transform -1 0 4224 0 1 9828
box -48 -56 432 834
use sg13g2_inv_1  _1654_
timestamp 1747056038
transform 1 0 2304 0 1 9828
box -48 -56 336 834
use sg13g2_xnor2_1  _1655_
timestamp 1747056038
transform -1 0 5664 0 -1 9828
box -48 -56 816 834
use sg13g2_xnor2_1  _1656_
timestamp 1747056038
transform 1 0 4128 0 -1 9828
box -48 -56 816 834
use sg13g2_nand2_1  _1657_
timestamp 1747056038
transform -1 0 6048 0 1 9828
box -48 -56 432 834
use sg13g2_nand2_1  _1658_
timestamp 1747056038
transform 1 0 1344 0 -1 8316
box -48 -56 432 834
use sg13g2_xnor2_1  _1659_
timestamp 1747056038
transform -1 0 4128 0 1 8316
box -48 -56 816 834
use sg13g2_xor2_1  _1660_
timestamp 1747056038
transform 1 0 3360 0 -1 9828
box -48 -56 816 834
use sg13g2_a21oi_1  _1661_
timestamp 1747056038
transform -1 0 5664 0 1 8316
box -48 -56 528 834
use sg13g2_o21ai_1  _1662_
timestamp 1747056038
transform 1 0 4608 0 1 9828
box -48 -56 538 834
use sg13g2_a221oi_1  _1663_
timestamp 1747056038
transform 1 0 4704 0 -1 14364
box -48 -56 816 834
use sg13g2_o21ai_1  _1664_
timestamp 1747056038
transform -1 0 4608 0 1 18900
box -48 -56 538 834
use sg13g2_o21ai_1  _1665_
timestamp 1747056038
transform -1 0 5088 0 1 18900
box -48 -56 538 834
use sg13g2_a21oi_1  _1666_
timestamp 1747056038
transform -1 0 6912 0 -1 21924
box -48 -56 528 834
use sg13g2_o21ai_1  _1667_
timestamp 1747056038
transform 1 0 6912 0 1 20412
box -48 -56 538 834
use sg13g2_a21oi_1  _1668_
timestamp 1747056038
transform 1 0 6336 0 1 21924
box -48 -56 528 834
use sg13g2_a22oi_1  _1669_
timestamp 1747056038
transform 1 0 6336 0 -1 18900
box -48 -56 624 834
use sg13g2_o21ai_1  _1670_
timestamp 1747056038
transform -1 0 6912 0 1 18900
box -48 -56 538 834
use sg13g2_a22oi_1  _1671_
timestamp 1747056038
transform -1 0 5664 0 1 9828
box -48 -56 624 834
use sg13g2_xor2_1  _1672_
timestamp 1747056038
transform 1 0 6240 0 -1 8316
box -48 -56 816 834
use sg13g2_xor2_1  _1673_
timestamp 1747056038
transform -1 0 6240 0 -1 8316
box -48 -56 816 834
use sg13g2_and2_1  _1674_
timestamp 1747056038
transform 1 0 3936 0 1 6804
box -48 -56 528 834
use sg13g2_xor2_1  _1675_
timestamp 1747056038
transform 1 0 4416 0 1 8316
box -48 -56 816 834
use sg13g2_o21ai_1  _1676_
timestamp 1747056038
transform 1 0 3456 0 1 6804
box -48 -56 538 834
use sg13g2_xnor2_1  _1677_
timestamp 1747056038
transform 1 0 4800 0 1 6804
box -48 -56 816 834
use sg13g2_a21oi_1  _1678_
timestamp 1747056038
transform 1 0 4992 0 -1 8316
box -48 -56 528 834
use sg13g2_o21ai_1  _1679_
timestamp 1747056038
transform 1 0 5952 0 1 6804
box -48 -56 538 834
use sg13g2_a21oi_1  _1680_
timestamp 1747056038
transform 1 0 6144 0 -1 12852
box -48 -56 528 834
use sg13g2_o21ai_1  _1681_
timestamp 1747056038
transform 1 0 5664 0 1 12852
box -48 -56 538 834
use sg13g2_o21ai_1  _1682_
timestamp 1747056038
transform -1 0 6336 0 1 18900
box -48 -56 538 834
use sg13g2_a22oi_1  _1683_
timestamp 1747056038
transform 1 0 5760 0 -1 20412
box -48 -56 624 834
use sg13g2_inv_1  _1684_
timestamp 1747056038
transform 1 0 3840 0 -1 20412
box -48 -56 336 834
use sg13g2_a21oi_1  _1685_
timestamp 1747056038
transform -1 0 5760 0 -1 21924
box -48 -56 528 834
use sg13g2_o21ai_1  _1686_
timestamp 1747056038
transform 1 0 4032 0 1 21924
box -48 -56 538 834
use sg13g2_a21oi_1  _1687_
timestamp 1747056038
transform -1 0 5280 0 -1 21924
box -48 -56 528 834
use sg13g2_a22oi_1  _1688_
timestamp 1747056038
transform 1 0 7872 0 1 15876
box -48 -56 624 834
use sg13g2_o21ai_1  _1689_
timestamp 1747056038
transform -1 0 7584 0 -1 15876
box -48 -56 538 834
use sg13g2_nand2_1  _1690_
timestamp 1747056038
transform 1 0 5280 0 -1 15876
box -48 -56 432 834
use sg13g2_nand2_1  _1691_
timestamp 1747056038
transform -1 0 10272 0 1 3780
box -48 -56 432 834
use sg13g2_xnor2_1  _1692_
timestamp 1747056038
transform -1 0 10176 0 -1 6804
box -48 -56 816 834
use sg13g2_a21oi_1  _1693_
timestamp 1747056038
transform -1 0 6144 0 1 8316
box -48 -56 528 834
use sg13g2_xnor2_1  _1694_
timestamp 1747056038
transform -1 0 10176 0 1 6804
box -48 -56 816 834
use sg13g2_or2_1  _1695_
timestamp 1747056038
transform 1 0 7200 0 -1 8316
box -48 -56 528 834
use sg13g2_o21ai_1  _1696_
timestamp 1747056038
transform 1 0 7392 0 1 6804
box -48 -56 538 834
use sg13g2_and2_1  _1697_
timestamp 1747056038
transform 1 0 10176 0 -1 6804
box -48 -56 528 834
use sg13g2_xnor2_1  _1698_
timestamp 1747056038
transform 1 0 9312 0 1 8316
box -48 -56 816 834
use sg13g2_xor2_1  _1699_
timestamp 1747056038
transform -1 0 10368 0 -1 8316
box -48 -56 816 834
use sg13g2_o21ai_1  _1700_
timestamp 1747056038
transform -1 0 9312 0 1 8316
box -48 -56 538 834
use sg13g2_a21oi_1  _1701_
timestamp 1747056038
transform -1 0 9120 0 -1 9828
box -48 -56 528 834
use sg13g2_nor2_1  _1702_
timestamp 1747056038
transform 1 0 3744 0 1 14364
box -48 -56 432 834
use sg13g2_o21ai_1  _1703_
timestamp 1747056038
transform -1 0 10368 0 -1 15876
box -48 -56 538 834
use sg13g2_o21ai_1  _1704_
timestamp 1747056038
transform 1 0 5280 0 1 14364
box -48 -56 538 834
use sg13g2_nand2_1  _1705_
timestamp 1747056038
transform -1 0 5280 0 1 14364
box -48 -56 432 834
use sg13g2_o21ai_1  _1706_
timestamp 1747056038
transform -1 0 5280 0 -1 15876
box -48 -56 538 834
use sg13g2_a21oi_1  _1707_
timestamp 1747056038
transform 1 0 3552 0 1 18900
box -48 -56 528 834
use sg13g2_o21ai_1  _1708_
timestamp 1747056038
transform -1 0 3360 0 -1 20412
box -48 -56 538 834
use sg13g2_a21oi_1  _1709_
timestamp 1747056038
transform 1 0 3072 0 -1 18900
box -48 -56 528 834
use sg13g2_a21oi_2  _1710_
timestamp 1747056038
transform 1 0 10080 0 1 8316
box -48 -56 816 834
use sg13g2_xnor2_1  _1711_
timestamp 1747056038
transform -1 0 16800 0 1 8316
box -48 -56 816 834
use sg13g2_xnor2_1  _1712_
timestamp 1747056038
transform -1 0 16032 0 1 8316
box -48 -56 816 834
use sg13g2_and2_1  _1713_
timestamp 1747056038
transform 1 0 18144 0 -1 6804
box -48 -56 528 834
use sg13g2_xor2_1  _1714_
timestamp 1747056038
transform 1 0 17280 0 1 6804
box -48 -56 816 834
use sg13g2_o21ai_1  _1715_
timestamp 1747056038
transform -1 0 9408 0 1 6804
box -48 -56 538 834
use sg13g2_xor2_1  _1716_
timestamp 1747056038
transform -1 0 18240 0 -1 8316
box -48 -56 816 834
use sg13g2_a21oi_1  _1717_
timestamp 1747056038
transform 1 0 14592 0 -1 8316
box -48 -56 528 834
use sg13g2_o21ai_1  _1718_
timestamp 1747056038
transform -1 0 15552 0 -1 8316
box -48 -56 538 834
use sg13g2_nand2b_1  _1719_
timestamp 1747056038
transform -1 0 9408 0 1 14364
box -48 -56 528 834
use sg13g2_o21ai_1  _1720_
timestamp 1747056038
transform 1 0 8640 0 -1 15876
box -48 -56 538 834
use sg13g2_a21oi_2  _1721_
timestamp 1747056038
transform -1 0 9888 0 -1 15876
box -48 -56 816 834
use sg13g2_a22oi_1  _1722_
timestamp 1747056038
transform 1 0 10752 0 1 14364
box -48 -56 624 834
use sg13g2_o21ai_1  _1723_
timestamp 1747056038
transform -1 0 10752 0 1 14364
box -48 -56 538 834
use sg13g2_o21ai_1  _1724_
timestamp 1747056038
transform -1 0 4416 0 1 15876
box -48 -56 538 834
use sg13g2_a21oi_1  _1725_
timestamp 1747056038
transform 1 0 3168 0 -1 15876
box -48 -56 528 834
use sg13g2_nor2_1  _1726_
timestamp 1747056038
transform 1 0 2112 0 -1 6804
box -48 -56 432 834
use sg13g2_o21ai_1  _1727_
timestamp 1747056038
transform 1 0 1248 0 -1 20412
box -48 -56 538 834
use sg13g2_a21oi_1  _1728_
timestamp 1747056038
transform 1 0 3360 0 -1 20412
box -48 -56 528 834
use sg13g2_nand2b_1  _1729_
timestamp 1747056038
transform -1 0 17472 0 -1 9828
box -48 -56 528 834
use sg13g2_o21ai_1  _1730_
timestamp 1747056038
transform 1 0 16800 0 1 8316
box -48 -56 538 834
use sg13g2_nor2_1  _1731_
timestamp 1747056038
transform 1 0 17472 0 -1 9828
box -48 -56 432 834
use sg13g2_xor2_1  _1732_
timestamp 1747056038
transform 1 0 17856 0 -1 9828
box -48 -56 816 834
use sg13g2_xnor2_1  _1733_
timestamp 1747056038
transform 1 0 18048 0 1 8316
box -48 -56 816 834
use sg13g2_a21oi_1  _1734_
timestamp 1747056038
transform 1 0 18624 0 -1 6804
box -48 -56 528 834
use sg13g2_nor2_1  _1735_
timestamp 1747056038
transform 1 0 19008 0 -1 8316
box -48 -56 432 834
use sg13g2_xor2_1  _1736_
timestamp 1747056038
transform 1 0 18048 0 1 6804
box -48 -56 816 834
use sg13g2_xnor2_1  _1737_
timestamp 1747056038
transform 1 0 18240 0 -1 8316
box -48 -56 816 834
use sg13g2_xnor2_1  _1738_
timestamp 1747056038
transform -1 0 20256 0 -1 9828
box -48 -56 816 834
use sg13g2_o21ai_1  _1739_
timestamp 1747056038
transform -1 0 13824 0 -1 12852
box -48 -56 538 834
use sg13g2_a21oi_1  _1740_
timestamp 1747056038
transform 1 0 12288 0 1 12852
box -48 -56 528 834
use sg13g2_a22oi_1  _1741_
timestamp 1747056038
transform 1 0 10944 0 1 15876
box -48 -56 624 834
use sg13g2_o21ai_1  _1742_
timestamp 1747056038
transform 1 0 11328 0 -1 17388
box -48 -56 538 834
use sg13g2_inv_1  _1743_
timestamp 1747056038
transform -1 0 13248 0 -1 18900
box -48 -56 336 834
use sg13g2_o21ai_1  _1744_
timestamp 1747056038
transform -1 0 12480 0 1 17388
box -48 -56 538 834
use sg13g2_a221oi_1  _1745_
timestamp 1747056038
transform 1 0 11904 0 -1 17388
box -48 -56 816 834
use sg13g2_a21oi_1  _1746_
timestamp 1747056038
transform 1 0 11520 0 1 17388
box -48 -56 528 834
use sg13g2_a21oi_1  _1747_
timestamp 1747056038
transform 1 0 3264 0 1 17388
box -48 -56 528 834
use sg13g2_o21ai_1  _1748_
timestamp 1747056038
transform -1 0 3072 0 -1 18900
box -48 -56 538 834
use sg13g2_a21oi_1  _1749_
timestamp 1747056038
transform 1 0 672 0 1 17388
box -48 -56 528 834
use sg13g2_a21oi_2  _1750_
timestamp 1747056038
transform -1 0 19584 0 1 8316
box -48 -56 816 834
use sg13g2_nor2b_1  _1751_
timestamp 1747056038
transform 1 0 22464 0 1 6804
box -54 -56 528 834
use sg13g2_xnor2_1  _1752_
timestamp 1747056038
transform -1 0 22272 0 -1 8316
box -48 -56 816 834
use sg13g2_nand2b_1  _1753_
timestamp 1747056038
transform 1 0 22656 0 1 8316
box -48 -56 528 834
use sg13g2_xor2_1  _1754_
timestamp 1747056038
transform 1 0 20544 0 1 8316
box -48 -56 816 834
use sg13g2_xnor2_1  _1755_
timestamp 1747056038
transform 1 0 20064 0 -1 8316
box -48 -56 816 834
use sg13g2_a221oi_1  _1756_
timestamp 1747056038
transform 1 0 18816 0 1 6804
box -48 -56 816 834
use sg13g2_nor3_1  _1757_
timestamp 1747056038
transform 1 0 20160 0 1 6804
box -48 -56 528 834
use sg13g2_o21ai_1  _1758_
timestamp 1747056038
transform 1 0 20640 0 1 6804
box -48 -56 538 834
use sg13g2_nand2b_1  _1759_
timestamp 1747056038
transform 1 0 20832 0 -1 8316
box -48 -56 528 834
use sg13g2_xnor2_1  _1760_
timestamp 1747056038
transform -1 0 21792 0 -1 9828
box -48 -56 816 834
use sg13g2_a21oi_1  _1761_
timestamp 1747056038
transform 1 0 16128 0 -1 12852
box -48 -56 528 834
use sg13g2_o21ai_1  _1762_
timestamp 1747056038
transform -1 0 14208 0 1 14364
box -48 -56 538 834
use sg13g2_nand2_1  _1763_
timestamp 1747056038
transform 1 0 13344 0 -1 15876
box -48 -56 432 834
use sg13g2_a22oi_1  _1764_
timestamp 1747056038
transform -1 0 13344 0 1 15876
box -48 -56 624 834
use sg13g2_nand2_2  _1765_
timestamp 1747056038
transform 1 0 13152 0 -1 17388
box -48 -56 624 834
use sg13g2_o21ai_1  _1766_
timestamp 1747056038
transform -1 0 13344 0 1 17388
box -48 -56 538 834
use sg13g2_a21oi_1  _1767_
timestamp 1747056038
transform -1 0 13152 0 -1 17388
box -48 -56 528 834
use sg13g2_o21ai_1  _1768_
timestamp 1747056038
transform -1 0 13824 0 1 12852
box -48 -56 538 834
use sg13g2_o21ai_1  _1769_
timestamp 1747056038
transform 1 0 3456 0 1 15876
box -48 -56 538 834
use sg13g2_inv_1  _1770_
timestamp 1747056038
transform -1 0 4032 0 -1 17388
box -48 -56 336 834
use sg13g2_a21oi_1  _1771_
timestamp 1747056038
transform 1 0 2496 0 1 15876
box -48 -56 528 834
use sg13g2_o21ai_1  _1772_
timestamp 1747056038
transform 1 0 2304 0 -1 15876
box -48 -56 538 834
use sg13g2_a21oi_1  _1773_
timestamp 1747056038
transform 1 0 1344 0 -1 15876
box -48 -56 528 834
use sg13g2_nor3_1  _1774_
timestamp 1747056038
transform 1 0 22944 0 -1 5292
box -48 -56 528 834
use sg13g2_or3_1  _1775_
timestamp 1747056038
transform 1 0 22272 0 -1 8316
box -48 -56 720 834
use sg13g2_o21ai_1  _1776_
timestamp 1747056038
transform 1 0 26592 0 -1 8316
box -48 -56 538 834
use sg13g2_a21oi_1  _1777_
timestamp 1747056038
transform 1 0 25632 0 -1 8316
box -48 -56 528 834
use sg13g2_nand3_1  _1778_
timestamp 1747056038
transform 1 0 22944 0 1 6804
box -48 -56 528 834
use sg13g2_nand3_1  _1779_
timestamp 1747056038
transform 1 0 21120 0 1 6804
box -48 -56 528 834
use sg13g2_o21ai_1  _1780_
timestamp 1747056038
transform -1 0 24096 0 -1 8316
box -48 -56 538 834
use sg13g2_a21oi_1  _1781_
timestamp 1747056038
transform 1 0 23136 0 -1 8316
box -48 -56 528 834
use sg13g2_nand2_1  _1782_
timestamp 1747056038
transform -1 0 27552 0 1 8316
box -48 -56 432 834
use sg13g2_nor2_1  _1783_
timestamp 1747056038
transform -1 0 27168 0 1 8316
box -48 -56 432 834
use sg13g2_xnor2_1  _1784_
timestamp 1747056038
transform -1 0 26304 0 1 8316
box -48 -56 816 834
use sg13g2_a21oi_1  _1785_
timestamp 1747056038
transform 1 0 21312 0 1 8316
box -48 -56 528 834
use sg13g2_xnor2_1  _1786_
timestamp 1747056038
transform -1 0 24000 0 1 8316
box -48 -56 816 834
use sg13g2_xnor2_1  _1787_
timestamp 1747056038
transform -1 0 23520 0 -1 9828
box -48 -56 816 834
use sg13g2_o21ai_1  _1788_
timestamp 1747056038
transform 1 0 15072 0 1 11340
box -48 -56 538 834
use sg13g2_a21oi_1  _1789_
timestamp 1747056038
transform 1 0 16032 0 1 14364
box -48 -56 528 834
use sg13g2_nor2_1  _1790_
timestamp 1747056038
transform -1 0 18240 0 1 17388
box -48 -56 432 834
use sg13g2_a221oi_1  _1791_
timestamp 1747056038
transform -1 0 16032 0 1 17388
box -48 -56 816 834
use sg13g2_a21oi_1  _1792_
timestamp 1747056038
transform 1 0 15168 0 1 18900
box -48 -56 528 834
use sg13g2_o21ai_1  _1793_
timestamp 1747056038
transform 1 0 14688 0 1 18900
box -48 -56 538 834
use sg13g2_a21o_1  _1794_
timestamp 1747056038
transform 1 0 15360 0 1 14364
box -48 -56 720 834
use sg13g2_a21oi_1  _1795_
timestamp 1747056038
transform 1 0 15072 0 -1 20412
box -48 -56 528 834
use sg13g2_a21oi_1  _1796_
timestamp 1747056038
transform 1 0 14208 0 1 18900
box -48 -56 528 834
use sg13g2_o21ai_1  _1797_
timestamp 1747056038
transform 1 0 14976 0 1 20412
box -48 -56 538 834
use sg13g2_a21oi_2  _1798_
timestamp 1747056038
transform -1 0 15648 0 -1 21924
box -48 -56 816 834
use sg13g2_xor2_1  _1799_
timestamp 1747056038
transform -1 0 19680 0 -1 12852
box -48 -56 816 834
use sg13g2_a21oi_1  _1800_
timestamp 1747056038
transform 1 0 17376 0 -1 12852
box -48 -56 528 834
use sg13g2_o21ai_1  _1801_
timestamp 1747056038
transform -1 0 26784 0 1 8316
box -48 -56 538 834
use sg13g2_xnor2_1  _1802_
timestamp 1747056038
transform 1 0 24000 0 1 8316
box -48 -56 816 834
use sg13g2_xnor2_1  _1803_
timestamp 1747056038
transform -1 0 25536 0 1 8316
box -48 -56 816 834
use sg13g2_xnor2_1  _1804_
timestamp 1747056038
transform 1 0 23136 0 1 9828
box -48 -56 816 834
use sg13g2_a21oi_1  _1805_
timestamp 1747056038
transform 1 0 26112 0 -1 8316
box -48 -56 528 834
use sg13g2_o21ai_1  _1806_
timestamp 1747056038
transform 1 0 24096 0 -1 8316
box -48 -56 538 834
use sg13g2_xnor2_1  _1807_
timestamp 1747056038
transform 1 0 23520 0 -1 9828
box -48 -56 816 834
use sg13g2_xnor2_1  _1808_
timestamp 1747056038
transform -1 0 24672 0 1 9828
box -48 -56 816 834
use sg13g2_a21oi_1  _1809_
timestamp 1747056038
transform 1 0 17376 0 1 11340
box -48 -56 528 834
use sg13g2_o21ai_1  _1810_
timestamp 1747056038
transform -1 0 17280 0 -1 12852
box -48 -56 538 834
use sg13g2_nor2_1  _1811_
timestamp 1747056038
transform 1 0 16032 0 1 17388
box -48 -56 432 834
use sg13g2_a221oi_1  _1812_
timestamp 1747056038
transform 1 0 16320 0 1 15876
box -48 -56 816 834
use sg13g2_nor2_1  _1813_
timestamp 1747056038
transform -1 0 17280 0 -1 17388
box -48 -56 432 834
use sg13g2_a221oi_1  _1814_
timestamp 1747056038
transform -1 0 16992 0 -1 18900
box -48 -56 816 834
use sg13g2_o21ai_1  _1815_
timestamp 1747056038
transform -1 0 17376 0 1 12852
box -48 -56 538 834
use sg13g2_a21oi_1  _1816_
timestamp 1747056038
transform 1 0 16128 0 1 18900
box -48 -56 528 834
use sg13g2_a21oi_1  _1817_
timestamp 1747056038
transform -1 0 17568 0 1 18900
box -48 -56 528 834
use sg13g2_o21ai_1  _1818_
timestamp 1747056038
transform 1 0 15840 0 -1 20412
box -48 -56 538 834
use sg13g2_a21oi_2  _1819_
timestamp 1747056038
transform 1 0 17568 0 -1 20412
box -48 -56 816 834
use sg13g2_a21o_1  _1820_
timestamp 1747056038
transform 1 0 25152 0 1 21924
box -48 -56 720 834
use sg13g2_nand3_1  _1821_
timestamp 1747056038
transform -1 0 23904 0 1 14364
box -48 -56 528 834
use sg13g2_o21ai_1  _1822_
timestamp 1747056038
transform -1 0 22560 0 1 14364
box -48 -56 538 834
use sg13g2_nand2_1  _1823_
timestamp 1747056038
transform -1 0 22752 0 -1 14364
box -48 -56 432 834
use sg13g2_nor4_1  _1824_
timestamp 1747056038
transform 1 0 21408 0 -1 15876
box -48 -56 624 834
use sg13g2_nand3_1  _1825_
timestamp 1747056038
transform 1 0 21600 0 1 14364
box -48 -56 528 834
use sg13g2_o21ai_1  _1826_
timestamp 1747056038
transform 1 0 21984 0 -1 15876
box -48 -56 538 834
use sg13g2_and3_2  _1827_
timestamp 1747056038
transform -1 0 22368 0 1 15876
box -48 -56 720 834
use sg13g2_nand3_1  _1828_
timestamp 1747056038
transform -1 0 22848 0 1 15876
box -48 -56 528 834
use sg13g2_nor2_2  _1829_
timestamp 1747056038
transform -1 0 22752 0 -1 18900
box -48 -56 624 834
use sg13g2_nand2_2  _1830_
timestamp 1747056038
transform -1 0 20352 0 1 15876
box -48 -56 624 834
use sg13g2_and2_1  _1831_
timestamp 1747056038
transform -1 0 18432 0 -1 18900
box -48 -56 528 834
use sg13g2_nor3_1  _1832_
timestamp 1747056038
transform 1 0 21024 0 1 12852
box -48 -56 528 834
use sg13g2_xnor2_1  _1833_
timestamp 1747056038
transform -1 0 20736 0 -1 11340
box -48 -56 816 834
use sg13g2_nor2_1  _1834_
timestamp 1747056038
transform 1 0 18144 0 1 9828
box -48 -56 432 834
use sg13g2_nor2_1  _1835_
timestamp 1747056038
transform -1 0 20448 0 -1 12852
box -48 -56 432 834
use sg13g2_xnor2_1  _1836_
timestamp 1747056038
transform 1 0 19776 0 1 11340
box -48 -56 816 834
use sg13g2_nor2_1  _1837_
timestamp 1747056038
transform -1 0 22176 0 1 8316
box -48 -56 432 834
use sg13g2_xnor2_1  _1838_
timestamp 1747056038
transform 1 0 24768 0 1 12852
box -48 -56 816 834
use sg13g2_nor2_1  _1839_
timestamp 1747056038
transform -1 0 28416 0 -1 12852
box -48 -56 432 834
use sg13g2_nand2_1  _1840_
timestamp 1747056038
transform 1 0 27456 0 -1 11340
box -48 -56 432 834
use sg13g2_nor2_2  _1841_
timestamp 1747056038
transform 1 0 24768 0 -1 12852
box -48 -56 624 834
use sg13g2_a21oi_1  _1842_
timestamp 1747056038
transform -1 0 25824 0 -1 12852
box -48 -56 528 834
use sg13g2_nor3_1  _1843_
timestamp 1747056038
transform 1 0 24288 0 1 12852
box -48 -56 528 834
use sg13g2_o21ai_1  _1844_
timestamp 1747056038
transform 1 0 27072 0 -1 12852
box -48 -56 538 834
use sg13g2_a21oi_1  _1845_
timestamp 1747056038
transform 1 0 27552 0 -1 12852
box -48 -56 528 834
use sg13g2_nor3_1  _1846_
timestamp 1747056038
transform -1 0 28032 0 1 11340
box -48 -56 528 834
use sg13g2_xnor2_1  _1847_
timestamp 1747056038
transform 1 0 24384 0 -1 9828
box -48 -56 816 834
use sg13g2_nor2_1  _1848_
timestamp 1747056038
transform 1 0 26016 0 -1 9828
box -48 -56 432 834
use sg13g2_nand3_1  _1849_
timestamp 1747056038
transform -1 0 24480 0 1 15876
box -48 -56 528 834
use sg13g2_xor2_1  _1850_
timestamp 1747056038
transform -1 0 25824 0 -1 15876
box -48 -56 816 834
use sg13g2_nor2_1  _1851_
timestamp 1747056038
transform 1 0 23328 0 1 17388
box -48 -56 432 834
use sg13g2_nor2_1  _1852_
timestamp 1747056038
transform -1 0 28992 0 1 15876
box -48 -56 432 834
use sg13g2_xnor2_1  _1853_
timestamp 1747056038
transform 1 0 24288 0 -1 15876
box -48 -56 816 834
use sg13g2_nor2_1  _1854_
timestamp 1747056038
transform -1 0 27552 0 1 17388
box -48 -56 432 834
use sg13g2_nand3_1  _1855_
timestamp 1747056038
transform 1 0 17184 0 1 26460
box -48 -56 528 834
use sg13g2_nor4_1  _1856_
timestamp 1747056038
transform 1 0 18912 0 -1 26460
box -48 -56 624 834
use sg13g2_nor2_1  _1857_
timestamp 1747056038
transform -1 0 29568 0 1 24948
box -48 -56 432 834
use sg13g2_and3_1  _1858_
timestamp 1747056038
transform 1 0 14880 0 1 26460
box -48 -56 720 834
use sg13g2_nand3_1  _1859_
timestamp 1747056038
transform 1 0 19680 0 1 24948
box -48 -56 528 834
use sg13g2_and2_1  _1860_
timestamp 1747056038
transform 1 0 18720 0 1 24948
box -48 -56 528 834
use sg13g2_nor4_2  _1861_
timestamp 1747056038
transform 1 0 18624 0 -1 24948
box -48 -56 1200 834
use sg13g2_or4_1  _1862_
timestamp 1747056038
transform 1 0 18720 0 1 26460
box -48 -56 816 834
use sg13g2_nand4_1  _1863_
timestamp 1747056038
transform 1 0 18144 0 1 26460
box -48 -56 624 834
use sg13g2_o21ai_1  _1864_
timestamp 1747056038
transform 1 0 19200 0 1 24948
box -48 -56 538 834
use sg13g2_inv_1  _1865_
timestamp 1747056038
transform -1 0 20448 0 1 24948
box -48 -56 336 834
use sg13g2_nor3_1  _1866_
timestamp 1747056038
transform 1 0 17664 0 -1 24948
box -48 -56 528 834
use sg13g2_nor2b_2  _1867_
timestamp 1747056038
transform -1 0 17664 0 -1 24948
box -54 -56 720 834
use sg13g2_nor2_1  _1868_
timestamp 1747056038
transform -1 0 30816 0 1 20412
box -48 -56 432 834
use sg13g2_nor2b_1  _1869_
timestamp 1747056038
transform 1 0 1920 0 -1 26460
box -54 -56 528 834
use sg13g2_nor3_1  _1870_
timestamp 1747056038
transform 1 0 768 0 1 24948
box -48 -56 528 834
use sg13g2_a21oi_1  _1871_
timestamp 1747056038
transform 1 0 1056 0 1 23436
box -48 -56 528 834
use sg13g2_and4_1  _1872_
timestamp 1747056038
transform 1 0 5952 0 1 23436
box -48 -56 816 834
use sg13g2_and3_1  _1873_
timestamp 1747056038
transform -1 0 2208 0 1 21924
box -48 -56 720 834
use sg13g2_nor3_1  _1874_
timestamp 1747056038
transform -1 0 1056 0 1 23436
box -48 -56 528 834
use sg13g2_nor2_1  _1875_
timestamp 1747056038
transform 1 0 576 0 -1 11340
box -48 -56 432 834
use sg13g2_and2_1  _1876_
timestamp 1747056038
transform 1 0 672 0 -1 14364
box -48 -56 528 834
use sg13g2_nor3_1  _1877_
timestamp 1747056038
transform -1 0 3552 0 1 14364
box -48 -56 528 834
use sg13g2_nor2b_1  _1878_
timestamp 1747056038
transform 1 0 864 0 -1 15876
box -54 -56 528 834
use sg13g2_a21oi_1  _1879_
timestamp 1747056038
transform -1 0 1824 0 -1 9828
box -48 -56 528 834
use sg13g2_o21ai_1  _1880_
timestamp 1747056038
transform 1 0 1824 0 -1 9828
box -48 -56 538 834
use sg13g2_inv_1  _1881_
timestamp 1747056038
transform 1 0 576 0 -1 9828
box -48 -56 336 834
use sg13g2_nand2_1  _1882_
timestamp 1747056038
transform 1 0 2016 0 -1 8316
box -48 -56 432 834
use sg13g2_xor2_1  _1883_
timestamp 1747056038
transform 1 0 2880 0 -1 6804
box -48 -56 816 834
use sg13g2_nor2_1  _1884_
timestamp 1747056038
transform -1 0 3840 0 1 5292
box -48 -56 432 834
use sg13g2_nor2_1  _1885_
timestamp 1747056038
transform -1 0 5952 0 1 6804
box -48 -56 432 834
use sg13g2_a21oi_1  _1886_
timestamp 1747056038
transform 1 0 5472 0 1 5292
box -48 -56 528 834
use sg13g2_o21ai_1  _1887_
timestamp 1747056038
transform 1 0 4992 0 1 5292
box -48 -56 538 834
use sg13g2_inv_1  _1888_
timestamp 1747056038
transform 1 0 6144 0 -1 5292
box -48 -56 336 834
use sg13g2_and4_2  _1889_
timestamp 1747056038
transform 1 0 4128 0 -1 8316
box -48 -56 912 834
use sg13g2_xnor2_1  _1890_
timestamp 1747056038
transform 1 0 9408 0 -1 5292
box -48 -56 816 834
use sg13g2_nor2_1  _1891_
timestamp 1747056038
transform -1 0 11040 0 -1 5292
box -48 -56 432 834
use sg13g2_a21oi_1  _1892_
timestamp 1747056038
transform -1 0 14112 0 -1 5292
box -48 -56 528 834
use sg13g2_and3_1  _1893_
timestamp 1747056038
transform -1 0 13440 0 1 5292
box -48 -56 720 834
use sg13g2_nor3_1  _1894_
timestamp 1747056038
transform 1 0 12672 0 -1 5292
box -48 -56 528 834
use sg13g2_nand3_1  _1895_
timestamp 1747056038
transform 1 0 13152 0 -1 5292
box -48 -56 528 834
use sg13g2_xnor2_1  _1896_
timestamp 1747056038
transform 1 0 19392 0 -1 5292
box -48 -56 816 834
use sg13g2_nor2_1  _1897_
timestamp 1747056038
transform 1 0 19584 0 1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _1898_
timestamp 1747056038
transform 1 0 19008 0 -1 5292
box -48 -56 432 834
use sg13g2_nor2_1  _1899_
timestamp 1747056038
transform -1 0 20640 0 1 3780
box -48 -56 432 834
use sg13g2_a21oi_1  _1900_
timestamp 1747056038
transform -1 0 21600 0 1 5292
box -48 -56 528 834
use sg13g2_nor2b_1  _1901_
timestamp 1747056038
transform 1 0 19776 0 -1 6804
box -54 -56 528 834
use sg13g2_or3_1  _1902_
timestamp 1747056038
transform 1 0 20160 0 -1 5292
box -48 -56 720 834
use sg13g2_xor2_1  _1903_
timestamp 1747056038
transform -1 0 23808 0 -1 6804
box -48 -56 816 834
use sg13g2_nor2_1  _1904_
timestamp 1747056038
transform -1 0 23808 0 -1 5292
box -48 -56 432 834
use sg13g2_nor2_1  _1905_
timestamp 1747056038
transform 1 0 22560 0 -1 5292
box -48 -56 432 834
use sg13g2_nor2_1  _1906_
timestamp 1747056038
transform -1 0 24192 0 -1 6804
box -48 -56 432 834
use sg13g2_a21oi_1  _1907_
timestamp 1747056038
transform 1 0 23808 0 -1 5292
box -48 -56 528 834
use sg13g2_nor2b_1  _1908_
timestamp 1747056038
transform 1 0 24768 0 1 5292
box -54 -56 528 834
use sg13g2_xor2_1  _1909_
timestamp 1747056038
transform 1 0 12768 0 -1 21924
box -48 -56 816 834
use sg13g2_xor2_1  _1910_
timestamp 1747056038
transform 1 0 3936 0 -1 24948
box -48 -56 816 834
use sg13g2_xor2_1  _1911_
timestamp 1747056038
transform 1 0 3360 0 -1 23436
box -48 -56 816 834
use sg13g2_nor3_1  _1912_
timestamp 1747056038
transform -1 0 13248 0 -1 24948
box -48 -56 528 834
use sg13g2_nor3_1  _1913_
timestamp 1747056038
transform 1 0 15456 0 1 21924
box -48 -56 528 834
use sg13g2_nor2_1  _1914_
timestamp 1747056038
transform -1 0 16416 0 -1 21924
box -48 -56 432 834
use sg13g2_nand2_2  _1915_
timestamp 1747056038
transform -1 0 14880 0 1 14364
box -48 -56 624 834
use sg13g2_and2_1  _1916_
timestamp 1747056038
transform -1 0 23136 0 -1 24948
box -48 -56 528 834
use sg13g2_a221oi_1  _1917_
timestamp 1747056038
transform -1 0 14496 0 -1 23436
box -48 -56 816 834
use sg13g2_a21oi_1  _1918_
timestamp 1747056038
transform 1 0 8736 0 -1 24948
box -48 -56 528 834
use sg13g2_and2_1  _1919_
timestamp 1747056038
transform 1 0 29184 0 1 23436
box -48 -56 528 834
use sg13g2_a221oi_1  _1920_
timestamp 1747056038
transform -1 0 25824 0 1 23436
box -48 -56 816 834
use sg13g2_a21oi_1  _1921_
timestamp 1747056038
transform 1 0 28704 0 1 24948
box -48 -56 528 834
use sg13g2_nand3_1  _1922_
timestamp 1747056038
transform -1 0 24192 0 -1 23436
box -48 -56 528 834
use sg13g2_a21oi_1  _1923_
timestamp 1747056038
transform 1 0 13248 0 1 24948
box -48 -56 528 834
use sg13g2_a22oi_1  _1924_
timestamp 1747056038
transform 1 0 12672 0 1 24948
box -48 -56 624 834
use sg13g2_and2_1  _1925_
timestamp 1747056038
transform 1 0 28224 0 1 23436
box -48 -56 528 834
use sg13g2_a221oi_1  _1926_
timestamp 1747056038
transform -1 0 16704 0 1 23436
box -48 -56 816 834
use sg13g2_a21oi_1  _1927_
timestamp 1747056038
transform 1 0 16128 0 1 24948
box -48 -56 528 834
use sg13g2_nand2_1  _1928_
timestamp 1747056038
transform 1 0 17856 0 -1 23436
box -48 -56 432 834
use sg13g2_nand3_1  _1929_
timestamp 1747056038
transform 1 0 15936 0 1 21924
box -48 -56 528 834
use sg13g2_nand3_1  _1930_
timestamp 1747056038
transform 1 0 18240 0 -1 23436
box -48 -56 528 834
use sg13g2_and2_1  _1931_
timestamp 1747056038
transform -1 0 25152 0 1 21924
box -48 -56 528 834
use sg13g2_a22oi_1  _1932_
timestamp 1747056038
transform 1 0 23904 0 -1 21924
box -48 -56 624 834
use sg13g2_nand2_1  _1933_
timestamp 1747056038
transform -1 0 30336 0 -1 23436
box -48 -56 432 834
use sg13g2_o21ai_1  _1934_
timestamp 1747056038
transform 1 0 22464 0 1 23436
box -48 -56 538 834
use sg13g2_nand3_1  _1935_
timestamp 1747056038
transform 1 0 23616 0 -1 20412
box -48 -56 528 834
use sg13g2_o21ai_1  _1936_
timestamp 1747056038
transform 1 0 24096 0 -1 20412
box -48 -56 538 834
use sg13g2_mux2_1  _1937_
timestamp 1747056038
transform 1 0 24576 0 -1 20412
box -48 -56 1008 834
use sg13g2_nand3_1  _1938_
timestamp 1747056038
transform 1 0 26688 0 1 21924
box -48 -56 528 834
use sg13g2_o21ai_1  _1939_
timestamp 1747056038
transform 1 0 21216 0 1 21924
box -48 -56 538 834
use sg13g2_mux2_1  _1940_
timestamp 1747056038
transform 1 0 20064 0 -1 21924
box -48 -56 1008 834
use sg13g2_nor2_1  _1941_
timestamp 1747056038
transform 1 0 20640 0 1 12852
box -48 -56 432 834
use sg13g2_nand4_1  _1942_
timestamp 1747056038
transform -1 0 21888 0 -1 14364
box -48 -56 624 834
use sg13g2_nor4_1  _1943_
timestamp 1747056038
transform 1 0 20736 0 -1 14364
box -48 -56 624 834
use sg13g2_nand2_2  _1944_
timestamp 1747056038
transform 1 0 20352 0 1 18900
box -48 -56 624 834
use sg13g2_nand3_1  _1945_
timestamp 1747056038
transform 1 0 22176 0 1 12852
box -48 -56 528 834
use sg13g2_nor2_1  _1946_
timestamp 1747056038
transform -1 0 29088 0 1 12852
box -48 -56 432 834
use sg13g2_nand2_1  _1947_
timestamp 1747056038
transform -1 0 23040 0 1 12852
box -48 -56 432 834
use sg13g2_nor2_1  _1948_
timestamp 1747056038
transform -1 0 27072 0 -1 14364
box -48 -56 432 834
use sg13g2_and2_1  _1949_
timestamp 1747056038
transform 1 0 21888 0 -1 14364
box -48 -56 528 834
use sg13g2_nor4_1  _1950_
timestamp 1747056038
transform 1 0 22848 0 1 14364
box -48 -56 624 834
use sg13g2_a21oi_1  _1951_
timestamp 1747056038
transform -1 0 23520 0 1 12852
box -48 -56 528 834
use sg13g2_nor4_1  _1952_
timestamp 1747056038
transform 1 0 23328 0 -1 14364
box -48 -56 624 834
use sg13g2_a21oi_1  _1953_
timestamp 1747056038
transform 1 0 24480 0 -1 14364
box -48 -56 528 834
use sg13g2_a22oi_1  _1954_
timestamp 1747056038
transform 1 0 22752 0 -1 14364
box -48 -56 624 834
use sg13g2_nor2_1  _1955_
timestamp 1747056038
transform -1 0 29184 0 -1 15876
box -48 -56 432 834
use sg13g2_nand2b_1  _1956_
timestamp 1747056038
transform 1 0 23520 0 1 12852
box -48 -56 528 834
use sg13g2_a21oi_1  _1957_
timestamp 1747056038
transform -1 0 27072 0 -1 12852
box -48 -56 528 834
use sg13g2_nor2_1  _1958_
timestamp 1747056038
transform -1 0 21600 0 1 24948
box -48 -56 432 834
use sg13g2_o21ai_1  _1959_
timestamp 1747056038
transform -1 0 11616 0 -1 26460
box -48 -56 538 834
use sg13g2_a21oi_1  _1960_
timestamp 1747056038
transform -1 0 4800 0 1 24948
box -48 -56 528 834
use sg13g2_a21oi_1  _1961_
timestamp 1747056038
transform 1 0 6336 0 -1 27972
box -48 -56 528 834
use sg13g2_and3_1  _1962_
timestamp 1747056038
transform -1 0 8928 0 1 26460
box -48 -56 720 834
use sg13g2_nor3_1  _1963_
timestamp 1747056038
transform 1 0 5856 0 -1 26460
box -48 -56 528 834
use sg13g2_nand2b_2  _1964_
timestamp 1747056038
transform -1 0 17760 0 1 23436
box -48 -56 816 834
use sg13g2_nand2_1  _1965_
timestamp 1747056038
transform 1 0 3840 0 -1 27972
box -48 -56 432 834
use sg13g2_nand3_1  _1966_
timestamp 1747056038
transform 1 0 14208 0 1 24948
box -48 -56 528 834
use sg13g2_xnor2_1  _1967_
timestamp 1747056038
transform -1 0 9792 0 -1 26460
box -48 -56 816 834
use sg13g2_nor2_1  _1968_
timestamp 1747056038
transform 1 0 1728 0 1 26460
box -48 -56 432 834
use sg13g2_nand2_1  _1969_
timestamp 1747056038
transform -1 0 28704 0 1 26460
box -48 -56 432 834
use sg13g2_nand2_2  _1970_
timestamp 1747056038
transform 1 0 16608 0 1 24948
box -48 -56 624 834
use sg13g2_inv_1  _1971_
timestamp 1747056038
transform -1 0 21984 0 1 21924
box -48 -56 336 834
use sg13g2_nor2_1  _1972_
timestamp 1747056038
transform 1 0 14496 0 1 26460
box -48 -56 432 834
use sg13g2_xnor2_1  _1973_
timestamp 1747056038
transform 1 0 15360 0 1 24948
box -48 -56 816 834
use sg13g2_o21ai_1  _1974_
timestamp 1747056038
transform 1 0 17184 0 1 24948
box -48 -56 538 834
use sg13g2_a21oi_1  _1975_
timestamp 1747056038
transform 1 0 25824 0 1 23436
box -48 -56 528 834
use sg13g2_and3_1  _1976_
timestamp 1747056038
transform 1 0 22464 0 1 24948
box -48 -56 720 834
use sg13g2_nand2_1  _1977_
timestamp 1747056038
transform -1 0 30240 0 1 26460
box -48 -56 432 834
use sg13g2_nor3_1  _1978_
timestamp 1747056038
transform -1 0 26208 0 -1 27972
box -48 -56 528 834
use sg13g2_nand2_1  _1979_
timestamp 1747056038
transform 1 0 30240 0 1 26460
box -48 -56 432 834
use sg13g2_xnor2_1  _1980_
timestamp 1747056038
transform 1 0 21888 0 -1 26460
box -48 -56 816 834
use sg13g2_o21ai_1  _1981_
timestamp 1747056038
transform 1 0 27264 0 -1 26460
box -48 -56 538 834
use sg13g2_a21oi_1  _1982_
timestamp 1747056038
transform 1 0 27744 0 -1 26460
box -48 -56 528 834
use sg13g2_nor2b_1  _1983_
timestamp 1747056038
transform 1 0 27360 0 1 26460
box -54 -56 528 834
use sg13g2_nor2_1  _1984_
timestamp 1747056038
transform -1 0 29760 0 -1 26460
box -48 -56 432 834
use sg13g2_nor3_1  _1985_
timestamp 1747056038
transform -1 0 27360 0 1 26460
box -48 -56 528 834
use sg13g2_xnor2_1  _1986_
timestamp 1747056038
transform 1 0 23136 0 -1 26460
box -48 -56 816 834
use sg13g2_nor2_1  _1987_
timestamp 1747056038
transform -1 0 30528 0 -1 26460
box -48 -56 432 834
use sg13g2_nand2_1  _1988_
timestamp 1747056038
transform -1 0 29856 0 1 26460
box -48 -56 432 834
use sg13g2_a22oi_1  _1989_
timestamp 1747056038
transform -1 0 21792 0 -1 26460
box -48 -56 624 834
use sg13g2_a21oi_1  _1990_
timestamp 1747056038
transform 1 0 20544 0 -1 23436
box -48 -56 528 834
use sg13g2_nor2_1  _1991_
timestamp 1747056038
transform -1 0 28992 0 -1 26460
box -48 -56 432 834
use sg13g2_nand2_1  _1992_
timestamp 1747056038
transform -1 0 29376 0 -1 26460
box -48 -56 432 834
use sg13g2_xnor2_1  _1993_
timestamp 1747056038
transform 1 0 20448 0 1 24948
box -48 -56 816 834
use sg13g2_o21ai_1  _1994_
timestamp 1747056038
transform 1 0 22656 0 -1 26460
box -48 -56 538 834
use sg13g2_o21ai_1  _1995_
timestamp 1747056038
transform -1 0 13632 0 1 26460
box -48 -56 538 834
use sg13g2_nor3_1  _1996_
timestamp 1747056038
transform 1 0 13728 0 1 24948
box -48 -56 528 834
use sg13g2_nand3_1  _1997_
timestamp 1747056038
transform 1 0 14304 0 -1 26460
box -48 -56 528 834
use sg13g2_nor2_1  _1998_
timestamp 1747056038
transform 1 0 2400 0 -1 26460
box -48 -56 432 834
use sg13g2_nor4_1  _1999_
timestamp 1747056038
transform -1 0 14304 0 -1 26460
box -48 -56 624 834
use sg13g2_nor2_1  _2000_
timestamp 1747056038
transform 1 0 8352 0 -1 24948
box -48 -56 432 834
use sg13g2_nand4_1  _2001_
timestamp 1747056038
transform 1 0 13632 0 1 26460
box -48 -56 624 834
use sg13g2_a21oi_1  _2002_
timestamp 1747056038
transform -1 0 15264 0 -1 26460
box -48 -56 528 834
use sg13g2_a22oi_1  _2003_
timestamp 1747056038
transform -1 0 13632 0 -1 26460
box -48 -56 624 834
use sg13g2_nor2_1  _2004_
timestamp 1747056038
transform 1 0 1920 0 -1 27972
box -48 -56 432 834
use sg13g2_nand2b_1  _2005_
timestamp 1747056038
transform 1 0 13152 0 -1 27972
box -48 -56 528 834
use sg13g2_a21oi_1  _2006_
timestamp 1747056038
transform 1 0 13632 0 -1 27972
box -48 -56 528 834
use sg13g2_nor2_1  _2007_
timestamp 1747056038
transform -1 0 31200 0 1 23436
box -48 -56 432 834
use sg13g2_nor2_1  _2008_
timestamp 1747056038
transform 1 0 2112 0 1 26460
box -48 -56 432 834
use sg13g2_a21oi_1  _2009_
timestamp 1747056038
transform 1 0 6720 0 1 23436
box -48 -56 528 834
use sg13g2_o21ai_1  _2010_
timestamp 1747056038
transform 1 0 8928 0 -1 23436
box -48 -56 538 834
use sg13g2_nand2_1  _2011_
timestamp 1747056038
transform -1 0 28704 0 1 18900
box -48 -56 432 834
use sg13g2_o21ai_1  _2012_
timestamp 1747056038
transform -1 0 24384 0 1 18900
box -48 -56 538 834
use sg13g2_nand2_1  _2013_
timestamp 1747056038
transform -1 0 26496 0 1 18900
box -48 -56 432 834
use sg13g2_o21ai_1  _2014_
timestamp 1747056038
transform -1 0 23424 0 1 18900
box -48 -56 538 834
use sg13g2_mux2_1  _2015_
timestamp 1747056038
transform 1 0 2496 0 1 23436
box -48 -56 1008 834
use sg13g2_mux2_1  _2016_
timestamp 1747056038
transform -1 0 3360 0 1 24948
box -48 -56 1008 834
use sg13g2_mux2_1  _2017_
timestamp 1747056038
transform -1 0 13728 0 1 21924
box -48 -56 1008 834
use sg13g2_o21ai_1  _2018_
timestamp 1747056038
transform -1 0 17376 0 -1 21924
box -48 -56 538 834
use sg13g2_tiehi  _2019__26
timestamp 1747056038
transform -1 0 30336 0 1 24948
box -48 -56 432 834
use sg13g2_dfrbp_1  _2019_
timestamp 1747056038
transform -1 0 29664 0 1 21924
box -60 -56 2556 834
use sg13g2_tiehi  _2020__18
timestamp 1747056038
transform -1 0 30528 0 -1 24948
box -48 -56 432 834
use sg13g2_dfrbp_1  _2020_
timestamp 1747056038
transform 1 0 26016 0 -1 24948
box -60 -56 2556 834
use sg13g2_tiehi  _2021__58
timestamp 1747056038
transform -1 0 29760 0 -1 24948
box -48 -56 432 834
use sg13g2_dfrbp_1  _2021_
timestamp 1747056038
transform -1 0 26688 0 -1 23436
box -60 -56 2556 834
use sg13g2_tiehi  _2022__57
timestamp 1747056038
transform -1 0 30912 0 1 21924
box -48 -56 432 834
use sg13g2_dfrbp_1  _2022_
timestamp 1747056038
transform -1 0 27936 0 -1 21924
box -60 -56 2556 834
use sg13g2_dfrbp_1  _2023_
timestamp 1747056038
transform -1 0 29664 0 1 20412
box -60 -56 2556 834
use sg13g2_tiehi  _2023__56
timestamp 1747056038
transform -1 0 29856 0 -1 20412
box -48 -56 432 834
use sg13g2_tiehi  _2024__55
timestamp 1747056038
transform -1 0 21312 0 -1 20412
box -48 -56 432 834
use sg13g2_dfrbp_1  _2024_
timestamp 1747056038
transform 1 0 18432 0 -1 18900
box -60 -56 2556 834
use sg13g2_dfrbp_1  _2025_
timestamp 1747056038
transform 1 0 21408 0 -1 12852
box -60 -56 2556 834
use sg13g2_tiehi  _2025__54
timestamp 1747056038
transform -1 0 28416 0 1 11340
box -48 -56 432 834
use sg13g2_tiehi  _2026__53
timestamp 1747056038
transform 1 0 19104 0 -1 11340
box -48 -56 432 834
use sg13g2_dfrbp_1  _2026_
timestamp 1747056038
transform 1 0 19488 0 1 9828
box -60 -56 2556 834
use sg13g2_dfrbp_1  _2027_
timestamp 1747056038
transform 1 0 20736 0 1 11340
box -60 -56 2556 834
use sg13g2_tiehi  _2027__52
timestamp 1747056038
transform -1 0 22176 0 1 5292
box -48 -56 432 834
use sg13g2_dfrbp_1  _2028_
timestamp 1747056038
transform -1 0 28032 0 1 12852
box -60 -56 2556 834
use sg13g2_tiehi  _2028__51
timestamp 1747056038
transform -1 0 28800 0 -1 12852
box -48 -56 432 834
use sg13g2_dfrbp_1  _2029_
timestamp 1747056038
transform 1 0 24576 0 1 14364
box -60 -56 2556 834
use sg13g2_tiehi  _2029__50
timestamp 1747056038
transform -1 0 29952 0 -1 14364
box -48 -56 432 834
use sg13g2_tiehi  _2030__49
timestamp 1747056038
transform -1 0 29184 0 -1 12852
box -48 -56 432 834
use sg13g2_dfrbp_1  _2030_
timestamp 1747056038
transform -1 0 27552 0 1 11340
box -60 -56 2556 834
use sg13g2_dfrbp_1  _2031_
timestamp 1747056038
transform -1 0 27456 0 -1 11340
box -60 -56 2556 834
use sg13g2_tiehi  _2031__48
timestamp 1747056038
transform -1 0 27456 0 1 9828
box -48 -56 432 834
use sg13g2_tiehi  _2032__47
timestamp 1747056038
transform -1 0 29376 0 1 15876
box -48 -56 432 834
use sg13g2_dfrbp_1  _2032_
timestamp 1747056038
transform -1 0 28320 0 -1 15876
box -60 -56 2556 834
use sg13g2_tiehi  _2033__46
timestamp 1747056038
transform -1 0 27936 0 1 17388
box -48 -56 432 834
use sg13g2_dfrbp_1  _2033_
timestamp 1747056038
transform -1 0 28224 0 -1 17388
box -60 -56 2556 834
use sg13g2_dfrbp_1  _2034_
timestamp 1747056038
transform 1 0 576 0 -1 24948
box -60 -56 2556 834
use sg13g2_tiehi  _2034__45
timestamp 1747056038
transform -1 0 19776 0 1 14364
box -48 -56 432 834
use sg13g2_dfrbp_1  _2035_
timestamp 1747056038
transform 1 0 576 0 -1 23436
box -60 -56 2556 834
use sg13g2_tiehi  _2035__43
timestamp 1747056038
transform -1 0 30240 0 -1 20412
box -48 -56 432 834
use sg13g2_dfrbp_1  _2036_
timestamp 1747056038
transform -1 0 3072 0 1 14364
box -60 -56 2556 834
use sg13g2_tiehi  _2036__41
timestamp 1747056038
transform -1 0 2400 0 -1 14364
box -48 -56 432 834
use sg13g2_dfrbp_1  _2037_
timestamp 1747056038
transform 1 0 864 0 1 8316
box -60 -56 2556 834
use sg13g2_tiehi  _2037__39
timestamp 1747056038
transform -1 0 2880 0 -1 6804
box -48 -56 432 834
use sg13g2_dfrbp_1  _2038_
timestamp 1747056038
transform 1 0 3648 0 -1 6804
box -60 -56 2556 834
use sg13g2_tiehi  _2038__37
timestamp 1747056038
transform -1 0 4992 0 1 5292
box -48 -56 432 834
use sg13g2_dfrbp_1  _2039_
timestamp 1747056038
transform 1 0 6432 0 1 5292
box -60 -56 2556 834
use sg13g2_tiehi  _2039__35
timestamp 1747056038
transform -1 0 7872 0 -1 5292
box -48 -56 432 834
use sg13g2_dfrbp_1  _2040_
timestamp 1747056038
transform 1 0 10176 0 1 5292
box -60 -56 2556 834
use sg13g2_tiehi  _2040__33
timestamp 1747056038
transform -1 0 11424 0 -1 5292
box -48 -56 432 834
use sg13g2_dfrbp_1  _2041_
timestamp 1747056038
transform 1 0 13728 0 1 5292
box -60 -56 2556 834
use sg13g2_tiehi  _2041__31
timestamp 1747056038
transform -1 0 15360 0 -1 5292
box -48 -56 432 834
use sg13g2_dfrbp_1  _2042_
timestamp 1747056038
transform -1 0 19392 0 1 5292
box -60 -56 2556 834
use sg13g2_tiehi  _2042__29
timestamp 1747056038
transform 1 0 17952 0 -1 5292
box -48 -56 432 834
use sg13g2_dfrbp_1  _2043_
timestamp 1747056038
transform 1 0 20256 0 -1 6804
box -60 -56 2556 834
use sg13g2_tiehi  _2043__27
timestamp 1747056038
transform -1 0 21888 0 -1 5292
box -48 -56 432 834
use sg13g2_tiehi  _2044__25
timestamp 1747056038
transform -1 0 26304 0 -1 6804
box -48 -56 432 834
use sg13g2_dfrbp_1  _2044_
timestamp 1747056038
transform 1 0 22272 0 1 5292
box -60 -56 2556 834
use sg13g2_tiehi  _2045__23
timestamp 1747056038
transform -1 0 27456 0 -1 8316
box -48 -56 432 834
use sg13g2_dfrbp_1  _2045_
timestamp 1747056038
transform 1 0 23712 0 1 6804
box -60 -56 2556 834
use sg13g2_tiehi  _2046__21
timestamp 1747056038
transform -1 0 30720 0 -1 27972
box -48 -56 432 834
use sg13g2_dfrbp_1  _2046_
timestamp 1747056038
transform -1 0 7296 0 1 24948
box -60 -56 2556 834
use sg13g2_tiehi  _2047__20
timestamp 1747056038
transform -1 0 31104 0 1 24948
box -48 -56 432 834
use sg13g2_dfrbp_1  _2047_
timestamp 1747056038
transform -1 0 27840 0 1 24948
box -60 -56 2556 834
use sg13g2_tiehi  _2048__19
timestamp 1747056038
transform 1 0 3648 0 1 26460
box -48 -56 432 834
use sg13g2_dfrbp_1  _2048_
timestamp 1747056038
transform -1 0 11904 0 -1 24948
box -60 -56 2556 834
use sg13g2_dfrbp_1  _2049_
timestamp 1747056038
transform -1 0 15264 0 1 23436
box -60 -56 2556 834
use sg13g2_tiehi  _2049__17
timestamp 1747056038
transform 1 0 8544 0 -1 23436
box -48 -56 432 834
use sg13g2_tiehi  _2050__73
timestamp 1747056038
transform -1 0 29568 0 -1 23436
box -48 -56 432 834
use sg13g2_dfrbp_1  _2050_
timestamp 1747056038
transform 1 0 18720 0 1 21924
box -60 -56 2556 834
use sg13g2_tiehi  _2051__72
timestamp 1747056038
transform -1 0 31104 0 -1 23436
box -48 -56 432 834
use sg13g2_dfrbp_1  _2051_
timestamp 1747056038
transform 1 0 21984 0 1 21924
box -60 -56 2556 834
use sg13g2_dfrbp_1  _2052_
timestamp 1747056038
transform -1 0 28128 0 -1 20412
box -60 -56 2556 834
use sg13g2_tiehi  _2052__71
timestamp 1747056038
transform -1 0 28512 0 -1 18900
box -48 -56 432 834
use sg13g2_tiehi  _2053__70
timestamp 1747056038
transform -1 0 30720 0 -1 23436
box -48 -56 432 834
use sg13g2_dfrbp_1  _2053_
timestamp 1747056038
transform 1 0 21024 0 -1 21924
box -60 -56 2556 834
use sg13g2_tiehi  _2054__69
timestamp 1747056038
transform -1 0 30144 0 1 14364
box -48 -56 432 834
use sg13g2_dfrbp_1  _2054_
timestamp 1747056038
transform 1 0 27072 0 -1 14364
box -60 -56 2556 834
use sg13g2_dfrbp_1  _2055_
timestamp 1747056038
transform 1 0 4896 0 1 26460
box -60 -56 2556 834
use sg13g2_tiehi  _2055__68
timestamp 1747056038
transform -1 0 31200 0 1 20412
box -48 -56 432 834
use sg13g2_dfrbp_1  _2056_
timestamp 1747056038
transform 1 0 6816 0 -1 27972
box -60 -56 2556 834
use sg13g2_tiehi  _2056__66
timestamp 1747056038
transform -1 0 31296 0 -1 24948
box -48 -56 432 834
use sg13g2_tiehi  _2057__64
timestamp 1747056038
transform 1 0 3456 0 -1 27972
box -48 -56 432 834
use sg13g2_dfrbp_1  _2057_
timestamp 1747056038
transform 1 0 9792 0 1 26460
box -60 -56 2556 834
use sg13g2_dfrbp_1  _2058_
timestamp 1747056038
transform -1 0 16800 0 -1 27972
box -60 -56 2556 834
use sg13g2_tiehi  _2058__62
timestamp 1747056038
transform 1 0 4608 0 -1 27972
box -48 -56 432 834
use sg13g2_tiehi  _2059__60
timestamp 1747056038
transform -1 0 30720 0 1 24948
box -48 -56 432 834
use sg13g2_dfrbp_1  _2059_
timestamp 1747056038
transform -1 0 25632 0 -1 24948
box -60 -56 2556 834
use sg13g2_tiehi  _2060__44
timestamp 1747056038
transform -1 0 30336 0 -1 27972
box -48 -56 432 834
use sg13g2_dfrbp_1  _2060_
timestamp 1747056038
transform -1 0 24864 0 -1 27972
box -60 -56 2556 834
use sg13g2_tiehi  _2061__40
timestamp 1747056038
transform -1 0 31392 0 1 26460
box -48 -56 432 834
use sg13g2_dfrbp_1  _2061_
timestamp 1747056038
transform -1 0 27264 0 -1 26460
box -60 -56 2556 834
use sg13g2_dfrbp_1  _2062_
timestamp 1747056038
transform -1 0 26880 0 1 26460
box -60 -56 2556 834
use sg13g2_tiehi  _2062__36
timestamp 1747056038
transform -1 0 30816 0 -1 21924
box -48 -56 432 834
use sg13g2_dfrbp_1  _2063_
timestamp 1747056038
transform -1 0 22368 0 -1 27972
box -60 -56 2556 834
use sg13g2_tiehi  _2063__32
timestamp 1747056038
transform -1 0 29088 0 1 26460
box -48 -56 432 834
use sg13g2_dfrbp_1  _2064_
timestamp 1747056038
transform -1 0 22368 0 -1 24948
box -60 -56 2556 834
use sg13g2_tiehi  _2064__28
timestamp 1747056038
transform -1 0 29952 0 -1 23436
box -48 -56 432 834
use sg13g2_dfrbp_1  _2065_
timestamp 1747056038
transform -1 0 12384 0 -1 27972
box -60 -56 2556 834
use sg13g2_tiehi  _2065__24
timestamp 1747056038
transform 1 0 1536 0 -1 26460
box -48 -56 432 834
use sg13g2_tiehi  _2066__22
timestamp 1747056038
transform -1 0 31296 0 1 21924
box -48 -56 432 834
use sg13g2_dfrbp_1  _2066_
timestamp 1747056038
transform -1 0 30432 0 -1 21924
box -60 -56 2556 834
use sg13g2_tiehi  _2067__67
timestamp 1747056038
transform -1 0 30912 0 -1 24948
box -48 -56 432 834
use sg13g2_dfrbp_1  _2067_
timestamp 1747056038
transform -1 0 29184 0 -1 23436
box -60 -56 2556 834
use sg13g2_tiehi  _2068__65
timestamp 1747056038
transform 1 0 1152 0 -1 27972
box -48 -56 432 834
use sg13g2_dfrbp_1  _2068_
timestamp 1747056038
transform 1 0 5088 0 -1 24948
box -60 -56 2556 834
use sg13g2_tiehi  _2069__63
timestamp 1747056038
transform 1 0 3264 0 1 26460
box -48 -56 432 834
use sg13g2_dfrbp_1  _2069_
timestamp 1747056038
transform 1 0 9408 0 -1 23436
box -60 -56 2556 834
use sg13g2_tiehi  _2070__61
timestamp 1747056038
transform -1 0 29088 0 1 18900
box -48 -56 432 834
use sg13g2_dfrbp_1  _2070_
timestamp 1747056038
transform 1 0 25248 0 -1 18900
box -60 -56 2556 834
use sg13g2_dfrbp_1  _2071_
timestamp 1747056038
transform 1 0 22752 0 -1 18900
box -60 -56 2556 834
use sg13g2_tiehi  _2071__59
timestamp 1747056038
transform -1 0 27168 0 1 17388
box -48 -56 432 834
use sg13g2_dfrbp_1  _2072_
timestamp 1747056038
transform 1 0 3456 0 1 23436
box -60 -56 2556 834
use sg13g2_tiehi  _2072__42
timestamp 1747056038
transform -1 0 4800 0 1 6804
box -48 -56 432 834
use sg13g2_dfrbp_1  _2073_
timestamp 1747056038
transform 1 0 2784 0 -1 26460
box -60 -56 2556 834
use sg13g2_tiehi  _2073__38
timestamp 1747056038
transform -1 0 20736 0 1 15876
box -48 -56 432 834
use sg13g2_dfrbp_1  _2074_
timestamp 1747056038
transform -1 0 12768 0 1 21924
box -60 -56 2556 834
use sg13g2_tiehi  _2074__34
timestamp 1747056038
transform 1 0 4800 0 1 20412
box -48 -56 432 834
use sg13g2_tiehi  _2075__30
timestamp 1747056038
transform -1 0 29952 0 -1 27972
box -48 -56 432 834
use sg13g2_dfrbp_1  _2075_
timestamp 1747056038
transform 1 0 16800 0 -1 27972
box -60 -56 2556 834
use sg13g2_buf_2  _2141_
timestamp 1747056038
transform 1 0 11232 0 -1 21924
box -48 -56 528 834
use sg13g2_buf_2  _2142_
timestamp 1747056038
transform -1 0 19200 0 1 20412
box -48 -56 528 834
use sg13g2_buf_2  _2143_
timestamp 1747056038
transform -1 0 15168 0 1 21924
box -48 -56 528 834
use sg13g2_buf_2  _2144_
timestamp 1747056038
transform -1 0 18336 0 -1 21924
box -48 -56 528 834
use sg13g2_buf_1  _2145_
timestamp 1747056038
transform -1 0 18720 0 -1 21924
box -48 -56 432 834
use sg13g2_buf_1  _2146_
timestamp 1747056038
transform -1 0 20448 0 -1 23436
box -48 -56 432 834
use sg13g2_buf_2  clkbuf_0_clk
timestamp 1747056038
transform 1 0 16032 0 -1 17388
box -48 -56 528 834
use sg13g2_buf_2  clkbuf_4_0_0_clk
timestamp 1747056038
transform -1 0 8448 0 1 14364
box -48 -56 528 834
use sg13g2_buf_2  clkbuf_4_1_0_clk
timestamp 1747056038
transform 1 0 8640 0 1 17388
box -48 -56 528 834
use sg13g2_buf_2  clkbuf_4_2_0_clk
timestamp 1747056038
transform 1 0 15648 0 1 18900
box -48 -56 528 834
use sg13g2_buf_2  clkbuf_4_3_0_clk
timestamp 1747056038
transform 1 0 12768 0 -1 20412
box -48 -56 528 834
use sg13g2_buf_2  clkbuf_4_4_0_clk
timestamp 1747056038
transform 1 0 5376 0 -1 26460
box -48 -56 528 834
use sg13g2_buf_2  clkbuf_4_5_0_clk
timestamp 1747056038
transform 1 0 5376 0 -1 27972
box -48 -56 528 834
use sg13g2_buf_2  clkbuf_4_6_0_clk
timestamp 1747056038
transform -1 0 16992 0 -1 24948
box -48 -56 528 834
use sg13g2_buf_2  clkbuf_4_7_0_clk
timestamp 1747056038
transform 1 0 12576 0 -1 26460
box -48 -56 528 834
use sg13g2_buf_2  clkbuf_4_8_0_clk
timestamp 1747056038
transform -1 0 22656 0 1 8316
box -48 -56 528 834
use sg13g2_buf_2  clkbuf_4_9_0_clk
timestamp 1747056038
transform -1 0 19968 0 -1 11340
box -48 -56 528 834
use sg13g2_buf_2  clkbuf_4_10_0_clk
timestamp 1747056038
transform 1 0 28224 0 1 12852
box -48 -56 528 834
use sg13g2_buf_2  clkbuf_4_11_0_clk
timestamp 1747056038
transform -1 0 28608 0 1 14364
box -48 -56 528 834
use sg13g2_buf_2  clkbuf_4_12_0_clk
timestamp 1747056038
transform -1 0 27936 0 1 18900
box -48 -56 528 834
use sg13g2_buf_2  clkbuf_4_13_0_clk
timestamp 1747056038
transform -1 0 29184 0 1 23436
box -48 -56 528 834
use sg13g2_buf_2  clkbuf_4_14_0_clk
timestamp 1747056038
transform -1 0 29472 0 -1 20412
box -48 -56 528 834
use sg13g2_buf_2  clkbuf_4_15_0_clk
timestamp 1747056038
transform 1 0 28512 0 -1 24948
box -48 -56 528 834
use sg13g2_inv_1  clkload0
timestamp 1747056038
transform 1 0 13920 0 1 18900
box -48 -56 336 834
use sg13g2_inv_1  clkload1
timestamp 1747056038
transform -1 0 4416 0 -1 23436
box -48 -56 336 834
use sg13g2_inv_1  clkload2
timestamp 1747056038
transform 1 0 14208 0 1 26460
box -48 -56 336 834
use sg13g2_inv_1  clkload3
timestamp 1747056038
transform 1 0 21984 0 1 9828
box -48 -56 336 834
use sg13g2_inv_1  clkload4
timestamp 1747056038
transform 1 0 29184 0 -1 15876
box -48 -56 336 834
use sg13g2_inv_1  clkload5
timestamp 1747056038
transform 1 0 23904 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  clkload6
timestamp 1747056038
transform 1 0 31104 0 -1 23436
box -48 -56 336 834
use sg13g2_tielo  controller_11
timestamp 1747056038
transform -1 0 31296 0 -1 26460
box -48 -56 432 834
use sg13g2_tielo  controller_12
timestamp 1747056038
transform -1 0 20160 0 1 14364
box -48 -56 432 834
use sg13g2_tielo  controller_13
timestamp 1747056038
transform -1 0 8064 0 -1 8316
box -48 -56 432 834
use sg13g2_tielo  controller_14
timestamp 1747056038
transform -1 0 29472 0 1 18900
box -48 -56 432 834
use sg13g2_tielo  controller_15
timestamp 1747056038
transform -1 0 30912 0 -1 26460
box -48 -56 432 834
use sg13g2_tielo  controller_16
timestamp 1747056038
transform -1 0 29856 0 1 18900
box -48 -56 432 834
use sg13g2_tiehi  controller_74
timestamp 1747056038
transform -1 0 28320 0 1 17388
box -48 -56 432 834
use sg13g2_tiehi  controller_75
timestamp 1747056038
transform -1 0 31200 0 -1 21924
box -48 -56 432 834
use sg13g2_buf_2  fanout314
timestamp 1747056038
transform 1 0 14976 0 -1 24948
box -48 -56 528 834
use sg13g2_buf_2  fanout315
timestamp 1747056038
transform -1 0 16704 0 -1 23436
box -48 -56 528 834
use sg13g2_buf_2  fanout316
timestamp 1747056038
transform 1 0 18624 0 -1 11340
box -48 -56 528 834
use sg13g2_buf_2  fanout317
timestamp 1747056038
transform 1 0 18624 0 1 15876
box -48 -56 528 834
use sg13g2_buf_2  fanout318
timestamp 1747056038
transform 1 0 17280 0 -1 17388
box -48 -56 528 834
use sg13g2_buf_2  fanout319
timestamp 1747056038
transform 1 0 21696 0 -1 18900
box -48 -56 528 834
use sg13g2_buf_4  fanout320
timestamp 1747056038
transform 1 0 17952 0 1 11340
box -48 -56 816 834
use sg13g2_buf_2  fanout321
timestamp 1747056038
transform 1 0 18144 0 1 15876
box -48 -56 528 834
use sg13g2_buf_2  fanout322
timestamp 1747056038
transform 1 0 10752 0 -1 11340
box -48 -56 528 834
use sg13g2_buf_4  fanout323
timestamp 1747056038
transform 1 0 11712 0 1 23436
box -48 -56 816 834
use sg13g2_buf_2  fanout324
timestamp 1747056038
transform 1 0 12480 0 -1 18900
box -48 -56 528 834
use sg13g2_buf_2  fanout325
timestamp 1747056038
transform 1 0 16896 0 1 17388
box -48 -56 528 834
use sg13g2_buf_2  fanout326
timestamp 1747056038
transform -1 0 17856 0 1 17388
box -48 -56 528 834
use sg13g2_buf_2  fanout327
timestamp 1747056038
transform -1 0 6240 0 1 14364
box -48 -56 528 834
use sg13g2_buf_2  fanout328
timestamp 1747056038
transform 1 0 576 0 -1 18900
box -48 -56 528 834
use sg13g2_buf_2  fanout329
timestamp 1747056038
transform 1 0 2784 0 1 20412
box -48 -56 528 834
use sg13g2_buf_2  fanout330
timestamp 1747056038
transform 1 0 5184 0 1 20412
box -48 -56 528 834
use sg13g2_buf_2  fanout331
timestamp 1747056038
transform 1 0 15744 0 1 20412
box -48 -56 528 834
use sg13g2_buf_4  fanout332
timestamp 1747056038
transform -1 0 2400 0 -1 21924
box -48 -56 816 834
use sg13g2_buf_2  fanout333
timestamp 1747056038
transform 1 0 672 0 -1 21924
box -48 -56 528 834
use sg13g2_buf_2  fanout334
timestamp 1747056038
transform -1 0 6528 0 -1 23436
box -48 -56 528 834
use sg13g2_buf_4  fanout335
timestamp 1747056038
transform -1 0 14592 0 1 21924
box -48 -56 816 834
use sg13g2_buf_2  fanout336
timestamp 1747056038
transform -1 0 9408 0 1 21924
box -48 -56 528 834
use sg13g2_buf_2  fanout337
timestamp 1747056038
transform -1 0 9792 0 1 15876
box -48 -56 528 834
use sg13g2_buf_1  fanout338
timestamp 1747056038
transform 1 0 8928 0 1 15876
box -48 -56 432 834
use sg13g2_buf_2  fanout339
timestamp 1747056038
transform -1 0 11520 0 1 9828
box -48 -56 528 834
use sg13g2_buf_1  fanout340
timestamp 1747056038
transform 1 0 11232 0 -1 11340
box -48 -56 432 834
use sg13g2_buf_2  fanout341
timestamp 1747056038
transform 1 0 8448 0 1 14364
box -48 -56 528 834
use sg13g2_buf_2  fanout342
timestamp 1747056038
transform 1 0 11808 0 1 12852
box -48 -56 528 834
use sg13g2_buf_1  fanout343
timestamp 1747056038
transform -1 0 12768 0 1 14364
box -48 -56 432 834
use sg13g2_buf_2  fanout344
timestamp 1747056038
transform -1 0 13344 0 1 12852
box -48 -56 528 834
use sg13g2_buf_2  fanout345
timestamp 1747056038
transform -1 0 11232 0 -1 14364
box -48 -56 528 834
use sg13g2_buf_2  fanout346
timestamp 1747056038
transform -1 0 10272 0 -1 21924
box -48 -56 528 834
use sg13g2_buf_2  fanout347
timestamp 1747056038
transform 1 0 4320 0 1 17388
box -48 -56 528 834
use sg13g2_buf_1  fanout348
timestamp 1747056038
transform 1 0 672 0 1 21924
box -48 -56 432 834
use sg13g2_buf_2  fanout349
timestamp 1747056038
transform 1 0 11328 0 1 20412
box -48 -56 528 834
use sg13g2_buf_2  fanout350
timestamp 1747056038
transform -1 0 12768 0 1 20412
box -48 -56 528 834
use sg13g2_buf_2  fanout351
timestamp 1747056038
transform -1 0 12288 0 1 20412
box -48 -56 528 834
use sg13g2_buf_2  fanout352
timestamp 1747056038
transform 1 0 11328 0 1 12852
box -48 -56 528 834
use sg13g2_buf_2  fanout353
timestamp 1747056038
transform -1 0 12096 0 1 18900
box -48 -56 528 834
use sg13g2_buf_2  fanout354
timestamp 1747056038
transform -1 0 11520 0 1 17388
box -48 -56 528 834
use sg13g2_buf_2  fanout355
timestamp 1747056038
transform 1 0 3360 0 -1 12852
box -48 -56 528 834
use sg13g2_buf_2  fanout356
timestamp 1747056038
transform -1 0 10656 0 1 24948
box -48 -56 528 834
use sg13g2_buf_2  fanout357
timestamp 1747056038
transform 1 0 2976 0 1 15876
box -48 -56 528 834
use sg13g2_buf_1  fanout358
timestamp 1747056038
transform 1 0 1344 0 1 26460
box -48 -56 432 834
use sg13g2_buf_2  fanout359
timestamp 1747056038
transform 1 0 8832 0 -1 21924
box -48 -56 528 834
use sg13g2_buf_2  fanout360
timestamp 1747056038
transform -1 0 9792 0 -1 21924
box -48 -56 528 834
use sg13g2_buf_2  fanout361
timestamp 1747056038
transform 1 0 8352 0 -1 21924
box -48 -56 528 834
use sg13g2_buf_2  fanout362
timestamp 1747056038
transform -1 0 10752 0 -1 21924
box -48 -56 528 834
use sg13g2_buf_2  fanout363
timestamp 1747056038
transform 1 0 10272 0 -1 17388
box -48 -56 528 834
use sg13g2_buf_4  fanout364
timestamp 1747056038
transform 1 0 7200 0 1 23436
box -48 -56 816 834
use sg13g2_buf_4  fanout365
timestamp 1747056038
transform 1 0 19584 0 -1 26460
box -48 -56 816 834
use sg13g2_buf_1  fanout366
timestamp 1747056038
transform -1 0 29472 0 1 26460
box -48 -56 432 834
use sg13g2_buf_2  fanout367
timestamp 1747056038
transform 1 0 10752 0 -1 21924
box -48 -56 528 834
use sg13g2_buf_4  fanout368
timestamp 1747056038
transform -1 0 25344 0 1 17388
box -48 -56 816 834
use sg13g2_buf_2  fanout369
timestamp 1747056038
transform 1 0 25344 0 1 17388
box -48 -56 528 834
use sg13g2_buf_4  fanout370
timestamp 1747056038
transform 1 0 11424 0 -1 20412
box -48 -56 816 834
use sg13g2_buf_1  fanout371
timestamp 1747056038
transform -1 0 9504 0 1 20412
box -48 -56 432 834
use sg13g2_buf_2  fanout372
timestamp 1747056038
transform 1 0 9312 0 -1 18900
box -48 -56 528 834
use sg13g2_buf_2  fanout373
timestamp 1747056038
transform -1 0 8640 0 1 17388
box -48 -56 528 834
use sg13g2_buf_1  fanout374
timestamp 1747056038
transform 1 0 576 0 1 26460
box -48 -56 432 834
use sg13g2_buf_2  fanout375
timestamp 1747056038
transform 1 0 17664 0 1 26460
box -48 -56 528 834
use sg13g2_buf_2  fanout376
timestamp 1747056038
transform -1 0 26688 0 -1 27972
box -48 -56 528 834
use sg13g2_buf_1  fanout377
timestamp 1747056038
transform -1 0 31008 0 1 26460
box -48 -56 432 834
use sg13g2_buf_2  fanout378
timestamp 1747056038
transform 1 0 10656 0 -1 26460
box -48 -56 528 834
use sg13g2_buf_2  fanout379
timestamp 1747056038
transform 1 0 9312 0 -1 27972
box -48 -56 528 834
use sg13g2_buf_2  fanout380
timestamp 1747056038
transform 1 0 5856 0 -1 27972
box -48 -56 528 834
use sg13g2_buf_1  fanout381
timestamp 1747056038
transform -1 0 19488 0 1 15876
box -48 -56 432 834
use sg13g2_buf_2  fanout382
timestamp 1747056038
transform 1 0 14880 0 -1 12852
box -48 -56 528 834
use sg13g2_buf_2  fanout383
timestamp 1747056038
transform 1 0 16224 0 1 5292
box -48 -56 528 834
use sg13g2_buf_4  fanout384
timestamp 1747056038
transform -1 0 16224 0 -1 5292
box -48 -56 816 834
use sg13g2_buf_2  fanout385
timestamp 1747056038
transform 1 0 8928 0 -1 5292
box -48 -56 528 834
use sg13g2_buf_2  fanout386
timestamp 1747056038
transform -1 0 9408 0 -1 6804
box -48 -56 528 834
use sg13g2_buf_2  fanout387
timestamp 1747056038
transform 1 0 6336 0 -1 6804
box -48 -56 528 834
use sg13g2_buf_2  fanout388
timestamp 1747056038
transform -1 0 6432 0 1 5292
box -48 -56 528 834
use sg13g2_buf_2  fanout389
timestamp 1747056038
transform 1 0 2400 0 -1 8316
box -48 -56 528 834
use sg13g2_buf_2  fanout390
timestamp 1747056038
transform -1 0 4128 0 -1 8316
box -48 -56 528 834
use sg13g2_buf_2  fanout391
timestamp 1747056038
transform 1 0 768 0 1 11340
box -48 -56 528 834
use sg13g2_buf_2  fanout392
timestamp 1747056038
transform 1 0 1056 0 1 21924
box -48 -56 528 834
use sg13g2_buf_4  fanout393
timestamp 1747056038
transform -1 0 26016 0 -1 9828
box -48 -56 816 834
use sg13g2_buf_1  fanout394
timestamp 1747056038
transform 1 0 26400 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_4  fanout395
timestamp 1747056038
transform 1 0 23616 0 -1 11340
box -48 -56 816 834
use sg13g2_buf_2  fanout396
timestamp 1747056038
transform 1 0 24672 0 1 9828
box -48 -56 528 834
use sg13g2_buf_2  fanout397
timestamp 1747056038
transform 1 0 19392 0 -1 8316
box -48 -56 528 834
use sg13g2_buf_2  fanout398
timestamp 1747056038
transform -1 0 28800 0 -1 15876
box -48 -56 528 834
use sg13g2_buf_2  fanout399
timestamp 1747056038
transform -1 0 26304 0 -1 12852
box -48 -56 528 834
use sg13g2_buf_4  fanout400
timestamp 1747056038
transform 1 0 18240 0 1 12852
box -48 -56 816 834
use sg13g2_buf_4  fanout401
timestamp 1747056038
transform 1 0 11616 0 -1 12852
box -48 -56 816 834
use sg13g2_buf_2  fanout402
timestamp 1747056038
transform -1 0 24864 0 -1 11340
box -48 -56 528 834
use sg13g2_buf_4  fanout403
timestamp 1747056038
transform 1 0 21984 0 -1 9828
box -48 -56 816 834
use sg13g2_buf_2  fanout404
timestamp 1747056038
transform -1 0 23616 0 -1 11340
box -48 -56 528 834
use sg13g2_buf_2  fanout405
timestamp 1747056038
transform 1 0 2496 0 1 11340
box -48 -56 528 834
use sg13g2_buf_2  fanout406
timestamp 1747056038
transform 1 0 10656 0 -1 12852
box -48 -56 528 834
use sg13g2_buf_2  fanout407
timestamp 1747056038
transform 1 0 23232 0 1 11340
box -48 -56 528 834
use sg13g2_buf_4  fanout408
timestamp 1747056038
transform -1 0 21696 0 -1 18900
box -48 -56 816 834
use sg13g2_buf_1  fanout409
timestamp 1747056038
transform -1 0 20928 0 1 17388
box -48 -56 432 834
use sg13g2_buf_2  fanout410
timestamp 1747056038
transform 1 0 960 0 -1 26460
box -48 -56 528 834
use sg13g2_buf_4  fanout411
timestamp 1747056038
transform 1 0 12768 0 -1 23436
box -48 -56 816 834
use sg13g2_buf_2  fanout412
timestamp 1747056038
transform -1 0 24960 0 -1 21924
box -48 -56 528 834
use sg13g2_buf_2  fanout413
timestamp 1747056038
transform -1 0 24096 0 1 20412
box -48 -56 528 834
use sg13g2_buf_2  fanout414
timestamp 1747056038
transform 1 0 22848 0 1 17388
box -48 -56 528 834
use sg13g2_buf_2  fanout415
timestamp 1747056038
transform -1 0 19680 0 1 20412
box -48 -56 528 834
use sg13g2_buf_2  fanout416
timestamp 1747056038
transform 1 0 18240 0 1 21924
box -48 -56 528 834
use sg13g2_buf_4  fanout417
timestamp 1747056038
transform 1 0 19296 0 -1 21924
box -48 -56 816 834
use sg13g2_buf_4  fanout418
timestamp 1747056038
transform 1 0 22848 0 1 20412
box -48 -56 816 834
use sg13g2_decap_8  FILLER_0_0
timestamp 1747056097
transform 1 0 576 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_7
timestamp 1747056097
transform 1 0 1248 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_14
timestamp 1747056097
transform 1 0 1920 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_21
timestamp 1747056097
transform 1 0 2592 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_28
timestamp 1747056097
transform 1 0 3264 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_35
timestamp 1747056097
transform 1 0 3936 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_42
timestamp 1747056097
transform 1 0 4608 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_49
timestamp 1747056097
transform 1 0 5280 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_56
timestamp 1747056097
transform 1 0 5952 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_63
timestamp 1747056097
transform 1 0 6624 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_70
timestamp 1747056097
transform 1 0 7296 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_77
timestamp 1747056097
transform 1 0 7968 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_84
timestamp 1747056097
transform 1 0 8640 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_91
timestamp 1747056097
transform 1 0 9312 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_98
timestamp 1747056097
transform 1 0 9984 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_105
timestamp 1747056097
transform 1 0 10656 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_112
timestamp 1747056097
transform 1 0 11328 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_119
timestamp 1747056097
transform 1 0 12000 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_126
timestamp 1747056097
transform 1 0 12672 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_133
timestamp 1747056097
transform 1 0 13344 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_140
timestamp 1747056097
transform 1 0 14016 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_147
timestamp 1747056097
transform 1 0 14688 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_154
timestamp 1747056097
transform 1 0 15360 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_161
timestamp 1747056097
transform 1 0 16032 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_168
timestamp 1747056097
transform 1 0 16704 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_175
timestamp 1747056097
transform 1 0 17376 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_182
timestamp 1747056097
transform 1 0 18048 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_189
timestamp 1747056097
transform 1 0 18720 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_196
timestamp 1747056097
transform 1 0 19392 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_203
timestamp 1747056097
transform 1 0 20064 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_210
timestamp 1747056097
transform 1 0 20736 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_217
timestamp 1747056097
transform 1 0 21408 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_224
timestamp 1747056097
transform 1 0 22080 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_231
timestamp 1747056097
transform 1 0 22752 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_238
timestamp 1747056097
transform 1 0 23424 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_245
timestamp 1747056097
transform 1 0 24096 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_252
timestamp 1747056097
transform 1 0 24768 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_259
timestamp 1747056097
transform 1 0 25440 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_266
timestamp 1747056097
transform 1 0 26112 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_273
timestamp 1747056097
transform 1 0 26784 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_280
timestamp 1747056097
transform 1 0 27456 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_287
timestamp 1747056097
transform 1 0 28128 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_294
timestamp 1747056097
transform 1 0 28800 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_301
timestamp 1747056097
transform 1 0 29472 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_308
timestamp 1747056097
transform 1 0 30144 0 1 756
box -48 -56 720 834
use sg13g2_decap_4  FILLER_0_315
timestamp 1747056038
transform 1 0 30816 0 1 756
box -48 -56 432 834
use sg13g2_fill_2  FILLER_0_319
timestamp 1747056038
transform 1 0 31200 0 1 756
box -48 -56 240 834
use sg13g2_decap_8  FILLER_1_0
timestamp 1747056097
transform 1 0 576 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_7
timestamp 1747056097
transform 1 0 1248 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_14
timestamp 1747056097
transform 1 0 1920 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_21
timestamp 1747056097
transform 1 0 2592 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_28
timestamp 1747056097
transform 1 0 3264 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_35
timestamp 1747056097
transform 1 0 3936 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_42
timestamp 1747056097
transform 1 0 4608 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_49
timestamp 1747056097
transform 1 0 5280 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_56
timestamp 1747056097
transform 1 0 5952 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_63
timestamp 1747056097
transform 1 0 6624 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_70
timestamp 1747056097
transform 1 0 7296 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_77
timestamp 1747056097
transform 1 0 7968 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_84
timestamp 1747056097
transform 1 0 8640 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_91
timestamp 1747056097
transform 1 0 9312 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_98
timestamp 1747056097
transform 1 0 9984 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_105
timestamp 1747056097
transform 1 0 10656 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_112
timestamp 1747056097
transform 1 0 11328 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_119
timestamp 1747056097
transform 1 0 12000 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_126
timestamp 1747056097
transform 1 0 12672 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_133
timestamp 1747056097
transform 1 0 13344 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_140
timestamp 1747056097
transform 1 0 14016 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_147
timestamp 1747056097
transform 1 0 14688 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_154
timestamp 1747056097
transform 1 0 15360 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_161
timestamp 1747056097
transform 1 0 16032 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_168
timestamp 1747056097
transform 1 0 16704 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_175
timestamp 1747056097
transform 1 0 17376 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_182
timestamp 1747056097
transform 1 0 18048 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_189
timestamp 1747056097
transform 1 0 18720 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_196
timestamp 1747056097
transform 1 0 19392 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_203
timestamp 1747056097
transform 1 0 20064 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_210
timestamp 1747056097
transform 1 0 20736 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_217
timestamp 1747056097
transform 1 0 21408 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_224
timestamp 1747056097
transform 1 0 22080 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_231
timestamp 1747056097
transform 1 0 22752 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_238
timestamp 1747056097
transform 1 0 23424 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_245
timestamp 1747056097
transform 1 0 24096 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_252
timestamp 1747056097
transform 1 0 24768 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_259
timestamp 1747056097
transform 1 0 25440 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_266
timestamp 1747056097
transform 1 0 26112 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_273
timestamp 1747056097
transform 1 0 26784 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_280
timestamp 1747056097
transform 1 0 27456 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_287
timestamp 1747056097
transform 1 0 28128 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_294
timestamp 1747056097
transform 1 0 28800 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_301
timestamp 1747056097
transform 1 0 29472 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_308
timestamp 1747056097
transform 1 0 30144 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_1_315
timestamp 1747056038
transform 1 0 30816 0 -1 2268
box -48 -56 432 834
use sg13g2_fill_2  FILLER_1_319
timestamp 1747056038
transform 1 0 31200 0 -1 2268
box -48 -56 240 834
use sg13g2_decap_8  FILLER_2_0
timestamp 1747056097
transform 1 0 576 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_7
timestamp 1747056097
transform 1 0 1248 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_14
timestamp 1747056097
transform 1 0 1920 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_21
timestamp 1747056097
transform 1 0 2592 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_28
timestamp 1747056097
transform 1 0 3264 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_35
timestamp 1747056097
transform 1 0 3936 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_42
timestamp 1747056097
transform 1 0 4608 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_49
timestamp 1747056097
transform 1 0 5280 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_56
timestamp 1747056097
transform 1 0 5952 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_63
timestamp 1747056097
transform 1 0 6624 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_70
timestamp 1747056097
transform 1 0 7296 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_77
timestamp 1747056097
transform 1 0 7968 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_84
timestamp 1747056097
transform 1 0 8640 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_91
timestamp 1747056097
transform 1 0 9312 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_98
timestamp 1747056097
transform 1 0 9984 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_105
timestamp 1747056097
transform 1 0 10656 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_112
timestamp 1747056097
transform 1 0 11328 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_119
timestamp 1747056097
transform 1 0 12000 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_126
timestamp 1747056097
transform 1 0 12672 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_133
timestamp 1747056097
transform 1 0 13344 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_140
timestamp 1747056097
transform 1 0 14016 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_147
timestamp 1747056097
transform 1 0 14688 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_154
timestamp 1747056097
transform 1 0 15360 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_161
timestamp 1747056097
transform 1 0 16032 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_168
timestamp 1747056097
transform 1 0 16704 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_175
timestamp 1747056097
transform 1 0 17376 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_182
timestamp 1747056097
transform 1 0 18048 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_189
timestamp 1747056097
transform 1 0 18720 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_196
timestamp 1747056097
transform 1 0 19392 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_203
timestamp 1747056097
transform 1 0 20064 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_210
timestamp 1747056097
transform 1 0 20736 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_217
timestamp 1747056097
transform 1 0 21408 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_224
timestamp 1747056097
transform 1 0 22080 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_231
timestamp 1747056097
transform 1 0 22752 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_238
timestamp 1747056097
transform 1 0 23424 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_245
timestamp 1747056097
transform 1 0 24096 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_252
timestamp 1747056097
transform 1 0 24768 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_259
timestamp 1747056097
transform 1 0 25440 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_266
timestamp 1747056097
transform 1 0 26112 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_273
timestamp 1747056097
transform 1 0 26784 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_280
timestamp 1747056097
transform 1 0 27456 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_287
timestamp 1747056097
transform 1 0 28128 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_294
timestamp 1747056097
transform 1 0 28800 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_301
timestamp 1747056097
transform 1 0 29472 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_308
timestamp 1747056097
transform 1 0 30144 0 1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_315
timestamp 1747056038
transform 1 0 30816 0 1 2268
box -48 -56 432 834
use sg13g2_fill_2  FILLER_2_319
timestamp 1747056038
transform 1 0 31200 0 1 2268
box -48 -56 240 834
use sg13g2_decap_8  FILLER_3_0
timestamp 1747056097
transform 1 0 576 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_7
timestamp 1747056097
transform 1 0 1248 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_14
timestamp 1747056097
transform 1 0 1920 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_21
timestamp 1747056097
transform 1 0 2592 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_28
timestamp 1747056097
transform 1 0 3264 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_35
timestamp 1747056097
transform 1 0 3936 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_42
timestamp 1747056097
transform 1 0 4608 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_49
timestamp 1747056097
transform 1 0 5280 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_56
timestamp 1747056097
transform 1 0 5952 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_63
timestamp 1747056097
transform 1 0 6624 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_70
timestamp 1747056097
transform 1 0 7296 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_77
timestamp 1747056097
transform 1 0 7968 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_84
timestamp 1747056097
transform 1 0 8640 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_91
timestamp 1747056097
transform 1 0 9312 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_98
timestamp 1747056097
transform 1 0 9984 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_105
timestamp 1747056097
transform 1 0 10656 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_112
timestamp 1747056097
transform 1 0 11328 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_119
timestamp 1747056097
transform 1 0 12000 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_126
timestamp 1747056097
transform 1 0 12672 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_133
timestamp 1747056097
transform 1 0 13344 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_140
timestamp 1747056097
transform 1 0 14016 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_147
timestamp 1747056097
transform 1 0 14688 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_154
timestamp 1747056097
transform 1 0 15360 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_161
timestamp 1747056097
transform 1 0 16032 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_168
timestamp 1747056097
transform 1 0 16704 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_175
timestamp 1747056097
transform 1 0 17376 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_182
timestamp 1747056097
transform 1 0 18048 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_189
timestamp 1747056097
transform 1 0 18720 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_196
timestamp 1747056097
transform 1 0 19392 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_203
timestamp 1747056097
transform 1 0 20064 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_210
timestamp 1747056097
transform 1 0 20736 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_217
timestamp 1747056097
transform 1 0 21408 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_224
timestamp 1747056097
transform 1 0 22080 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_231
timestamp 1747056097
transform 1 0 22752 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_238
timestamp 1747056097
transform 1 0 23424 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_245
timestamp 1747056097
transform 1 0 24096 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_252
timestamp 1747056097
transform 1 0 24768 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_259
timestamp 1747056097
transform 1 0 25440 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_266
timestamp 1747056097
transform 1 0 26112 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_273
timestamp 1747056097
transform 1 0 26784 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_280
timestamp 1747056097
transform 1 0 27456 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_287
timestamp 1747056097
transform 1 0 28128 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_294
timestamp 1747056097
transform 1 0 28800 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_301
timestamp 1747056097
transform 1 0 29472 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_308
timestamp 1747056097
transform 1 0 30144 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_315
timestamp 1747056038
transform 1 0 30816 0 -1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_3_319
timestamp 1747056038
transform 1 0 31200 0 -1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_4_0
timestamp 1747056097
transform 1 0 576 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_7
timestamp 1747056097
transform 1 0 1248 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_14
timestamp 1747056097
transform 1 0 1920 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_21
timestamp 1747056097
transform 1 0 2592 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_28
timestamp 1747056097
transform 1 0 3264 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_35
timestamp 1747056097
transform 1 0 3936 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_42
timestamp 1747056097
transform 1 0 4608 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_49
timestamp 1747056097
transform 1 0 5280 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_56
timestamp 1747056097
transform 1 0 5952 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_63
timestamp 1747056097
transform 1 0 6624 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_70
timestamp 1747056097
transform 1 0 7296 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_77
timestamp 1747056097
transform 1 0 7968 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_84
timestamp 1747056097
transform 1 0 8640 0 1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_91
timestamp 1747056038
transform 1 0 9312 0 1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_4_95
timestamp 1747056038
transform 1 0 9696 0 1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_4_101
timestamp 1747056097
transform 1 0 10272 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_108
timestamp 1747056097
transform 1 0 10944 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_115
timestamp 1747056097
transform 1 0 11616 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_122
timestamp 1747056097
transform 1 0 12288 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_129
timestamp 1747056097
transform 1 0 12960 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_136
timestamp 1747056097
transform 1 0 13632 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_143
timestamp 1747056097
transform 1 0 14304 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_150
timestamp 1747056097
transform 1 0 14976 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_157
timestamp 1747056097
transform 1 0 15648 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_164
timestamp 1747056097
transform 1 0 16320 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_171
timestamp 1747056097
transform 1 0 16992 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_178
timestamp 1747056097
transform 1 0 17664 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_185
timestamp 1747056097
transform 1 0 18336 0 1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_192
timestamp 1747056038
transform 1 0 19008 0 1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_4_196
timestamp 1747056038
transform 1 0 19392 0 1 3780
box -48 -56 240 834
use sg13g2_fill_2  FILLER_4_202
timestamp 1747056038
transform 1 0 19968 0 1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_204
timestamp 1747056097
transform 1 0 20160 0 1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_212
timestamp 1747056097
transform 1 0 20928 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_219
timestamp 1747056097
transform 1 0 21600 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_226
timestamp 1747056097
transform 1 0 22272 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_233
timestamp 1747056097
transform 1 0 22944 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_240
timestamp 1747056097
transform 1 0 23616 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_247
timestamp 1747056097
transform 1 0 24288 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_254
timestamp 1747056097
transform 1 0 24960 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_261
timestamp 1747056097
transform 1 0 25632 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_268
timestamp 1747056097
transform 1 0 26304 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_275
timestamp 1747056097
transform 1 0 26976 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_282
timestamp 1747056097
transform 1 0 27648 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_289
timestamp 1747056097
transform 1 0 28320 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_296
timestamp 1747056097
transform 1 0 28992 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_303
timestamp 1747056097
transform 1 0 29664 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_310
timestamp 1747056097
transform 1 0 30336 0 1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_317
timestamp 1747056038
transform 1 0 31008 0 1 3780
box -48 -56 432 834
use sg13g2_decap_8  FILLER_5_0
timestamp 1747056097
transform 1 0 576 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_7
timestamp 1747056097
transform 1 0 1248 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_14
timestamp 1747056097
transform 1 0 1920 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_21
timestamp 1747056097
transform 1 0 2592 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_28
timestamp 1747056097
transform 1 0 3264 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_35
timestamp 1747056097
transform 1 0 3936 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_42
timestamp 1747056097
transform 1 0 4608 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_49
timestamp 1747056097
transform 1 0 5280 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_56
timestamp 1747056038
transform 1 0 5952 0 -1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_5_61
timestamp 1747056097
transform 1 0 6432 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_68
timestamp 1747056038
transform 1 0 7104 0 -1 5292
box -48 -56 432 834
use sg13g2_decap_8  FILLER_5_76
timestamp 1747056097
transform 1 0 7872 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_83
timestamp 1747056038
transform 1 0 8544 0 -1 5292
box -48 -56 432 834
use sg13g2_fill_1  FILLER_5_100
timestamp 1747056097
transform 1 0 10176 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_4  FILLER_5_122
timestamp 1747056038
transform 1 0 12288 0 -1 5292
box -48 -56 432 834
use sg13g2_fill_1  FILLER_5_154
timestamp 1747056097
transform 1 0 15360 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_172
timestamp 1747056097
transform 1 0 17088 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_179
timestamp 1747056038
transform 1 0 17760 0 -1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_5_185
timestamp 1747056097
transform 1 0 18336 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_222
timestamp 1747056097
transform 1 0 21888 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_247
timestamp 1747056097
transform 1 0 24288 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_254
timestamp 1747056097
transform 1 0 24960 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_261
timestamp 1747056097
transform 1 0 25632 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_268
timestamp 1747056097
transform 1 0 26304 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_275
timestamp 1747056097
transform 1 0 26976 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_282
timestamp 1747056097
transform 1 0 27648 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_289
timestamp 1747056097
transform 1 0 28320 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_296
timestamp 1747056097
transform 1 0 28992 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_303
timestamp 1747056097
transform 1 0 29664 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_310
timestamp 1747056097
transform 1 0 30336 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_317
timestamp 1747056038
transform 1 0 31008 0 -1 5292
box -48 -56 432 834
use sg13g2_decap_8  FILLER_6_0
timestamp 1747056097
transform 1 0 576 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_7
timestamp 1747056097
transform 1 0 1248 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_14
timestamp 1747056097
transform 1 0 1920 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_21
timestamp 1747056097
transform 1 0 2592 0 1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_28
timestamp 1747056038
transform 1 0 3264 0 1 5292
box -48 -56 240 834
use sg13g2_fill_2  FILLER_6_39
timestamp 1747056038
transform 1 0 4320 0 1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_41
timestamp 1747056097
transform 1 0 4512 0 1 5292
box -48 -56 144 834
use sg13g2_fill_2  FILLER_6_87
timestamp 1747056038
transform 1 0 8928 0 1 5292
box -48 -56 240 834
use sg13g2_fill_2  FILLER_6_98
timestamp 1747056038
transform 1 0 9984 0 1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_126
timestamp 1747056097
transform 1 0 12672 0 1 5292
box -48 -56 144 834
use sg13g2_fill_2  FILLER_6_134
timestamp 1747056038
transform 1 0 13440 0 1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_136
timestamp 1747056097
transform 1 0 13632 0 1 5292
box -48 -56 144 834
use sg13g2_fill_2  FILLER_6_168
timestamp 1747056038
transform 1 0 16704 0 1 5292
box -48 -56 240 834
use sg13g2_fill_2  FILLER_6_219
timestamp 1747056038
transform 1 0 21600 0 1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_225
timestamp 1747056097
transform 1 0 22176 0 1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_257
timestamp 1747056097
transform 1 0 25248 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_264
timestamp 1747056097
transform 1 0 25920 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_271
timestamp 1747056097
transform 1 0 26592 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_278
timestamp 1747056097
transform 1 0 27264 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_285
timestamp 1747056097
transform 1 0 27936 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_292
timestamp 1747056097
transform 1 0 28608 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_299
timestamp 1747056097
transform 1 0 29280 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_306
timestamp 1747056097
transform 1 0 29952 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_313
timestamp 1747056097
transform 1 0 30624 0 1 5292
box -48 -56 720 834
use sg13g2_fill_1  FILLER_6_320
timestamp 1747056097
transform 1 0 31296 0 1 5292
box -48 -56 144 834
use sg13g2_decap_4  FILLER_7_0
timestamp 1747056038
transform 1 0 576 0 -1 6804
box -48 -56 432 834
use sg13g2_fill_1  FILLER_7_4
timestamp 1747056097
transform 1 0 960 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_7_13
timestamp 1747056038
transform 1 0 1824 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_15
timestamp 1747056097
transform 1 0 2016 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_7_58
timestamp 1747056038
transform 1 0 6144 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_78
timestamp 1747056097
transform 1 0 8064 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_7_121
timestamp 1747056038
transform 1 0 12192 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_2  FILLER_7_154
timestamp 1747056038
transform 1 0 15360 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_2  FILLER_7_164
timestamp 1747056038
transform 1 0 16320 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_166
timestamp 1747056097
transform 1 0 16512 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_7_193
timestamp 1747056097
transform 1 0 19104 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_7_198
timestamp 1747056038
transform 1 0 19584 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_2  FILLER_7_231
timestamp 1747056038
transform 1 0 22752 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_233
timestamp 1747056097
transform 1 0 22944 0 -1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_268
timestamp 1747056097
transform 1 0 26304 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_275
timestamp 1747056097
transform 1 0 26976 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_282
timestamp 1747056097
transform 1 0 27648 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_289
timestamp 1747056097
transform 1 0 28320 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_296
timestamp 1747056097
transform 1 0 28992 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_303
timestamp 1747056097
transform 1 0 29664 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_310
timestamp 1747056097
transform 1 0 30336 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_4  FILLER_7_317
timestamp 1747056038
transform 1 0 31008 0 -1 6804
box -48 -56 432 834
use sg13g2_fill_1  FILLER_8_29
timestamp 1747056097
transform 1 0 3360 0 1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_8_61
timestamp 1747056097
transform 1 0 6432 0 1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_8_76
timestamp 1747056038
transform 1 0 7872 0 1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_86
timestamp 1747056097
transform 1 0 8832 0 1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_8_100
timestamp 1747056097
transform 1 0 10176 0 1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_8_127
timestamp 1747056038
transform 1 0 12768 0 1 6804
box -48 -56 240 834
use sg13g2_fill_2  FILLER_8_150
timestamp 1747056038
transform 1 0 14976 0 1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_173
timestamp 1747056097
transform 1 0 17184 0 1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_8_203
timestamp 1747056097
transform 1 0 20064 0 1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_8_238
timestamp 1747056038
transform 1 0 23424 0 1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_240
timestamp 1747056097
transform 1 0 23616 0 1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_276
timestamp 1747056097
transform 1 0 27072 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_283
timestamp 1747056097
transform 1 0 27744 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_290
timestamp 1747056097
transform 1 0 28416 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_297
timestamp 1747056097
transform 1 0 29088 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_304
timestamp 1747056097
transform 1 0 29760 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_311
timestamp 1747056097
transform 1 0 30432 0 1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_8_318
timestamp 1747056038
transform 1 0 31104 0 1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_320
timestamp 1747056097
transform 1 0 31296 0 1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_9_12
timestamp 1747056038
transform 1 0 1728 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_14
timestamp 1747056097
transform 1 0 1920 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_9_67
timestamp 1747056038
transform 1 0 7008 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_2  FILLER_9_127
timestamp 1747056038
transform 1 0 12768 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_129
timestamp 1747056097
transform 1 0 12960 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_9_138
timestamp 1747056038
transform 1 0 13824 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_140
timestamp 1747056097
transform 1 0 14016 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_9_156
timestamp 1747056038
transform 1 0 15552 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_2  FILLER_9_174
timestamp 1747056038
transform 1 0 17280 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_2  FILLER_9_201
timestamp 1747056038
transform 1 0 19872 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_2  FILLER_9_216
timestamp 1747056038
transform 1 0 21312 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_2  FILLER_9_233
timestamp 1747056038
transform 1 0 22944 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_2  FILLER_9_250
timestamp 1747056038
transform 1 0 24576 0 -1 8316
box -48 -56 240 834
use sg13g2_decap_8  FILLER_9_280
timestamp 1747056097
transform 1 0 27456 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_287
timestamp 1747056097
transform 1 0 28128 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_294
timestamp 1747056097
transform 1 0 28800 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_301
timestamp 1747056097
transform 1 0 29472 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_308
timestamp 1747056097
transform 1 0 30144 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_4  FILLER_9_315
timestamp 1747056038
transform 1 0 30816 0 -1 8316
box -48 -56 432 834
use sg13g2_fill_2  FILLER_9_319
timestamp 1747056038
transform 1 0 31200 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_2  FILLER_10_0
timestamp 1747056038
transform 1 0 576 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_2
timestamp 1747056097
transform 1 0 768 0 1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_10_37
timestamp 1747056038
transform 1 0 4128 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_39
timestamp 1747056097
transform 1 0 4320 0 1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_10_119
timestamp 1747056038
transform 1 0 12000 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_121
timestamp 1747056097
transform 1 0 12192 0 1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_10_151
timestamp 1747056038
transform 1 0 15072 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_178
timestamp 1747056097
transform 1 0 17664 0 1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_10_206
timestamp 1747056038
transform 1 0 20352 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_235
timestamp 1747056097
transform 1 0 23136 0 1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_281
timestamp 1747056097
transform 1 0 27552 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_288
timestamp 1747056097
transform 1 0 28224 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_295
timestamp 1747056097
transform 1 0 28896 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_302
timestamp 1747056097
transform 1 0 29568 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_309
timestamp 1747056097
transform 1 0 30240 0 1 8316
box -48 -56 720 834
use sg13g2_decap_4  FILLER_10_316
timestamp 1747056038
transform 1 0 30912 0 1 8316
box -48 -56 432 834
use sg13g2_fill_1  FILLER_10_320
timestamp 1747056097
transform 1 0 31296 0 1 8316
box -48 -56 144 834
use sg13g2_fill_1  FILLER_11_7
timestamp 1747056097
transform 1 0 1248 0 -1 9828
box -48 -56 144 834
use sg13g2_fill_2  FILLER_11_27
timestamp 1747056038
transform 1 0 3168 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_53
timestamp 1747056097
transform 1 0 5664 0 -1 9828
box -48 -56 144 834
use sg13g2_fill_2  FILLER_11_75
timestamp 1747056038
transform 1 0 7776 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_2  FILLER_11_82
timestamp 1747056038
transform 1 0 8448 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_94
timestamp 1747056097
transform 1 0 9600 0 -1 9828
box -48 -56 144 834
use sg13g2_fill_2  FILLER_11_100
timestamp 1747056038
transform 1 0 10176 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_107
timestamp 1747056097
transform 1 0 10848 0 -1 9828
box -48 -56 144 834
use sg13g2_fill_1  FILLER_11_135
timestamp 1747056097
transform 1 0 13536 0 -1 9828
box -48 -56 144 834
use sg13g2_fill_1  FILLER_11_157
timestamp 1747056097
transform 1 0 15648 0 -1 9828
box -48 -56 144 834
use sg13g2_fill_1  FILLER_11_188
timestamp 1747056097
transform 1 0 18624 0 -1 9828
box -48 -56 144 834
use sg13g2_fill_2  FILLER_11_221
timestamp 1747056038
transform 1 0 21792 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_247
timestamp 1747056097
transform 1 0 24288 0 -1 9828
box -48 -56 144 834
use sg13g2_fill_1  FILLER_11_256
timestamp 1747056097
transform 1 0 25152 0 -1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_273
timestamp 1747056097
transform 1 0 26784 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_280
timestamp 1747056097
transform 1 0 27456 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_287
timestamp 1747056097
transform 1 0 28128 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_294
timestamp 1747056097
transform 1 0 28800 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_301
timestamp 1747056097
transform 1 0 29472 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_308
timestamp 1747056097
transform 1 0 30144 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_11_315
timestamp 1747056038
transform 1 0 30816 0 -1 9828
box -48 -56 432 834
use sg13g2_fill_2  FILLER_11_319
timestamp 1747056038
transform 1 0 31200 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_12_0
timestamp 1747056097
transform 1 0 576 0 1 9828
box -48 -56 144 834
use sg13g2_fill_1  FILLER_12_33
timestamp 1747056097
transform 1 0 3744 0 1 9828
box -48 -56 144 834
use sg13g2_fill_1  FILLER_12_65
timestamp 1747056097
transform 1 0 6816 0 1 9828
box -48 -56 144 834
use sg13g2_fill_2  FILLER_12_129
timestamp 1747056038
transform 1 0 12960 0 1 9828
box -48 -56 240 834
use sg13g2_fill_2  FILLER_12_195
timestamp 1747056038
transform 1 0 19296 0 1 9828
box -48 -56 240 834
use sg13g2_fill_2  FILLER_12_256
timestamp 1747056038
transform 1 0 25152 0 1 9828
box -48 -56 240 834
use sg13g2_decap_8  FILLER_12_280
timestamp 1747056097
transform 1 0 27456 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_287
timestamp 1747056097
transform 1 0 28128 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_294
timestamp 1747056097
transform 1 0 28800 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_301
timestamp 1747056097
transform 1 0 29472 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_308
timestamp 1747056097
transform 1 0 30144 0 1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_12_315
timestamp 1747056038
transform 1 0 30816 0 1 9828
box -48 -56 432 834
use sg13g2_fill_2  FILLER_12_319
timestamp 1747056038
transform 1 0 31200 0 1 9828
box -48 -56 240 834
use sg13g2_fill_2  FILLER_13_20
timestamp 1747056038
transform 1 0 2496 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_2  FILLER_13_58
timestamp 1747056038
transform 1 0 6144 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_13_95
timestamp 1747056097
transform 1 0 9696 0 -1 11340
box -48 -56 144 834
use sg13g2_fill_1  FILLER_13_124
timestamp 1747056097
transform 1 0 12480 0 -1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_13_154
timestamp 1747056038
transform 1 0 15360 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_13_156
timestamp 1747056097
transform 1 0 15552 0 -1 11340
box -48 -56 144 834
use sg13g2_fill_1  FILLER_13_210
timestamp 1747056097
transform 1 0 20736 0 -1 11340
box -48 -56 144 834
use sg13g2_fill_1  FILLER_13_253
timestamp 1747056097
transform 1 0 24864 0 -1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_13_284
timestamp 1747056097
transform 1 0 27840 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_291
timestamp 1747056097
transform 1 0 28512 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_298
timestamp 1747056097
transform 1 0 29184 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_305
timestamp 1747056097
transform 1 0 29856 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_312
timestamp 1747056097
transform 1 0 30528 0 -1 11340
box -48 -56 720 834
use sg13g2_fill_2  FILLER_13_319
timestamp 1747056038
transform 1 0 31200 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_2  FILLER_14_0
timestamp 1747056038
transform 1 0 576 0 1 11340
box -48 -56 240 834
use sg13g2_fill_2  FILLER_14_35
timestamp 1747056038
transform 1 0 3936 0 1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_14_50
timestamp 1747056097
transform 1 0 5376 0 1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_14_56
timestamp 1747056038
transform 1 0 5952 0 1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_14_124
timestamp 1747056097
transform 1 0 12480 0 1 11340
box -48 -56 144 834
use sg13g2_fill_1  FILLER_14_169
timestamp 1747056097
transform 1 0 16800 0 1 11340
box -48 -56 144 834
use sg13g2_fill_1  FILLER_14_180
timestamp 1747056097
transform 1 0 17856 0 1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_14_198
timestamp 1747056038
transform 1 0 19584 0 1 11340
box -48 -56 240 834
use sg13g2_fill_2  FILLER_14_208
timestamp 1747056038
transform 1 0 20544 0 1 11340
box -48 -56 240 834
use sg13g2_decap_8  FILLER_14_290
timestamp 1747056097
transform 1 0 28416 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_297
timestamp 1747056097
transform 1 0 29088 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_304
timestamp 1747056097
transform 1 0 29760 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_311
timestamp 1747056097
transform 1 0 30432 0 1 11340
box -48 -56 720 834
use sg13g2_fill_2  FILLER_14_318
timestamp 1747056038
transform 1 0 31104 0 1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_14_320
timestamp 1747056097
transform 1 0 31296 0 1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_15_0
timestamp 1747056038
transform 1 0 576 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_2  FILLER_15_27
timestamp 1747056038
transform 1 0 3168 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_15_34
timestamp 1747056097
transform 1 0 3840 0 -1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_15_48
timestamp 1747056038
transform 1 0 5184 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_2  FILLER_15_72
timestamp 1747056038
transform 1 0 7488 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_15_74
timestamp 1747056097
transform 1 0 7680 0 -1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_15_103
timestamp 1747056038
transform 1 0 10464 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_15_123
timestamp 1747056097
transform 1 0 12384 0 -1 12852
box -48 -56 144 834
use sg13g2_fill_1  FILLER_15_132
timestamp 1747056097
transform 1 0 13248 0 -1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_15_146
timestamp 1747056038
transform 1 0 14592 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_15_148
timestamp 1747056097
transform 1 0 14784 0 -1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_15_167
timestamp 1747056038
transform 1 0 16608 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_15_174
timestamp 1747056097
transform 1 0 17280 0 -1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_15_180
timestamp 1747056038
transform 1 0 17856 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_15_182
timestamp 1747056097
transform 1 0 18048 0 -1 12852
box -48 -56 144 834
use sg13g2_fill_1  FILLER_15_207
timestamp 1747056097
transform 1 0 20448 0 -1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_15_268
timestamp 1747056038
transform 1 0 26304 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_15_270
timestamp 1747056097
transform 1 0 26496 0 -1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_15_298
timestamp 1747056097
transform 1 0 29184 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_305
timestamp 1747056097
transform 1 0 29856 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_312
timestamp 1747056097
transform 1 0 30528 0 -1 12852
box -48 -56 720 834
use sg13g2_fill_2  FILLER_15_319
timestamp 1747056038
transform 1 0 31200 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_2  FILLER_16_0
timestamp 1747056038
transform 1 0 576 0 1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_16_2
timestamp 1747056097
transform 1 0 768 0 1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_16_12
timestamp 1747056038
transform 1 0 1728 0 1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_16_14
timestamp 1747056097
transform 1 0 1920 0 1 12852
box -48 -56 144 834
use sg13g2_fill_1  FILLER_16_23
timestamp 1747056097
transform 1 0 2784 0 1 12852
box -48 -56 144 834
use sg13g2_fill_1  FILLER_16_29
timestamp 1747056097
transform 1 0 3360 0 1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_16_35
timestamp 1747056038
transform 1 0 3936 0 1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_16_37
timestamp 1747056097
transform 1 0 4128 0 1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_16_46
timestamp 1747056038
transform 1 0 4992 0 1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_16_68
timestamp 1747056097
transform 1 0 7104 0 1 12852
box -48 -56 144 834
use sg13g2_fill_1  FILLER_16_90
timestamp 1747056097
transform 1 0 9216 0 1 12852
box -48 -56 144 834
use sg13g2_fill_1  FILLER_16_111
timestamp 1747056097
transform 1 0 11232 0 1 12852
box -48 -56 144 834
use sg13g2_fill_1  FILLER_16_127
timestamp 1747056097
transform 1 0 12768 0 1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_16_138
timestamp 1747056038
transform 1 0 13824 0 1 12852
box -48 -56 240 834
use sg13g2_fill_2  FILLER_16_145
timestamp 1747056038
transform 1 0 14496 0 1 12852
box -48 -56 240 834
use sg13g2_fill_2  FILLER_16_167
timestamp 1747056038
transform 1 0 16608 0 1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_16_169
timestamp 1747056097
transform 1 0 16800 0 1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_16_175
timestamp 1747056038
transform 1 0 17376 0 1 12852
box -48 -56 240 834
use sg13g2_fill_2  FILLER_16_286
timestamp 1747056038
transform 1 0 28032 0 1 12852
box -48 -56 240 834
use sg13g2_decap_8  FILLER_16_297
timestamp 1747056097
transform 1 0 29088 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_304
timestamp 1747056097
transform 1 0 29760 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_311
timestamp 1747056097
transform 1 0 30432 0 1 12852
box -48 -56 720 834
use sg13g2_fill_2  FILLER_16_318
timestamp 1747056038
transform 1 0 31104 0 1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_16_320
timestamp 1747056097
transform 1 0 31296 0 1 12852
box -48 -56 144 834
use sg13g2_fill_1  FILLER_17_0
timestamp 1747056097
transform 1 0 576 0 -1 14364
box -48 -56 144 834
use sg13g2_fill_1  FILLER_17_111
timestamp 1747056097
transform 1 0 11232 0 -1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_17_147
timestamp 1747056038
transform 1 0 14688 0 -1 14364
box -48 -56 240 834
use sg13g2_fill_2  FILLER_17_164
timestamp 1747056038
transform 1 0 16320 0 -1 14364
box -48 -56 240 834
use sg13g2_fill_2  FILLER_17_182
timestamp 1747056038
transform 1 0 18048 0 -1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_17_243
timestamp 1747056097
transform 1 0 23904 0 -1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_17_306
timestamp 1747056097
transform 1 0 29952 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_313
timestamp 1747056097
transform 1 0 30624 0 -1 14364
box -48 -56 720 834
use sg13g2_fill_1  FILLER_17_320
timestamp 1747056097
transform 1 0 31296 0 -1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_18_31
timestamp 1747056038
transform 1 0 3552 0 1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_18_112
timestamp 1747056097
transform 1 0 11328 0 1 14364
box -48 -56 144 834
use sg13g2_fill_1  FILLER_18_122
timestamp 1747056097
transform 1 0 12288 0 1 14364
box -48 -56 144 834
use sg13g2_fill_1  FILLER_18_142
timestamp 1747056097
transform 1 0 14208 0 1 14364
box -48 -56 144 834
use sg13g2_fill_1  FILLER_18_153
timestamp 1747056097
transform 1 0 15264 0 1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_18_170
timestamp 1747056038
transform 1 0 16896 0 1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_18_172
timestamp 1747056097
transform 1 0 17088 0 1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_18_177
timestamp 1747056038
transform 1 0 17568 0 1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_18_179
timestamp 1747056097
transform 1 0 17760 0 1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_18_276
timestamp 1747056038
transform 1 0 27072 0 1 14364
box -48 -56 240 834
use sg13g2_fill_2  FILLER_18_292
timestamp 1747056038
transform 1 0 28608 0 1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_18_294
timestamp 1747056097
transform 1 0 28800 0 1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_18_308
timestamp 1747056097
transform 1 0 30144 0 1 14364
box -48 -56 720 834
use sg13g2_decap_4  FILLER_18_315
timestamp 1747056038
transform 1 0 30816 0 1 14364
box -48 -56 432 834
use sg13g2_fill_2  FILLER_18_319
timestamp 1747056038
transform 1 0 31200 0 1 14364
box -48 -56 240 834
use sg13g2_fill_2  FILLER_19_0
timestamp 1747056038
transform 1 0 576 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_19_2
timestamp 1747056097
transform 1 0 768 0 -1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_19_42
timestamp 1747056038
transform 1 0 4608 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_19_63
timestamp 1747056097
transform 1 0 6624 0 -1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_19_102
timestamp 1747056097
transform 1 0 10368 0 -1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_19_111
timestamp 1747056038
transform 1 0 11232 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_2  FILLER_19_153
timestamp 1747056038
transform 1 0 15264 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_2  FILLER_19_163
timestamp 1747056038
transform 1 0 16224 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_19_165
timestamp 1747056097
transform 1 0 16416 0 -1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_19_171
timestamp 1747056038
transform 1 0 16992 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_19_188
timestamp 1747056097
transform 1 0 18624 0 -1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_19_215
timestamp 1747056038
transform 1 0 21216 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_2  FILLER_19_233
timestamp 1747056038
transform 1 0 22944 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_19_246
timestamp 1747056097
transform 1 0 24192 0 -1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_19_301
timestamp 1747056097
transform 1 0 29472 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_308
timestamp 1747056097
transform 1 0 30144 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_4  FILLER_19_315
timestamp 1747056038
transform 1 0 30816 0 -1 15876
box -48 -56 432 834
use sg13g2_fill_2  FILLER_19_319
timestamp 1747056038
transform 1 0 31200 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_2  FILLER_20_0
timestamp 1747056038
transform 1 0 576 0 1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_20_56
timestamp 1747056097
transform 1 0 5952 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_82
timestamp 1747056097
transform 1 0 8448 0 1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_20_96
timestamp 1747056038
transform 1 0 9792 0 1 15876
box -48 -56 240 834
use sg13g2_fill_2  FILLER_20_120
timestamp 1747056038
transform 1 0 12096 0 1 15876
box -48 -56 240 834
use sg13g2_fill_2  FILLER_20_145
timestamp 1747056038
transform 1 0 14496 0 1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_20_147
timestamp 1747056097
transform 1 0 14688 0 1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_20_232
timestamp 1747056038
transform 1 0 22848 0 1 15876
box -48 -56 240 834
use sg13g2_decap_8  FILLER_20_300
timestamp 1747056097
transform 1 0 29376 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_307
timestamp 1747056097
transform 1 0 30048 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_314
timestamp 1747056097
transform 1 0 30720 0 1 15876
box -48 -56 720 834
use sg13g2_fill_2  FILLER_21_0
timestamp 1747056038
transform 1 0 576 0 -1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_21_2
timestamp 1747056097
transform 1 0 768 0 -1 17388
box -48 -56 144 834
use sg13g2_fill_2  FILLER_21_23
timestamp 1747056038
transform 1 0 2784 0 -1 17388
box -48 -56 240 834
use sg13g2_fill_2  FILLER_21_40
timestamp 1747056038
transform 1 0 4416 0 -1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_21_42
timestamp 1747056097
transform 1 0 4608 0 -1 17388
box -48 -56 144 834
use sg13g2_fill_2  FILLER_21_64
timestamp 1747056038
transform 1 0 6720 0 -1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_21_66
timestamp 1747056097
transform 1 0 6912 0 -1 17388
box -48 -56 144 834
use sg13g2_fill_2  FILLER_21_72
timestamp 1747056038
transform 1 0 7488 0 -1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_21_80
timestamp 1747056097
transform 1 0 8256 0 -1 17388
box -48 -56 144 834
use sg13g2_fill_2  FILLER_21_99
timestamp 1747056038
transform 1 0 10080 0 -1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_21_106
timestamp 1747056097
transform 1 0 10752 0 -1 17388
box -48 -56 144 834
use sg13g2_fill_1  FILLER_21_117
timestamp 1747056097
transform 1 0 11808 0 -1 17388
box -48 -56 144 834
use sg13g2_fill_1  FILLER_21_146
timestamp 1747056097
transform 1 0 14592 0 -1 17388
box -48 -56 144 834
use sg13g2_fill_1  FILLER_21_179
timestamp 1747056097
transform 1 0 17760 0 -1 17388
box -48 -56 144 834
use sg13g2_fill_2  FILLER_21_205
timestamp 1747056038
transform 1 0 20256 0 -1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_21_217
timestamp 1747056097
transform 1 0 21408 0 -1 17388
box -48 -56 144 834
use sg13g2_fill_1  FILLER_21_240
timestamp 1747056097
transform 1 0 23616 0 -1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_21_288
timestamp 1747056097
transform 1 0 28224 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_295
timestamp 1747056097
transform 1 0 28896 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_302
timestamp 1747056097
transform 1 0 29568 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_309
timestamp 1747056097
transform 1 0 30240 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_21_316
timestamp 1747056038
transform 1 0 30912 0 -1 17388
box -48 -56 432 834
use sg13g2_fill_1  FILLER_21_320
timestamp 1747056097
transform 1 0 31296 0 -1 17388
box -48 -56 144 834
use sg13g2_fill_1  FILLER_22_0
timestamp 1747056097
transform 1 0 576 0 1 17388
box -48 -56 144 834
use sg13g2_fill_1  FILLER_22_38
timestamp 1747056097
transform 1 0 4224 0 1 17388
box -48 -56 144 834
use sg13g2_fill_2  FILLER_22_77
timestamp 1747056038
transform 1 0 7968 0 1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_22_102
timestamp 1747056097
transform 1 0 10368 0 1 17388
box -48 -56 144 834
use sg13g2_fill_2  FILLER_22_107
timestamp 1747056038
transform 1 0 10848 0 1 17388
box -48 -56 240 834
use sg13g2_fill_2  FILLER_22_151
timestamp 1747056038
transform 1 0 15072 0 1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_22_165
timestamp 1747056097
transform 1 0 16416 0 1 17388
box -48 -56 144 834
use sg13g2_fill_1  FILLER_22_212
timestamp 1747056097
transform 1 0 20928 0 1 17388
box -48 -56 144 834
use sg13g2_fill_2  FILLER_22_229
timestamp 1747056038
transform 1 0 22560 0 1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_22_231
timestamp 1747056097
transform 1 0 22752 0 1 17388
box -48 -56 144 834
use sg13g2_fill_1  FILLER_22_249
timestamp 1747056097
transform 1 0 24480 0 1 17388
box -48 -56 144 834
use sg13g2_fill_1  FILLER_22_263
timestamp 1747056097
transform 1 0 25824 0 1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_22_289
timestamp 1747056097
transform 1 0 28320 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_296
timestamp 1747056097
transform 1 0 28992 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_303
timestamp 1747056097
transform 1 0 29664 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_310
timestamp 1747056097
transform 1 0 30336 0 1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_22_317
timestamp 1747056038
transform 1 0 31008 0 1 17388
box -48 -56 432 834
use sg13g2_fill_1  FILLER_23_15
timestamp 1747056097
transform 1 0 2016 0 -1 18900
box -48 -56 144 834
use sg13g2_fill_1  FILLER_23_35
timestamp 1747056097
transform 1 0 3936 0 -1 18900
box -48 -56 144 834
use sg13g2_fill_2  FILLER_23_40
timestamp 1747056038
transform 1 0 4416 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_23_42
timestamp 1747056097
transform 1 0 4608 0 -1 18900
box -48 -56 144 834
use sg13g2_fill_2  FILLER_23_121
timestamp 1747056038
transform 1 0 12192 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_23_123
timestamp 1747056097
transform 1 0 12384 0 -1 18900
box -48 -56 144 834
use sg13g2_fill_1  FILLER_23_150
timestamp 1747056097
transform 1 0 14976 0 -1 18900
box -48 -56 144 834
use sg13g2_fill_1  FILLER_23_157
timestamp 1747056097
transform 1 0 15648 0 -1 18900
box -48 -56 144 834
use sg13g2_fill_2  FILLER_23_179
timestamp 1747056038
transform 1 0 17760 0 -1 18900
box -48 -56 240 834
use sg13g2_decap_8  FILLER_23_298
timestamp 1747056097
transform 1 0 29184 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_305
timestamp 1747056097
transform 1 0 29856 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_312
timestamp 1747056097
transform 1 0 30528 0 -1 18900
box -48 -56 720 834
use sg13g2_fill_2  FILLER_23_319
timestamp 1747056038
transform 1 0 31200 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_2  FILLER_24_0
timestamp 1747056038
transform 1 0 576 0 1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_24_2
timestamp 1747056097
transform 1 0 768 0 1 18900
box -48 -56 144 834
use sg13g2_fill_1  FILLER_24_36
timestamp 1747056097
transform 1 0 4032 0 1 18900
box -48 -56 144 834
use sg13g2_fill_2  FILLER_24_53
timestamp 1747056038
transform 1 0 5664 0 1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_24_60
timestamp 1747056097
transform 1 0 6336 0 1 18900
box -48 -56 144 834
use sg13g2_fill_1  FILLER_24_82
timestamp 1747056097
transform 1 0 8448 0 1 18900
box -48 -56 144 834
use sg13g2_fill_2  FILLER_24_120
timestamp 1747056038
transform 1 0 12096 0 1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_24_122
timestamp 1747056097
transform 1 0 12288 0 1 18900
box -48 -56 144 834
use sg13g2_fill_1  FILLER_24_128
timestamp 1747056097
transform 1 0 12864 0 1 18900
box -48 -56 144 834
use sg13g2_fill_2  FILLER_24_216
timestamp 1747056038
transform 1 0 21312 0 1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_24_242
timestamp 1747056097
transform 1 0 23808 0 1 18900
box -48 -56 144 834
use sg13g2_fill_1  FILLER_24_270
timestamp 1747056097
transform 1 0 26496 0 1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_24_305
timestamp 1747056097
transform 1 0 29856 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_312
timestamp 1747056097
transform 1 0 30528 0 1 18900
box -48 -56 720 834
use sg13g2_fill_2  FILLER_24_319
timestamp 1747056038
transform 1 0 31200 0 1 18900
box -48 -56 240 834
use sg13g2_fill_2  FILLER_25_0
timestamp 1747056038
transform 1 0 576 0 -1 20412
box -48 -56 240 834
use sg13g2_fill_2  FILLER_25_22
timestamp 1747056038
transform 1 0 2688 0 -1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_25_112
timestamp 1747056097
transform 1 0 11328 0 -1 20412
box -48 -56 144 834
use sg13g2_fill_1  FILLER_25_121
timestamp 1747056097
transform 1 0 12192 0 -1 20412
box -48 -56 144 834
use sg13g2_fill_2  FILLER_25_149
timestamp 1747056038
transform 1 0 14880 0 -1 20412
box -48 -56 240 834
use sg13g2_fill_2  FILLER_25_156
timestamp 1747056038
transform 1 0 15552 0 -1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_25_158
timestamp 1747056097
transform 1 0 15744 0 -1 20412
box -48 -56 144 834
use sg13g2_fill_2  FILLER_25_190
timestamp 1747056038
transform 1 0 18816 0 -1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_25_239
timestamp 1747056097
transform 1 0 23520 0 -1 20412
box -48 -56 144 834
use sg13g2_fill_1  FILLER_25_260
timestamp 1747056097
transform 1 0 25536 0 -1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_25_312
timestamp 1747056097
transform 1 0 30528 0 -1 20412
box -48 -56 720 834
use sg13g2_fill_2  FILLER_25_319
timestamp 1747056038
transform 1 0 31200 0 -1 20412
box -48 -56 240 834
use sg13g2_fill_2  FILLER_26_0
timestamp 1747056038
transform 1 0 576 0 1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_26_28
timestamp 1747056097
transform 1 0 3264 0 1 20412
box -48 -56 144 834
use sg13g2_fill_2  FILLER_26_42
timestamp 1747056038
transform 1 0 4608 0 1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_26_53
timestamp 1747056097
transform 1 0 5664 0 1 20412
box -48 -56 144 834
use sg13g2_fill_1  FILLER_26_93
timestamp 1747056097
transform 1 0 9504 0 1 20412
box -48 -56 144 834
use sg13g2_fill_2  FILLER_26_104
timestamp 1747056038
transform 1 0 10560 0 1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_26_106
timestamp 1747056097
transform 1 0 10752 0 1 20412
box -48 -56 144 834
use sg13g2_fill_2  FILLER_26_155
timestamp 1747056038
transform 1 0 15456 0 1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_26_157
timestamp 1747056097
transform 1 0 15648 0 1 20412
box -48 -56 144 834
use sg13g2_fill_1  FILLER_26_167
timestamp 1747056097
transform 1 0 16608 0 1 20412
box -48 -56 144 834
use sg13g2_fill_2  FILLER_26_199
timestamp 1747056038
transform 1 0 19680 0 1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_26_201
timestamp 1747056097
transform 1 0 19872 0 1 20412
box -48 -56 144 834
use sg13g2_fill_2  FILLER_26_230
timestamp 1747056038
transform 1 0 22656 0 1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_26_245
timestamp 1747056097
transform 1 0 24096 0 1 20412
box -48 -56 144 834
use sg13g2_fill_2  FILLER_26_251
timestamp 1747056038
transform 1 0 24672 0 1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_26_267
timestamp 1747056097
transform 1 0 26208 0 1 20412
box -48 -56 144 834
use sg13g2_fill_2  FILLER_26_319
timestamp 1747056038
transform 1 0 31200 0 1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_27_0
timestamp 1747056097
transform 1 0 576 0 -1 21924
box -48 -56 144 834
use sg13g2_fill_2  FILLER_27_36
timestamp 1747056038
transform 1 0 4032 0 -1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_27_38
timestamp 1747056097
transform 1 0 4224 0 -1 21924
box -48 -56 144 834
use sg13g2_fill_2  FILLER_27_59
timestamp 1747056038
transform 1 0 6240 0 -1 21924
box -48 -56 240 834
use sg13g2_fill_2  FILLER_27_125
timestamp 1747056038
transform 1 0 12576 0 -1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_27_135
timestamp 1747056097
transform 1 0 13536 0 -1 21924
box -48 -56 144 834
use sg13g2_fill_1  FILLER_27_165
timestamp 1747056097
transform 1 0 16416 0 -1 21924
box -48 -56 144 834
use sg13g2_fill_1  FILLER_27_194
timestamp 1747056097
transform 1 0 19200 0 -1 21924
box -48 -56 144 834
use sg13g2_fill_2  FILLER_27_319
timestamp 1747056038
transform 1 0 31200 0 -1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_28_0
timestamp 1747056097
transform 1 0 576 0 1 21924
box -48 -56 144 834
use sg13g2_fill_2  FILLER_28_17
timestamp 1747056038
transform 1 0 2208 0 1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_28_19
timestamp 1747056097
transform 1 0 2400 0 1 21924
box -48 -56 144 834
use sg13g2_fill_1  FILLER_28_59
timestamp 1747056097
transform 1 0 6240 0 1 21924
box -48 -56 144 834
use sg13g2_fill_1  FILLER_28_86
timestamp 1747056097
transform 1 0 8832 0 1 21924
box -48 -56 144 834
use sg13g2_fill_2  FILLER_28_92
timestamp 1747056038
transform 1 0 9408 0 1 21924
box -48 -56 240 834
use sg13g2_fill_2  FILLER_28_99
timestamp 1747056038
transform 1 0 10080 0 1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_28_137
timestamp 1747056097
transform 1 0 13728 0 1 21924
box -48 -56 144 834
use sg13g2_fill_1  FILLER_28_146
timestamp 1747056097
transform 1 0 14592 0 1 21924
box -48 -56 144 834
use sg13g2_fill_2  FILLER_28_249
timestamp 1747056038
transform 1 0 24480 0 1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_28_320
timestamp 1747056097
transform 1 0 31296 0 1 21924
box -48 -56 144 834
use sg13g2_fill_2  FILLER_29_26
timestamp 1747056038
transform 1 0 3072 0 -1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_29_28
timestamp 1747056097
transform 1 0 3264 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_29_62
timestamp 1747056097
transform 1 0 6528 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_29_135
timestamp 1747056038
transform 1 0 13536 0 -1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_29_154
timestamp 1747056097
transform 1 0 15360 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_29_168
timestamp 1747056038
transform 1 0 16704 0 -1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_29_179
timestamp 1747056097
transform 1 0 17760 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_29_207
timestamp 1747056097
transform 1 0 20448 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_29_222
timestamp 1747056097
transform 1 0 21888 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_19
timestamp 1747056097
transform 1 0 2400 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_85
timestamp 1747056097
transform 1 0 8736 0 1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_30_106
timestamp 1747056038
transform 1 0 10752 0 1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_30_153
timestamp 1747056097
transform 1 0 15264 0 1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_30_179
timestamp 1747056038
transform 1 0 17760 0 1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_30_233
timestamp 1747056097
transform 1 0 22944 0 1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_30_268
timestamp 1747056038
transform 1 0 26304 0 1 23436
box -48 -56 240 834
use sg13g2_fill_2  FILLER_30_319
timestamp 1747056038
transform 1 0 31200 0 1 23436
box -48 -56 240 834
use sg13g2_fill_2  FILLER_31_90
timestamp 1747056038
transform 1 0 9216 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_31_149
timestamp 1747056097
transform 1 0 14880 0 -1 24948
box -48 -56 144 834
use sg13g2_fill_2  FILLER_31_155
timestamp 1747056038
transform 1 0 15456 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_31_200
timestamp 1747056097
transform 1 0 19776 0 -1 24948
box -48 -56 144 834
use sg13g2_fill_1  FILLER_31_320
timestamp 1747056097
transform 1 0 31296 0 -1 24948
box -48 -56 144 834
use sg13g2_fill_2  FILLER_32_0
timestamp 1747056038
transform 1 0 576 0 1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_32_38
timestamp 1747056097
transform 1 0 4224 0 1 24948
box -48 -56 144 834
use sg13g2_fill_1  FILLER_32_105
timestamp 1747056097
transform 1 0 10656 0 1 24948
box -48 -56 144 834
use sg13g2_fill_2  FILLER_32_152
timestamp 1747056038
transform 1 0 15168 0 1 24948
box -48 -56 240 834
use sg13g2_fill_2  FILLER_32_178
timestamp 1747056038
transform 1 0 17664 0 1 24948
box -48 -56 240 834
use sg13g2_fill_2  FILLER_32_318
timestamp 1747056038
transform 1 0 31104 0 1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_32_320
timestamp 1747056097
transform 1 0 31296 0 1 24948
box -48 -56 144 834
use sg13g2_fill_1  FILLER_33_9
timestamp 1747056097
transform 1 0 1440 0 -1 26460
box -48 -56 144 834
use sg13g2_fill_1  FILLER_33_49
timestamp 1747056097
transform 1 0 5280 0 -1 26460
box -48 -56 144 834
use sg13g2_fill_2  FILLER_33_86
timestamp 1747056038
transform 1 0 8832 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_33_136
timestamp 1747056097
transform 1 0 13632 0 -1 26460
box -48 -56 144 834
use sg13g2_fill_2  FILLER_33_183
timestamp 1747056038
transform 1 0 18144 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_33_190
timestamp 1747056097
transform 1 0 18816 0 -1 26460
box -48 -56 144 834
use sg13g2_fill_1  FILLER_33_197
timestamp 1747056097
transform 1 0 19488 0 -1 26460
box -48 -56 144 834
use sg13g2_fill_1  FILLER_33_221
timestamp 1747056097
transform 1 0 21792 0 -1 26460
box -48 -56 144 834
use sg13g2_fill_1  FILLER_33_320
timestamp 1747056097
transform 1 0 31296 0 -1 26460
box -48 -56 144 834
use sg13g2_fill_1  FILLER_34_228
timestamp 1747056097
transform 1 0 22464 0 1 26460
box -48 -56 144 834
use sg13g2_fill_1  FILLER_34_247
timestamp 1747056097
transform 1 0 24288 0 1 26460
box -48 -56 144 834
use sg13g2_fill_2  FILLER_35_0
timestamp 1747056038
transform 1 0 576 0 -1 27972
box -48 -56 240 834
use sg13g2_fill_1  FILLER_35_96
timestamp 1747056097
transform 1 0 9792 0 -1 27972
box -48 -56 144 834
use sg13g2_fill_2  FILLER_35_141
timestamp 1747056038
transform 1 0 14112 0 -1 27972
box -48 -56 240 834
use sg13g2_fill_1  FILLER_35_314
timestamp 1747056097
transform 1 0 30720 0 -1 27972
box -48 -56 144 834
use sg13g2_fill_1  FILLER_35_320
timestamp 1747056097
transform 1 0 31296 0 -1 27972
box -48 -56 144 834
use sg13g2_dlygate4sd3_1  hold1
timestamp 1747056038
transform -1 0 29760 0 1 14364
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold2
timestamp 1747056038
transform -1 0 20352 0 1 18900
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold3
timestamp 1747056038
transform 1 0 23040 0 1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold4
timestamp 1747056038
transform -1 0 23712 0 -1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold5
timestamp 1747056038
transform -1 0 10656 0 -1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold6
timestamp 1747056038
transform 1 0 24384 0 1 18900
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold7
timestamp 1747056038
transform -1 0 27360 0 1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold8
timestamp 1747056038
transform -1 0 19584 0 -1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold9
timestamp 1747056038
transform 1 0 11904 0 -1 24948
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold10
timestamp 1747056038
transform -1 0 23424 0 1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold11
timestamp 1747056038
transform 1 0 24000 0 1 24948
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold12
timestamp 1747056038
transform -1 0 4224 0 1 24948
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold13
timestamp 1747056038
transform -1 0 2112 0 1 24948
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold14
timestamp 1747056038
transform 1 0 26592 0 1 18900
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold15
timestamp 1747056038
transform -1 0 22848 0 -1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold16
timestamp 1747056038
transform -1 0 21888 0 -1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold17
timestamp 1747056038
transform 1 0 28128 0 -1 20412
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold18
timestamp 1747056038
transform -1 0 28224 0 1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold19
timestamp 1747056038
transform -1 0 26208 0 1 20412
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold20
timestamp 1747056038
transform 1 0 26304 0 1 20412
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold21
timestamp 1747056038
transform -1 0 25056 0 1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold22
timestamp 1747056038
transform -1 0 28704 0 1 24948
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold23
timestamp 1747056038
transform -1 0 27072 0 1 6804
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold24
timestamp 1747056038
transform 1 0 24768 0 -1 8316
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold25
timestamp 1747056038
transform -1 0 25056 0 -1 6804
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold26
timestamp 1747056038
transform -1 0 7200 0 -1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold27
timestamp 1747056038
transform -1 0 8928 0 1 24948
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold28
timestamp 1747056038
transform 1 0 14016 0 -1 24948
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold29
timestamp 1747056038
transform -1 0 16512 0 -1 24948
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold30
timestamp 1747056038
transform 1 0 20352 0 -1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold31
timestamp 1747056038
transform -1 0 22464 0 1 24948
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold32
timestamp 1747056038
transform 1 0 24480 0 1 15876
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold33
timestamp 1747056038
transform 1 0 25920 0 1 17388
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold34
timestamp 1747056038
transform 1 0 25248 0 1 18900
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold35
timestamp 1747056038
transform 1 0 25824 0 1 21924
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold36
timestamp 1747056038
transform 1 0 14496 0 -1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold37
timestamp 1747056038
transform -1 0 5280 0 -1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold38
timestamp 1747056038
transform -1 0 22464 0 1 6804
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold39
timestamp 1747056038
transform -1 0 21120 0 1 5292
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold40
timestamp 1747056038
transform -1 0 25920 0 -1 6804
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold41
timestamp 1747056038
transform 1 0 11904 0 -1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold42
timestamp 1747056038
transform -1 0 26688 0 -1 14364
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold43
timestamp 1747056038
transform -1 0 3936 0 -1 24948
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold44
timestamp 1747056038
transform -1 0 2400 0 1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold45
timestamp 1747056038
transform -1 0 4896 0 1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold46
timestamp 1747056038
transform 1 0 24864 0 -1 27972
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold47
timestamp 1747056038
transform 1 0 23904 0 -1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold48
timestamp 1747056038
transform 1 0 23136 0 1 24948
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold49
timestamp 1747056038
transform -1 0 24288 0 1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold50
timestamp 1747056038
transform 1 0 20736 0 1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold51
timestamp 1747056038
transform -1 0 22464 0 1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold52
timestamp 1747056038
transform 1 0 15840 0 1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold53
timestamp 1747056038
transform 1 0 27264 0 1 14364
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold54
timestamp 1747056038
transform -1 0 25824 0 -1 14364
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold55
timestamp 1747056038
transform 1 0 24192 0 1 11340
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold56
timestamp 1747056038
transform -1 0 22560 0 -1 11340
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold57
timestamp 1747056038
transform 1 0 20832 0 -1 11340
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold58
timestamp 1747056038
transform 1 0 7392 0 1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold59
timestamp 1747056038
transform -1 0 8064 0 -1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold60
timestamp 1747056038
transform 1 0 8928 0 1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold61
timestamp 1747056038
transform -1 0 23136 0 1 9828
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold62
timestamp 1747056038
transform -1 0 26208 0 1 15876
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold63
timestamp 1747056038
transform 1 0 25344 0 1 9828
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold64
timestamp 1747056038
transform -1 0 27072 0 1 9828
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold65
timestamp 1747056038
transform -1 0 13152 0 1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold66
timestamp 1747056038
transform -1 0 2016 0 -1 14364
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold67
timestamp 1747056038
transform -1 0 3168 0 -1 9828
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold68
timestamp 1747056038
transform 1 0 11712 0 -1 21924
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold69
timestamp 1747056038
transform 1 0 6528 0 1 6804
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold70
timestamp 1747056038
transform 1 0 9120 0 1 5292
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold71
timestamp 1747056038
transform 1 0 19488 0 1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold72
timestamp 1747056038
transform -1 0 24768 0 -1 12852
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold73
timestamp 1747056038
transform 1 0 16224 0 -1 5292
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold74
timestamp 1747056038
transform 1 0 19392 0 1 5292
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold75
timestamp 1747056038
transform 1 0 864 0 1 12852
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold76
timestamp 1747056038
transform 1 0 14112 0 -1 5292
box -48 -56 912 834
use sg13g2_buf_2  input1
timestamp 1747056038
transform -1 0 31296 0 -1 27972
box -48 -56 528 834
use sg13g2_buf_1  input2
timestamp 1747056038
transform -1 0 30432 0 1 20412
box -48 -56 432 834
use sg13g2_buf_2  input3
timestamp 1747056038
transform -1 0 29568 0 -1 27972
box -48 -56 528 834
use sg13g2_buf_2  input4
timestamp 1747056038
transform -1 0 29088 0 -1 27972
box -48 -56 528 834
use sg13g2_buf_2  input5
timestamp 1747056038
transform -1 0 28320 0 1 26460
box -48 -56 528 834
use sg13g2_buf_2  input6
timestamp 1747056038
transform -1 0 28608 0 -1 27972
box -48 -56 528 834
use sg13g2_buf_2  input7
timestamp 1747056038
transform -1 0 28128 0 -1 27972
box -48 -56 528 834
use sg13g2_buf_2  input8
timestamp 1747056038
transform -1 0 27648 0 -1 27972
box -48 -56 528 834
use sg13g2_buf_2  input9
timestamp 1747056038
transform -1 0 27168 0 -1 27972
box -48 -56 528 834
use sg13g2_buf_1  input10
timestamp 1747056038
transform -1 0 30144 0 -1 26460
box -48 -56 432 834
<< labels >>
flabel metal5 s 27638 712 28078 28016 0 FreeSans 3200 90 0 0 VGND
port 1 nsew
flabel metal5 s 19864 712 20304 28016 0 FreeSans 3200 90 0 0 VGND
port 1 nsew
flabel metal5 s 12090 712 12530 28016 0 FreeSans 3200 90 0 0 VGND
port 1 nsew
flabel metal5 s 4316 712 4756 28016 0 FreeSans 3200 90 0 0 VGND
port 1 nsew
flabel metal5 s 26398 712 26838 28016 0 FreeSans 3200 90 0 0 VPWR
port 2 nsew
flabel metal5 s 18624 712 19064 28016 0 FreeSans 3200 90 0 0 VPWR
port 2 nsew
flabel metal5 s 10850 712 11290 28016 0 FreeSans 3200 90 0 0 VPWR
port 2 nsew
flabel metal5 s 3076 712 3516 28016 0 FreeSans 3200 90 0 0 VPWR
port 2 nsew
flabel metal3 s 11576 28600 11656 29000 0 FreeSans 400 90 0 0 b6
port 3 nsew
flabel metal3 s 14648 28600 14728 29000 0 FreeSans 400 90 0 0 b7
port 4 nsew
flabel metal3 s 30008 28600 30088 29000 0 FreeSans 400 90 0 0 clk
port 5 nsew
flabel metal2 s 0 8864 400 8944 0 FreeSans 400 0 0 0 db[0]
port 6 nsew
flabel metal2 s 0 8444 400 8524 0 FreeSans 400 0 0 0 db[1]
port 7 nsew
flabel metal2 s 0 8024 400 8104 0 FreeSans 400 0 0 0 db[2]
port 8 nsew
flabel metal2 s 0 7604 400 7684 0 FreeSans 400 0 0 0 db[3]
port 9 nsew
flabel metal2 s 0 7184 400 7264 0 FreeSans 400 0 0 0 db[4]
port 10 nsew
flabel metal2 s 0 6764 400 6844 0 FreeSans 400 0 0 0 db[5]
port 11 nsew
flabel metal2 s 0 6344 400 6424 0 FreeSans 400 0 0 0 db[6]
port 12 nsew
flabel metal2 s 0 5924 400 6004 0 FreeSans 400 0 0 0 db[7]
port 13 nsew
flabel metal2 s 0 15584 400 15664 0 FreeSans 400 0 0 0 dg[0]
port 14 nsew
flabel metal2 s 0 15164 400 15244 0 FreeSans 400 0 0 0 dg[1]
port 15 nsew
flabel metal2 s 0 14744 400 14824 0 FreeSans 400 0 0 0 dg[2]
port 16 nsew
flabel metal2 s 0 14324 400 14404 0 FreeSans 400 0 0 0 dg[3]
port 17 nsew
flabel metal2 s 0 13904 400 13984 0 FreeSans 400 0 0 0 dg[4]
port 18 nsew
flabel metal2 s 0 13484 400 13564 0 FreeSans 400 0 0 0 dg[5]
port 19 nsew
flabel metal2 s 0 13064 400 13144 0 FreeSans 400 0 0 0 dg[6]
port 20 nsew
flabel metal2 s 0 12644 400 12724 0 FreeSans 400 0 0 0 dg[7]
port 21 nsew
flabel metal2 s 0 22304 400 22384 0 FreeSans 400 0 0 0 dr[0]
port 22 nsew
flabel metal2 s 0 21884 400 21964 0 FreeSans 400 0 0 0 dr[1]
port 23 nsew
flabel metal2 s 0 21464 400 21544 0 FreeSans 400 0 0 0 dr[2]
port 24 nsew
flabel metal2 s 0 21044 400 21124 0 FreeSans 400 0 0 0 dr[3]
port 25 nsew
flabel metal2 s 0 20624 400 20704 0 FreeSans 400 0 0 0 dr[4]
port 26 nsew
flabel metal2 s 0 20204 400 20284 0 FreeSans 400 0 0 0 dr[5]
port 27 nsew
flabel metal2 s 0 19784 400 19864 0 FreeSans 400 0 0 0 dr[6]
port 28 nsew
flabel metal2 s 0 19364 400 19444 0 FreeSans 400 0 0 0 dr[7]
port 29 nsew
flabel metal3 s 30776 28600 30856 29000 0 FreeSans 400 90 0 0 ena
port 30 nsew
flabel metal3 s 12344 28600 12424 29000 0 FreeSans 400 90 0 0 g6
port 31 nsew
flabel metal3 s 15416 28600 15496 29000 0 FreeSans 400 90 0 0 g7
port 32 nsew
flabel metal3 s 9272 28600 9352 29000 0 FreeSans 400 90 0 0 hblank
port 33 nsew
flabel metal3 s 10808 28600 10888 29000 0 FreeSans 400 90 0 0 hsync
port 34 nsew
flabel metal3 s 13112 28600 13192 29000 0 FreeSans 400 90 0 0 r6
port 35 nsew
flabel metal3 s 16184 28600 16264 29000 0 FreeSans 400 90 0 0 r7
port 36 nsew
flabel metal3 s 29240 28600 29320 29000 0 FreeSans 400 90 0 0 rst_n
port 37 nsew
flabel metal3 s 28472 28600 28552 29000 0 FreeSans 400 90 0 0 ui_in[0]
port 38 nsew
flabel metal3 s 27704 28600 27784 29000 0 FreeSans 400 90 0 0 ui_in[1]
port 39 nsew
flabel metal3 s 26936 28600 27016 29000 0 FreeSans 400 90 0 0 ui_in[2]
port 40 nsew
flabel metal3 s 26168 28600 26248 29000 0 FreeSans 400 90 0 0 ui_in[3]
port 41 nsew
flabel metal3 s 25400 28600 25480 29000 0 FreeSans 400 90 0 0 ui_in[4]
port 42 nsew
flabel metal3 s 24632 28600 24712 29000 0 FreeSans 400 90 0 0 ui_in[5]
port 43 nsew
flabel metal3 s 23864 28600 23944 29000 0 FreeSans 400 90 0 0 ui_in[6]
port 44 nsew
flabel metal3 s 23096 28600 23176 29000 0 FreeSans 400 90 0 0 ui_in[7]
port 45 nsew
flabel metal3 s 3896 28600 3976 29000 0 FreeSans 400 90 0 0 uio_oe[0]
port 46 nsew
flabel metal3 s 3128 28600 3208 29000 0 FreeSans 400 90 0 0 uio_oe[1]
port 47 nsew
flabel metal3 s 8504 28600 8584 29000 0 FreeSans 400 90 0 0 uio_out2
port 48 nsew
flabel metal3 s 7736 28600 7816 29000 0 FreeSans 400 90 0 0 uio_out3
port 49 nsew
flabel metal3 s 6968 28600 7048 29000 0 FreeSans 400 90 0 0 uio_out4
port 50 nsew
flabel metal3 s 6200 28600 6280 29000 0 FreeSans 400 90 0 0 uio_out5
port 51 nsew
flabel metal3 s 5432 28600 5512 29000 0 FreeSans 400 90 0 0 uio_out6
port 52 nsew
flabel metal3 s 4664 28600 4744 29000 0 FreeSans 400 90 0 0 uio_out7
port 53 nsew
flabel metal3 s 10040 28600 10120 29000 0 FreeSans 400 90 0 0 vblank
port 54 nsew
flabel metal3 s 13880 28600 13960 29000 0 FreeSans 400 90 0 0 vsync
port 55 nsew
<< properties >>
string FIXED_BBOX 0 0 32000 29000
string GDS_END 2361606
string GDS_FILE ../gds/controller.gds
string GDS_START 261558
<< end >>
