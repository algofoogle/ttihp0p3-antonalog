magic
tech ihp-sg13g2
magscale 1 2
timestamp 1746869612
<< metal1 >>
rect 288 25724 2304 25748
rect 288 25684 1544 25724
rect 1912 25684 2304 25724
rect 288 25660 2304 25684
rect 268 24968 2304 24992
rect 268 24928 304 24968
rect 672 24928 2304 24968
rect 268 24904 2304 24928
rect 288 24212 2304 24236
rect 288 24172 1544 24212
rect 1912 24172 2304 24212
rect 288 24148 2304 24172
rect 730 24044 788 24045
rect 730 24004 739 24044
rect 779 24004 788 24044
rect 730 24003 788 24004
rect 1515 23876 1557 23885
rect 1515 23836 1516 23876
rect 1556 23836 1557 23876
rect 1515 23827 1557 23836
rect 268 23456 2304 23480
rect 268 23416 304 23456
rect 672 23416 2304 23456
rect 268 23392 2304 23416
rect 730 23204 788 23205
rect 730 23164 739 23204
rect 779 23164 788 23204
rect 730 23163 788 23164
rect 1515 23036 1557 23045
rect 1515 22996 1516 23036
rect 1556 22996 1557 23036
rect 1515 22987 1557 22996
rect 288 22700 2304 22724
rect 288 22660 1544 22700
rect 1912 22660 2304 22700
rect 288 22636 2304 22660
rect 538 22448 596 22449
rect 538 22408 547 22448
rect 587 22408 596 22448
rect 538 22407 596 22408
rect 1515 22364 1557 22373
rect 1515 22324 1516 22364
rect 1556 22324 1557 22364
rect 1515 22315 1557 22324
rect 268 21944 2304 21968
rect 268 21904 304 21944
rect 672 21904 2304 21944
rect 268 21880 2304 21904
rect 1114 21608 1172 21609
rect 1114 21568 1123 21608
rect 1163 21568 1172 21608
rect 1114 21567 1172 21568
rect 2091 21524 2133 21533
rect 2091 21484 2092 21524
rect 2132 21484 2133 21524
rect 2091 21475 2133 21484
rect 288 21188 2304 21212
rect 288 21148 1544 21188
rect 1912 21148 2304 21188
rect 288 21124 2304 21148
rect 1114 20936 1172 20937
rect 1114 20896 1123 20936
rect 1163 20896 1172 20936
rect 1114 20895 1172 20896
rect 2091 20852 2133 20861
rect 2091 20812 2092 20852
rect 2132 20812 2133 20852
rect 2091 20803 2133 20812
rect 268 20432 2304 20456
rect 268 20392 304 20432
rect 672 20392 2304 20432
rect 268 20368 2304 20392
rect 730 20264 788 20265
rect 730 20224 739 20264
rect 779 20224 788 20264
rect 730 20223 788 20224
rect 1515 20012 1557 20021
rect 1515 19972 1516 20012
rect 1556 19972 1557 20012
rect 1515 19963 1557 19972
rect 288 19676 2304 19700
rect 288 19636 1544 19676
rect 1912 19636 2304 19676
rect 288 19612 2304 19636
rect 730 19508 788 19509
rect 730 19468 739 19508
rect 779 19468 788 19508
rect 730 19467 788 19468
rect 1515 19340 1557 19349
rect 1515 19300 1516 19340
rect 1556 19300 1557 19340
rect 1515 19291 1557 19300
rect 268 18920 2304 18944
rect 268 18880 304 18920
rect 672 18880 2304 18920
rect 268 18856 2304 18880
rect 538 18584 596 18585
rect 538 18544 547 18584
rect 587 18544 596 18584
rect 538 18543 596 18544
rect 1515 18500 1557 18509
rect 1515 18460 1516 18500
rect 1556 18460 1557 18500
rect 1515 18451 1557 18460
rect 288 18164 2304 18188
rect 288 18124 1544 18164
rect 1912 18124 2304 18164
rect 288 18100 2304 18124
rect 268 17408 2304 17432
rect 268 17368 304 17408
rect 672 17368 2304 17408
rect 268 17344 2304 17368
rect 288 16652 2304 16676
rect 288 16612 1544 16652
rect 1912 16612 2304 16652
rect 288 16588 2304 16612
rect 268 15896 2304 15920
rect 268 15856 304 15896
rect 672 15856 2304 15896
rect 268 15832 2304 15856
rect 730 15728 788 15729
rect 730 15688 739 15728
rect 779 15688 788 15728
rect 730 15687 788 15688
rect 1515 15476 1557 15485
rect 1515 15436 1516 15476
rect 1556 15436 1557 15476
rect 1515 15427 1557 15436
rect 288 15140 2304 15164
rect 288 15100 1544 15140
rect 1912 15100 2304 15140
rect 288 15076 2304 15100
rect 538 14888 596 14889
rect 538 14848 547 14888
rect 587 14848 596 14888
rect 538 14847 596 14848
rect 1515 14804 1557 14813
rect 1515 14764 1516 14804
rect 1556 14764 1557 14804
rect 1515 14755 1557 14764
rect 268 14384 2304 14408
rect 268 14344 304 14384
rect 672 14344 2304 14384
rect 268 14320 2304 14344
rect 538 13964 596 13965
rect 538 13924 547 13964
rect 587 13924 596 13964
rect 538 13923 596 13924
rect 1515 13964 1557 13973
rect 1515 13924 1516 13964
rect 1556 13924 1557 13964
rect 1515 13915 1557 13924
rect 288 13628 2304 13652
rect 288 13588 1544 13628
rect 1912 13588 2304 13628
rect 288 13564 2304 13588
rect 2091 13292 2133 13301
rect 2091 13252 2092 13292
rect 2132 13252 2133 13292
rect 2091 13243 2133 13252
rect 1306 13040 1364 13041
rect 1306 13000 1315 13040
rect 1355 13000 1364 13040
rect 1306 12999 1364 13000
rect 268 12872 2304 12896
rect 268 12832 304 12872
rect 672 12832 2304 12872
rect 268 12808 2304 12832
rect 2091 12452 2133 12461
rect 2091 12412 2092 12452
rect 2132 12412 2133 12452
rect 2091 12403 2133 12412
rect 1306 12284 1364 12285
rect 1306 12244 1315 12284
rect 1355 12244 1364 12284
rect 1306 12243 1364 12244
rect 288 12116 2304 12140
rect 288 12076 1544 12116
rect 1912 12076 2304 12116
rect 288 12052 2304 12076
rect 1515 11780 1557 11789
rect 1515 11740 1516 11780
rect 1556 11740 1557 11780
rect 1515 11731 1557 11740
rect 730 11528 788 11529
rect 730 11488 739 11528
rect 779 11488 788 11528
rect 730 11487 788 11488
rect 268 11360 2304 11384
rect 268 11320 304 11360
rect 672 11320 2304 11360
rect 268 11296 2304 11320
rect 1515 10940 1557 10949
rect 1515 10900 1516 10940
rect 1556 10900 1557 10940
rect 1515 10891 1557 10900
rect 538 10856 596 10857
rect 538 10816 547 10856
rect 587 10816 596 10856
rect 538 10815 596 10816
rect 288 10604 2304 10628
rect 288 10564 1544 10604
rect 1912 10564 2304 10604
rect 288 10540 2304 10564
rect 2091 10268 2133 10277
rect 2091 10228 2092 10268
rect 2132 10228 2133 10268
rect 2091 10219 2133 10228
rect 1114 10184 1172 10185
rect 1114 10144 1123 10184
rect 1163 10144 1172 10184
rect 1114 10143 1172 10144
rect 268 9848 2304 9872
rect 268 9808 304 9848
rect 672 9808 2304 9848
rect 268 9784 2304 9808
rect 288 9092 2304 9116
rect 288 9052 1544 9092
rect 1912 9052 2304 9092
rect 288 9028 2304 9052
rect 268 8336 2304 8360
rect 268 8296 304 8336
rect 672 8296 2304 8336
rect 268 8272 2304 8296
rect 288 7580 2304 7604
rect 288 7540 1544 7580
rect 1912 7540 2304 7580
rect 288 7516 2304 7540
rect 1515 7244 1557 7253
rect 1515 7204 1516 7244
rect 1556 7204 1557 7244
rect 1515 7195 1557 7204
rect 730 6992 788 6993
rect 730 6952 739 6992
rect 779 6952 788 6992
rect 730 6951 788 6952
rect 268 6824 2304 6848
rect 268 6784 304 6824
rect 672 6784 2304 6824
rect 268 6760 2304 6784
rect 1515 6404 1557 6413
rect 1515 6364 1516 6404
rect 1556 6364 1557 6404
rect 1515 6355 1557 6364
rect 538 6320 596 6321
rect 538 6280 547 6320
rect 587 6280 596 6320
rect 538 6279 596 6280
rect 288 6068 2304 6092
rect 288 6028 1544 6068
rect 1912 6028 2304 6068
rect 288 6004 2304 6028
rect 1515 5732 1557 5741
rect 1515 5692 1516 5732
rect 1556 5692 1557 5732
rect 1515 5683 1557 5692
rect 730 5480 788 5481
rect 730 5440 739 5480
rect 779 5440 788 5480
rect 730 5439 788 5440
rect 268 5312 2304 5336
rect 268 5272 304 5312
rect 672 5272 2304 5312
rect 268 5248 2304 5272
rect 2091 4892 2133 4901
rect 2091 4852 2092 4892
rect 2132 4852 2133 4892
rect 2091 4843 2133 4852
rect 1114 4808 1172 4809
rect 1114 4768 1123 4808
rect 1163 4768 1172 4808
rect 1114 4767 1172 4768
rect 288 4556 2304 4580
rect 288 4516 1544 4556
rect 1912 4516 2304 4556
rect 288 4492 2304 4516
rect 2091 4220 2133 4229
rect 2091 4180 2092 4220
rect 2132 4180 2133 4220
rect 2091 4171 2133 4180
rect 1306 3968 1364 3969
rect 1306 3928 1315 3968
rect 1355 3928 1364 3968
rect 1306 3927 1364 3928
rect 268 3800 2304 3824
rect 268 3760 304 3800
rect 672 3760 2304 3800
rect 268 3736 2304 3760
rect 2091 3380 2133 3389
rect 2091 3340 2092 3380
rect 2132 3340 2133 3380
rect 2091 3331 2133 3340
rect 1114 3296 1172 3297
rect 1114 3256 1123 3296
rect 1163 3256 1172 3296
rect 1114 3255 1172 3256
rect 288 3044 2304 3068
rect 288 3004 1544 3044
rect 1912 3004 2304 3044
rect 288 2980 2304 3004
rect 730 2876 788 2877
rect 730 2836 739 2876
rect 779 2836 788 2876
rect 730 2835 788 2836
rect 1515 2708 1557 2717
rect 1515 2668 1516 2708
rect 1556 2668 1557 2708
rect 1515 2659 1557 2668
rect 268 2288 2304 2312
rect 268 2248 304 2288
rect 672 2248 2304 2288
rect 268 2224 2304 2248
rect 1515 1868 1557 1877
rect 1515 1828 1516 1868
rect 1556 1828 1557 1868
rect 1515 1819 1557 1828
rect 538 1784 596 1785
rect 538 1744 547 1784
rect 587 1744 596 1784
rect 538 1743 596 1744
rect 288 1532 2304 1556
rect 288 1492 1544 1532
rect 1912 1492 2304 1532
rect 288 1468 2304 1492
rect 268 776 2304 800
rect 268 736 304 776
rect 672 736 2304 776
rect 268 712 2304 736
rect 288 20 2304 44
rect 288 -20 1544 20
rect 1912 -20 2304 20
rect 288 -44 2304 -20
<< via1 >>
rect 1544 25684 1912 25724
rect 304 24928 672 24968
rect 1544 24172 1912 24212
rect 739 24004 779 24044
rect 1516 23836 1556 23876
rect 304 23416 672 23456
rect 739 23164 779 23204
rect 1516 22996 1556 23036
rect 1544 22660 1912 22700
rect 547 22408 587 22448
rect 1516 22324 1556 22364
rect 304 21904 672 21944
rect 1123 21568 1163 21608
rect 2092 21484 2132 21524
rect 1544 21148 1912 21188
rect 1123 20896 1163 20936
rect 2092 20812 2132 20852
rect 304 20392 672 20432
rect 739 20224 779 20264
rect 1516 19972 1556 20012
rect 1544 19636 1912 19676
rect 739 19468 779 19508
rect 1516 19300 1556 19340
rect 304 18880 672 18920
rect 547 18544 587 18584
rect 1516 18460 1556 18500
rect 1544 18124 1912 18164
rect 304 17368 672 17408
rect 1544 16612 1912 16652
rect 304 15856 672 15896
rect 739 15688 779 15728
rect 1516 15436 1556 15476
rect 1544 15100 1912 15140
rect 547 14848 587 14888
rect 1516 14764 1556 14804
rect 304 14344 672 14384
rect 547 13924 587 13964
rect 1516 13924 1556 13964
rect 1544 13588 1912 13628
rect 2092 13252 2132 13292
rect 1315 13000 1355 13040
rect 304 12832 672 12872
rect 2092 12412 2132 12452
rect 1315 12244 1355 12284
rect 1544 12076 1912 12116
rect 1516 11740 1556 11780
rect 739 11488 779 11528
rect 304 11320 672 11360
rect 1516 10900 1556 10940
rect 547 10816 587 10856
rect 1544 10564 1912 10604
rect 2092 10228 2132 10268
rect 1123 10144 1163 10184
rect 304 9808 672 9848
rect 1544 9052 1912 9092
rect 304 8296 672 8336
rect 1544 7540 1912 7580
rect 1516 7204 1556 7244
rect 739 6952 779 6992
rect 304 6784 672 6824
rect 1516 6364 1556 6404
rect 547 6280 587 6320
rect 1544 6028 1912 6068
rect 1516 5692 1556 5732
rect 739 5440 779 5480
rect 304 5272 672 5312
rect 2092 4852 2132 4892
rect 1123 4768 1163 4808
rect 1544 4516 1912 4556
rect 2092 4180 2132 4220
rect 1315 3928 1355 3968
rect 304 3760 672 3800
rect 2092 3340 2132 3380
rect 1123 3256 1163 3296
rect 1544 3004 1912 3044
rect 739 2836 779 2876
rect 1516 2668 1556 2708
rect 304 2248 672 2288
rect 1516 1828 1556 1868
rect 547 1744 587 1784
rect 1544 1492 1912 1532
rect 304 736 672 776
rect 1544 -20 1912 20
<< metal2 >>
rect 1535 25684 1544 25724
rect 1912 25684 1921 25724
rect 0 25052 100 25072
rect 0 25012 172 25052
rect 212 25012 221 25052
rect 0 24992 100 25012
rect 295 24928 304 24968
rect 672 24928 681 24968
rect 1535 24172 1544 24212
rect 1912 24172 1921 24212
rect 0 24128 100 24148
rect 0 24088 788 24128
rect 0 24068 100 24088
rect 748 24044 788 24088
rect 730 24004 739 24044
rect 779 24004 788 24044
rect 1507 23836 1516 23876
rect 1556 23836 2380 23876
rect 2420 23836 2429 23876
rect 295 23416 304 23456
rect 672 23416 681 23456
rect 0 23204 100 23224
rect 0 23164 739 23204
rect 779 23164 788 23204
rect 0 23144 100 23164
rect 1507 22996 1516 23036
rect 1556 22996 2284 23036
rect 2324 22996 2333 23036
rect 1535 22660 1544 22700
rect 1912 22660 1921 22700
rect 163 22408 172 22448
rect 212 22408 547 22448
rect 587 22408 596 22448
rect 1507 22324 1516 22364
rect 1556 22324 1996 22364
rect 2036 22324 2045 22364
rect 0 22280 100 22300
rect 0 22240 1132 22280
rect 1172 22240 1181 22280
rect 0 22220 100 22240
rect 295 21904 304 21944
rect 672 21904 681 21944
rect 1001 21568 1123 21608
rect 1172 21568 1181 21608
rect 2057 21484 2092 21524
rect 2132 21484 2188 21524
rect 2228 21484 2237 21524
rect 0 21356 100 21376
rect 0 21316 1132 21356
rect 1172 21316 1181 21356
rect 0 21296 100 21316
rect 1535 21148 1544 21188
rect 1912 21148 1921 21188
rect 2500 21104 2600 21124
rect 1987 21064 1996 21104
rect 2036 21064 2600 21104
rect 2500 21044 2600 21064
rect 1001 20896 1123 20936
rect 1172 20896 1181 20936
rect 1961 20812 2092 20852
rect 2132 20812 2141 20852
rect 2500 20684 2600 20704
rect 2371 20644 2380 20684
rect 2420 20644 2600 20684
rect 2500 20624 2600 20644
rect 0 20432 100 20452
rect 0 20392 212 20432
rect 295 20392 304 20432
rect 672 20392 681 20432
rect 0 20372 100 20392
rect 172 20264 212 20392
rect 2500 20264 2600 20284
rect 172 20224 739 20264
rect 779 20224 788 20264
rect 2275 20224 2284 20264
rect 2324 20224 2600 20264
rect 2500 20204 2600 20224
rect 1507 19972 1516 20012
rect 1556 19972 1996 20012
rect 2036 19972 2045 20012
rect 2500 19844 2600 19864
rect 2179 19804 2188 19844
rect 2228 19804 2600 19844
rect 2500 19784 2600 19804
rect 1535 19636 1544 19676
rect 1912 19636 1921 19676
rect 0 19508 100 19528
rect 0 19468 739 19508
rect 779 19468 788 19508
rect 0 19448 100 19468
rect 2500 19424 2600 19444
rect 2083 19384 2092 19424
rect 2132 19384 2600 19424
rect 2500 19364 2600 19384
rect 1385 19300 1516 19340
rect 1556 19300 1565 19340
rect 2500 19004 2600 19024
rect 1987 18964 1996 19004
rect 2036 18964 2600 19004
rect 2500 18944 2600 18964
rect 295 18880 304 18920
rect 672 18880 681 18920
rect 0 18584 100 18604
rect 2500 18584 2600 18604
rect 0 18544 547 18584
rect 587 18544 596 18584
rect 1507 18544 1516 18584
rect 1556 18544 2600 18584
rect 0 18524 100 18544
rect 2500 18524 2600 18544
rect 1507 18460 1516 18500
rect 1556 18460 2036 18500
rect 1996 18164 2036 18460
rect 2500 18164 2600 18184
rect 1535 18124 1544 18164
rect 1912 18124 1921 18164
rect 1996 18124 2600 18164
rect 2500 18104 2600 18124
rect 295 17368 304 17408
rect 672 17368 681 17408
rect 1535 16612 1544 16652
rect 1912 16612 1921 16652
rect 295 15856 304 15896
rect 672 15856 681 15896
rect 0 15812 100 15832
rect 0 15772 788 15812
rect 0 15752 100 15772
rect 748 15728 788 15772
rect 730 15688 739 15728
rect 779 15688 788 15728
rect 1507 15436 1516 15476
rect 1556 15436 1996 15476
rect 2036 15436 2045 15476
rect 1535 15100 1544 15140
rect 1912 15100 1921 15140
rect 0 14888 100 14908
rect 0 14848 547 14888
rect 587 14848 596 14888
rect 0 14828 100 14848
rect 1507 14764 1516 14804
rect 1556 14764 1708 14804
rect 1748 14764 1757 14804
rect 2500 14384 2600 14404
rect 295 14344 304 14384
rect 672 14344 681 14384
rect 1987 14344 1996 14384
rect 2036 14344 2600 14384
rect 2500 14324 2600 14344
rect 0 13964 100 13984
rect 2500 13964 2600 13984
rect 0 13924 547 13964
rect 587 13924 596 13964
rect 1507 13924 1516 13964
rect 1556 13924 1565 13964
rect 1699 13924 1708 13964
rect 1748 13924 2600 13964
rect 0 13904 100 13924
rect 1516 13880 1556 13924
rect 2500 13904 2600 13924
rect 1516 13840 2036 13880
rect 1535 13588 1544 13628
rect 1912 13588 1921 13628
rect 1996 13544 2036 13840
rect 2500 13544 2600 13564
rect 1996 13504 2600 13544
rect 2500 13484 2600 13504
rect 2083 13252 2092 13292
rect 2132 13252 2141 13292
rect 2092 13124 2132 13252
rect 2500 13124 2600 13144
rect 2092 13084 2600 13124
rect 2500 13064 2600 13084
rect 0 13040 100 13060
rect 0 13000 1315 13040
rect 1355 13000 1364 13040
rect 0 12980 100 13000
rect 295 12832 304 12872
rect 672 12832 681 12872
rect 2500 12704 2600 12724
rect 2092 12664 2600 12704
rect 2092 12452 2132 12664
rect 2500 12644 2600 12664
rect 2083 12412 2092 12452
rect 2132 12412 2141 12452
rect 2500 12284 2600 12304
rect 1306 12244 1315 12284
rect 1355 12244 1364 12284
rect 1987 12244 1996 12284
rect 2036 12244 2600 12284
rect 0 12116 100 12136
rect 1324 12116 1364 12244
rect 2500 12224 2600 12244
rect 0 12076 1364 12116
rect 1535 12076 1544 12116
rect 1912 12076 1921 12116
rect 0 12056 100 12076
rect 2500 11864 2600 11884
rect 1507 11824 1516 11864
rect 1556 11824 2600 11864
rect 2500 11804 2600 11824
rect 1507 11740 1516 11780
rect 1556 11740 1996 11780
rect 2036 11740 2045 11780
rect 730 11488 739 11528
rect 779 11488 788 11528
rect 295 11320 304 11360
rect 672 11320 681 11360
rect 0 11192 100 11212
rect 748 11192 788 11488
rect 2500 11444 2600 11464
rect 2083 11404 2092 11444
rect 2132 11404 2600 11444
rect 2500 11384 2600 11404
rect 0 11152 788 11192
rect 0 11132 100 11152
rect 1385 10900 1516 10940
rect 1556 10900 1565 10940
rect 425 10816 547 10856
rect 596 10816 605 10856
rect 1535 10564 1544 10604
rect 1912 10564 1921 10604
rect 0 10268 100 10288
rect 0 10228 556 10268
rect 596 10228 605 10268
rect 1961 10228 2092 10268
rect 2132 10228 2141 10268
rect 0 10208 100 10228
rect 1001 10144 1123 10184
rect 1172 10144 1181 10184
rect 295 9808 304 9848
rect 672 9808 681 9848
rect 0 9344 100 9364
rect 0 9304 1132 9344
rect 1172 9304 1181 9344
rect 0 9284 100 9304
rect 1535 9052 1544 9092
rect 1912 9052 1921 9092
rect 295 8296 304 8336
rect 672 8296 681 8336
rect 2500 7664 2600 7684
rect 1996 7624 2600 7664
rect 1535 7540 1544 7580
rect 1912 7540 1921 7580
rect 1996 7244 2036 7624
rect 2500 7604 2600 7624
rect 2500 7244 2600 7264
rect 1507 7204 1516 7244
rect 1556 7204 2036 7244
rect 2083 7204 2092 7244
rect 2132 7204 2600 7244
rect 2500 7184 2600 7204
rect 30 6952 739 6992
rect 779 6952 788 6992
rect 30 6740 70 6952
rect 2500 6824 2600 6844
rect 295 6784 304 6824
rect 672 6784 681 6824
rect 1987 6784 1996 6824
rect 2036 6784 2600 6824
rect 2500 6764 2600 6784
rect 30 6700 212 6740
rect 0 6572 100 6592
rect 172 6572 212 6700
rect 0 6532 212 6572
rect 0 6512 100 6532
rect 2500 6404 2600 6424
rect 1507 6364 1516 6404
rect 1556 6364 2092 6404
rect 2132 6364 2141 6404
rect 2275 6364 2284 6404
rect 2324 6364 2600 6404
rect 2500 6344 2600 6364
rect 259 6280 268 6320
rect 308 6280 547 6320
rect 587 6280 596 6320
rect 1535 6028 1544 6068
rect 1912 6028 1921 6068
rect 2500 5984 2600 6004
rect 2371 5944 2380 5984
rect 2420 5944 2600 5984
rect 2500 5924 2600 5944
rect 1507 5692 1516 5732
rect 1556 5692 1996 5732
rect 2036 5692 2045 5732
rect 0 5648 100 5668
rect 0 5608 268 5648
rect 308 5608 317 5648
rect 0 5588 100 5608
rect 2500 5564 2600 5584
rect 2083 5524 2092 5564
rect 2132 5524 2600 5564
rect 2500 5504 2600 5524
rect 617 5440 739 5480
rect 788 5440 797 5480
rect 295 5272 304 5312
rect 672 5272 681 5312
rect 2500 5144 2600 5164
rect 2179 5104 2188 5144
rect 2228 5104 2600 5144
rect 2500 5084 2600 5104
rect 1961 4852 2092 4892
rect 2132 4852 2141 4892
rect 835 4768 844 4808
rect 884 4768 1123 4808
rect 1163 4768 1172 4808
rect 0 4724 100 4744
rect 2500 4724 2600 4744
rect 0 4684 748 4724
rect 788 4684 797 4724
rect 1987 4684 1996 4724
rect 2036 4684 2600 4724
rect 0 4664 100 4684
rect 2500 4664 2600 4684
rect 1535 4516 1544 4556
rect 1912 4516 1921 4556
rect 2083 4180 2092 4220
rect 2132 4180 2284 4220
rect 2324 4180 2333 4220
rect 1306 3928 1315 3968
rect 1355 3928 1364 3968
rect 1324 3884 1364 3928
rect 172 3844 1364 3884
rect 0 3800 100 3820
rect 172 3800 212 3844
rect 0 3760 212 3800
rect 295 3760 304 3800
rect 672 3760 681 3800
rect 0 3740 100 3760
rect 2057 3340 2092 3380
rect 2132 3340 2188 3380
rect 2228 3340 2237 3380
rect 1001 3256 1123 3296
rect 1172 3256 1181 3296
rect 1535 3004 1544 3044
rect 1912 3004 1921 3044
rect 0 2876 100 2896
rect 0 2836 739 2876
rect 779 2836 788 2876
rect 0 2816 100 2836
rect 1507 2668 1516 2708
rect 1556 2668 2380 2708
rect 2420 2668 2429 2708
rect 295 2248 304 2288
rect 672 2248 681 2288
rect 0 1952 100 1972
rect 0 1912 844 1952
rect 884 1912 893 1952
rect 0 1892 100 1912
rect 1507 1828 1516 1868
rect 1556 1828 1996 1868
rect 2036 1828 2045 1868
rect 163 1744 172 1784
rect 212 1744 547 1784
rect 587 1744 596 1784
rect 1535 1492 1544 1532
rect 1912 1492 1921 1532
rect 0 1028 100 1048
rect 0 988 1132 1028
rect 1172 988 1181 1028
rect 0 968 100 988
rect 295 736 304 776
rect 672 736 681 776
rect 0 104 100 124
rect 0 64 172 104
rect 212 64 221 104
rect 0 44 100 64
rect 1535 -20 1544 20
rect 1912 -20 1921 20
<< via2 >>
rect 1544 25684 1912 25724
rect 172 25012 212 25052
rect 304 24928 672 24968
rect 1544 24172 1912 24212
rect 2380 23836 2420 23876
rect 304 23416 672 23456
rect 2284 22996 2324 23036
rect 1544 22660 1912 22700
rect 172 22408 212 22448
rect 1996 22324 2036 22364
rect 1132 22240 1172 22280
rect 304 21904 672 21944
rect 1132 21568 1163 21608
rect 1163 21568 1172 21608
rect 2188 21484 2228 21524
rect 1132 21316 1172 21356
rect 1544 21148 1912 21188
rect 1996 21064 2036 21104
rect 1132 20896 1163 20936
rect 1163 20896 1172 20936
rect 2092 20812 2132 20852
rect 2380 20644 2420 20684
rect 304 20392 672 20432
rect 2284 20224 2324 20264
rect 1996 19972 2036 20012
rect 2188 19804 2228 19844
rect 1544 19636 1912 19676
rect 2092 19384 2132 19424
rect 1516 19300 1556 19340
rect 1996 18964 2036 19004
rect 304 18880 672 18920
rect 1516 18544 1556 18584
rect 1544 18124 1912 18164
rect 304 17368 672 17408
rect 1544 16612 1912 16652
rect 304 15856 672 15896
rect 1996 15436 2036 15476
rect 1544 15100 1912 15140
rect 1708 14764 1748 14804
rect 304 14344 672 14384
rect 1996 14344 2036 14384
rect 1708 13924 1748 13964
rect 1544 13588 1912 13628
rect 304 12832 672 12872
rect 1996 12244 2036 12284
rect 1544 12076 1912 12116
rect 1516 11824 1556 11864
rect 1996 11740 2036 11780
rect 304 11320 672 11360
rect 2092 11404 2132 11444
rect 1516 10900 1556 10940
rect 556 10816 587 10856
rect 587 10816 596 10856
rect 1544 10564 1912 10604
rect 556 10228 596 10268
rect 2092 10228 2132 10268
rect 1132 10144 1163 10184
rect 1163 10144 1172 10184
rect 304 9808 672 9848
rect 1132 9304 1172 9344
rect 1544 9052 1912 9092
rect 304 8296 672 8336
rect 1544 7540 1912 7580
rect 2092 7204 2132 7244
rect 304 6784 672 6824
rect 1996 6784 2036 6824
rect 2092 6364 2132 6404
rect 2284 6364 2324 6404
rect 268 6280 308 6320
rect 1544 6028 1912 6068
rect 2380 5944 2420 5984
rect 1996 5692 2036 5732
rect 268 5608 308 5648
rect 2092 5524 2132 5564
rect 748 5440 779 5480
rect 779 5440 788 5480
rect 304 5272 672 5312
rect 2188 5104 2228 5144
rect 2092 4852 2132 4892
rect 844 4768 884 4808
rect 748 4684 788 4724
rect 1996 4684 2036 4724
rect 1544 4516 1912 4556
rect 2284 4180 2324 4220
rect 304 3760 672 3800
rect 2188 3340 2228 3380
rect 1132 3256 1163 3296
rect 1163 3256 1172 3296
rect 1544 3004 1912 3044
rect 2380 2668 2420 2708
rect 304 2248 672 2288
rect 844 1912 884 1952
rect 1996 1828 2036 1868
rect 172 1744 212 1784
rect 1544 1492 1912 1532
rect 1132 988 1172 1028
rect 304 736 672 776
rect 172 64 212 104
rect 1544 -20 1912 20
<< metal3 >>
rect 1544 25724 1912 25733
rect 1544 25675 1912 25684
rect 172 25052 212 25061
rect 172 22448 212 25012
rect 304 24968 672 24977
rect 304 24919 672 24928
rect 1544 24212 1912 24221
rect 1544 24163 1912 24172
rect 2380 23876 2420 23885
rect 304 23456 672 23465
rect 304 23407 672 23416
rect 2284 23036 2324 23045
rect 1544 22700 1912 22709
rect 1544 22651 1912 22660
rect 172 22399 212 22408
rect 1996 22364 2036 22373
rect 1132 22280 1172 22289
rect 304 21944 672 21953
rect 304 21895 672 21904
rect 1132 21608 1172 22240
rect 1132 21559 1172 21568
rect 1132 21356 1172 21365
rect 1132 20936 1172 21316
rect 1544 21188 1912 21197
rect 1544 21139 1912 21148
rect 1996 21104 2036 22324
rect 1996 21055 2036 21064
rect 2188 21524 2228 21533
rect 1132 20887 1172 20896
rect 2092 20852 2132 20861
rect 304 20432 672 20441
rect 304 20383 672 20392
rect 1996 20012 2036 20021
rect 1544 19676 1912 19685
rect 1544 19627 1912 19636
rect 1516 19340 1556 19349
rect 304 18920 672 18929
rect 304 18871 672 18880
rect 1516 18584 1556 19300
rect 1996 19004 2036 19972
rect 2092 19424 2132 20812
rect 2188 19844 2228 21484
rect 2284 20264 2324 22996
rect 2380 20684 2420 23836
rect 2380 20635 2420 20644
rect 2284 20215 2324 20224
rect 2188 19795 2228 19804
rect 2092 19375 2132 19384
rect 1996 18955 2036 18964
rect 1516 18535 1556 18544
rect 1544 18164 1912 18173
rect 1544 18115 1912 18124
rect 304 17408 672 17417
rect 304 17359 672 17368
rect 1544 16652 1912 16661
rect 1544 16603 1912 16612
rect 304 15896 672 15905
rect 304 15847 672 15856
rect 1996 15476 2036 15485
rect 1544 15140 1912 15149
rect 1544 15091 1912 15100
rect 1708 14804 1748 14813
rect 304 14384 672 14393
rect 304 14335 672 14344
rect 1708 13964 1748 14764
rect 1996 14384 2036 15436
rect 1996 14335 2036 14344
rect 1708 13915 1748 13924
rect 1544 13628 1912 13637
rect 1544 13579 1912 13588
rect 304 12872 672 12881
rect 304 12823 672 12832
rect 1996 12284 2036 12293
rect 1544 12116 1912 12125
rect 1544 12067 1912 12076
rect 1516 11864 1556 11873
rect 304 11360 672 11369
rect 304 11311 672 11320
rect 1516 10940 1556 11824
rect 1996 11780 2036 12244
rect 1996 11731 2036 11740
rect 1516 10891 1556 10900
rect 2092 11444 2132 11453
rect 556 10856 596 10865
rect 556 10268 596 10816
rect 1544 10604 1912 10613
rect 1544 10555 1912 10564
rect 556 10219 596 10228
rect 2092 10268 2132 11404
rect 2092 10219 2132 10228
rect 1132 10184 1172 10193
rect 304 9848 672 9857
rect 304 9799 672 9808
rect 1132 9344 1172 10144
rect 1132 9295 1172 9304
rect 1544 9092 1912 9101
rect 1544 9043 1912 9052
rect 304 8336 672 8345
rect 304 8287 672 8296
rect 1544 7580 1912 7589
rect 1544 7531 1912 7540
rect 2092 7244 2132 7253
rect 304 6824 672 6833
rect 304 6775 672 6784
rect 1996 6824 2036 6833
rect 268 6320 308 6329
rect 268 5648 308 6280
rect 1544 6068 1912 6077
rect 1544 6019 1912 6028
rect 1996 5732 2036 6784
rect 2092 6404 2132 7204
rect 2092 6355 2132 6364
rect 2284 6404 2324 6413
rect 1996 5683 2036 5692
rect 268 5599 308 5608
rect 2092 5564 2132 5573
rect 748 5480 788 5489
rect 304 5312 672 5321
rect 304 5263 672 5272
rect 748 4724 788 5440
rect 2092 4892 2132 5524
rect 2092 4843 2132 4852
rect 2188 5144 2228 5153
rect 748 4675 788 4684
rect 844 4808 884 4817
rect 304 3800 672 3809
rect 304 3751 672 3760
rect 304 2288 672 2297
rect 304 2239 672 2248
rect 844 1952 884 4768
rect 1996 4724 2036 4733
rect 1544 4556 1912 4565
rect 1544 4507 1912 4516
rect 844 1903 884 1912
rect 1132 3296 1172 3305
rect 172 1784 212 1793
rect 172 104 212 1744
rect 1132 1028 1172 3256
rect 1544 3044 1912 3053
rect 1544 2995 1912 3004
rect 1996 1868 2036 4684
rect 2188 3380 2228 5104
rect 2284 4220 2324 6364
rect 2284 4171 2324 4180
rect 2380 5984 2420 5993
rect 2188 3331 2228 3340
rect 2380 2708 2420 5944
rect 2380 2659 2420 2668
rect 1996 1819 2036 1828
rect 1544 1532 1912 1541
rect 1544 1483 1912 1492
rect 1132 979 1172 988
rect 304 776 672 785
rect 304 727 672 736
rect 172 55 212 64
rect 1544 20 1912 29
rect 1544 -29 1912 -20
<< via3 >>
rect 1544 25684 1912 25724
rect 304 24928 672 24968
rect 1544 24172 1912 24212
rect 304 23416 672 23456
rect 1544 22660 1912 22700
rect 304 21904 672 21944
rect 1544 21148 1912 21188
rect 304 20392 672 20432
rect 1544 19636 1912 19676
rect 304 18880 672 18920
rect 1544 18124 1912 18164
rect 304 17368 672 17408
rect 1544 16612 1912 16652
rect 304 15856 672 15896
rect 1544 15100 1912 15140
rect 304 14344 672 14384
rect 1544 13588 1912 13628
rect 304 12832 672 12872
rect 1544 12076 1912 12116
rect 304 11320 672 11360
rect 1544 10564 1912 10604
rect 304 9808 672 9848
rect 1544 9052 1912 9092
rect 304 8296 672 8336
rect 1544 7540 1912 7580
rect 304 6784 672 6824
rect 1544 6028 1912 6068
rect 304 5272 672 5312
rect 304 3760 672 3800
rect 304 2248 672 2288
rect 1544 4516 1912 4556
rect 1544 3004 1912 3044
rect 1544 1492 1912 1532
rect 304 736 672 776
rect 1544 -20 1912 20
<< metal4 >>
rect 1535 25684 1544 25724
rect 1912 25684 1921 25724
rect 295 24928 304 24968
rect 672 24928 681 24968
rect 1535 24172 1544 24212
rect 1912 24172 1921 24212
rect 295 23416 304 23456
rect 672 23416 681 23456
rect 1535 22660 1544 22700
rect 1912 22660 1921 22700
rect 295 21904 304 21944
rect 672 21904 681 21944
rect 1535 21148 1544 21188
rect 1912 21148 1921 21188
rect 295 20392 304 20432
rect 672 20392 681 20432
rect 1535 19636 1544 19676
rect 1912 19636 1921 19676
rect 295 18880 304 18920
rect 672 18880 681 18920
rect 1535 18124 1544 18164
rect 1912 18124 1921 18164
rect 295 17368 304 17408
rect 672 17368 681 17408
rect 1535 16612 1544 16652
rect 1912 16612 1921 16652
rect 295 15856 304 15896
rect 672 15856 681 15896
rect 1535 15100 1544 15140
rect 1912 15100 1921 15140
rect 295 14344 304 14384
rect 672 14344 681 14384
rect 1535 13588 1544 13628
rect 1912 13588 1921 13628
rect 295 12832 304 12872
rect 672 12832 681 12872
rect 1535 12076 1544 12116
rect 1912 12076 1921 12116
rect 295 11320 304 11360
rect 672 11320 681 11360
rect 1535 10564 1544 10604
rect 1912 10564 1921 10604
rect 295 9808 304 9848
rect 672 9808 681 9848
rect 1535 9052 1544 9092
rect 1912 9052 1921 9092
rect 295 8296 304 8336
rect 672 8296 681 8336
rect 1535 7540 1544 7580
rect 1912 7540 1921 7580
rect 295 6784 304 6824
rect 672 6784 681 6824
rect 1535 6028 1544 6068
rect 1912 6028 1921 6068
rect 295 5272 304 5312
rect 672 5272 681 5312
rect 1535 4516 1544 4556
rect 1912 4516 1921 4556
rect 295 3760 304 3800
rect 672 3760 681 3800
rect 1535 3004 1544 3044
rect 1912 3004 1921 3044
rect 295 2248 304 2288
rect 672 2248 681 2288
rect 1535 1492 1544 1532
rect 1912 1492 1921 1532
rect 295 736 304 776
rect 672 736 681 776
rect 1535 -20 1544 20
rect 1912 -20 1921 20
<< via4 >>
rect 1544 25684 1912 25724
rect 304 24928 672 24968
rect 1544 24172 1912 24212
rect 304 23416 672 23456
rect 1544 22660 1912 22700
rect 304 21904 672 21944
rect 1544 21148 1912 21188
rect 304 20392 672 20432
rect 1544 19636 1912 19676
rect 304 18880 672 18920
rect 1544 18124 1912 18164
rect 304 17368 672 17408
rect 1544 16612 1912 16652
rect 304 15856 672 15896
rect 1544 15100 1912 15140
rect 304 14344 672 14384
rect 1544 13588 1912 13628
rect 304 12832 672 12872
rect 1544 12076 1912 12116
rect 304 11320 672 11360
rect 1544 10564 1912 10604
rect 304 9808 672 9848
rect 1544 9052 1912 9092
rect 304 8296 672 8336
rect 1544 7540 1912 7580
rect 304 6784 672 6824
rect 1544 6028 1912 6068
rect 304 5272 672 5312
rect 1544 4516 1912 4556
rect 304 3760 672 3800
rect 1544 3004 1912 3044
rect 304 2248 672 2288
rect 1544 1492 1912 1532
rect 304 736 672 776
rect 1544 -20 1912 20
<< metal5 >>
rect 268 24968 708 25748
rect 268 24928 304 24968
rect 672 24928 708 24968
rect 268 23456 708 24928
rect 268 23416 304 23456
rect 672 23416 708 23456
rect 268 21944 708 23416
rect 268 21904 304 21944
rect 672 21904 708 21944
rect 268 20432 708 21904
rect 268 20392 304 20432
rect 672 20392 708 20432
rect 268 18920 708 20392
rect 268 18880 304 18920
rect 672 18880 708 18920
rect 268 17408 708 18880
rect 268 17368 304 17408
rect 672 17368 708 17408
rect 268 15896 708 17368
rect 268 15856 304 15896
rect 672 15856 708 15896
rect 268 14384 708 15856
rect 268 14344 304 14384
rect 672 14344 708 14384
rect 268 12872 708 14344
rect 268 12832 304 12872
rect 672 12832 708 12872
rect 268 11360 708 12832
rect 268 11320 304 11360
rect 672 11320 708 11360
rect 268 9848 708 11320
rect 268 9808 304 9848
rect 672 9808 708 9848
rect 268 8336 708 9808
rect 268 8296 304 8336
rect 672 8296 708 8336
rect 268 6824 708 8296
rect 268 6784 304 6824
rect 672 6784 708 6824
rect 268 5312 708 6784
rect 268 5272 304 5312
rect 672 5272 708 5312
rect 268 3800 708 5272
rect 268 3760 304 3800
rect 672 3760 708 3800
rect 268 2288 708 3760
rect 268 2248 304 2288
rect 672 2248 708 2288
rect 268 776 708 2248
rect 268 736 304 776
rect 672 736 708 776
rect 268 -44 708 736
rect 1508 25724 1948 25748
rect 1508 25684 1544 25724
rect 1912 25684 1948 25724
rect 1508 24212 1948 25684
rect 1508 24172 1544 24212
rect 1912 24172 1948 24212
rect 1508 22700 1948 24172
rect 1508 22660 1544 22700
rect 1912 22660 1948 22700
rect 1508 21188 1948 22660
rect 1508 21148 1544 21188
rect 1912 21148 1948 21188
rect 1508 19676 1948 21148
rect 1508 19636 1544 19676
rect 1912 19636 1948 19676
rect 1508 18164 1948 19636
rect 1508 18124 1544 18164
rect 1912 18124 1948 18164
rect 1508 16652 1948 18124
rect 1508 16612 1544 16652
rect 1912 16612 1948 16652
rect 1508 15140 1948 16612
rect 1508 15100 1544 15140
rect 1912 15100 1948 15140
rect 1508 13628 1948 15100
rect 1508 13588 1544 13628
rect 1912 13588 1948 13628
rect 1508 12116 1948 13588
rect 1508 12076 1544 12116
rect 1912 12076 1948 12116
rect 1508 10604 1948 12076
rect 1508 10564 1544 10604
rect 1912 10564 1948 10604
rect 1508 9092 1948 10564
rect 1508 9052 1544 9092
rect 1912 9052 1948 9092
rect 1508 7580 1948 9052
rect 1508 7540 1544 7580
rect 1912 7540 1948 7580
rect 1508 6068 1948 7540
rect 1508 6028 1544 6068
rect 1912 6028 1948 6068
rect 1508 4556 1948 6028
rect 1508 4516 1544 4556
rect 1912 4516 1948 4556
rect 1508 3044 1948 4516
rect 1508 3004 1544 3044
rect 1912 3004 1948 3044
rect 1508 1532 1948 3004
rect 1508 1492 1544 1532
rect 1912 1492 1948 1532
rect 1508 20 1948 1492
rect 1508 -20 1544 20
rect 1912 -20 1948 20
rect 1508 -44 1948 -20
use sg13g2_decap_8  FILLER_0_0
timestamp 1746816402
transform 1 0 288 0 1 0
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_7
timestamp 1746816402
transform 1 0 960 0 1 0
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_14
timestamp 1746816402
transform 1 0 1632 0 1 0
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_0
timestamp 1746816402
transform 1 0 288 0 -1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_7
timestamp 1746816402
transform 1 0 960 0 -1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_14
timestamp 1746816402
transform 1 0 1632 0 -1 1512
box -48 -56 720 834
use sg13g2_fill_1  FILLER_2_0
timestamp 1746816402
transform 1 0 288 0 1 1512
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_14
timestamp 1746816402
transform 1 0 1632 0 1 1512
box -48 -56 720 834
use sg13g2_fill_1  FILLER_3_0
timestamp 1746816402
transform 1 0 288 0 -1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_14
timestamp 1746816402
transform 1 0 1632 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_0
timestamp 1746816402
transform 1 0 288 0 1 3024
box -48 -56 720 834
use sg13g2_fill_1  FILLER_4_20
timestamp 1746816402
transform 1 0 2208 0 1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_0
timestamp 1746816402
transform 1 0 288 0 -1 4536
box -48 -56 720 834
use sg13g2_fill_1  FILLER_5_20
timestamp 1746816402
transform 1 0 2208 0 -1 4536
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_0
timestamp 1746816402
transform 1 0 288 0 1 4536
box -48 -56 720 834
use sg13g2_fill_1  FILLER_6_20
timestamp 1746816402
transform 1 0 2208 0 1 4536
box -48 -56 144 834
use sg13g2_fill_1  FILLER_7_0
timestamp 1746816402
transform 1 0 288 0 -1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_14
timestamp 1746816402
transform 1 0 1632 0 -1 6048
box -48 -56 720 834
use sg13g2_fill_1  FILLER_8_0
timestamp 1746816402
transform 1 0 288 0 1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_14
timestamp 1746816402
transform 1 0 1632 0 1 6048
box -48 -56 720 834
use sg13g2_fill_1  FILLER_9_0
timestamp 1746816402
transform 1 0 288 0 -1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_14
timestamp 1746816402
transform 1 0 1632 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_0
timestamp 1746816402
transform 1 0 288 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_7
timestamp 1746816402
transform 1 0 960 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_14
timestamp 1746816402
transform 1 0 1632 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_0
timestamp 1746816402
transform 1 0 288 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_7
timestamp 1746816402
transform 1 0 960 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_14
timestamp 1746816402
transform 1 0 1632 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_0
timestamp 1746816402
transform 1 0 288 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_7
timestamp 1746816402
transform 1 0 960 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_14
timestamp 1746816402
transform 1 0 1632 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_0
timestamp 1746816402
transform 1 0 288 0 -1 10584
box -48 -56 720 834
use sg13g2_fill_1  FILLER_13_20
timestamp 1746816402
transform 1 0 2208 0 -1 10584
box -48 -56 144 834
use sg13g2_fill_1  FILLER_14_0
timestamp 1746816402
transform 1 0 288 0 1 10584
box -48 -56 144 834
use sg13g2_decap_8  FILLER_14_14
timestamp 1746816402
transform 1 0 1632 0 1 10584
box -48 -56 720 834
use sg13g2_fill_1  FILLER_15_0
timestamp 1746816402
transform 1 0 288 0 -1 12096
box -48 -56 144 834
use sg13g2_decap_8  FILLER_15_14
timestamp 1746816402
transform 1 0 1632 0 -1 12096
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_0
timestamp 1746816402
transform 1 0 288 0 1 12096
box -48 -56 720 834
use sg13g2_fill_1  FILLER_16_20
timestamp 1746816402
transform 1 0 2208 0 1 12096
box -48 -56 144 834
use sg13g2_decap_8  FILLER_17_0
timestamp 1746816402
transform 1 0 288 0 -1 13608
box -48 -56 720 834
use sg13g2_fill_1  FILLER_17_20
timestamp 1746816402
transform 1 0 2208 0 -1 13608
box -48 -56 144 834
use sg13g2_fill_1  FILLER_18_0
timestamp 1746816402
transform 1 0 288 0 1 13608
box -48 -56 144 834
use sg13g2_decap_8  FILLER_18_14
timestamp 1746816402
transform 1 0 1632 0 1 13608
box -48 -56 720 834
use sg13g2_fill_1  FILLER_19_0
timestamp 1746816402
transform 1 0 288 0 -1 15120
box -48 -56 144 834
use sg13g2_decap_8  FILLER_19_14
timestamp 1746816402
transform 1 0 1632 0 -1 15120
box -48 -56 720 834
use sg13g2_fill_1  FILLER_20_0
timestamp 1746816402
transform 1 0 288 0 1 15120
box -48 -56 144 834
use sg13g2_decap_8  FILLER_20_14
timestamp 1746816402
transform 1 0 1632 0 1 15120
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_0
timestamp 1746816402
transform 1 0 288 0 -1 16632
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_7
timestamp 1746816402
transform 1 0 960 0 -1 16632
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_14
timestamp 1746816402
transform 1 0 1632 0 -1 16632
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_0
timestamp 1746816402
transform 1 0 288 0 1 16632
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_7
timestamp 1746816402
transform 1 0 960 0 1 16632
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_14
timestamp 1746816402
transform 1 0 1632 0 1 16632
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_0
timestamp 1746816402
transform 1 0 288 0 -1 18144
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_7
timestamp 1746816402
transform 1 0 960 0 -1 18144
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_14
timestamp 1746816402
transform 1 0 1632 0 -1 18144
box -48 -56 720 834
use sg13g2_fill_1  FILLER_24_0
timestamp 1746816402
transform 1 0 288 0 1 18144
box -48 -56 144 834
use sg13g2_decap_8  FILLER_24_14
timestamp 1746816402
transform 1 0 1632 0 1 18144
box -48 -56 720 834
use sg13g2_fill_1  FILLER_25_0
timestamp 1746816402
transform 1 0 288 0 -1 19656
box -48 -56 144 834
use sg13g2_decap_8  FILLER_25_14
timestamp 1746816402
transform 1 0 1632 0 -1 19656
box -48 -56 720 834
use sg13g2_fill_1  FILLER_26_0
timestamp 1746816402
transform 1 0 288 0 1 19656
box -48 -56 144 834
use sg13g2_decap_8  FILLER_26_14
timestamp 1746816402
transform 1 0 1632 0 1 19656
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_0
timestamp 1746816402
transform 1 0 288 0 -1 21168
box -48 -56 720 834
use sg13g2_fill_1  FILLER_27_20
timestamp 1746816402
transform 1 0 2208 0 -1 21168
box -48 -56 144 834
use sg13g2_decap_8  FILLER_28_0
timestamp 1746816402
transform 1 0 288 0 1 21168
box -48 -56 720 834
use sg13g2_fill_1  FILLER_28_20
timestamp 1746816402
transform 1 0 2208 0 1 21168
box -48 -56 144 834
use sg13g2_fill_1  FILLER_29_0
timestamp 1746816402
transform 1 0 288 0 -1 22680
box -48 -56 144 834
use sg13g2_decap_8  FILLER_29_14
timestamp 1746816402
transform 1 0 1632 0 -1 22680
box -48 -56 720 834
use sg13g2_fill_1  FILLER_30_0
timestamp 1746816402
transform 1 0 288 0 1 22680
box -48 -56 144 834
use sg13g2_decap_8  FILLER_30_14
timestamp 1746816402
transform 1 0 1632 0 1 22680
box -48 -56 720 834
use sg13g2_fill_1  FILLER_31_0
timestamp 1746816402
transform 1 0 288 0 -1 24192
box -48 -56 144 834
use sg13g2_decap_8  FILLER_31_14
timestamp 1746816402
transform 1 0 1632 0 -1 24192
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_0
timestamp 1746816402
transform 1 0 288 0 1 24192
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_7
timestamp 1746816402
transform 1 0 960 0 1 24192
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_14
timestamp 1746816402
transform 1 0 1632 0 1 24192
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_0
timestamp 1746816402
transform 1 0 288 0 -1 25704
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_7
timestamp 1746816402
transform 1 0 960 0 -1 25704
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_14
timestamp 1746816402
transform 1 0 1632 0 -1 25704
box -48 -56 720 834
use sg13g2_buf_8  rgb_buffer_cell\[0\]
timestamp 1746816402
transform -1 0 1632 0 -1 7560
box -48 -56 1296 834
use sg13g2_buf_8  rgb_buffer_cell\[1\]
timestamp 1746816402
transform -1 0 1632 0 1 6048
box -48 -56 1296 834
use sg13g2_buf_8  rgb_buffer_cell\[2\]
timestamp 1746816402
transform -1 0 1632 0 -1 6048
box -48 -56 1296 834
use sg13g2_buf_8  rgb_buffer_cell\[3\]
timestamp 1746816402
transform -1 0 2208 0 -1 4536
box -48 -56 1296 834
use sg13g2_buf_8  rgb_buffer_cell\[4\]
timestamp 1746816402
transform -1 0 1632 0 -1 3024
box -48 -56 1296 834
use sg13g2_buf_8  rgb_buffer_cell\[5\]
timestamp 1746816402
transform -1 0 2208 0 1 4536
box -48 -56 1296 834
use sg13g2_buf_8  rgb_buffer_cell\[6\]
timestamp 1746816402
transform -1 0 2208 0 1 3024
box -48 -56 1296 834
use sg13g2_buf_8  rgb_buffer_cell\[7\]
timestamp 1746816402
transform -1 0 1632 0 1 1512
box -48 -56 1296 834
use sg13g2_buf_8  rgb_buffer_cell\[8\]
timestamp 1746816402
transform -1 0 1632 0 1 15120
box -48 -56 1296 834
use sg13g2_buf_8  rgb_buffer_cell\[9\]
timestamp 1746816402
transform -1 0 1632 0 -1 15120
box -48 -56 1296 834
use sg13g2_buf_8  rgb_buffer_cell\[10\]
timestamp 1746816402
transform -1 0 1632 0 1 13608
box -48 -56 1296 834
use sg13g2_buf_8  rgb_buffer_cell\[11\]
timestamp 1746816402
transform -1 0 2208 0 -1 13608
box -48 -56 1296 834
use sg13g2_buf_8  rgb_buffer_cell\[12\]
timestamp 1746816402
transform -1 0 2208 0 1 12096
box -48 -56 1296 834
use sg13g2_buf_8  rgb_buffer_cell\[13\]
timestamp 1746816402
transform -1 0 1632 0 -1 12096
box -48 -56 1296 834
use sg13g2_buf_8  rgb_buffer_cell\[14\]
timestamp 1746816402
transform -1 0 1632 0 1 10584
box -48 -56 1296 834
use sg13g2_buf_8  rgb_buffer_cell\[15\]
timestamp 1746816402
transform -1 0 2208 0 -1 10584
box -48 -56 1296 834
use sg13g2_buf_8  rgb_buffer_cell\[16\]
timestamp 1746816402
transform -1 0 1632 0 -1 22680
box -48 -56 1296 834
use sg13g2_buf_8  rgb_buffer_cell\[17\]
timestamp 1746816402
transform -1 0 1632 0 -1 24192
box -48 -56 1296 834
use sg13g2_buf_8  rgb_buffer_cell\[18\]
timestamp 1746816402
transform -1 0 1632 0 1 22680
box -48 -56 1296 834
use sg13g2_buf_8  rgb_buffer_cell\[19\]
timestamp 1746816402
transform -1 0 2208 0 1 21168
box -48 -56 1296 834
use sg13g2_buf_8  rgb_buffer_cell\[20\]
timestamp 1746816402
transform -1 0 2208 0 -1 21168
box -48 -56 1296 834
use sg13g2_buf_8  rgb_buffer_cell\[21\]
timestamp 1746816402
transform -1 0 1632 0 1 19656
box -48 -56 1296 834
use sg13g2_buf_8  rgb_buffer_cell\[22\]
timestamp 1746816402
transform -1 0 1632 0 -1 19656
box -48 -56 1296 834
use sg13g2_buf_8  rgb_buffer_cell\[23\]
timestamp 1746816402
transform -1 0 1632 0 1 18144
box -48 -56 1296 834
<< labels >>
flabel metal5 s 1508 -44 1948 25748 0 FreeSans 3200 90 0 0 VGND
port 1 nsew
flabel metal5 s 268 -44 708 25748 0 FreeSans 3200 90 0 0 VPWR
port 2 nsew
flabel metal2 s 0 6512 100 6592 0 FreeSans 400 0 0 0 b[0]
port 3 nsew
flabel metal2 s 0 5588 100 5668 0 FreeSans 400 0 0 0 b[1]
port 4 nsew
flabel metal2 s 0 4664 100 4744 0 FreeSans 400 0 0 0 b[2]
port 5 nsew
flabel metal2 s 0 3740 100 3820 0 FreeSans 400 0 0 0 b[3]
port 6 nsew
flabel metal2 s 0 2816 100 2896 0 FreeSans 400 0 0 0 b[4]
port 7 nsew
flabel metal2 s 0 1892 100 1972 0 FreeSans 400 0 0 0 b[5]
port 8 nsew
flabel metal2 s 0 968 100 1048 0 FreeSans 400 0 0 0 b[6]
port 9 nsew
flabel metal2 s 0 44 100 124 0 FreeSans 400 0 0 0 b[7]
port 10 nsew
flabel metal2 s 2500 7604 2600 7684 0 FreeSans 400 0 0 0 db[0]
port 11 nsew
flabel metal2 s 2500 7184 2600 7264 0 FreeSans 400 0 0 0 db[1]
port 12 nsew
flabel metal2 s 2500 6764 2600 6844 0 FreeSans 400 0 0 0 db[2]
port 13 nsew
flabel metal2 s 2500 6344 2600 6424 0 FreeSans 400 0 0 0 db[3]
port 14 nsew
flabel metal2 s 2500 5924 2600 6004 0 FreeSans 400 0 0 0 db[4]
port 15 nsew
flabel metal2 s 2500 5504 2600 5584 0 FreeSans 400 0 0 0 db[5]
port 16 nsew
flabel metal2 s 2500 5084 2600 5164 0 FreeSans 400 0 0 0 db[6]
port 17 nsew
flabel metal2 s 2500 4664 2600 4744 0 FreeSans 400 0 0 0 db[7]
port 18 nsew
flabel metal2 s 2500 14324 2600 14404 0 FreeSans 400 0 0 0 dg[0]
port 19 nsew
flabel metal2 s 2500 13904 2600 13984 0 FreeSans 400 0 0 0 dg[1]
port 20 nsew
flabel metal2 s 2500 13484 2600 13564 0 FreeSans 400 0 0 0 dg[2]
port 21 nsew
flabel metal2 s 2500 13064 2600 13144 0 FreeSans 400 0 0 0 dg[3]
port 22 nsew
flabel metal2 s 2500 12644 2600 12724 0 FreeSans 400 0 0 0 dg[4]
port 23 nsew
flabel metal2 s 2500 12224 2600 12304 0 FreeSans 400 0 0 0 dg[5]
port 24 nsew
flabel metal2 s 2500 11804 2600 11884 0 FreeSans 400 0 0 0 dg[6]
port 25 nsew
flabel metal2 s 2500 11384 2600 11464 0 FreeSans 400 0 0 0 dg[7]
port 26 nsew
flabel metal2 s 2500 21044 2600 21124 0 FreeSans 400 0 0 0 dr[0]
port 27 nsew
flabel metal2 s 2500 20624 2600 20704 0 FreeSans 400 0 0 0 dr[1]
port 28 nsew
flabel metal2 s 2500 20204 2600 20284 0 FreeSans 400 0 0 0 dr[2]
port 29 nsew
flabel metal2 s 2500 19784 2600 19864 0 FreeSans 400 0 0 0 dr[3]
port 30 nsew
flabel metal2 s 2500 19364 2600 19444 0 FreeSans 400 0 0 0 dr[4]
port 31 nsew
flabel metal2 s 2500 18944 2600 19024 0 FreeSans 400 0 0 0 dr[5]
port 32 nsew
flabel metal2 s 2500 18524 2600 18604 0 FreeSans 400 0 0 0 dr[6]
port 33 nsew
flabel metal2 s 2500 18104 2600 18184 0 FreeSans 400 0 0 0 dr[7]
port 34 nsew
flabel metal2 s 0 15752 100 15832 0 FreeSans 400 0 0 0 g[0]
port 35 nsew
flabel metal2 s 0 14828 100 14908 0 FreeSans 400 0 0 0 g[1]
port 36 nsew
flabel metal2 s 0 13904 100 13984 0 FreeSans 400 0 0 0 g[2]
port 37 nsew
flabel metal2 s 0 12980 100 13060 0 FreeSans 400 0 0 0 g[3]
port 38 nsew
flabel metal2 s 0 12056 100 12136 0 FreeSans 400 0 0 0 g[4]
port 39 nsew
flabel metal2 s 0 11132 100 11212 0 FreeSans 400 0 0 0 g[5]
port 40 nsew
flabel metal2 s 0 10208 100 10288 0 FreeSans 400 0 0 0 g[6]
port 41 nsew
flabel metal2 s 0 9284 100 9364 0 FreeSans 400 0 0 0 g[7]
port 42 nsew
flabel metal2 s 0 24992 100 25072 0 FreeSans 400 0 0 0 r[0]
port 43 nsew
flabel metal2 s 0 24068 100 24148 0 FreeSans 400 0 0 0 r[1]
port 44 nsew
flabel metal2 s 0 23144 100 23224 0 FreeSans 400 0 0 0 r[2]
port 45 nsew
flabel metal2 s 0 22220 100 22300 0 FreeSans 400 0 0 0 r[3]
port 46 nsew
flabel metal2 s 0 21296 100 21376 0 FreeSans 400 0 0 0 r[4]
port 47 nsew
flabel metal2 s 0 20372 100 20452 0 FreeSans 400 0 0 0 r[5]
port 48 nsew
flabel metal2 s 0 19448 100 19528 0 FreeSans 400 0 0 0 r[6]
port 49 nsew
flabel metal2 s 0 18524 100 18604 0 FreeSans 400 0 0 0 r[7]
port 50 nsew
<< properties >>
string FIXED_BBOX 0 0 2600 26000
string GDS_END 107254
string GDS_FILE ../gds/rgb_buffers.gds
string GDS_START 14954
<< end >>
