magic
tech ihp-sg13g2
timestamp 1747537721
<< nwell >>
rect -24 175 600 417
<< pwell >>
rect 9 28 576 157
rect -13 -28 589 28
<< nmos >>
rect 57 70 70 144
rect 108 70 121 144
rect 210 70 223 144
rect 261 70 274 144
rect 312 70 325 144
rect 363 70 376 144
rect 465 70 478 144
rect 516 70 529 144
<< pmos >>
rect 57 206 70 318
rect 108 206 121 318
rect 210 206 223 318
rect 261 206 274 318
rect 312 206 325 318
rect 363 206 376 318
rect 465 206 478 318
rect 516 206 529 318
<< ndiff >>
rect 22 137 57 144
rect 22 121 30 137
rect 46 121 57 137
rect 22 93 57 121
rect 22 77 30 93
rect 46 77 57 93
rect 22 70 57 77
rect 70 137 108 144
rect 70 121 81 137
rect 97 121 108 137
rect 70 93 108 121
rect 70 77 81 93
rect 97 77 108 93
rect 70 70 108 77
rect 121 93 210 144
rect 121 77 132 93
rect 148 77 183 93
rect 199 77 210 93
rect 121 70 210 77
rect 223 137 261 144
rect 223 121 234 137
rect 250 121 261 137
rect 223 93 261 121
rect 223 77 234 93
rect 250 77 261 93
rect 223 70 261 77
rect 274 93 312 144
rect 274 77 285 93
rect 301 77 312 93
rect 274 70 312 77
rect 325 137 363 144
rect 325 121 336 137
rect 352 121 363 137
rect 325 93 363 121
rect 325 77 336 93
rect 352 77 363 93
rect 325 70 363 77
rect 376 93 465 144
rect 376 77 387 93
rect 403 77 438 93
rect 454 77 465 93
rect 376 70 465 77
rect 478 137 516 144
rect 478 121 489 137
rect 505 121 516 137
rect 478 93 516 121
rect 478 77 489 93
rect 505 77 516 93
rect 478 70 516 77
rect 529 137 563 144
rect 529 121 540 137
rect 556 121 563 137
rect 529 93 563 121
rect 529 77 540 93
rect 556 77 563 93
rect 529 70 563 77
<< pdiff >>
rect 22 311 57 318
rect 22 295 30 311
rect 46 295 57 311
rect 22 271 57 295
rect 22 255 30 271
rect 46 255 57 271
rect 22 229 57 255
rect 22 213 30 229
rect 46 213 57 229
rect 22 206 57 213
rect 70 311 108 318
rect 70 295 81 311
rect 97 295 108 311
rect 70 271 108 295
rect 70 255 81 271
rect 97 255 108 271
rect 70 229 108 255
rect 70 213 81 229
rect 97 213 108 229
rect 70 206 108 213
rect 121 311 155 318
rect 121 295 132 311
rect 148 295 155 311
rect 121 271 155 295
rect 121 255 132 271
rect 148 255 155 271
rect 121 206 155 255
rect 176 311 210 318
rect 176 295 183 311
rect 199 295 210 311
rect 176 271 210 295
rect 176 255 183 271
rect 199 255 210 271
rect 176 206 210 255
rect 223 271 261 318
rect 223 255 234 271
rect 250 255 261 271
rect 223 229 261 255
rect 223 213 234 229
rect 250 213 261 229
rect 223 206 261 213
rect 274 311 312 318
rect 274 295 285 311
rect 301 295 312 311
rect 274 271 312 295
rect 274 255 285 271
rect 301 255 312 271
rect 274 229 312 255
rect 274 213 285 229
rect 301 213 312 229
rect 274 206 312 213
rect 325 271 363 318
rect 325 255 336 271
rect 352 255 363 271
rect 325 229 363 255
rect 325 213 336 229
rect 352 213 363 229
rect 325 206 363 213
rect 376 311 410 318
rect 376 295 387 311
rect 403 295 410 311
rect 376 271 410 295
rect 376 255 387 271
rect 403 255 410 271
rect 376 206 410 255
rect 431 311 465 318
rect 431 295 438 311
rect 454 295 465 311
rect 431 271 465 295
rect 431 255 438 271
rect 454 255 465 271
rect 431 229 465 255
rect 431 213 438 229
rect 454 213 465 229
rect 431 206 465 213
rect 478 271 516 318
rect 478 255 489 271
rect 505 255 516 271
rect 478 229 516 255
rect 478 213 489 229
rect 505 213 516 229
rect 478 206 516 213
rect 529 311 563 318
rect 529 295 540 311
rect 556 295 563 311
rect 529 271 563 295
rect 529 255 540 271
rect 556 255 563 271
rect 529 229 563 255
rect 529 213 540 229
rect 556 213 563 229
rect 529 206 563 213
<< ndiffc >>
rect 30 121 46 137
rect 30 77 46 93
rect 81 121 97 137
rect 81 77 97 93
rect 132 77 148 93
rect 183 77 199 93
rect 234 121 250 137
rect 234 77 250 93
rect 285 77 301 93
rect 336 121 352 137
rect 336 77 352 93
rect 387 77 403 93
rect 438 77 454 93
rect 489 121 505 137
rect 489 77 505 93
rect 540 121 556 137
rect 540 77 556 93
<< pdiffc >>
rect 30 295 46 311
rect 30 255 46 271
rect 30 213 46 229
rect 81 295 97 311
rect 81 255 97 271
rect 81 213 97 229
rect 132 295 148 311
rect 132 255 148 271
rect 183 295 199 311
rect 183 255 199 271
rect 234 255 250 271
rect 234 213 250 229
rect 285 295 301 311
rect 285 255 301 271
rect 285 213 301 229
rect 336 255 352 271
rect 336 213 352 229
rect 387 295 403 311
rect 387 255 403 271
rect 438 295 454 311
rect 438 255 454 271
rect 438 213 454 229
rect 489 255 505 271
rect 489 213 505 229
rect 540 295 556 311
rect 540 255 556 271
rect 540 213 556 229
<< psubdiff >>
rect 0 8 576 15
rect 0 -8 16 8
rect 32 -8 64 8
rect 80 -8 112 8
rect 128 -8 160 8
rect 176 -8 208 8
rect 224 -8 256 8
rect 272 -8 304 8
rect 320 -8 352 8
rect 368 -8 400 8
rect 416 -8 448 8
rect 464 -8 496 8
rect 512 -8 544 8
rect 560 -8 576 8
rect 0 -15 576 -8
<< nsubdiff >>
rect 0 386 576 393
rect 0 370 16 386
rect 32 370 64 386
rect 80 370 112 386
rect 128 370 160 386
rect 176 370 208 386
rect 224 370 256 386
rect 272 370 304 386
rect 320 370 352 386
rect 368 370 400 386
rect 416 370 448 386
rect 464 370 496 386
rect 512 370 544 386
rect 560 370 576 386
rect 0 363 576 370
<< psubdiffcont >>
rect 16 -8 32 8
rect 64 -8 80 8
rect 112 -8 128 8
rect 160 -8 176 8
rect 208 -8 224 8
rect 256 -8 272 8
rect 304 -8 320 8
rect 352 -8 368 8
rect 400 -8 416 8
rect 448 -8 464 8
rect 496 -8 512 8
rect 544 -8 560 8
<< nsubdiffcont >>
rect 16 370 32 386
rect 64 370 80 386
rect 112 370 128 386
rect 160 370 176 386
rect 208 370 224 386
rect 256 370 272 386
rect 304 370 320 386
rect 352 370 368 386
rect 400 370 416 386
rect 448 370 464 386
rect 496 370 512 386
rect 544 370 560 386
<< poly >>
rect 57 318 70 336
rect 108 318 121 336
rect 210 318 223 336
rect 261 318 274 336
rect 312 318 325 336
rect 363 318 376 336
rect 465 318 478 336
rect 516 318 529 336
rect 57 190 70 206
rect 108 190 121 206
rect 210 190 223 206
rect 261 190 274 206
rect 312 190 325 206
rect 363 190 376 206
rect 465 190 478 206
rect 516 190 529 206
rect 48 183 129 190
rect 48 167 55 183
rect 71 167 106 183
rect 122 167 129 183
rect 48 160 129 167
rect 201 183 282 190
rect 201 167 208 183
rect 224 167 259 183
rect 275 167 282 183
rect 201 160 282 167
rect 303 183 384 190
rect 303 167 310 183
rect 326 167 361 183
rect 377 167 384 183
rect 303 160 384 167
rect 436 183 537 190
rect 436 167 443 183
rect 459 167 537 183
rect 436 160 537 167
rect 57 144 70 160
rect 108 144 121 160
rect 210 144 223 160
rect 261 144 274 160
rect 312 144 325 160
rect 363 144 376 160
rect 465 144 478 160
rect 516 144 529 160
rect 57 52 70 70
rect 108 52 121 70
rect 210 52 223 70
rect 261 52 274 70
rect 312 52 325 70
rect 363 52 376 70
rect 465 52 478 70
rect 516 52 529 70
<< polycont >>
rect 55 167 71 183
rect 106 167 122 183
rect 208 167 224 183
rect 259 167 275 183
rect 310 167 326 183
rect 361 167 377 183
rect 443 167 459 183
<< metal1 >>
rect 0 386 576 400
rect 0 370 16 386
rect 32 370 64 386
rect 80 370 112 386
rect 128 370 160 386
rect 176 370 208 386
rect 224 370 256 386
rect 272 370 304 386
rect 320 370 352 386
rect 368 370 400 386
rect 416 370 448 386
rect 464 370 496 386
rect 512 370 544 386
rect 560 370 576 386
rect 0 356 576 370
rect 25 311 51 356
rect 25 295 30 311
rect 46 295 51 311
rect 25 271 51 295
rect 25 255 30 271
rect 46 255 51 271
rect 25 229 51 255
rect 25 213 30 229
rect 46 213 51 229
rect 25 208 51 213
rect 76 311 102 316
rect 76 295 81 311
rect 97 295 102 311
rect 76 271 102 295
rect 76 255 81 271
rect 97 255 102 271
rect 76 234 102 255
rect 127 311 153 356
rect 127 295 132 311
rect 148 295 153 311
rect 127 271 153 295
rect 127 255 132 271
rect 148 255 153 271
rect 127 252 153 255
rect 178 311 408 320
rect 178 295 183 311
rect 199 295 285 311
rect 301 295 387 311
rect 403 295 408 311
rect 178 294 408 295
rect 178 271 204 294
rect 178 255 183 271
rect 199 255 204 271
rect 178 252 204 255
rect 229 271 255 276
rect 229 255 234 271
rect 250 255 255 271
rect 229 234 255 255
rect 76 229 255 234
rect 76 213 81 229
rect 97 213 234 229
rect 250 213 255 229
rect 76 212 255 213
rect 280 271 306 294
rect 280 255 285 271
rect 301 255 306 271
rect 280 229 306 255
rect 280 213 285 229
rect 301 213 306 229
rect 280 208 306 213
rect 331 271 357 276
rect 331 255 336 271
rect 352 255 357 271
rect 331 230 357 255
rect 382 271 408 294
rect 382 255 387 271
rect 403 255 408 271
rect 382 250 408 255
rect 433 311 561 320
rect 433 295 438 311
rect 454 295 540 311
rect 556 295 561 311
rect 433 294 561 295
rect 433 271 459 294
rect 433 255 438 271
rect 454 255 459 271
rect 433 230 459 255
rect 331 229 459 230
rect 331 213 336 229
rect 352 213 438 229
rect 454 213 459 229
rect 331 212 459 213
rect 484 271 510 276
rect 484 255 489 271
rect 505 255 510 271
rect 484 229 510 255
rect 484 213 489 229
rect 505 213 510 229
rect 48 183 129 190
rect 48 167 55 183
rect 71 167 106 183
rect 122 167 129 183
rect 48 157 129 167
rect 201 183 282 190
rect 201 167 208 183
rect 224 167 259 183
rect 275 167 282 183
rect 201 157 282 167
rect 303 183 384 190
rect 303 167 310 183
rect 326 167 361 183
rect 377 167 384 183
rect 303 157 384 167
rect 402 183 466 190
rect 402 167 443 183
rect 459 167 466 183
rect 402 157 466 167
rect 484 137 510 213
rect 535 271 561 294
rect 535 255 540 271
rect 556 255 561 271
rect 535 229 561 255
rect 535 213 540 229
rect 556 213 561 229
rect 535 208 561 213
rect 25 121 30 137
rect 46 121 51 137
rect 25 93 51 121
rect 25 77 30 93
rect 46 77 51 93
rect 25 22 51 77
rect 76 121 81 137
rect 97 121 234 137
rect 250 121 336 137
rect 352 121 489 137
rect 505 121 510 137
rect 76 117 510 121
rect 76 93 102 117
rect 76 77 81 93
rect 97 77 102 93
rect 76 72 102 77
rect 127 93 204 98
rect 127 77 132 93
rect 148 77 183 93
rect 199 77 204 93
rect 127 22 204 77
rect 229 93 255 117
rect 229 77 234 93
rect 250 77 255 93
rect 229 72 255 77
rect 280 93 306 98
rect 280 77 285 93
rect 301 77 306 93
rect 280 22 306 77
rect 331 93 357 117
rect 331 77 336 93
rect 352 77 357 93
rect 331 72 357 77
rect 382 93 459 98
rect 382 77 387 93
rect 403 77 438 93
rect 454 77 459 93
rect 382 22 459 77
rect 484 93 510 117
rect 484 77 489 93
rect 505 77 510 93
rect 484 72 510 77
rect 535 137 561 142
rect 535 121 540 137
rect 556 121 561 137
rect 535 93 561 121
rect 535 77 540 93
rect 556 77 561 93
rect 535 22 561 77
rect 0 8 576 22
rect 0 -8 16 8
rect 32 -8 64 8
rect 80 -8 112 8
rect 128 -8 160 8
rect 176 -8 208 8
rect 224 -8 256 8
rect 272 -8 304 8
rect 320 -8 352 8
rect 368 -8 400 8
rect 416 -8 448 8
rect 464 -8 496 8
rect 512 -8 544 8
rect 560 -8 576 8
rect 0 -22 576 -8
<< labels >>
flabel metal1 s 484 72 510 276 0 FreeSans 250 0 0 0 Y
port 4 nsew
flabel metal1 s 402 158 466 190 0 FreeSans 250 0 0 0 D
port 1 nsew
flabel metal1 s 0 356 576 400 0 FreeSans 250 0 0 0 VDD
port 5 nsew
flabel metal1 s 201 158 282 190 0 FreeSans 250 0 0 0 B
port 2 nsew
flabel metal1 s 48 158 129 190 0 FreeSans 250 0 0 0 A
port 7 nsew
flabel metal1 s 0 -22 576 22 0 FreeSans 250 0 0 0 VSS
port 6 nsew
flabel metal1 s 303 158 384 190 0 FreeSans 250 0 0 0 C
port 3 nsew
<< properties >>
string FIXED_BBOX 0 0 576 378
string GDS_END 244964
string GDS_FILE ../gds/controller.gds
string GDS_START 236706
<< end >>
