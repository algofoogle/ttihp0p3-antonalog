magic
tech ihp-sg13g2
timestamp 1747537721
<< nwell >>
rect -24 175 360 417
<< pwell >>
rect 34 28 320 148
rect -13 -28 349 28
<< nmos >>
rect 81 80 94 135
rect 145 61 158 135
rect 205 61 218 135
rect 248 61 261 135
<< pmos >>
rect 92 206 105 290
rect 146 206 159 318
rect 197 206 210 318
rect 248 206 261 318
<< ndiff >>
rect 47 115 81 135
rect 47 99 54 115
rect 70 99 81 115
rect 47 80 81 99
rect 94 91 145 135
rect 94 80 113 91
rect 101 75 113 80
rect 129 75 145 91
rect 101 61 145 75
rect 158 61 205 135
rect 218 61 248 135
rect 261 126 307 135
rect 261 110 282 126
rect 298 110 307 126
rect 261 85 307 110
rect 261 69 272 85
rect 288 69 307 85
rect 261 61 307 69
<< pdiff >>
rect 112 310 146 318
rect 112 294 119 310
rect 135 294 146 310
rect 112 290 146 294
rect 58 283 92 290
rect 58 267 65 283
rect 81 267 92 283
rect 58 241 92 267
rect 58 225 65 241
rect 81 225 92 241
rect 58 206 92 225
rect 105 275 146 290
rect 105 259 119 275
rect 135 259 146 275
rect 105 233 146 259
rect 105 217 119 233
rect 135 217 146 233
rect 105 206 146 217
rect 159 310 197 318
rect 159 294 170 310
rect 186 294 197 310
rect 159 276 197 294
rect 159 260 170 276
rect 186 260 197 276
rect 159 241 197 260
rect 159 225 170 241
rect 186 225 197 241
rect 159 206 197 225
rect 210 310 248 318
rect 210 294 221 310
rect 237 294 248 310
rect 210 275 248 294
rect 210 259 221 275
rect 237 259 248 275
rect 210 206 248 259
rect 261 310 295 318
rect 261 294 272 310
rect 288 294 295 310
rect 261 270 295 294
rect 261 254 272 270
rect 288 254 295 270
rect 261 230 295 254
rect 261 214 272 230
rect 288 214 295 230
rect 261 206 295 214
<< ndiffc >>
rect 54 99 70 115
rect 113 75 129 91
rect 282 110 298 126
rect 272 69 288 85
<< pdiffc >>
rect 119 294 135 310
rect 65 267 81 283
rect 65 225 81 241
rect 119 259 135 275
rect 119 217 135 233
rect 170 294 186 310
rect 170 260 186 276
rect 170 225 186 241
rect 221 294 237 310
rect 221 259 237 275
rect 272 294 288 310
rect 272 254 288 270
rect 272 214 288 230
<< psubdiff >>
rect 0 8 336 15
rect 0 -8 16 8
rect 32 -8 64 8
rect 80 -8 112 8
rect 128 -8 160 8
rect 176 -8 208 8
rect 224 -8 256 8
rect 272 -8 304 8
rect 320 -8 336 8
rect 0 -15 336 -8
<< nsubdiff >>
rect 0 386 336 393
rect 0 370 16 386
rect 32 370 64 386
rect 80 370 112 386
rect 128 370 160 386
rect 176 370 208 386
rect 224 370 256 386
rect 272 370 304 386
rect 320 370 336 386
rect 0 363 336 370
<< psubdiffcont >>
rect 16 -8 32 8
rect 64 -8 80 8
rect 112 -8 128 8
rect 160 -8 176 8
rect 208 -8 224 8
rect 256 -8 272 8
rect 304 -8 320 8
<< nsubdiffcont >>
rect 16 370 32 386
rect 64 370 80 386
rect 112 370 128 386
rect 160 370 176 386
rect 208 370 224 386
rect 256 370 272 386
rect 304 370 320 386
<< poly >>
rect 146 318 159 336
rect 197 318 210 336
rect 248 318 261 336
rect 92 290 105 308
rect 92 187 105 206
rect 146 187 159 206
rect 197 190 210 206
rect 75 180 105 187
rect 75 164 82 180
rect 98 164 105 180
rect 75 157 105 164
rect 135 180 165 187
rect 135 164 142 180
rect 158 164 165 180
rect 135 157 165 164
rect 196 181 226 190
rect 248 185 261 206
rect 196 165 203 181
rect 219 165 226 181
rect 196 158 226 165
rect 247 178 277 185
rect 247 162 254 178
rect 270 162 277 178
rect 81 135 94 157
rect 145 135 158 157
rect 205 135 218 158
rect 247 155 277 162
rect 248 135 261 155
rect 81 62 94 80
rect 145 43 158 61
rect 205 43 218 61
rect 248 43 261 61
<< polycont >>
rect 82 164 98 180
rect 142 164 158 180
rect 203 165 219 181
rect 254 162 270 178
<< metal1 >>
rect 0 386 336 400
rect 0 370 16 386
rect 32 370 64 386
rect 80 370 112 386
rect 128 370 160 386
rect 176 370 208 386
rect 224 370 256 386
rect 272 370 304 386
rect 320 370 336 386
rect 0 356 336 370
rect 114 310 140 356
rect 114 294 119 310
rect 135 294 140 310
rect 44 283 86 286
rect 44 267 65 283
rect 81 267 86 283
rect 44 241 86 267
rect 44 225 65 241
rect 81 225 86 241
rect 44 223 86 225
rect 114 275 140 294
rect 114 259 119 275
rect 135 259 140 275
rect 114 233 140 259
rect 44 137 61 223
rect 114 217 119 233
rect 135 217 140 233
rect 165 310 191 313
rect 165 294 170 310
rect 186 294 191 310
rect 165 276 191 294
rect 165 260 170 276
rect 186 260 191 276
rect 165 241 191 260
rect 216 310 242 356
rect 216 294 221 310
rect 237 294 242 310
rect 216 275 242 294
rect 216 259 221 275
rect 237 259 242 275
rect 216 257 242 259
rect 264 310 313 320
rect 264 294 272 310
rect 288 294 313 310
rect 264 270 313 294
rect 165 225 170 241
rect 186 239 191 241
rect 264 254 272 270
rect 288 254 313 270
rect 264 239 313 254
rect 186 230 313 239
rect 186 225 272 230
rect 165 220 272 225
rect 264 214 272 220
rect 288 214 313 230
rect 264 210 313 214
rect 79 180 117 198
rect 79 164 82 180
rect 98 164 117 180
rect 79 157 117 164
rect 135 180 168 198
rect 135 164 142 180
rect 158 164 168 180
rect 135 157 168 164
rect 190 181 225 200
rect 190 165 203 181
rect 219 165 225 181
rect 190 157 225 165
rect 243 178 278 187
rect 243 162 254 178
rect 270 162 278 178
rect 243 154 278 162
rect 243 137 259 154
rect 44 120 259 137
rect 296 136 313 210
rect 277 126 313 136
rect 44 115 71 120
rect 44 99 54 115
rect 70 99 71 115
rect 277 110 282 126
rect 298 110 313 126
rect 277 101 313 110
rect 44 88 71 99
rect 108 91 135 96
rect 108 75 113 91
rect 129 75 135 91
rect 108 22 135 75
rect 263 85 313 101
rect 263 69 272 85
rect 288 69 313 85
rect 263 62 313 69
rect 0 8 336 22
rect 0 -8 16 8
rect 32 -8 64 8
rect 80 -8 112 8
rect 128 -8 160 8
rect 176 -8 208 8
rect 224 -8 256 8
rect 272 -8 304 8
rect 320 -8 336 8
rect 0 -22 336 -8
<< labels >>
flabel metal1 s 79 157 117 198 0 FreeSans 200 0 0 0 A_N
port 2 nsew
flabel metal1 s 264 210 313 320 0 FreeSans 200 0 0 0 Y
port 3 nsew
flabel metal1 s 0 356 336 400 0 FreeSans 200 0 0 0 VDD
port 4 nsew
flabel metal1 s 0 -22 336 22 0 FreeSans 200 0 0 0 VSS
port 5 nsew
flabel metal1 s 190 157 225 200 0 FreeSans 200 0 0 0 B
port 6 nsew
flabel metal1 s 135 157 168 198 0 FreeSans 200 0 0 0 C
port 7 nsew
<< properties >>
string FIXED_BBOX 0 0 336 378
string GDS_END 159590
string GDS_FILE ../gds/controller.gds
string GDS_START 153760
<< end >>
