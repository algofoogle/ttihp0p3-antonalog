magic
tech ihp-sg13g2
timestamp 1747485648
<< pwell >>
rect -1401 -512 1941 528
<< psubdiff >>
rect -1370 490 1910 497
rect -1370 474 -1324 490
rect 1864 474 1910 490
rect -1370 467 1910 474
rect -1370 451 -1340 467
rect -1370 -435 -1363 451
rect -1347 -435 -1340 451
rect -1370 -451 -1340 -435
rect 1880 451 1910 467
rect 1880 -435 1887 451
rect 1903 -435 1910 451
rect 1880 -451 1910 -435
rect -1370 -458 1910 -451
rect -1370 -474 -1324 -458
rect 1864 -474 1910 -458
rect -1370 -481 1910 -474
<< psubdiffcont >>
rect -1324 474 1864 490
rect -1363 -435 -1347 451
rect 1887 -435 1903 451
rect -1324 -474 1864 -458
<< metal1 >>
rect -1363 474 -1324 490
rect 1864 474 1903 490
rect -1363 451 -1347 474
rect -1363 -458 -1347 -435
rect 1887 451 1903 474
rect 1887 -458 1903 -435
rect -1363 -474 -1324 -458
rect 1864 -474 1903 -458
<< end >>
