magic
tech ihp-sg13g2
magscale 1 2
timestamp 1746816455
<< metal1 >>
rect 2687 27560 3127 27569
rect 2687 27120 2688 27560
rect 3126 27120 3824 27560
rect 2687 27111 3127 27120
rect 3705 26378 3785 26387
rect 3705 26298 3706 26378
rect 3784 26298 3785 26378
rect 3705 26289 3785 26298
rect 5265 25482 5345 25491
rect 5265 25402 5266 25482
rect 5344 25402 5345 25482
rect 5265 25393 5345 25402
rect 3703 24596 3783 24605
rect 3703 24516 3704 24596
rect 3782 24516 3783 24596
rect 3703 24507 3783 24516
rect 5265 23708 5345 23717
rect 5265 23628 5266 23708
rect 5344 23628 5345 23708
rect 5265 23619 5345 23628
rect 3695 22820 3775 22829
rect 3695 22740 3696 22820
rect 3774 22740 3775 22820
rect 3695 22731 3775 22740
rect 5249 21940 5329 21949
rect 5249 21860 5250 21940
rect 5328 21860 5329 21940
rect 5249 21851 5329 21860
rect 3695 21020 3775 21029
rect 3695 20940 3696 21020
rect 3774 20940 3775 21020
rect 3695 20931 3775 20940
rect 5227 20646 5407 20655
rect 5227 20466 5228 20646
rect 5406 20466 5407 20646
rect 5227 20457 5407 20466
rect 2657 20324 3097 20333
rect 2657 19884 2658 20324
rect 3096 19924 3662 20324
rect 5249 20150 5329 20159
rect 5249 20070 5250 20150
rect 5328 20070 5329 20150
rect 5249 20061 5329 20070
rect 3096 19884 5642 19924
rect 2657 19875 3097 19884
rect 3222 19680 5642 19884
rect 3218 19628 5642 19680
rect 3218 19174 5712 19628
rect 3218 18784 3936 19174
rect 3719 18054 3799 18063
rect 3719 17974 3720 18054
rect 3798 17974 3799 18054
rect 3719 17965 3799 17974
rect 5275 17158 5355 17167
rect 5275 17078 5276 17158
rect 5354 17078 5355 17158
rect 5275 17069 5355 17078
rect 3713 16276 3793 16285
rect 3713 16196 3714 16276
rect 3792 16196 3793 16276
rect 3713 16187 3793 16196
rect 5285 15388 5383 15389
rect 5285 15310 5294 15388
rect 5374 15310 5383 15388
rect 5285 15309 5383 15310
rect 3719 14484 3799 14493
rect 3719 14404 3720 14484
rect 3798 14404 3799 14484
rect 3719 14395 3799 14404
rect 5265 13612 5345 13621
rect 5265 13532 5266 13612
rect 5344 13532 5345 13612
rect 5265 13523 5345 13532
rect 3709 12720 3789 12729
rect 3709 12640 3710 12720
rect 3788 12640 3789 12720
rect 3709 12631 3789 12640
rect 5219 12338 5399 12347
rect 5219 12158 5220 12338
rect 5398 12158 5399 12338
rect 5219 12149 5399 12158
rect 5269 11834 5349 11843
rect 2621 11752 3061 11761
rect 5269 11754 5270 11834
rect 5348 11754 5349 11834
rect 2621 11312 2622 11752
rect 3060 11746 3152 11752
rect 3060 11584 3680 11746
rect 5269 11745 5349 11754
rect 3060 11320 5664 11584
rect 3060 11318 5696 11320
rect 3060 11312 3152 11318
rect 2621 11303 3061 11312
rect 3428 11006 5696 11318
rect 3462 10842 5696 11006
rect 3462 10452 3900 10842
rect 3723 9720 3803 9729
rect 3723 9640 3724 9720
rect 3802 9640 3803 9720
rect 3723 9631 3803 9640
rect 5281 8842 5361 8851
rect 5281 8762 5282 8842
rect 5360 8762 5361 8842
rect 5281 8753 5361 8762
rect 3729 7948 3809 7957
rect 3729 7868 3730 7948
rect 3808 7868 3809 7948
rect 3729 7859 3809 7868
rect 5285 7054 5365 7063
rect 5285 6974 5286 7054
rect 5364 6974 5365 7054
rect 5285 6965 5365 6974
rect 3729 6176 3809 6185
rect 3729 6096 3730 6176
rect 3808 6096 3809 6176
rect 3729 6087 3809 6096
rect 5271 5286 5351 5295
rect 5271 5206 5272 5286
rect 5350 5206 5351 5286
rect 5271 5197 5351 5206
rect 3713 4398 3793 4407
rect 3713 4318 3714 4398
rect 3792 4318 3793 4398
rect 3713 4309 3793 4318
rect 5223 4010 5403 4019
rect 5223 3830 5224 4010
rect 5402 3830 5403 4010
rect 5223 3821 5403 3830
rect 5271 3504 5351 3513
rect 5271 3424 5272 3504
rect 5350 3424 5351 3504
rect 5271 3415 5351 3424
rect 2581 3334 3021 3343
rect 2581 2894 2582 3334
rect 3020 3328 3112 3334
rect 3020 3312 3226 3328
rect 3020 3299 3370 3312
rect 3020 2949 5639 3299
rect 3020 2906 3370 2949
rect 3020 2900 3226 2906
rect 3020 2894 3112 2900
rect 2581 2885 3021 2894
<< via1 >>
rect 2688 27120 3126 27560
rect 3706 26298 3784 26378
rect 5266 25402 5344 25482
rect 3704 24516 3782 24596
rect 5266 23628 5344 23708
rect 3696 22740 3774 22820
rect 5250 21860 5328 21940
rect 3696 20940 3774 21020
rect 5228 20466 5406 20646
rect 2658 19884 3096 20324
rect 5250 20070 5328 20150
rect 3720 17974 3798 18054
rect 5276 17078 5354 17158
rect 3714 16196 3792 16276
rect 5294 15310 5374 15388
rect 3720 14404 3798 14484
rect 5266 13532 5344 13612
rect 3710 12640 3788 12720
rect 5220 12158 5398 12338
rect 5270 11754 5348 11834
rect 2622 11312 3060 11752
rect 3724 9640 3802 9720
rect 5282 8762 5360 8842
rect 3730 7868 3808 7948
rect 5286 6974 5364 7054
rect 3730 6096 3808 6176
rect 5272 5206 5350 5286
rect 3714 4318 3792 4398
rect 5224 3830 5402 4010
rect 5272 3424 5350 3504
rect 2582 2894 3020 3334
<< metal2 >>
rect 2686 27560 3126 27569
rect 2679 27120 2686 27560
rect 3126 27120 3135 27560
rect 2686 27111 3126 27120
rect 3697 26298 3706 26378
rect 3784 26298 7298 26378
rect 5257 25402 5266 25482
rect 5344 25402 7106 25482
rect 3695 24516 3704 24596
rect 3782 24516 6900 24596
rect 5257 23628 5266 23708
rect 5344 23628 6650 23708
rect 3687 22740 3696 22820
rect 3774 22740 6422 22820
rect 5241 21860 5250 21940
rect 5328 21860 6188 21940
rect 3007 21600 3016 21780
rect 3196 21600 3205 21780
rect 3016 20646 3196 21600
rect 6108 21440 6188 21860
rect 6342 21860 6422 22740
rect 6570 22280 6650 23628
rect 6820 22700 6900 24516
rect 7026 23120 7106 25402
rect 7218 23540 7298 26298
rect 7218 23460 7726 23540
rect 7026 23040 7682 23120
rect 6820 22620 7698 22700
rect 6570 22200 7690 22280
rect 6342 21780 7674 21860
rect 6108 21360 7682 21440
rect 3687 20940 3696 21020
rect 3774 20940 7690 21020
rect 3016 20466 5228 20646
rect 5406 20466 5415 20646
rect 7116 20520 7690 20600
rect 2656 20324 3096 20333
rect 2649 19884 2656 20324
rect 3096 19884 3105 20324
rect 7116 20150 7196 20520
rect 5241 20070 5250 20150
rect 5328 20070 7196 20150
rect 2656 19875 3096 19884
rect 3711 17974 3720 18054
rect 3798 17974 7262 18054
rect 5267 17078 5276 17158
rect 5354 17078 7020 17158
rect 6940 16400 7020 17078
rect 7182 16820 7262 17974
rect 7182 16740 7686 16820
rect 6940 16320 7586 16400
rect 3705 16196 3714 16276
rect 3792 16196 6784 16276
rect 6704 15980 6784 16196
rect 6704 15900 7592 15980
rect 5294 15480 7680 15560
rect 5294 15388 5374 15480
rect 5294 15301 5374 15310
rect 5860 15060 7672 15140
rect 5860 14484 5940 15060
rect 3711 14404 3720 14484
rect 3798 14404 5940 14484
rect 6276 14640 7596 14720
rect 6276 13612 6356 14640
rect 5257 13532 5266 13612
rect 5344 13532 6356 13612
rect 6676 14220 7596 14300
rect 6676 12720 6756 14220
rect 3701 12640 3710 12720
rect 3788 12640 6756 12720
rect 7064 13800 7600 13880
rect 2707 12158 2716 12338
rect 2896 12158 5220 12338
rect 5398 12158 5407 12338
rect 7064 11834 7144 13800
rect 2620 11752 3060 11761
rect 5261 11754 5270 11834
rect 5348 11754 7144 11834
rect 2613 11312 2620 11752
rect 3060 11312 3069 11752
rect 2620 11303 3060 11312
rect 5326 10020 7680 10100
rect 5326 9720 5406 10020
rect 3715 9640 3724 9720
rect 3802 9640 5406 9720
rect 5598 9600 7590 9680
rect 5598 8842 5678 9600
rect 5273 8762 5282 8842
rect 5360 8762 5678 8842
rect 5814 9180 7586 9260
rect 5814 7948 5894 9180
rect 3721 7868 3730 7948
rect 3808 7868 5894 7948
rect 6030 8760 7580 8840
rect 6030 7054 6110 8760
rect 5277 6974 5286 7054
rect 5364 6974 6110 7054
rect 6240 8340 7596 8420
rect 6240 6176 6320 8340
rect 3721 6096 3730 6176
rect 3808 6096 6320 6176
rect 6440 7920 7586 8000
rect 6440 5286 6520 7920
rect 5263 5206 5272 5286
rect 5350 5206 6520 5286
rect 6646 7500 7590 7580
rect 6646 4398 6726 7500
rect 3705 4318 3714 4398
rect 3792 4318 6726 4398
rect 6888 7080 7616 7160
rect 1634 4010 1814 4019
rect 1814 3830 5224 4010
rect 5402 3830 5411 4010
rect 1634 3821 1814 3830
rect 6888 3504 6968 7080
rect 5263 3424 5272 3504
rect 5350 3424 6968 3504
rect 2580 3334 3020 3343
rect 2573 2894 2580 3334
rect 3020 2894 3029 3334
rect 2580 2885 3020 2894
<< via2 >>
rect 2686 27120 2688 27560
rect 2688 27120 3126 27560
rect 3016 21600 3196 21780
rect 2656 19884 2658 20324
rect 2658 19884 3096 20324
rect 2716 12158 2896 12338
rect 2620 11312 2622 11752
rect 2622 11312 3060 11752
rect 1634 3830 1814 4010
rect 2580 2894 2582 3334
rect 2582 2894 3020 3334
<< metal3 >>
rect 10502 30465 10621 30479
rect 10502 30373 10515 30465
rect 10607 30373 10621 30465
rect 10502 30019 10621 30373
rect 11270 30465 11389 30479
rect 11270 30373 11283 30465
rect 11375 30373 11389 30465
rect 11270 30019 11389 30373
rect 12038 30465 12157 30479
rect 12038 30373 12051 30465
rect 12143 30373 12157 30465
rect 12038 30019 12157 30373
rect 12806 30465 12925 30479
rect 12806 30373 12819 30465
rect 12911 30373 12925 30465
rect 12806 30019 12925 30373
rect 13574 30465 13693 30479
rect 13574 30373 13587 30465
rect 13679 30373 13693 30465
rect 13574 30019 13693 30373
rect 14342 30465 14461 30479
rect 14342 30373 14355 30465
rect 14447 30373 14461 30465
rect 14342 30019 14461 30373
rect 15110 30465 15229 30479
rect 15110 30373 15123 30465
rect 15215 30373 15229 30465
rect 15110 30019 15229 30373
rect 15878 30465 15997 30479
rect 15878 30373 15891 30465
rect 15983 30373 15997 30465
rect 15878 30019 15997 30373
rect 16646 30465 16765 30479
rect 16646 30373 16659 30465
rect 16751 30373 16765 30465
rect 16646 30019 16765 30373
rect 17414 30465 17533 30479
rect 17414 30373 17427 30465
rect 17519 30373 17533 30465
rect 17414 30019 17533 30373
rect 18182 30465 18301 30479
rect 18182 30373 18195 30465
rect 18287 30373 18301 30465
rect 18182 30019 18301 30373
rect 18950 30465 19069 30479
rect 18950 30373 18963 30465
rect 19055 30373 19069 30465
rect 18950 30019 19069 30373
rect 19718 30465 19837 30479
rect 19718 30373 19731 30465
rect 19823 30373 19837 30465
rect 19718 30019 19837 30373
rect 20486 30465 20605 30479
rect 20486 30373 20499 30465
rect 20591 30373 20605 30465
rect 20486 30019 20605 30373
rect 21254 30465 21373 30479
rect 21254 30373 21267 30465
rect 21359 30373 21373 30465
rect 21254 30019 21373 30373
rect 22022 30465 22141 30479
rect 22022 30373 22035 30465
rect 22127 30373 22141 30465
rect 22022 30019 22141 30373
rect 22790 30465 22909 30479
rect 22790 30373 22803 30465
rect 22895 30373 22909 30465
rect 22790 30019 22909 30373
rect 23558 30465 23677 30479
rect 23558 30373 23571 30465
rect 23663 30373 23677 30465
rect 23558 30019 23677 30373
rect 30471 30362 30480 30458
rect 30576 30362 30585 30458
rect 31239 30362 31248 30458
rect 31344 30362 31353 30458
rect 32007 30362 32016 30458
rect 32112 30362 32121 30458
rect 32775 30362 32784 30458
rect 32880 30362 32889 30458
rect 33543 30362 33552 30458
rect 33648 30362 33657 30458
rect 34311 30362 34320 30458
rect 34416 30362 34425 30458
rect 35079 30362 35088 30458
rect 35184 30362 35193 30458
rect 35847 30362 35856 30458
rect 35952 30362 35961 30458
rect 36615 30362 36624 30458
rect 36720 30362 36729 30458
rect 37383 30362 37392 30458
rect 37488 30362 37497 30458
rect 38151 30362 38160 30458
rect 38256 30362 38265 30458
rect 30480 30010 30576 30362
rect 31248 30010 31344 30362
rect 32016 30010 32112 30362
rect 32784 30010 32880 30362
rect 33552 30010 33648 30362
rect 34320 30010 34416 30362
rect 35088 30010 35184 30362
rect 35856 30010 35952 30362
rect 36624 30010 36720 30362
rect 37392 30010 37488 30362
rect 38160 30010 38256 30362
rect 2677 27120 2686 27560
rect 3126 27120 3135 27560
rect 3007 24596 3016 24776
rect 3196 24596 3205 24776
rect 3016 21780 3196 24596
rect 3016 21591 3196 21600
rect 2181 21396 2190 21576
rect 2370 21396 2379 21576
rect 2190 19098 2370 21396
rect 2647 19884 2656 20324
rect 3096 19884 3105 20324
rect 2190 18918 2896 19098
rect 1625 18196 1634 18376
rect 1814 18196 1823 18376
rect 1634 4010 1814 18196
rect 2716 12338 2896 18918
rect 2716 12149 2896 12158
rect 2611 11312 2620 11752
rect 3060 11312 3069 11752
rect 1625 3830 1634 4010
rect 1814 3830 1823 4010
rect 2571 2894 2580 3334
rect 3020 2894 3029 3334
<< via3 >>
rect 10515 30373 10607 30465
rect 11283 30373 11375 30465
rect 12051 30373 12143 30465
rect 12819 30373 12911 30465
rect 13587 30373 13679 30465
rect 14355 30373 14447 30465
rect 15123 30373 15215 30465
rect 15891 30373 15983 30465
rect 16659 30373 16751 30465
rect 17427 30373 17519 30465
rect 18195 30373 18287 30465
rect 18963 30373 19055 30465
rect 19731 30373 19823 30465
rect 20499 30373 20591 30465
rect 21267 30373 21359 30465
rect 22035 30373 22127 30465
rect 22803 30373 22895 30465
rect 23571 30373 23663 30465
rect 30480 30362 30576 30458
rect 31248 30362 31344 30458
rect 32016 30362 32112 30458
rect 32784 30362 32880 30458
rect 33552 30362 33648 30458
rect 34320 30362 34416 30458
rect 35088 30362 35184 30458
rect 35856 30362 35952 30458
rect 36624 30362 36720 30458
rect 37392 30362 37488 30458
rect 38160 30362 38256 30458
rect 2686 27120 3126 27560
rect 3016 24596 3196 24776
rect 2190 21396 2370 21576
rect 2656 19884 3096 20324
rect 1634 18196 1814 18376
rect 2620 11312 3060 11752
rect 2580 2894 3020 3334
<< metal4 >>
rect 10515 30465 10607 30474
rect 11283 30465 11375 30474
rect 12051 30465 12143 30474
rect 12819 30465 12911 30474
rect 13587 30465 13679 30474
rect 14355 30465 14447 30474
rect 15123 30465 15215 30474
rect 15891 30465 15983 30474
rect 16659 30465 16751 30474
rect 17427 30465 17519 30474
rect 18195 30465 18287 30474
rect 18963 30465 19055 30474
rect 19731 30465 19823 30474
rect 20499 30465 20591 30474
rect 21267 30465 21359 30474
rect 22035 30465 22127 30474
rect 22803 30465 22895 30474
rect 23571 30465 23663 30474
rect 10508 30375 10515 30462
rect 10607 30375 10613 30462
rect 11276 30375 11283 30462
rect 11375 30375 11381 30462
rect 12044 30375 12051 30462
rect 12143 30375 12149 30462
rect 12812 30375 12819 30462
rect 12911 30375 12917 30462
rect 13580 30375 13587 30462
rect 13679 30375 13685 30462
rect 14348 30375 14355 30462
rect 14447 30375 14453 30462
rect 15116 30375 15123 30462
rect 15215 30375 15221 30462
rect 15884 30375 15891 30462
rect 15983 30375 15989 30462
rect 16652 30375 16659 30462
rect 16751 30375 16757 30462
rect 17420 30375 17427 30462
rect 17519 30375 17525 30462
rect 18188 30375 18195 30462
rect 18287 30375 18293 30462
rect 18956 30375 18963 30462
rect 19055 30375 19061 30462
rect 19724 30375 19731 30462
rect 19823 30375 19829 30462
rect 20492 30375 20499 30462
rect 20591 30375 20597 30462
rect 21260 30375 21267 30462
rect 21359 30375 21365 30462
rect 22028 30375 22035 30462
rect 22127 30375 22133 30462
rect 22796 30375 22803 30462
rect 22895 30375 22901 30462
rect 23564 30375 23571 30462
rect 23663 30375 23669 30462
rect 30480 30458 30576 30467
rect 31248 30458 31344 30467
rect 32016 30458 32112 30467
rect 32784 30458 32880 30467
rect 33552 30458 33648 30467
rect 34320 30458 34416 30467
rect 35088 30458 35184 30467
rect 35856 30458 35952 30467
rect 36624 30458 36720 30467
rect 37392 30458 37488 30467
rect 38160 30458 38256 30467
rect 10515 30364 10607 30373
rect 11283 30364 11375 30373
rect 12051 30364 12143 30373
rect 12819 30364 12911 30373
rect 13587 30364 13679 30373
rect 14355 30364 14447 30373
rect 15123 30364 15215 30373
rect 15891 30364 15983 30373
rect 16659 30364 16751 30373
rect 17427 30364 17519 30373
rect 18195 30364 18287 30373
rect 18963 30364 19055 30373
rect 19731 30364 19823 30373
rect 20499 30364 20591 30373
rect 21267 30364 21359 30373
rect 22035 30364 22127 30373
rect 22803 30364 22895 30373
rect 23571 30364 23663 30373
rect 30471 30362 30480 30458
rect 30576 30362 30585 30458
rect 31239 30362 31248 30458
rect 31344 30362 31353 30458
rect 32007 30362 32016 30458
rect 32112 30362 32121 30458
rect 32775 30362 32784 30458
rect 32880 30362 32889 30458
rect 33543 30362 33552 30458
rect 33648 30362 33657 30458
rect 34311 30362 34320 30458
rect 34416 30362 34425 30458
rect 35079 30362 35088 30458
rect 35184 30362 35193 30458
rect 35847 30362 35856 30458
rect 35952 30362 35961 30458
rect 36615 30362 36624 30458
rect 36720 30362 36729 30458
rect 37383 30362 37392 30458
rect 37488 30362 37497 30458
rect 38151 30362 38160 30458
rect 38256 30362 38265 30458
rect 30480 30353 30576 30362
rect 31248 30353 31344 30362
rect 32016 30353 32112 30362
rect 32784 30353 32880 30362
rect 33552 30353 33648 30362
rect 34320 30353 34416 30362
rect 35088 30353 35184 30362
rect 35856 30353 35952 30362
rect 36624 30353 36720 30362
rect 37392 30353 37488 30362
rect 38160 30353 38256 30362
rect 2686 27560 3126 27569
rect 2686 27111 3126 27120
rect 416 24776 596 24785
rect 3016 24776 3196 24785
rect 596 24596 3016 24776
rect 416 24587 596 24596
rect 3016 24587 3196 24596
rect 418 21576 598 21585
rect 2190 21576 2370 21585
rect 598 21396 2190 21576
rect 418 21387 598 21396
rect 2190 21387 2370 21396
rect 2656 20324 3096 20333
rect 2656 19875 3096 19884
rect 392 18376 572 18385
rect 1634 18376 1814 18385
rect 572 18196 1634 18376
rect 392 18187 572 18196
rect 1634 18187 1814 18196
rect 2620 11752 3060 11761
rect 2620 11303 3060 11312
rect 2580 3334 3020 3343
rect 2580 2885 3020 2894
rect 7113 1659 7718 1668
rect 7718 1584 38332 1659
rect 7718 1144 11718 1584
rect 12158 1144 19492 1584
rect 19932 1578 38332 1584
rect 19932 1144 27266 1578
rect 7718 1138 27266 1144
rect 27706 1570 38332 1578
rect 27706 1138 35040 1570
rect 7718 1130 35040 1138
rect 35480 1130 38332 1570
rect 7718 1054 38332 1130
rect 7113 1045 7718 1054
<< via4 >>
rect 10517 30375 10604 30462
rect 11285 30375 11372 30462
rect 12053 30375 12140 30462
rect 12821 30375 12908 30462
rect 13589 30375 13676 30462
rect 14357 30375 14444 30462
rect 15125 30375 15212 30462
rect 15893 30375 15980 30462
rect 16661 30375 16748 30462
rect 17429 30375 17516 30462
rect 18197 30375 18284 30462
rect 18965 30375 19052 30462
rect 19733 30375 19820 30462
rect 20501 30375 20588 30462
rect 21269 30375 21356 30462
rect 22037 30375 22124 30462
rect 22805 30375 22892 30462
rect 23573 30375 23660 30462
rect 30480 30362 30576 30458
rect 31248 30362 31344 30458
rect 32016 30362 32112 30458
rect 32784 30362 32880 30458
rect 33552 30362 33648 30458
rect 34320 30362 34416 30458
rect 35088 30362 35184 30458
rect 35856 30362 35952 30458
rect 36624 30362 36720 30458
rect 37392 30362 37488 30458
rect 38160 30362 38256 30458
rect 2686 27120 3126 27560
rect 416 24596 596 24776
rect 418 21396 598 21576
rect 2656 19884 3096 20324
rect 392 18196 572 18376
rect 2620 11312 3060 11752
rect 2580 2894 3020 3334
rect 7113 1054 7718 1659
rect 11718 1144 12158 1584
rect 19492 1144 19932 1584
rect 27266 1138 27706 1578
rect 35040 1130 35480 1570
<< metal5 >>
rect 958 30596 1732 30678
rect 791 30592 1732 30596
rect 5922 30592 5982 30996
rect 6690 30592 6750 30996
rect 7458 30592 7518 30996
rect 8226 30592 8286 30996
rect 8994 30592 9054 30996
rect 9762 30592 9822 30996
rect 791 30532 9822 30592
rect 791 30456 1732 30532
rect 10530 30522 10590 30996
rect 11298 30522 11358 30996
rect 12066 30522 12126 30996
rect 12834 30522 12894 30996
rect 13602 30522 13662 30996
rect 14370 30522 14430 30996
rect 15138 30522 15198 30996
rect 15906 30522 15966 30996
rect 16674 30522 16734 30996
rect 17442 30522 17502 30996
rect 18210 30522 18270 30996
rect 18978 30522 19038 30996
rect 19746 30522 19806 30996
rect 20514 30522 20574 30996
rect 21282 30522 21342 30996
rect 22050 30522 22110 30996
rect 22818 30522 22878 30996
rect 23586 30522 23646 30996
rect 24354 30796 24414 30996
rect 25122 30796 25182 30996
rect 25890 30796 25950 30996
rect 26658 30796 26718 30996
rect 27426 30796 27486 30996
rect 28194 30796 28254 30996
rect 28962 30796 29022 30996
rect 29730 30796 29790 30996
rect 30498 30522 30558 30996
rect 31266 30522 31326 30996
rect 32034 30522 32094 30996
rect 32802 30522 32862 30996
rect 33570 30522 33630 30996
rect 34338 30522 34398 30996
rect 35106 30522 35166 30996
rect 35874 30522 35934 30996
rect 36642 30522 36702 30996
rect 37410 30522 37470 30996
rect 38178 30522 38238 30996
rect 800 30446 1732 30456
rect 10517 30462 10604 30522
rect 800 27560 1240 30446
rect 10517 30366 10604 30375
rect 11285 30462 11372 30522
rect 11285 30366 11372 30375
rect 12053 30462 12140 30522
rect 12053 30366 12140 30375
rect 12821 30462 12908 30522
rect 12821 30366 12908 30375
rect 13589 30462 13676 30522
rect 13589 30366 13676 30375
rect 14357 30462 14444 30522
rect 14357 30366 14444 30375
rect 15125 30462 15212 30522
rect 15125 30366 15212 30375
rect 15893 30462 15980 30522
rect 15893 30366 15980 30375
rect 16661 30462 16748 30522
rect 16661 30366 16748 30375
rect 17429 30462 17516 30522
rect 17429 30366 17516 30375
rect 18197 30462 18284 30522
rect 18197 30366 18284 30375
rect 18965 30462 19052 30522
rect 18965 30366 19052 30375
rect 19733 30462 19820 30522
rect 19733 30366 19820 30375
rect 20501 30462 20588 30522
rect 20501 30366 20588 30375
rect 21269 30462 21356 30522
rect 21269 30366 21356 30375
rect 22037 30462 22124 30522
rect 22037 30366 22124 30375
rect 22805 30462 22892 30522
rect 22805 30366 22892 30375
rect 23573 30462 23660 30522
rect 23573 30366 23660 30375
rect 30480 30458 30576 30522
rect 30480 30353 30576 30362
rect 31248 30458 31344 30522
rect 31248 30353 31344 30362
rect 32016 30458 32112 30522
rect 32016 30353 32112 30362
rect 32784 30458 32880 30522
rect 32784 30353 32880 30362
rect 33552 30458 33648 30522
rect 33552 30353 33648 30362
rect 34320 30458 34416 30522
rect 34320 30353 34416 30362
rect 35088 30458 35184 30522
rect 35088 30353 35184 30362
rect 35856 30458 35952 30522
rect 35856 30353 35952 30362
rect 36624 30458 36720 30522
rect 36624 30353 36720 30362
rect 37392 30458 37488 30522
rect 37392 30353 37488 30362
rect 38160 30458 38256 30522
rect 38160 30353 38256 30362
rect 800 27120 2686 27560
rect 3126 27120 3135 27560
rect 0 24596 416 24776
rect 596 24596 605 24776
rect 0 21396 418 21576
rect 598 21396 607 21576
rect 800 20324 1240 27120
rect 800 19884 2656 20324
rect 3096 19884 3105 20324
rect 0 18196 392 18376
rect 572 18196 581 18376
rect 0 14996 200 15176
rect 800 11752 1240 19884
rect 800 11312 2620 11752
rect 3060 11312 3069 11752
rect 800 3334 1240 11312
rect 800 2894 2580 3334
rect 3020 2894 3029 3334
rect 800 1576 1240 2894
rect 6420 1576 7113 1659
rect 800 1136 7113 1576
rect 800 0 1240 1136
rect 6420 1054 7113 1136
rect 7718 1054 7727 1659
rect 10448 796 10968 2534
rect 11718 1584 12158 2488
rect 11718 1135 12158 1144
rect 18214 796 18734 2540
rect 19492 1584 19932 2372
rect 19492 1135 19932 1144
rect 25998 796 26518 2556
rect 27266 1578 27706 2372
rect 27266 1129 27706 1138
rect 33750 796 34270 2482
rect 35040 1570 35480 2372
rect 35040 1121 35480 1130
rect 39800 796 40240 30596
rect 7168 356 40240 796
rect 7254 276 40240 356
rect 39800 0 40240 276
use r2r_dac  blue_dac
timestamp 1746810912
transform 0 1 3516 -1 0 10920
box -142 -18 7922 2062
use controller  controller_0
timestamp 1746816402
transform 1 0 7402 0 1 1156
box 0 700 31805 29000
use r2r_dac  green_dac
timestamp 1746810912
transform 0 1 3512 -1 0 19246
box -142 -18 7922 2062
use r2r_dac  red_dac
timestamp 1746810912
transform 0 1 3492 -1 0 27566
box -142 -18 7922 2062
<< labels >>
flabel metal5 s 37410 30796 37470 30996 4 FreeSans 320 0 0 0 clk
port 2 nsew
flabel metal5 s 38178 30796 38238 30996 4 FreeSans 320 0 0 0 ena
port 3 nsew
flabel metal5 s 36642 30796 36702 30996 4 FreeSans 320 0 0 0 rst_n
port 4 nsew
flabel metal5 s 35874 30796 35934 30996 4 FreeSans 320 0 0 0 ui_in[0]
port 5 nsew
flabel metal5 s 35106 30796 35166 30996 4 FreeSans 320 0 0 0 ui_in[1]
port 6 nsew
flabel metal5 s 34338 30796 34398 30996 4 FreeSans 320 0 0 0 ui_in[2]
port 7 nsew
flabel metal5 s 33570 30796 33630 30996 4 FreeSans 320 0 0 0 ui_in[3]
port 8 nsew
flabel metal5 s 32802 30796 32862 30996 4 FreeSans 320 0 0 0 ui_in[4]
port 9 nsew
flabel metal5 s 32034 30796 32094 30996 4 FreeSans 320 0 0 0 ui_in[5]
port 10 nsew
flabel metal5 s 31266 30796 31326 30996 4 FreeSans 320 0 0 0 ui_in[6]
port 11 nsew
flabel metal5 s 30498 30796 30558 30996 4 FreeSans 320 0 0 0 ui_in[7]
port 12 nsew
flabel metal5 s 29730 30796 29790 30996 4 FreeSans 320 0 0 0 uio_in[0]
port 13 nsew
flabel metal5 s 28962 30796 29022 30996 4 FreeSans 320 0 0 0 uio_in[1]
port 14 nsew
flabel metal5 s 28194 30796 28254 30996 4 FreeSans 320 0 0 0 uio_in[2]
port 15 nsew
flabel metal5 s 27426 30796 27486 30996 4 FreeSans 320 0 0 0 uio_in[3]
port 16 nsew
flabel metal5 s 26658 30796 26718 30996 4 FreeSans 320 0 0 0 uio_in[4]
port 17 nsew
flabel metal5 s 25890 30796 25950 30996 4 FreeSans 320 0 0 0 uio_in[5]
port 18 nsew
flabel metal5 s 25122 30796 25182 30996 4 FreeSans 320 0 0 0 uio_in[6]
port 19 nsew
flabel metal5 s 24354 30796 24414 30996 4 FreeSans 320 0 0 0 uio_in[7]
port 20 nsew
flabel metal5 s 11298 30796 11358 30996 4 FreeSans 320 0 0 0 uio_oe[0]
port 21 nsew
flabel metal5 s 10530 30796 10590 30996 4 FreeSans 320 0 0 0 uio_oe[1]
port 22 nsew
flabel metal5 s 9762 30796 9822 30996 4 FreeSans 320 0 0 0 uio_oe[2]
port 23 nsew
flabel metal5 s 8994 30796 9054 30996 4 FreeSans 320 0 0 0 uio_oe[3]
port 24 nsew
flabel metal5 s 8226 30796 8286 30996 4 FreeSans 320 0 0 0 uio_oe[4]
port 25 nsew
flabel metal5 s 7458 30796 7518 30996 4 FreeSans 320 0 0 0 uio_oe[5]
port 26 nsew
flabel metal5 s 6690 30796 6750 30996 4 FreeSans 320 0 0 0 uio_oe[6]
port 27 nsew
flabel metal5 s 5922 30796 5982 30996 4 FreeSans 320 0 0 0 uio_oe[7]
port 28 nsew
flabel metal5 s 17442 30796 17502 30996 4 FreeSans 320 0 0 0 uio_out[0]
port 29 nsew
flabel metal5 s 16674 30796 16734 30996 4 FreeSans 320 0 0 0 uio_out[1]
port 30 nsew
flabel metal5 s 15906 30796 15966 30996 4 FreeSans 320 0 0 0 uio_out[2]
port 31 nsew
flabel metal5 s 15138 30796 15198 30996 4 FreeSans 320 0 0 0 uio_out[3]
port 32 nsew
flabel metal5 s 14370 30796 14430 30996 4 FreeSans 320 0 0 0 uio_out[4]
port 33 nsew
flabel metal5 s 13602 30796 13662 30996 4 FreeSans 320 0 0 0 uio_out[5]
port 34 nsew
flabel metal5 s 12834 30796 12894 30996 4 FreeSans 320 0 0 0 uio_out[6]
port 35 nsew
flabel metal5 s 12066 30796 12126 30996 4 FreeSans 320 0 0 0 uio_out[7]
port 36 nsew
flabel metal5 s 23586 30796 23646 30996 4 FreeSans 320 0 0 0 uo_out[0]
port 37 nsew
flabel metal5 s 22818 30796 22878 30996 4 FreeSans 320 0 0 0 uo_out[1]
port 38 nsew
flabel metal5 s 22050 30796 22110 30996 4 FreeSans 320 0 0 0 uo_out[2]
port 39 nsew
flabel metal5 s 21282 30796 21342 30996 4 FreeSans 320 0 0 0 uo_out[3]
port 40 nsew
flabel metal5 s 20514 30796 20574 30996 4 FreeSans 320 0 0 0 uo_out[4]
port 41 nsew
flabel metal5 s 19746 30796 19806 30996 4 FreeSans 320 0 0 0 uo_out[5]
port 42 nsew
flabel metal5 s 18978 30796 19038 30996 4 FreeSans 320 0 0 0 uo_out[6]
port 43 nsew
flabel metal5 s 18210 30796 18270 30996 4 FreeSans 320 0 0 0 uo_out[7]
port 44 nsew
flabel metal5 s 0 24596 200 24776 0 FreeSans 320 0 0 0 ua[0]
port 45 nsew
flabel metal5 s 0 21396 200 21576 0 FreeSans 320 0 0 0 ua[1]
port 46 nsew
flabel metal5 s 0 18196 200 18376 0 FreeSans 320 0 0 0 ua[2]
port 47 nsew
flabel metal5 s 0 14996 200 15176 0 FreeSans 320 0 0 0 ua[3]
port 48 nsew
flabel metal5 s 800 0 1240 30596 0 FreeSans 320 0 0 0 VGND
port 49 nsew
flabel metal5 s 39800 0 40240 30596 0 FreeSans 320 0 0 0 VPWR
port 50 nsew
<< properties >>
string FIXED_BBOX 0 0 40416 30996
<< end >>
