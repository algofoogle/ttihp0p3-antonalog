magic
tech ihp-sg13g2
magscale 1 2
timestamp 1747056038
<< nwell >>
rect -48 350 624 834
<< pwell >>
rect 16 56 546 296
rect -26 -56 602 56
<< nmos >>
rect 120 122 146 270
rect 221 122 247 270
rect 324 122 350 270
rect 426 122 452 270
<< pmos >>
rect 120 426 146 650
rect 222 426 248 650
rect 324 426 350 650
rect 426 426 452 650
<< ndiff >>
rect 42 256 120 270
rect 42 224 56 256
rect 88 224 120 256
rect 42 168 120 224
rect 42 136 56 168
rect 88 136 120 168
rect 42 122 120 136
rect 146 122 221 270
rect 247 122 324 270
rect 350 122 426 270
rect 452 256 520 270
rect 452 224 474 256
rect 506 224 520 256
rect 452 168 520 224
rect 452 136 474 168
rect 506 136 520 168
rect 452 122 520 136
<< pdiff >>
rect 52 635 120 650
rect 52 603 66 635
rect 98 603 120 635
rect 52 556 120 603
rect 52 524 66 556
rect 98 524 120 556
rect 52 472 120 524
rect 52 440 66 472
rect 98 440 120 472
rect 52 426 120 440
rect 146 635 222 650
rect 146 603 168 635
rect 200 603 222 635
rect 146 556 222 603
rect 146 524 168 556
rect 200 524 222 556
rect 146 472 222 524
rect 146 440 168 472
rect 200 440 222 472
rect 146 426 222 440
rect 248 635 324 650
rect 248 603 270 635
rect 302 603 324 635
rect 248 556 324 603
rect 248 524 270 556
rect 302 524 324 556
rect 248 426 324 524
rect 350 635 426 650
rect 350 603 372 635
rect 404 603 426 635
rect 350 556 426 603
rect 350 524 372 556
rect 404 524 426 556
rect 350 472 426 524
rect 350 440 372 472
rect 404 440 426 472
rect 350 426 426 440
rect 452 635 520 650
rect 452 603 474 635
rect 506 603 520 635
rect 452 556 520 603
rect 452 524 474 556
rect 506 524 520 556
rect 452 426 520 524
<< ndiffc >>
rect 56 224 88 256
rect 56 136 88 168
rect 474 224 506 256
rect 474 136 506 168
<< pdiffc >>
rect 66 603 98 635
rect 66 524 98 556
rect 66 440 98 472
rect 168 603 200 635
rect 168 524 200 556
rect 168 440 200 472
rect 270 603 302 635
rect 270 524 302 556
rect 372 603 404 635
rect 372 524 404 556
rect 372 440 404 472
rect 474 603 506 635
rect 474 524 506 556
<< psubdiff >>
rect 0 16 576 30
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 576 16
rect 0 -30 576 -16
<< nsubdiff >>
rect 0 772 576 786
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 576 772
rect 0 726 576 740
<< psubdiffcont >>
rect 32 -16 64 16
rect 128 -16 160 16
rect 224 -16 256 16
rect 320 -16 352 16
rect 416 -16 448 16
rect 512 -16 544 16
<< nsubdiffcont >>
rect 32 740 64 772
rect 128 740 160 772
rect 224 740 256 772
rect 320 740 352 772
rect 416 740 448 772
rect 512 740 544 772
<< poly >>
rect 120 650 146 686
rect 222 650 248 686
rect 324 650 350 686
rect 426 650 452 686
rect 120 374 146 426
rect 222 380 248 426
rect 72 360 146 374
rect 72 328 86 360
rect 118 328 146 360
rect 72 314 146 328
rect 205 363 265 380
rect 324 371 350 426
rect 426 393 452 426
rect 409 379 469 393
rect 205 331 219 363
rect 251 331 265 363
rect 205 317 265 331
rect 307 357 367 371
rect 307 325 321 357
rect 353 325 367 357
rect 409 347 423 379
rect 455 347 469 379
rect 409 333 469 347
rect 120 270 146 314
rect 221 270 247 317
rect 307 311 367 325
rect 324 270 350 311
rect 426 270 452 333
rect 120 86 146 122
rect 221 86 247 122
rect 324 86 350 122
rect 426 86 452 122
<< polycont >>
rect 86 328 118 360
rect 219 331 251 363
rect 321 325 353 357
rect 423 347 455 379
<< metal1 >>
rect 0 772 576 800
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 576 772
rect 0 712 576 740
rect 56 635 108 712
rect 56 603 66 635
rect 98 603 108 635
rect 56 556 108 603
rect 56 524 66 556
rect 98 524 108 556
rect 56 472 108 524
rect 56 440 66 472
rect 98 440 108 472
rect 56 436 108 440
rect 158 635 210 645
rect 158 603 168 635
rect 200 603 210 635
rect 158 556 210 603
rect 158 524 168 556
rect 200 524 210 556
rect 158 479 210 524
rect 260 635 312 712
rect 260 603 270 635
rect 302 603 312 635
rect 260 556 312 603
rect 260 524 270 556
rect 302 524 312 556
rect 260 515 312 524
rect 362 635 414 645
rect 362 603 372 635
rect 404 603 414 635
rect 362 556 414 603
rect 362 524 372 556
rect 404 524 414 556
rect 362 479 414 524
rect 464 635 516 712
rect 464 603 474 635
rect 506 603 516 635
rect 464 556 516 603
rect 464 524 474 556
rect 506 524 516 556
rect 464 515 516 524
rect 158 472 540 479
rect 158 440 168 472
rect 200 440 372 472
rect 404 440 540 472
rect 158 436 540 440
rect 72 360 138 400
rect 72 328 86 360
rect 118 328 138 360
rect 72 310 138 328
rect 190 363 264 400
rect 190 331 219 363
rect 251 331 264 363
rect 190 310 264 331
rect 300 357 366 400
rect 300 325 321 357
rect 353 325 366 357
rect 300 310 366 325
rect 402 379 456 400
rect 402 347 423 379
rect 455 347 456 379
rect 402 310 456 347
rect 492 266 540 436
rect 45 256 99 266
rect 45 224 56 256
rect 88 224 99 256
rect 45 168 99 224
rect 45 136 56 168
rect 88 136 99 168
rect 45 44 99 136
rect 464 256 540 266
rect 464 224 474 256
rect 506 224 540 256
rect 464 168 540 224
rect 464 136 474 168
rect 506 136 540 168
rect 464 126 540 136
rect 0 16 576 44
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 576 16
rect 0 -44 576 -16
<< labels >>
flabel metal1 s 0 712 576 800 0 FreeSans 400 0 0 0 VDD
port 2 nsew
flabel metal1 s 492 126 540 479 0 FreeSans 400 0 0 0 Y
port 3 nsew
flabel metal1 s 300 310 366 400 0 FreeSans 400 0 0 0 B
port 4 nsew
flabel metal1 s 190 310 264 400 0 FreeSans 400 0 0 0 C
port 5 nsew
flabel metal1 s 0 -44 576 44 0 FreeSans 400 0 0 0 VSS
port 6 nsew
flabel metal1 s 402 310 456 400 0 FreeSans 400 0 0 0 A
port 7 nsew
flabel metal1 s 72 310 138 400 0 FreeSans 500 0 0 0 D
port 8 nsew
<< properties >>
string FIXED_BBOX 0 0 576 756
string GDS_END 195444
string GDS_FILE ../gds/controller.gds
string GDS_START 190770
<< end >>
