magic
tech ihp-sg13g2
timestamp 1747537721
<< nwell >>
rect -24 175 456 417
<< pwell >>
rect 247 136 427 146
rect 54 28 427 136
rect -13 -28 445 28
<< nmos >>
rect 101 59 114 123
rect 140 59 153 123
rect 179 59 192 123
rect 236 59 249 123
rect 287 59 300 133
rect 352 59 365 133
<< pmos >>
rect 74 234 87 318
rect 125 234 138 318
rect 176 234 189 318
rect 233 234 246 318
rect 287 206 300 318
rect 352 206 365 318
<< ndiff >>
rect 260 123 287 133
rect 67 116 101 123
rect 67 100 74 116
rect 90 100 101 116
rect 67 82 101 100
rect 67 66 74 82
rect 90 66 101 82
rect 67 59 101 66
rect 114 59 140 123
rect 153 59 179 123
rect 192 59 236 123
rect 249 116 287 123
rect 249 100 260 116
rect 276 100 287 116
rect 249 82 287 100
rect 249 66 260 82
rect 276 66 287 82
rect 249 59 287 66
rect 300 126 352 133
rect 300 110 325 126
rect 341 110 352 126
rect 300 82 352 110
rect 300 66 325 82
rect 341 66 352 82
rect 300 59 352 66
rect 365 126 414 133
rect 365 110 391 126
rect 407 110 414 126
rect 365 82 414 110
rect 365 66 391 82
rect 407 66 414 82
rect 365 59 414 66
<< pdiff >>
rect 40 311 74 318
rect 40 295 47 311
rect 63 295 74 311
rect 40 273 74 295
rect 40 257 47 273
rect 63 257 74 273
rect 40 234 74 257
rect 87 311 125 318
rect 87 295 98 311
rect 114 295 125 311
rect 87 257 125 295
rect 87 241 98 257
rect 114 241 125 257
rect 87 234 125 241
rect 138 311 176 318
rect 138 295 149 311
rect 165 295 176 311
rect 138 273 176 295
rect 138 257 149 273
rect 165 257 176 273
rect 138 234 176 257
rect 189 311 233 318
rect 189 295 203 311
rect 219 295 233 311
rect 189 257 233 295
rect 189 241 203 257
rect 219 241 233 257
rect 189 234 233 241
rect 246 311 287 318
rect 246 295 259 311
rect 275 295 287 311
rect 246 276 287 295
rect 246 260 259 276
rect 275 260 287 276
rect 246 234 287 260
rect 264 206 287 234
rect 300 311 352 318
rect 300 295 325 311
rect 341 295 352 311
rect 300 271 352 295
rect 300 255 325 271
rect 341 255 352 271
rect 300 229 352 255
rect 300 213 325 229
rect 341 213 352 229
rect 300 206 352 213
rect 365 311 414 318
rect 365 295 391 311
rect 407 295 414 311
rect 365 271 414 295
rect 365 255 391 271
rect 407 255 414 271
rect 365 229 414 255
rect 365 213 391 229
rect 407 213 414 229
rect 365 206 414 213
<< ndiffc >>
rect 74 100 90 116
rect 74 66 90 82
rect 260 100 276 116
rect 260 66 276 82
rect 325 110 341 126
rect 325 66 341 82
rect 391 110 407 126
rect 391 66 407 82
<< pdiffc >>
rect 47 295 63 311
rect 47 257 63 273
rect 98 295 114 311
rect 98 241 114 257
rect 149 295 165 311
rect 149 257 165 273
rect 203 295 219 311
rect 203 241 219 257
rect 259 295 275 311
rect 259 260 275 276
rect 325 295 341 311
rect 325 255 341 271
rect 325 213 341 229
rect 391 295 407 311
rect 391 255 407 271
rect 391 213 407 229
<< psubdiff >>
rect 0 8 432 15
rect 0 -8 16 8
rect 32 -8 64 8
rect 80 -8 112 8
rect 128 -8 160 8
rect 176 -8 208 8
rect 224 -8 256 8
rect 272 -8 304 8
rect 320 -8 352 8
rect 368 -8 400 8
rect 416 -8 432 8
rect 0 -15 432 -8
<< nsubdiff >>
rect 0 386 432 393
rect 0 370 16 386
rect 32 370 64 386
rect 80 370 112 386
rect 128 370 160 386
rect 176 370 208 386
rect 224 370 256 386
rect 272 370 304 386
rect 320 370 352 386
rect 368 370 400 386
rect 416 370 432 386
rect 0 363 432 370
<< psubdiffcont >>
rect 16 -8 32 8
rect 64 -8 80 8
rect 112 -8 128 8
rect 160 -8 176 8
rect 208 -8 224 8
rect 256 -8 272 8
rect 304 -8 320 8
rect 352 -8 368 8
rect 400 -8 416 8
<< nsubdiffcont >>
rect 16 370 32 386
rect 64 370 80 386
rect 112 370 128 386
rect 160 370 176 386
rect 208 370 224 386
rect 256 370 272 386
rect 304 370 320 386
rect 352 370 368 386
rect 400 370 416 386
<< poly >>
rect 74 318 87 336
rect 125 318 138 336
rect 176 318 189 336
rect 233 318 246 336
rect 287 318 300 336
rect 352 318 365 336
rect 74 226 87 234
rect 125 226 138 234
rect 73 201 91 226
rect 123 202 141 226
rect 176 213 189 234
rect 69 192 102 201
rect 69 176 77 192
rect 93 176 102 192
rect 69 158 102 176
rect 123 193 158 202
rect 176 201 212 213
rect 123 177 133 193
rect 149 177 158 193
rect 123 169 158 177
rect 179 192 212 201
rect 179 176 187 192
rect 203 176 212 192
rect 69 142 77 158
rect 93 145 102 158
rect 93 142 114 145
rect 69 130 114 142
rect 101 123 114 130
rect 140 123 153 169
rect 179 158 212 176
rect 179 142 187 158
rect 203 142 212 158
rect 233 190 246 234
rect 287 190 300 206
rect 352 190 365 206
rect 233 181 266 190
rect 233 165 241 181
rect 257 165 266 181
rect 233 157 266 165
rect 287 178 365 190
rect 287 162 295 178
rect 311 162 365 178
rect 179 134 212 142
rect 179 123 192 134
rect 236 123 249 157
rect 287 154 365 162
rect 287 133 300 154
rect 352 133 365 154
rect 101 41 114 59
rect 140 41 153 59
rect 179 41 192 59
rect 236 41 249 59
rect 287 41 300 59
rect 352 41 365 59
<< polycont >>
rect 77 176 93 192
rect 133 177 149 193
rect 187 176 203 192
rect 77 142 93 158
rect 187 142 203 158
rect 241 165 257 181
rect 295 162 311 178
<< metal1 >>
rect 0 386 432 400
rect 0 370 16 386
rect 32 370 64 386
rect 80 370 112 386
rect 128 370 160 386
rect 176 370 208 386
rect 224 370 256 386
rect 272 370 304 386
rect 320 370 352 386
rect 368 370 400 386
rect 416 370 432 386
rect 0 356 432 370
rect 42 311 68 356
rect 42 295 47 311
rect 63 295 68 311
rect 42 273 68 295
rect 42 257 47 273
rect 63 257 68 273
rect 42 256 68 257
rect 93 311 119 312
rect 93 295 98 311
rect 114 295 119 311
rect 93 257 119 295
rect 93 241 98 257
rect 114 241 119 257
rect 144 311 170 356
rect 144 295 149 311
rect 165 295 170 311
rect 144 273 170 295
rect 144 257 149 273
rect 165 257 170 273
rect 144 256 170 257
rect 198 311 224 312
rect 198 295 203 311
rect 219 295 224 311
rect 198 257 224 295
rect 254 311 280 356
rect 254 295 259 311
rect 275 295 280 311
rect 254 276 280 295
rect 254 260 259 276
rect 275 260 280 276
rect 254 258 280 260
rect 320 311 368 312
rect 320 295 325 311
rect 341 295 368 311
rect 320 271 368 295
rect 93 238 119 241
rect 198 241 203 257
rect 219 241 224 257
rect 198 238 224 241
rect 320 255 325 271
rect 341 255 368 271
rect 35 222 301 238
rect 35 117 52 222
rect 70 192 107 201
rect 70 176 77 192
rect 93 176 107 192
rect 70 158 107 176
rect 70 142 77 158
rect 93 142 107 158
rect 70 135 107 142
rect 125 193 156 202
rect 125 177 133 193
rect 149 177 156 193
rect 35 116 99 117
rect 35 100 74 116
rect 90 100 99 116
rect 35 82 99 100
rect 35 66 74 82
rect 90 66 99 82
rect 125 66 156 177
rect 179 192 212 201
rect 179 176 187 192
rect 203 176 212 192
rect 179 158 212 176
rect 179 142 187 158
rect 203 142 212 158
rect 231 181 266 200
rect 231 165 241 181
rect 257 165 266 181
rect 231 157 266 165
rect 285 187 301 222
rect 320 229 368 255
rect 320 213 325 229
rect 341 213 368 229
rect 386 311 412 356
rect 386 295 391 311
rect 407 295 412 311
rect 386 271 412 295
rect 386 255 391 271
rect 407 255 412 271
rect 386 229 412 255
rect 386 213 391 229
rect 407 213 412 229
rect 320 207 368 213
rect 285 178 320 187
rect 285 162 295 178
rect 311 162 320 178
rect 285 154 320 162
rect 179 66 212 142
rect 352 126 368 207
rect 255 116 281 121
rect 255 100 260 116
rect 276 100 281 116
rect 255 82 281 100
rect 255 66 260 82
rect 276 66 281 82
rect 35 64 99 66
rect 255 22 281 66
rect 320 110 325 126
rect 341 110 368 126
rect 320 82 368 110
rect 320 66 325 82
rect 341 66 368 82
rect 320 64 368 66
rect 386 110 391 126
rect 407 110 412 126
rect 386 82 412 110
rect 386 66 391 82
rect 407 66 412 82
rect 386 22 412 66
rect 0 8 432 22
rect 0 -8 16 8
rect 32 -8 64 8
rect 80 -8 112 8
rect 128 -8 160 8
rect 176 -8 208 8
rect 224 -8 256 8
rect 272 -8 304 8
rect 320 -8 352 8
rect 368 -8 400 8
rect 416 -8 432 8
rect 0 -22 432 -8
<< labels >>
flabel metal1 s 320 207 368 312 0 FreeSans 200 0 0 0 X
port 2 nsew
flabel metal1 s 125 66 156 202 0 FreeSans 200 0 0 0 B
port 3 nsew
flabel metal1 s 70 135 107 201 0 FreeSans 200 0 0 0 A
port 4 nsew
flabel metal1 s 0 356 432 400 0 FreeSans 200 0 0 0 VDD
port 5 nsew
flabel metal1 s 0 -22 432 22 0 FreeSans 200 0 0 0 VSS
port 6 nsew
flabel metal1 s 179 66 212 201 0 FreeSans 200 0 0 0 C
port 7 nsew
flabel metal1 s 231 157 266 200 0 FreeSans 200 0 0 0 D
port 8 nsew
<< properties >>
string FIXED_BBOX 0 0 432 378
string GDS_END 113568
string GDS_FILE ../gds/controller.gds
string GDS_START 107454
<< end >>
