magic
tech ihp-sg13g2
magscale 1 2
timestamp 1746816402
<< nwell >>
rect -48 350 528 834
<< pwell >>
rect 63 56 481 292
rect -26 -56 506 56
<< nmos >>
rect 157 118 183 266
rect 259 118 285 266
rect 361 138 387 266
<< pmos >>
rect 157 412 183 636
rect 259 412 285 636
rect 361 427 387 627
<< ndiff >>
rect 89 251 157 266
rect 89 219 103 251
rect 135 219 157 251
rect 89 164 157 219
rect 89 132 103 164
rect 135 132 157 164
rect 89 118 157 132
rect 183 251 259 266
rect 183 219 205 251
rect 237 219 259 251
rect 183 164 259 219
rect 183 132 205 164
rect 237 132 259 164
rect 183 118 259 132
rect 285 195 361 266
rect 285 163 307 195
rect 339 163 361 195
rect 285 138 361 163
rect 387 252 455 266
rect 387 220 409 252
rect 441 220 455 252
rect 387 184 455 220
rect 387 152 409 184
rect 441 152 455 184
rect 387 138 455 152
rect 285 118 347 138
<< pdiff >>
rect 26 621 157 636
rect 26 589 40 621
rect 72 589 157 621
rect 26 534 157 589
rect 26 502 40 534
rect 72 502 157 534
rect 26 459 157 502
rect 26 427 40 459
rect 72 427 157 459
rect 26 412 157 427
rect 183 458 259 636
rect 183 426 205 458
rect 237 426 259 458
rect 183 412 259 426
rect 285 627 347 636
rect 285 613 361 627
rect 285 581 307 613
rect 339 581 361 613
rect 285 427 361 581
rect 387 609 455 627
rect 387 577 409 609
rect 441 577 455 609
rect 387 541 455 577
rect 387 509 409 541
rect 441 509 455 541
rect 387 473 455 509
rect 387 441 409 473
rect 441 441 455 473
rect 387 427 455 441
rect 285 412 347 427
<< ndiffc >>
rect 103 219 135 251
rect 103 132 135 164
rect 205 219 237 251
rect 205 132 237 164
rect 307 163 339 195
rect 409 220 441 252
rect 409 152 441 184
<< pdiffc >>
rect 40 589 72 621
rect 40 502 72 534
rect 40 427 72 459
rect 205 426 237 458
rect 307 581 339 613
rect 409 577 441 609
rect 409 509 441 541
rect 409 441 441 473
<< psubdiff >>
rect 0 16 480 30
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 480 16
rect 0 -30 480 -16
<< nsubdiff >>
rect 0 772 480 786
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 480 772
rect 0 726 480 740
<< psubdiffcont >>
rect 32 -16 64 16
rect 128 -16 160 16
rect 224 -16 256 16
rect 320 -16 352 16
rect 416 -16 448 16
<< nsubdiffcont >>
rect 32 740 64 772
rect 128 740 160 772
rect 224 740 256 772
rect 320 740 352 772
rect 416 740 448 772
<< poly >>
rect 157 636 183 672
rect 259 636 285 672
rect 361 627 387 663
rect 157 370 183 412
rect 259 370 285 412
rect 21 353 285 370
rect 21 321 38 353
rect 70 321 106 353
rect 138 321 285 353
rect 21 304 285 321
rect 157 266 183 304
rect 259 266 285 304
rect 361 380 387 427
rect 361 363 431 380
rect 361 331 382 363
rect 414 331 431 363
rect 361 314 431 331
rect 361 266 387 314
rect 157 82 183 118
rect 259 82 285 118
rect 361 102 387 138
<< polycont >>
rect 38 321 70 353
rect 106 321 138 353
rect 382 331 414 363
<< metal1 >>
rect 0 772 480 800
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 480 772
rect 0 712 480 740
rect 30 621 82 712
rect 30 589 40 621
rect 72 589 82 621
rect 30 534 82 589
rect 297 613 349 712
rect 297 581 307 613
rect 339 581 349 613
rect 297 579 349 581
rect 394 609 452 620
rect 394 577 409 609
rect 441 577 452 609
rect 394 542 452 577
rect 30 502 40 534
rect 72 502 82 534
rect 30 459 82 502
rect 30 427 40 459
rect 72 427 82 459
rect 30 424 82 427
rect 121 541 452 542
rect 121 510 409 541
rect 121 370 153 510
rect 21 353 153 370
rect 21 321 38 353
rect 70 321 106 353
rect 138 321 153 353
rect 21 304 153 321
rect 189 458 255 474
rect 189 426 205 458
rect 237 426 255 458
rect 93 251 145 255
rect 93 219 103 251
rect 135 219 145 251
rect 93 164 145 219
rect 93 132 103 164
rect 135 132 145 164
rect 93 44 145 132
rect 189 251 255 426
rect 189 219 205 251
rect 237 219 255 251
rect 299 278 331 510
rect 394 509 409 510
rect 441 509 452 541
rect 394 473 452 509
rect 394 441 409 473
rect 441 441 452 473
rect 394 436 452 441
rect 367 363 455 400
rect 367 331 382 363
rect 414 331 455 363
rect 367 314 455 331
rect 299 252 451 278
rect 299 246 409 252
rect 189 164 255 219
rect 399 220 409 246
rect 441 220 451 252
rect 189 132 205 164
rect 237 132 255 164
rect 189 127 255 132
rect 297 195 349 199
rect 297 163 307 195
rect 339 163 349 195
rect 297 44 349 163
rect 399 184 451 220
rect 399 152 409 184
rect 441 152 451 184
rect 399 144 451 152
rect 0 16 480 44
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 480 16
rect 0 -44 480 -16
<< labels >>
flabel metal1 s 0 -44 480 44 0 FreeSans 400 0 0 0 VSS
port 2 nsew
flabel metal1 s 0 712 480 800 0 FreeSans 400 0 0 0 VDD
port 3 nsew
flabel metal1 s 189 127 255 474 0 FreeSans 400 0 0 0 X
port 4 nsew
flabel metal1 s 367 314 455 400 0 FreeSans 400 0 0 0 A
port 5 nsew
<< properties >>
string FIXED_BBOX 0 0 480 756
string GDS_END 27744
string GDS_FILE ../gds/controller.gds
string GDS_START 23448
<< end >>
