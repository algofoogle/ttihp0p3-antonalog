magic
tech ihp-sg13g2
timestamp 1747537721
<< nwell >>
rect -24 175 360 417
<< pwell >>
rect 25 28 336 157
rect -13 -28 349 28
<< nmos >>
rect 72 80 85 144
rect 123 80 136 144
rect 174 80 187 144
rect 225 70 238 144
rect 276 70 289 144
<< pmos >>
rect 72 235 85 319
rect 123 235 136 319
rect 174 235 187 319
rect 225 217 238 329
rect 276 217 289 329
<< ndiff >>
rect 38 126 72 144
rect 38 110 45 126
rect 61 110 72 126
rect 38 80 72 110
rect 85 80 123 144
rect 136 80 174 144
rect 187 105 225 144
rect 187 89 198 105
rect 214 89 225 105
rect 187 80 225 89
rect 194 70 225 80
rect 238 131 276 144
rect 238 115 249 131
rect 265 115 276 131
rect 238 97 276 115
rect 238 81 249 97
rect 265 81 276 97
rect 238 70 276 81
rect 289 97 323 144
rect 289 81 300 97
rect 316 81 323 97
rect 289 70 323 81
<< pdiff >>
rect 194 319 225 329
rect 38 309 72 319
rect 38 293 45 309
rect 61 293 72 309
rect 38 263 72 293
rect 38 247 45 263
rect 61 247 72 263
rect 38 235 72 247
rect 85 290 123 319
rect 85 274 96 290
rect 112 274 123 290
rect 85 235 123 274
rect 136 306 174 319
rect 136 290 147 306
rect 163 290 174 306
rect 136 267 174 290
rect 136 251 147 267
rect 163 251 174 267
rect 136 235 174 251
rect 187 313 225 319
rect 187 297 198 313
rect 214 297 225 313
rect 187 279 225 297
rect 187 263 198 279
rect 214 263 225 279
rect 187 235 225 263
rect 202 217 225 235
rect 238 322 276 329
rect 238 306 249 322
rect 265 306 276 322
rect 238 286 276 306
rect 238 270 249 286
rect 265 270 276 286
rect 238 217 276 270
rect 289 322 324 329
rect 289 306 301 322
rect 317 306 324 322
rect 289 217 324 306
<< ndiffc >>
rect 45 110 61 126
rect 198 89 214 105
rect 249 115 265 131
rect 249 81 265 97
rect 300 81 316 97
<< pdiffc >>
rect 45 293 61 309
rect 45 247 61 263
rect 96 274 112 290
rect 147 290 163 306
rect 147 251 163 267
rect 198 297 214 313
rect 198 263 214 279
rect 249 306 265 322
rect 249 270 265 286
rect 301 306 317 322
<< psubdiff >>
rect 0 8 336 15
rect 0 -8 16 8
rect 32 -8 64 8
rect 80 -8 112 8
rect 128 -8 160 8
rect 176 -8 208 8
rect 224 -8 256 8
rect 272 -8 304 8
rect 320 -8 336 8
rect 0 -15 336 -8
<< nsubdiff >>
rect 0 386 336 393
rect 0 370 16 386
rect 32 370 64 386
rect 80 370 112 386
rect 128 370 160 386
rect 176 370 208 386
rect 224 370 256 386
rect 272 370 304 386
rect 320 370 336 386
rect 0 363 336 370
<< psubdiffcont >>
rect 16 -8 32 8
rect 64 -8 80 8
rect 112 -8 128 8
rect 160 -8 176 8
rect 208 -8 224 8
rect 256 -8 272 8
rect 304 -8 320 8
<< nsubdiffcont >>
rect 16 370 32 386
rect 64 370 80 386
rect 112 370 128 386
rect 160 370 176 386
rect 208 370 224 386
rect 256 370 272 386
rect 304 370 320 386
<< poly >>
rect 72 319 85 337
rect 123 319 136 337
rect 174 319 187 337
rect 225 329 238 350
rect 276 329 289 350
rect 72 144 85 235
rect 123 198 136 235
rect 174 200 187 235
rect 225 206 238 217
rect 276 206 289 217
rect 109 189 142 198
rect 109 173 117 189
rect 133 173 142 189
rect 109 165 142 173
rect 173 191 206 200
rect 173 175 181 191
rect 197 175 206 191
rect 173 167 206 175
rect 225 198 289 206
rect 225 182 240 198
rect 256 182 289 198
rect 225 173 289 182
rect 123 144 136 165
rect 174 144 187 167
rect 225 144 238 173
rect 276 144 289 173
rect 72 73 85 80
rect 35 66 102 73
rect 35 50 43 66
rect 59 50 77 66
rect 93 50 102 66
rect 123 54 136 80
rect 174 54 187 80
rect 225 52 238 70
rect 276 51 289 70
rect 35 39 102 50
<< polycont >>
rect 117 173 133 189
rect 181 175 197 191
rect 240 182 256 198
rect 43 50 59 66
rect 77 50 93 66
<< metal1 >>
rect 0 386 336 400
rect 0 370 16 386
rect 32 370 64 386
rect 80 370 112 386
rect 128 370 160 386
rect 176 370 208 386
rect 224 370 256 386
rect 272 370 304 386
rect 320 370 336 386
rect 0 356 336 370
rect 40 309 66 311
rect 40 293 45 309
rect 61 293 66 309
rect 40 263 66 293
rect 91 290 117 356
rect 193 313 219 356
rect 91 274 96 290
rect 112 274 117 290
rect 91 273 117 274
rect 142 306 168 308
rect 142 290 147 306
rect 163 290 168 306
rect 40 247 45 263
rect 61 247 66 263
rect 40 232 66 247
rect 142 267 168 290
rect 142 251 147 267
rect 163 251 168 267
rect 193 297 198 313
rect 214 297 219 313
rect 193 279 219 297
rect 193 263 198 279
rect 214 263 219 279
rect 193 261 219 263
rect 243 322 270 336
rect 243 306 249 322
rect 265 306 270 322
rect 243 286 270 306
rect 295 322 322 356
rect 295 306 301 322
rect 317 306 322 322
rect 295 287 322 306
rect 243 270 249 286
rect 265 270 270 286
rect 243 269 270 270
rect 243 251 306 269
rect 142 232 168 251
rect 40 216 240 232
rect 40 126 66 216
rect 224 206 240 216
rect 224 198 264 206
rect 109 189 154 198
rect 109 173 117 189
rect 133 173 154 189
rect 109 140 154 173
rect 173 191 206 195
rect 173 175 181 191
rect 197 175 206 191
rect 173 140 206 175
rect 224 182 240 198
rect 256 182 264 198
rect 224 173 264 182
rect 283 155 306 251
rect 40 110 45 126
rect 61 110 66 126
rect 244 131 306 155
rect 244 115 249 131
rect 265 129 306 131
rect 265 115 270 129
rect 40 109 66 110
rect 122 79 159 109
rect 35 66 159 79
rect 35 50 43 66
rect 59 50 77 66
rect 93 50 159 66
rect 35 47 159 50
rect 193 105 219 114
rect 193 89 198 105
rect 214 89 219 105
rect 193 22 219 89
rect 244 97 270 115
rect 244 81 249 97
rect 265 81 270 97
rect 244 77 270 81
rect 295 97 321 109
rect 295 81 300 97
rect 316 81 321 97
rect 295 22 321 81
rect 0 8 336 22
rect 0 -8 16 8
rect 32 -8 64 8
rect 80 -8 112 8
rect 128 -8 160 8
rect 176 -8 208 8
rect 224 -8 256 8
rect 272 -8 304 8
rect 320 -8 336 8
rect 0 -22 336 -8
<< labels >>
flabel metal1 s 244 129 306 155 0 FreeSans 200 0 0 0 X
port 2 nsew
flabel metal1 s 109 140 154 198 0 FreeSans 200 0 0 0 B
port 3 nsew
flabel metal1 s 0 356 336 400 0 FreeSans 200 0 0 0 VDD
port 4 nsew
flabel metal1 s 0 -22 336 22 0 FreeSans 200 0 0 0 VSS
port 5 nsew
flabel metal1 s 173 140 206 195 0 FreeSans 200 0 0 0 C
port 6 nsew
flabel metal1 s 122 47 159 109 0 FreeSans 200 0 0 0 A
port 7 nsew
<< properties >>
string FIXED_BBOX 0 0 336 378
string GDS_END 226730
string GDS_FILE ../gds/controller.gds
string GDS_START 220982
<< end >>
