magic
tech ihp-sg13g2
magscale 1 2
timestamp 1747537721
<< nwell >>
rect -48 350 720 834
<< pwell >>
rect 427 254 635 292
rect 47 56 635 254
rect -26 -56 698 56
<< nmos >>
rect 141 118 167 228
rect 243 118 269 228
rect 413 118 439 228
rect 515 118 541 266
<< pmos >>
rect 141 412 167 612
rect 218 412 244 612
rect 332 412 358 612
rect 502 412 528 636
<< ndiff >>
rect 453 228 515 266
rect 73 189 141 228
rect 73 157 87 189
rect 119 157 141 189
rect 73 118 141 157
rect 167 176 243 228
rect 167 144 189 176
rect 221 144 243 176
rect 167 118 243 144
rect 269 184 413 228
rect 269 152 291 184
rect 323 152 359 184
rect 391 152 413 184
rect 269 118 413 152
rect 439 176 515 228
rect 439 144 461 176
rect 493 144 515 176
rect 439 118 515 144
rect 541 251 609 266
rect 541 219 563 251
rect 595 219 609 251
rect 541 165 609 219
rect 541 133 563 165
rect 595 133 609 165
rect 541 118 609 133
<< pdiff >>
rect 428 612 502 636
rect 73 597 141 612
rect 73 565 87 597
rect 119 565 141 597
rect 73 483 141 565
rect 73 451 87 483
rect 119 451 141 483
rect 73 412 141 451
rect 167 412 218 612
rect 244 412 332 612
rect 358 598 502 612
rect 358 566 380 598
rect 412 566 448 598
rect 480 566 502 598
rect 358 530 502 566
rect 358 498 380 530
rect 412 498 448 530
rect 480 498 502 530
rect 358 412 502 498
rect 528 621 596 636
rect 528 589 550 621
rect 582 589 596 621
rect 528 540 596 589
rect 528 508 550 540
rect 582 508 596 540
rect 528 460 596 508
rect 528 428 550 460
rect 582 428 596 460
rect 528 412 596 428
<< ndiffc >>
rect 87 157 119 189
rect 189 144 221 176
rect 291 152 323 184
rect 359 152 391 184
rect 461 144 493 176
rect 563 219 595 251
rect 563 133 595 165
<< pdiffc >>
rect 87 565 119 597
rect 87 451 119 483
rect 380 566 412 598
rect 448 566 480 598
rect 380 498 412 530
rect 448 498 480 530
rect 550 589 582 621
rect 550 508 582 540
rect 550 428 582 460
<< psubdiff >>
rect 0 16 672 30
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 608 16
rect 640 -16 672 16
rect 0 -30 672 -16
<< nsubdiff >>
rect 0 772 672 786
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 608 772
rect 640 740 672 772
rect 0 726 672 740
<< psubdiffcont >>
rect 32 -16 64 16
rect 128 -16 160 16
rect 224 -16 256 16
rect 320 -16 352 16
rect 416 -16 448 16
rect 512 -16 544 16
rect 608 -16 640 16
<< nsubdiffcont >>
rect 32 740 64 772
rect 128 740 160 772
rect 224 740 256 772
rect 320 740 352 772
rect 416 740 448 772
rect 512 740 544 772
rect 608 740 640 772
<< poly >>
rect 141 612 167 648
rect 218 612 244 648
rect 332 612 358 648
rect 502 636 528 672
rect 141 380 167 412
rect 99 363 167 380
rect 99 331 116 363
rect 148 331 167 363
rect 99 314 167 331
rect 218 380 244 412
rect 332 380 358 412
rect 218 363 284 380
rect 218 331 235 363
rect 267 331 284 363
rect 218 314 284 331
rect 332 363 439 380
rect 502 367 528 412
rect 332 331 365 363
rect 397 331 439 363
rect 332 314 439 331
rect 141 228 167 314
rect 243 228 269 314
rect 413 228 439 314
rect 479 353 541 367
rect 479 321 493 353
rect 525 321 541 353
rect 479 307 541 321
rect 515 266 541 307
rect 141 82 167 118
rect 243 82 269 118
rect 413 82 439 118
rect 515 82 541 118
<< polycont >>
rect 116 331 148 363
rect 235 331 267 363
rect 365 331 397 363
rect 493 321 525 353
<< metal1 >>
rect 0 772 672 800
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 608 772
rect 640 740 672 772
rect 0 712 672 740
rect 77 597 129 599
rect 77 565 87 597
rect 119 565 129 597
rect 77 483 129 565
rect 370 598 490 712
rect 370 566 380 598
rect 412 566 448 598
rect 480 566 490 598
rect 370 530 490 566
rect 370 498 380 530
rect 412 498 448 530
rect 480 498 490 530
rect 370 495 490 498
rect 540 621 610 640
rect 540 589 550 621
rect 582 589 610 621
rect 540 540 610 589
rect 540 508 550 540
rect 582 508 610 540
rect 77 451 87 483
rect 119 459 129 483
rect 540 460 610 508
rect 119 451 503 459
rect 77 424 503 451
rect 59 363 167 387
rect 59 331 116 363
rect 148 331 167 363
rect 59 301 167 331
rect 218 363 312 387
rect 218 331 235 363
rect 267 331 312 363
rect 218 301 312 331
rect 348 363 414 387
rect 348 331 365 363
rect 397 331 414 363
rect 348 301 414 331
rect 469 370 503 424
rect 540 428 550 460
rect 582 428 610 460
rect 540 408 610 428
rect 469 353 542 370
rect 469 321 493 353
rect 525 321 542 353
rect 469 304 542 321
rect 469 265 503 304
rect 77 223 503 265
rect 578 261 610 408
rect 552 251 610 261
rect 77 222 393 223
rect 77 189 129 222
rect 77 157 87 189
rect 119 157 129 189
rect 289 184 393 222
rect 77 153 129 157
rect 179 176 231 178
rect 179 144 189 176
rect 221 144 231 176
rect 179 44 231 144
rect 289 152 291 184
rect 323 152 359 184
rect 391 152 393 184
rect 552 219 563 251
rect 595 219 610 251
rect 289 135 393 152
rect 451 176 503 178
rect 451 144 461 176
rect 493 144 503 176
rect 451 44 503 144
rect 552 165 610 219
rect 552 133 563 165
rect 595 133 610 165
rect 552 121 610 133
rect 0 16 672 44
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 608 16
rect 640 -16 672 16
rect 0 -44 672 -16
<< labels >>
flabel metal1 s 0 712 672 800 0 FreeSans 400 0 0 0 VDD
port 2 nsew
flabel metal1 s 0 -44 672 44 0 FreeSans 400 0 0 0 VSS
port 3 nsew
flabel metal1 s 59 301 167 387 0 FreeSans 400 0 0 0 C
port 4 nsew
flabel metal1 s 218 301 312 387 0 FreeSans 400 0 0 0 B
port 5 nsew
flabel metal1 s 348 301 414 387 0 FreeSans 400 0 0 0 A
port 6 nsew
flabel metal1 s 540 408 610 640 0 FreeSans 400 0 0 0 X
port 7 nsew
<< properties >>
string FIXED_BBOX 0 0 672 756
string GDS_END 128346
string GDS_FILE ../gds/controller.gds
string GDS_START 122822
<< end >>
