magic
tech ihp-sg13g2
magscale 1 2
timestamp 1746816402
<< nwell >>
rect -48 350 432 834
<< pwell >>
rect -3 56 342 281
rect -26 -56 410 56
<< nmos >>
rect 91 195 117 255
rect 221 96 247 255
<< pmos >>
rect 97 429 123 561
rect 222 429 248 660
<< ndiff >>
rect 23 241 91 255
rect 23 209 37 241
rect 69 209 91 241
rect 23 195 91 209
rect 117 195 221 255
rect 137 96 221 195
rect 247 239 316 255
rect 247 207 270 239
rect 302 207 316 239
rect 247 96 316 207
rect 137 36 202 96
<< pdiff >>
rect 23 660 204 720
rect 23 615 222 660
rect 141 561 222 615
rect 23 478 97 561
rect 23 446 37 478
rect 69 446 97 478
rect 23 429 97 446
rect 123 429 222 561
rect 248 563 316 660
rect 248 531 270 563
rect 302 531 316 563
rect 248 475 316 531
rect 248 443 270 475
rect 302 443 316 475
rect 248 429 316 443
<< ndiffc >>
rect 37 209 69 241
rect 270 207 302 239
<< pdiffc >>
rect 37 446 69 478
rect 270 531 302 563
rect 270 443 302 475
<< psubdiff >>
rect 137 30 202 36
rect 0 16 384 30
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 384 16
rect 0 -30 384 -16
<< nsubdiff >>
rect 0 772 384 786
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 384 772
rect 0 726 384 740
rect 23 720 204 726
<< psubdiffcont >>
rect 32 -16 64 16
rect 128 -16 160 16
rect 224 -16 256 16
rect 320 -16 352 16
<< nsubdiffcont >>
rect 32 740 64 772
rect 128 740 160 772
rect 224 740 256 772
rect 320 740 352 772
<< poly >>
rect 222 660 248 698
rect 97 561 123 599
rect 97 413 123 429
rect 91 387 123 413
rect 222 395 248 429
rect 91 331 117 387
rect 222 381 319 395
rect 222 366 273 381
rect 259 349 273 366
rect 305 349 319 381
rect 259 342 319 349
rect 260 341 319 342
rect 261 340 319 341
rect 262 339 319 340
rect 263 338 319 339
rect 264 337 319 338
rect 265 336 319 337
rect 266 335 319 336
rect 23 317 117 331
rect 23 285 37 317
rect 69 285 117 317
rect 23 271 117 285
rect 91 255 117 271
rect 169 328 222 329
rect 169 327 223 328
rect 169 326 224 327
rect 169 325 225 326
rect 169 324 226 325
rect 169 323 227 324
rect 169 322 228 323
rect 169 315 229 322
rect 169 283 183 315
rect 215 298 229 315
rect 215 283 247 298
rect 169 269 247 283
rect 221 255 247 269
rect 91 157 117 195
rect 221 60 247 96
<< polycont >>
rect 273 349 305 381
rect 37 285 69 317
rect 183 283 215 315
<< metal1 >>
rect 0 772 384 800
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 384 772
rect 0 712 384 740
rect 260 563 317 582
rect 260 531 270 563
rect 302 531 317 563
rect 27 478 79 490
rect 27 446 37 478
rect 69 446 79 478
rect 27 438 79 446
rect 39 406 79 438
rect 260 475 317 531
rect 260 443 270 475
rect 302 443 317 475
rect 260 426 317 443
rect 39 363 224 406
rect 27 317 79 327
rect 27 285 37 317
rect 69 285 79 317
rect 27 241 79 285
rect 174 315 224 363
rect 174 283 183 315
rect 215 283 224 315
rect 174 271 224 283
rect 260 381 315 390
rect 260 349 273 381
rect 305 349 315 381
rect 27 209 37 241
rect 69 209 79 241
rect 27 206 79 209
rect 260 239 315 349
rect 260 207 270 239
rect 302 207 315 239
rect 260 197 315 207
rect 0 16 384 44
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 384 16
rect 0 -44 384 -16
<< labels >>
flabel metal1 s 260 426 317 582 0 FreeSans 400 0 0 0 L_HI
port 2 nsew
flabel metal1 s 0 712 384 800 0 FreeSans 400 0 0 0 VDD
port 3 nsew
flabel metal1 s 0 -44 384 44 0 FreeSans 400 0 0 0 VSS
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 384 756
string GDS_END 20344
string GDS_FILE ../gds/controller.gds
string GDS_START 16892
<< end >>
