** sch_path: /home/anton/projects/ttihp0p3-antonalog/xschem/tb_r2r_dac.sch
**.subckt tb_r2r_dac
x1 IN[7] IN[6] IN[5] IN[4] IN[3] IN[2] IN[1] IN[0] net1 GND r2r_dac
V4 IN[3] GND pulse(0 1.2 8u 0 0 8u 16u)
V3 IN[2] GND pulse(0 1.2 4u 0 0 4u 8u)
V2 IN[1] GND pulse(0 1.2 2u 0 0 2u 4u)
V1 IN[0] GND pulse(0 1.2 1u 0 0 1u 2u)
R1 OUT net1 500R m=1
C1 OUT GND 10p m=1
V8 IN[7] GND pulse(0 1.2 128u 0 0 128u 256u)
V7 IN[6] GND pulse(0 1.2 64u 0 0 64u 128u)
V6 IN[5] GND pulse(0 1.2 32u 0 0 32u 64u)
V5 IN[4] GND pulse(0 1.2 16u 0 0 16u 32u)
**** begin user architecture code

.control
tran 10n 256u
write tb_r2r_dac.raw
.endc


.lib /home/anton/asic/IHP-Open-PDK/ihp-sg13g2/libs.tech/ngspice/models/cornerRES.lib res_typ

**** end user architecture code
**.ends

* expanding   symbol:  r2r_dac.sym # of pins=3
** sym_path: /home/anton/projects/ttihp0p3-antonalog/xschem/r2r_dac.sym
** sch_path: /home/anton/projects/ttihp0p3-antonalog/xschem/r2r_dac.sch
.subckt r2r_dac IN[7] IN[6] IN[5] IN[4] IN[3] IN[2] IN[1] IN[0] OUT GND
*.ipin IN[7],IN[6],IN[5],IN[4],IN[3],IN[2],IN[1],IN[0]
*.iopin GND
*.opin OUT
XR0a net1 IN[0] rhigh w=1.0e-6 l=6.0e-6 m=1 b=0
XR0b net3 net1 rhigh w=1.0e-6 l=6.0e-6 m=1 b=0
XR1c net3 net4 rhigh w=1.0e-6 l=6.0e-6 m=1 b=0
XR0c net2 net3 rhigh w=1.0e-6 l=6.0e-6 m=1 b=0
XR0d GND net2 rhigh w=1.0e-6 l=6.0e-6 m=1 b=0
XR1a net5 IN[1] rhigh w=1.0e-6 l=6.0e-6 m=1 b=0
XR1b net4 net5 rhigh w=1.0e-6 l=6.0e-6 m=1 b=0
XR2c net4 net6 rhigh w=1.0e-6 l=6.0e-6 m=1 b=0
XR2a net7 IN[2] rhigh w=1.0e-6 l=6.0e-6 m=1 b=0
XR2b net6 net7 rhigh w=1.0e-6 l=6.0e-6 m=1 b=0
XR3c net6 net8 rhigh w=1.0e-6 l=6.0e-6 m=1 b=0
XR3a net9 IN[3] rhigh w=1.0e-6 l=6.0e-6 m=1 b=0
XR3b net8 net9 rhigh w=1.0e-6 l=6.0e-6 m=1 b=0
XR4c net8 net10 rhigh w=1.0e-6 l=6.0e-6 m=1 b=0
XR4a net11 IN[4] rhigh w=1.0e-6 l=6.0e-6 m=1 b=0
XR4b net10 net11 rhigh w=1.0e-6 l=6.0e-6 m=1 b=0
XR5c net10 net12 rhigh w=1.0e-6 l=6.0e-6 m=1 b=0
XR5a net13 IN[5] rhigh w=1.0e-6 l=6.0e-6 m=1 b=0
XR5b net12 net13 rhigh w=1.0e-6 l=6.0e-6 m=1 b=0
XR6c net12 net14 rhigh w=1.0e-6 l=6.0e-6 m=1 b=0
XR6a net15 IN[6] rhigh w=1.0e-6 l=6.0e-6 m=1 b=0
XR6b net14 net15 rhigh w=1.0e-6 l=6.0e-6 m=1 b=0
XR7c net14 OUT rhigh w=1.0e-6 l=6.0e-6 m=1 b=0
XR7a net16 IN[7] rhigh w=1.0e-6 l=6.0e-6 m=1 b=0
XR7b OUT net16 rhigh w=1.0e-6 l=6.0e-6 m=1 b=0
.ends

.end
