magic
tech ihp-sg13g2
magscale 1 2
timestamp 1746816402
<< nwell >>
rect -48 350 816 834
<< pwell >>
rect 46 56 709 292
rect -26 -56 794 56
<< nmos >>
rect 140 156 166 266
rect 242 156 268 266
rect 385 156 411 266
rect 487 156 513 266
rect 589 118 615 266
<< pmos >>
rect 148 436 174 636
rect 234 436 260 636
rect 348 436 374 636
rect 462 436 488 636
rect 593 412 619 636
<< ndiff >>
rect 72 227 140 266
rect 72 195 86 227
rect 118 195 140 227
rect 72 156 140 195
rect 166 213 242 266
rect 166 181 188 213
rect 220 181 242 213
rect 166 156 242 181
rect 268 197 385 266
rect 268 165 301 197
rect 333 165 385 197
rect 268 156 385 165
rect 411 213 487 266
rect 411 181 433 213
rect 465 181 487 213
rect 411 156 487 181
rect 513 200 589 266
rect 513 168 535 200
rect 567 168 589 200
rect 513 156 589 168
rect 282 150 371 156
rect 527 118 589 156
rect 615 249 683 266
rect 615 217 637 249
rect 669 217 683 249
rect 615 166 683 217
rect 615 134 637 166
rect 669 134 683 166
rect 615 118 683 134
<< pdiff >>
rect 80 621 148 636
rect 80 589 94 621
rect 126 589 148 621
rect 80 553 148 589
rect 80 521 94 553
rect 126 521 148 553
rect 80 483 148 521
rect 80 451 94 483
rect 126 451 148 483
rect 80 436 148 451
rect 174 436 234 636
rect 260 436 348 636
rect 374 436 462 636
rect 488 619 593 636
rect 488 587 510 619
rect 542 587 593 619
rect 488 551 593 587
rect 488 519 510 551
rect 542 519 593 551
rect 488 436 593 519
rect 545 412 593 436
rect 619 619 687 636
rect 619 587 641 619
rect 673 587 687 619
rect 619 540 687 587
rect 619 508 641 540
rect 673 508 687 540
rect 619 461 687 508
rect 619 429 641 461
rect 673 429 687 461
rect 619 412 687 429
<< ndiffc >>
rect 86 195 118 227
rect 188 181 220 213
rect 301 165 333 197
rect 433 181 465 213
rect 535 168 567 200
rect 637 217 669 249
rect 637 134 669 166
<< pdiffc >>
rect 94 589 126 621
rect 94 521 126 553
rect 94 451 126 483
rect 510 587 542 619
rect 510 519 542 551
rect 641 587 673 619
rect 641 508 673 540
rect 641 429 673 461
<< psubdiff >>
rect 0 16 768 30
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 608 16
rect 640 -16 704 16
rect 736 -16 768 16
rect 0 -30 768 -16
<< nsubdiff >>
rect 0 772 768 786
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 608 772
rect 640 740 704 772
rect 736 740 768 772
rect 0 726 768 740
<< psubdiffcont >>
rect 32 -16 64 16
rect 128 -16 160 16
rect 224 -16 256 16
rect 320 -16 352 16
rect 416 -16 448 16
rect 512 -16 544 16
rect 608 -16 640 16
rect 704 -16 736 16
<< nsubdiffcont >>
rect 32 740 64 772
rect 128 740 160 772
rect 224 740 256 772
rect 320 740 352 772
rect 416 740 448 772
rect 512 740 544 772
rect 608 740 640 772
rect 704 740 736 772
<< poly >>
rect 148 636 174 672
rect 234 636 260 672
rect 348 636 374 672
rect 462 636 488 672
rect 593 636 619 672
rect 148 394 174 436
rect 234 394 260 436
rect 348 394 374 436
rect 109 377 175 394
rect 109 345 126 377
rect 158 345 175 377
rect 109 328 175 345
rect 229 377 295 394
rect 229 345 246 377
rect 278 345 295 377
rect 229 328 295 345
rect 343 377 409 394
rect 462 380 488 436
rect 343 345 360 377
rect 392 345 409 377
rect 343 328 409 345
rect 457 363 524 380
rect 593 370 619 412
rect 457 331 474 363
rect 506 331 524 363
rect 140 266 166 328
rect 242 266 268 328
rect 343 306 411 328
rect 457 314 524 331
rect 566 353 632 370
rect 566 321 583 353
rect 615 321 632 353
rect 385 266 411 306
rect 487 266 513 314
rect 566 304 632 321
rect 589 266 615 304
rect 140 120 166 156
rect 242 120 268 156
rect 385 120 411 156
rect 487 120 513 156
rect 589 82 615 118
<< polycont >>
rect 126 345 158 377
rect 246 345 278 377
rect 360 345 392 377
rect 474 331 506 363
rect 583 321 615 353
<< metal1 >>
rect 0 772 768 800
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 608 772
rect 640 740 704 772
rect 736 740 768 772
rect 0 712 768 740
rect 84 621 136 624
rect 84 589 94 621
rect 126 589 136 621
rect 84 553 136 589
rect 84 521 94 553
rect 126 521 136 553
rect 84 483 136 521
rect 500 619 552 712
rect 500 587 510 619
rect 542 587 552 619
rect 500 551 552 587
rect 500 519 510 551
rect 542 519 552 551
rect 500 517 552 519
rect 631 619 700 621
rect 631 587 641 619
rect 673 587 700 619
rect 631 540 700 587
rect 84 451 94 483
rect 126 476 136 483
rect 631 508 641 540
rect 673 508 700 540
rect 126 451 591 476
rect 84 438 591 451
rect 53 377 175 387
rect 53 345 126 377
rect 158 345 175 377
rect 53 309 175 345
rect 229 377 304 394
rect 229 345 246 377
rect 278 345 304 377
rect 229 309 304 345
rect 343 377 409 394
rect 343 345 360 377
rect 392 345 409 377
rect 343 309 409 345
rect 454 363 521 395
rect 454 331 474 363
rect 506 331 521 363
rect 454 309 521 331
rect 557 370 591 438
rect 631 461 700 508
rect 631 429 641 461
rect 673 429 700 461
rect 631 408 700 429
rect 557 353 632 370
rect 557 321 583 353
rect 615 321 632 353
rect 557 304 632 321
rect 557 273 599 304
rect 184 239 599 273
rect 668 259 700 408
rect 636 249 700 259
rect 76 227 128 229
rect 76 195 86 227
rect 118 195 128 227
rect 76 44 128 195
rect 184 213 224 239
rect 184 181 188 213
rect 220 181 224 213
rect 429 213 469 239
rect 184 171 224 181
rect 291 197 343 200
rect 291 165 301 197
rect 333 165 343 197
rect 429 181 433 213
rect 465 181 469 213
rect 636 217 637 249
rect 669 217 700 249
rect 429 171 469 181
rect 525 200 577 202
rect 291 44 343 165
rect 525 168 535 200
rect 567 168 577 200
rect 525 44 577 168
rect 636 166 700 217
rect 636 134 637 166
rect 669 134 700 166
rect 636 124 700 134
rect 0 16 768 44
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 608 16
rect 640 -16 704 16
rect 736 -16 768 16
rect 0 -44 768 -16
<< labels >>
flabel metal1 s 631 408 700 621 0 FreeSans 400 0 0 0 X
port 2 nsew
flabel metal1 s 229 309 304 394 0 FreeSans 400 0 0 0 C
port 3 nsew
flabel metal1 s 53 309 175 387 0 FreeSans 400 0 0 0 D
port 4 nsew
flabel metal1 s 0 712 768 800 0 FreeSans 400 0 0 0 VDD
port 5 nsew
flabel metal1 s 0 -44 768 44 0 FreeSans 400 0 0 0 VSS
port 6 nsew
flabel metal1 s 454 309 521 395 0 FreeSans 400 0 0 0 A
port 7 nsew
flabel metal1 s 343 309 409 394 0 FreeSans 400 0 0 0 B
port 8 nsew
<< properties >>
string FIXED_BBOX 0 0 768 756
string GDS_END 225682
string GDS_FILE ../gds/controller.gds
string GDS_START 219360
<< end >>
