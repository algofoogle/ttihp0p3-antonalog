magic
tech ihp-sg13g2
timestamp 1747537721
<< nwell >>
rect -24 175 408 417
<< pwell >>
rect 23 28 354 146
rect -13 -28 397 28
<< nmos >>
rect 70 78 83 133
rect 121 78 134 133
rect 192 78 205 133
rect 243 78 256 133
rect 294 59 307 133
<< pmos >>
rect 74 218 87 318
rect 117 218 130 318
rect 174 218 187 318
rect 231 218 244 318
rect 296 206 309 318
<< ndiff >>
rect 36 113 70 133
rect 36 97 43 113
rect 59 97 70 113
rect 36 78 70 97
rect 83 106 121 133
rect 83 90 94 106
rect 110 90 121 106
rect 83 78 121 90
rect 134 98 192 133
rect 134 82 150 98
rect 166 82 192 98
rect 134 78 192 82
rect 205 106 243 133
rect 205 90 216 106
rect 232 90 243 106
rect 205 78 243 90
rect 256 100 294 133
rect 256 84 267 100
rect 283 84 294 100
rect 256 78 294 84
rect 141 75 185 78
rect 263 59 294 78
rect 307 124 341 133
rect 307 108 318 124
rect 334 108 341 124
rect 307 83 341 108
rect 307 67 318 83
rect 334 67 341 83
rect 307 59 341 67
<< pdiff >>
rect 40 310 74 318
rect 40 294 47 310
rect 63 294 74 310
rect 40 276 74 294
rect 40 260 47 276
rect 63 260 74 276
rect 40 241 74 260
rect 40 225 47 241
rect 63 225 74 241
rect 40 218 74 225
rect 87 218 117 318
rect 130 218 174 318
rect 187 218 231 318
rect 244 309 296 318
rect 244 293 255 309
rect 271 293 296 309
rect 244 275 296 293
rect 244 259 255 275
rect 271 259 296 275
rect 244 218 296 259
rect 272 206 296 218
rect 309 309 343 318
rect 309 293 320 309
rect 336 293 343 309
rect 309 270 343 293
rect 309 254 320 270
rect 336 254 343 270
rect 309 230 343 254
rect 309 214 320 230
rect 336 214 343 230
rect 309 206 343 214
<< ndiffc >>
rect 43 97 59 113
rect 94 90 110 106
rect 150 82 166 98
rect 216 90 232 106
rect 267 84 283 100
rect 318 108 334 124
rect 318 67 334 83
<< pdiffc >>
rect 47 294 63 310
rect 47 260 63 276
rect 47 225 63 241
rect 255 293 271 309
rect 255 259 271 275
rect 320 293 336 309
rect 320 254 336 270
rect 320 214 336 230
<< psubdiff >>
rect 0 8 384 15
rect 0 -8 16 8
rect 32 -8 64 8
rect 80 -8 112 8
rect 128 -8 160 8
rect 176 -8 208 8
rect 224 -8 256 8
rect 272 -8 304 8
rect 320 -8 352 8
rect 368 -8 384 8
rect 0 -15 384 -8
<< nsubdiff >>
rect 0 386 384 393
rect 0 370 16 386
rect 32 370 64 386
rect 80 370 112 386
rect 128 370 160 386
rect 176 370 208 386
rect 224 370 256 386
rect 272 370 304 386
rect 320 370 352 386
rect 368 370 384 386
rect 0 363 384 370
<< psubdiffcont >>
rect 16 -8 32 8
rect 64 -8 80 8
rect 112 -8 128 8
rect 160 -8 176 8
rect 208 -8 224 8
rect 256 -8 272 8
rect 304 -8 320 8
rect 352 -8 368 8
<< nsubdiffcont >>
rect 16 370 32 386
rect 64 370 80 386
rect 112 370 128 386
rect 160 370 176 386
rect 208 370 224 386
rect 256 370 272 386
rect 304 370 320 386
rect 352 370 368 386
<< poly >>
rect 74 318 87 336
rect 117 318 130 336
rect 174 318 187 336
rect 231 318 244 336
rect 296 318 309 336
rect 74 197 87 218
rect 117 197 130 218
rect 174 197 187 218
rect 54 188 87 197
rect 54 172 63 188
rect 79 172 87 188
rect 54 164 87 172
rect 114 188 147 197
rect 114 172 123 188
rect 139 172 147 188
rect 114 164 147 172
rect 171 188 204 197
rect 231 190 244 218
rect 171 172 180 188
rect 196 172 204 188
rect 171 164 204 172
rect 228 181 262 190
rect 296 185 309 206
rect 228 165 237 181
rect 253 165 262 181
rect 70 133 83 164
rect 121 133 134 164
rect 171 153 205 164
rect 228 157 262 165
rect 283 176 316 185
rect 283 160 291 176
rect 307 160 316 176
rect 192 133 205 153
rect 243 133 256 157
rect 283 152 316 160
rect 294 133 307 152
rect 70 60 83 78
rect 121 60 134 78
rect 192 60 205 78
rect 243 60 256 78
rect 294 41 307 59
<< polycont >>
rect 63 172 79 188
rect 123 172 139 188
rect 180 172 196 188
rect 237 165 253 181
rect 291 160 307 176
<< metal1 >>
rect 0 386 384 400
rect 0 370 16 386
rect 32 370 64 386
rect 80 370 112 386
rect 128 370 160 386
rect 176 370 208 386
rect 224 370 256 386
rect 272 370 304 386
rect 320 370 352 386
rect 368 370 384 386
rect 0 356 384 370
rect 42 310 68 312
rect 42 294 47 310
rect 63 294 68 310
rect 42 276 68 294
rect 42 260 47 276
rect 63 260 68 276
rect 42 241 68 260
rect 250 309 276 356
rect 250 293 255 309
rect 271 293 276 309
rect 250 275 276 293
rect 250 259 255 275
rect 271 259 276 275
rect 250 258 276 259
rect 315 309 350 310
rect 315 293 320 309
rect 336 293 350 309
rect 315 270 350 293
rect 42 225 47 241
rect 63 238 68 241
rect 315 254 320 270
rect 336 254 350 270
rect 63 225 295 238
rect 42 219 295 225
rect 26 188 87 193
rect 26 172 63 188
rect 79 172 87 188
rect 26 154 87 172
rect 114 188 152 197
rect 114 172 123 188
rect 139 172 152 188
rect 114 154 152 172
rect 171 188 204 197
rect 171 172 180 188
rect 196 172 204 188
rect 171 154 204 172
rect 227 181 260 197
rect 227 165 237 181
rect 253 165 260 181
rect 227 154 260 165
rect 278 185 295 219
rect 315 230 350 254
rect 315 214 320 230
rect 336 214 350 230
rect 315 204 350 214
rect 278 176 316 185
rect 278 160 291 176
rect 307 160 316 176
rect 278 152 316 160
rect 278 136 299 152
rect 92 119 299 136
rect 334 129 350 204
rect 318 124 350 129
rect 38 113 64 114
rect 38 97 43 113
rect 59 97 64 113
rect 38 22 64 97
rect 92 106 112 119
rect 92 90 94 106
rect 110 90 112 106
rect 214 106 234 119
rect 92 85 112 90
rect 145 98 171 100
rect 145 82 150 98
rect 166 82 171 98
rect 214 90 216 106
rect 232 90 234 106
rect 334 108 350 124
rect 214 85 234 90
rect 262 100 288 101
rect 145 22 171 82
rect 262 84 267 100
rect 283 84 288 100
rect 262 22 288 84
rect 318 83 350 108
rect 334 67 350 83
rect 318 62 350 67
rect 0 8 384 22
rect 0 -8 16 8
rect 32 -8 64 8
rect 80 -8 112 8
rect 128 -8 160 8
rect 176 -8 208 8
rect 224 -8 256 8
rect 272 -8 304 8
rect 320 -8 352 8
rect 368 -8 384 8
rect 0 -22 384 -8
<< labels >>
flabel metal1 s 315 204 350 310 0 FreeSans 200 0 0 0 X
port 2 nsew
flabel metal1 s 114 154 152 197 0 FreeSans 200 0 0 0 C
port 3 nsew
flabel metal1 s 26 154 87 193 0 FreeSans 200 0 0 0 D
port 4 nsew
flabel metal1 s 0 356 384 400 0 FreeSans 200 0 0 0 VDD
port 5 nsew
flabel metal1 s 0 -22 384 22 0 FreeSans 200 0 0 0 VSS
port 6 nsew
flabel metal1 s 227 154 260 197 0 FreeSans 200 0 0 0 A
port 7 nsew
flabel metal1 s 171 154 204 197 0 FreeSans 200 0 0 0 B
port 8 nsew
<< properties >>
string FIXED_BBOX 0 0 384 378
string GDS_END 251330
string GDS_FILE ../gds/controller.gds
string GDS_START 245008
<< end >>
