magic
tech ihp-sg13g2
timestamp 1747537721
<< nwell >>
rect -24 175 264 417
<< pwell >>
rect 8 28 232 148
rect -13 -28 253 28
<< nmos >>
rect 60 61 73 135
rect 119 61 132 135
rect 162 61 175 135
<< pmos >>
rect 60 213 73 325
rect 111 213 124 325
rect 162 213 175 325
<< ndiff >>
rect 21 91 60 135
rect 21 75 28 91
rect 44 75 60 91
rect 21 61 60 75
rect 73 61 119 135
rect 132 61 162 135
rect 175 126 219 135
rect 175 110 192 126
rect 208 110 219 126
rect 175 85 219 110
rect 175 69 186 85
rect 202 69 219 85
rect 175 61 219 69
<< pdiff >>
rect 26 317 60 325
rect 26 301 33 317
rect 49 301 60 317
rect 26 282 60 301
rect 26 266 33 282
rect 49 266 60 282
rect 26 240 60 266
rect 26 224 33 240
rect 49 224 60 240
rect 26 213 60 224
rect 73 317 111 325
rect 73 301 84 317
rect 100 301 111 317
rect 73 283 111 301
rect 73 267 84 283
rect 100 267 111 283
rect 73 248 111 267
rect 73 232 84 248
rect 100 232 111 248
rect 73 213 111 232
rect 124 317 162 325
rect 124 301 135 317
rect 151 301 162 317
rect 124 282 162 301
rect 124 266 135 282
rect 151 266 162 282
rect 124 213 162 266
rect 175 317 209 325
rect 175 301 186 317
rect 202 301 209 317
rect 175 277 209 301
rect 175 261 186 277
rect 202 261 209 277
rect 175 237 209 261
rect 175 221 186 237
rect 202 221 209 237
rect 175 213 209 221
<< ndiffc >>
rect 28 75 44 91
rect 192 110 208 126
rect 186 69 202 85
<< pdiffc >>
rect 33 301 49 317
rect 33 266 49 282
rect 33 224 49 240
rect 84 301 100 317
rect 84 267 100 283
rect 84 232 100 248
rect 135 301 151 317
rect 135 266 151 282
rect 186 301 202 317
rect 186 261 202 277
rect 186 221 202 237
<< psubdiff >>
rect 0 8 240 15
rect 0 -8 16 8
rect 32 -8 64 8
rect 80 -8 112 8
rect 128 -8 160 8
rect 176 -8 208 8
rect 224 -8 240 8
rect 0 -15 240 -8
<< nsubdiff >>
rect 0 386 240 393
rect 0 370 16 386
rect 32 370 64 386
rect 80 370 112 386
rect 128 370 160 386
rect 176 370 208 386
rect 224 370 240 386
rect 0 363 240 370
<< psubdiffcont >>
rect 16 -8 32 8
rect 64 -8 80 8
rect 112 -8 128 8
rect 160 -8 176 8
rect 208 -8 224 8
<< nsubdiffcont >>
rect 16 370 32 386
rect 64 370 80 386
rect 112 370 128 386
rect 160 370 176 386
rect 208 370 224 386
<< poly >>
rect 60 325 73 343
rect 111 325 124 343
rect 162 325 175 343
rect 60 187 73 213
rect 111 190 124 213
rect 36 180 73 187
rect 36 164 43 180
rect 59 164 73 180
rect 36 157 73 164
rect 102 181 132 190
rect 162 185 175 213
rect 102 165 109 181
rect 125 165 132 181
rect 102 158 132 165
rect 60 135 73 157
rect 119 135 132 158
rect 150 178 187 185
rect 150 162 160 178
rect 176 162 187 178
rect 150 155 187 162
rect 162 135 175 155
rect 60 43 73 61
rect 119 43 132 61
rect 162 43 175 61
<< polycont >>
rect 43 164 59 180
rect 109 165 125 181
rect 160 162 176 178
<< metal1 >>
rect 0 386 240 400
rect 0 370 16 386
rect 32 370 64 386
rect 80 370 112 386
rect 128 370 160 386
rect 176 370 208 386
rect 224 370 240 386
rect 0 356 240 370
rect 28 317 54 356
rect 28 301 33 317
rect 49 301 54 317
rect 28 282 54 301
rect 28 266 33 282
rect 49 266 54 282
rect 28 240 54 266
rect 28 224 33 240
rect 49 224 54 240
rect 28 217 54 224
rect 79 317 105 320
rect 79 301 84 317
rect 100 301 105 317
rect 79 283 105 301
rect 79 267 84 283
rect 100 267 105 283
rect 79 248 105 267
rect 130 317 156 356
rect 130 301 135 317
rect 151 301 156 317
rect 130 282 156 301
rect 130 266 135 282
rect 151 266 156 282
rect 130 257 156 266
rect 178 317 226 327
rect 178 301 186 317
rect 202 301 226 317
rect 178 277 226 301
rect 178 261 186 277
rect 202 261 226 277
rect 79 232 84 248
rect 100 239 105 248
rect 178 239 226 261
rect 100 237 226 239
rect 100 232 186 237
rect 79 221 186 232
rect 202 221 226 237
rect 79 218 226 221
rect 178 217 226 218
rect 36 180 69 198
rect 36 164 43 180
rect 59 164 69 180
rect 36 157 69 164
rect 95 181 132 200
rect 95 165 109 181
rect 125 165 132 181
rect 95 157 132 165
rect 153 178 187 199
rect 153 162 160 178
rect 176 162 187 178
rect 153 155 187 162
rect 205 136 226 217
rect 187 126 226 136
rect 187 110 192 126
rect 208 110 226 126
rect 187 101 226 110
rect 22 91 49 96
rect 22 75 28 91
rect 44 75 49 91
rect 22 22 49 75
rect 177 85 226 101
rect 177 69 186 85
rect 202 69 226 85
rect 177 62 226 69
rect 0 8 240 22
rect 0 -8 16 8
rect 32 -8 64 8
rect 80 -8 112 8
rect 128 -8 160 8
rect 176 -8 208 8
rect 224 -8 240 8
rect 0 -22 240 -8
<< labels >>
flabel metal1 s 0 356 240 400 0 FreeSans 200 0 0 0 VDD
port 2 nsew
flabel metal1 s 178 217 226 327 0 FreeSans 200 0 0 0 Y
port 3 nsew
flabel metal1 s 95 157 132 200 0 FreeSans 200 0 0 0 B
port 4 nsew
flabel metal1 s 36 157 69 198 0 FreeSans 200 0 0 0 C
port 5 nsew
flabel metal1 s 0 -22 240 22 0 FreeSans 200 0 0 0 VSS
port 6 nsew
flabel metal1 s 153 155 187 199 0 FreeSans 200 0 0 0 A
port 7 nsew
<< properties >>
string FIXED_BBOX 0 0 240 378
string GDS_END 122778
string GDS_FILE ../gds/controller.gds
string GDS_START 118150
<< end >>
