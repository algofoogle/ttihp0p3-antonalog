magic
tech ihp-sg13g2
magscale 1 2
timestamp 1747056038
<< nwell >>
rect -48 350 432 834
<< pwell >>
rect 27 56 344 292
rect -26 -56 410 56
<< nmos >>
rect 121 118 147 266
rect 223 118 249 266
<< pmos >>
rect 119 412 145 636
rect 222 412 248 636
<< ndiff >>
rect 53 250 121 266
rect 53 218 67 250
rect 99 218 121 250
rect 53 167 121 218
rect 53 135 67 167
rect 99 135 121 167
rect 53 118 121 135
rect 147 250 223 266
rect 147 218 169 250
rect 201 218 223 250
rect 147 167 223 218
rect 147 135 169 167
rect 201 135 223 167
rect 147 118 223 135
rect 249 250 318 266
rect 249 218 272 250
rect 304 218 318 250
rect 249 167 318 218
rect 249 135 272 167
rect 304 135 318 167
rect 249 118 318 135
<< pdiff >>
rect 51 619 119 636
rect 51 587 65 619
rect 97 587 119 619
rect 51 550 119 587
rect 51 518 65 550
rect 97 518 119 550
rect 51 479 119 518
rect 51 447 65 479
rect 97 447 119 479
rect 51 412 119 447
rect 145 619 222 636
rect 145 587 168 619
rect 200 587 222 619
rect 145 540 222 587
rect 145 508 168 540
rect 200 508 222 540
rect 145 461 222 508
rect 145 429 168 461
rect 200 429 222 461
rect 145 412 222 429
rect 248 619 316 636
rect 248 587 270 619
rect 302 587 316 619
rect 248 540 316 587
rect 248 508 270 540
rect 302 508 316 540
rect 248 461 316 508
rect 248 429 270 461
rect 302 429 316 461
rect 248 412 316 429
<< ndiffc >>
rect 67 218 99 250
rect 67 135 99 167
rect 169 218 201 250
rect 169 135 201 167
rect 272 218 304 250
rect 272 135 304 167
<< pdiffc >>
rect 65 587 97 619
rect 65 518 97 550
rect 65 447 97 479
rect 168 587 200 619
rect 168 508 200 540
rect 168 429 200 461
rect 270 587 302 619
rect 270 508 302 540
rect 270 429 302 461
<< psubdiff >>
rect 0 16 384 30
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 384 16
rect 0 -30 384 -16
<< nsubdiff >>
rect 0 772 384 786
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 384 772
rect 0 726 384 740
<< psubdiffcont >>
rect 32 -16 64 16
rect 128 -16 160 16
rect 224 -16 256 16
rect 320 -16 352 16
<< nsubdiffcont >>
rect 32 740 64 772
rect 128 740 160 772
rect 224 740 256 772
rect 320 740 352 772
<< poly >>
rect 119 636 145 672
rect 222 636 248 672
rect 119 397 145 412
rect 222 397 248 412
rect 119 370 157 397
rect 61 353 157 370
rect 61 321 78 353
rect 110 334 157 353
rect 211 334 248 397
rect 110 321 248 334
rect 61 317 248 321
rect 61 304 249 317
rect 121 266 147 304
rect 223 266 249 304
rect 121 82 147 118
rect 223 82 249 118
<< polycont >>
rect 78 321 110 353
<< metal1 >>
rect 0 772 384 800
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 384 772
rect 0 712 384 740
rect 55 619 107 712
rect 55 587 65 619
rect 97 587 107 619
rect 55 550 107 587
rect 55 518 65 550
rect 97 518 107 550
rect 55 479 107 518
rect 55 447 65 479
rect 97 447 107 479
rect 55 437 107 447
rect 165 619 204 636
rect 165 587 168 619
rect 200 587 204 619
rect 165 540 204 587
rect 165 508 168 540
rect 200 508 204 540
rect 165 461 204 508
rect 165 429 168 461
rect 200 429 204 461
rect 36 353 127 400
rect 36 321 78 353
rect 110 321 127 353
rect 36 304 127 321
rect 57 250 109 260
rect 57 218 67 250
rect 99 218 109 250
rect 57 167 109 218
rect 57 135 67 167
rect 99 135 109 167
rect 57 44 109 135
rect 165 250 204 429
rect 264 619 307 712
rect 264 587 270 619
rect 302 587 307 619
rect 264 540 307 587
rect 264 508 270 540
rect 302 508 307 540
rect 264 461 307 508
rect 264 429 270 461
rect 302 429 307 461
rect 264 419 307 429
rect 165 218 169 250
rect 201 218 204 250
rect 165 167 204 218
rect 165 135 169 167
rect 201 135 204 167
rect 165 114 204 135
rect 268 250 308 261
rect 268 218 272 250
rect 304 218 308 250
rect 268 167 308 218
rect 268 135 272 167
rect 304 135 308 167
rect 268 44 308 135
rect 0 16 384 44
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 384 16
rect 0 -44 384 -16
<< labels >>
flabel metal1 s 0 -44 384 44 0 FreeSans 400 0 0 0 VSS
port 2 nsew
flabel metal1 s 0 712 384 800 0 FreeSans 400 0 0 0 VDD
port 3 nsew
flabel metal1 s 165 114 204 636 0 FreeSans 400 0 0 0 Y
port 4 nsew
flabel metal1 s 36 304 127 400 0 FreeSans 400 0 0 0 A
port 5 nsew
<< properties >>
string FIXED_BBOX 0 0 384 756
string GDS_END 26516
string GDS_FILE ../gds/controller.gds
string GDS_START 22828
<< end >>
