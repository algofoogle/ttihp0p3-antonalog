magic
tech ihp-sg13g2
magscale 1 2
timestamp 1747056038
<< nwell >>
rect -48 350 432 834
<< pwell >>
rect -2 56 386 239
rect -26 -56 410 56
<< nmos >>
rect 92 129 292 213
<< pmos >>
rect 92 436 292 636
<< ndiff >>
rect 24 176 92 213
rect 24 144 38 176
rect 70 144 92 176
rect 24 129 92 144
rect 292 176 360 213
rect 292 144 314 176
rect 346 144 360 176
rect 292 129 360 144
<< pdiff >>
rect 24 621 92 636
rect 24 589 38 621
rect 70 589 92 621
rect 24 551 92 589
rect 24 519 38 551
rect 70 519 92 551
rect 24 436 92 519
rect 292 621 360 636
rect 292 589 314 621
rect 346 589 360 621
rect 292 551 360 589
rect 292 519 314 551
rect 346 519 360 551
rect 292 436 360 519
<< ndiffc >>
rect 38 144 70 176
rect 314 144 346 176
<< pdiffc >>
rect 38 589 70 621
rect 38 519 70 551
rect 314 589 346 621
rect 314 519 346 551
<< psubdiff >>
rect 0 16 384 30
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 384 16
rect 0 -30 384 -16
<< nsubdiff >>
rect 0 772 384 786
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 384 772
rect 0 726 384 740
<< psubdiffcont >>
rect 32 -16 64 16
rect 128 -16 160 16
rect 224 -16 256 16
rect 320 -16 352 16
<< nsubdiffcont >>
rect 32 740 64 772
rect 128 740 160 772
rect 224 740 256 772
rect 320 740 352 772
<< poly >>
rect 92 636 292 672
rect 92 400 292 436
rect 92 344 171 400
rect 92 312 122 344
rect 154 312 171 344
rect 92 295 171 312
rect 213 343 292 360
rect 213 311 230 343
rect 262 311 292 343
rect 213 249 292 311
rect 92 213 292 249
rect 92 93 292 129
<< polycont >>
rect 122 312 154 344
rect 230 311 262 343
<< metal1 >>
rect 0 772 384 800
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 384 772
rect 0 712 384 740
rect 26 621 80 712
rect 26 589 38 621
rect 70 589 80 621
rect 26 551 80 589
rect 26 519 38 551
rect 70 519 80 551
rect 26 507 80 519
rect 213 621 358 712
rect 213 589 314 621
rect 346 589 358 621
rect 213 551 358 589
rect 213 519 314 551
rect 346 519 358 551
rect 213 508 358 519
rect 106 344 171 361
rect 106 312 122 344
rect 154 312 171 344
rect 106 187 171 312
rect 213 343 281 508
rect 213 311 230 343
rect 262 311 281 343
rect 213 294 281 311
rect 26 176 171 187
rect 26 144 38 176
rect 70 144 171 176
rect 26 44 171 144
rect 302 176 358 187
rect 302 144 314 176
rect 346 144 358 176
rect 302 44 358 144
rect 0 16 384 44
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 384 16
rect 0 -44 384 -16
<< labels >>
flabel metal1 s 0 712 384 800 0 FreeSans 400 0 0 0 VDD
port 1 nsew
flabel metal1 s 0 -44 384 44 0 FreeSans 400 0 0 0 VSS
port 2 nsew
<< properties >>
string FIXED_BBOX 0 0 384 756
string GDS_END 5784
string GDS_FILE ../gds/controller.gds
string GDS_START 3516
<< end >>
