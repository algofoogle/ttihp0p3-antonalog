magic
tech ihp-sg13g2
magscale 1 2
timestamp 1746816402
<< nwell >>
rect -48 350 2064 834
rect 148 323 912 350
<< pwell >>
rect 1276 302 1573 314
rect 1276 272 1999 302
rect 45 56 1999 272
rect -26 -56 2042 56
<< nmos >>
rect 139 118 165 246
rect 282 118 308 246
rect 356 118 382 246
rect 474 118 500 246
rect 644 118 670 246
rect 784 118 810 246
rect 860 118 886 246
rect 997 118 1023 246
rect 1071 118 1097 246
rect 1351 160 1377 288
rect 1453 160 1479 288
rect 1765 148 1791 276
rect 1879 128 1905 276
<< pmos >>
rect 159 412 185 612
rect 269 385 295 585
rect 461 385 487 585
rect 563 385 589 585
rect 653 385 679 585
rect 779 385 805 585
rect 880 431 906 631
rect 1083 431 1109 631
rect 1163 431 1189 631
rect 1367 436 1393 636
rect 1482 436 1508 636
rect 1726 431 1752 631
rect 1883 412 1909 636
<< ndiff >>
rect 71 232 139 246
rect 71 200 85 232
rect 117 200 139 232
rect 71 164 139 200
rect 71 132 85 164
rect 117 132 139 164
rect 71 118 139 132
rect 165 164 282 246
rect 165 132 207 164
rect 239 132 282 164
rect 165 118 282 132
rect 308 118 356 246
rect 382 222 474 246
rect 382 190 420 222
rect 452 190 474 222
rect 382 118 474 190
rect 500 118 644 246
rect 670 164 784 246
rect 670 132 712 164
rect 744 132 784 164
rect 670 118 784 132
rect 810 118 860 246
rect 886 164 997 246
rect 886 132 925 164
rect 957 132 997 164
rect 886 118 997 132
rect 1023 118 1071 246
rect 1097 182 1165 246
rect 1302 229 1351 288
rect 1097 150 1119 182
rect 1151 150 1165 182
rect 1097 118 1165 150
rect 1219 215 1351 229
rect 1219 183 1233 215
rect 1265 183 1351 215
rect 1219 160 1351 183
rect 1377 274 1453 288
rect 1377 242 1399 274
rect 1431 242 1453 274
rect 1377 160 1453 242
rect 1479 206 1547 288
rect 1479 174 1501 206
rect 1533 174 1547 206
rect 1479 160 1547 174
rect 1693 262 1765 276
rect 1693 230 1707 262
rect 1739 230 1765 262
rect 1693 194 1765 230
rect 1693 162 1707 194
rect 1739 162 1765 194
rect 1219 124 1337 160
rect 1219 92 1233 124
rect 1265 92 1337 124
rect 1219 78 1337 92
rect 1693 148 1765 162
rect 1791 262 1879 276
rect 1791 230 1817 262
rect 1849 230 1879 262
rect 1791 194 1879 230
rect 1791 162 1817 194
rect 1849 162 1879 194
rect 1791 148 1879 162
rect 1825 128 1879 148
rect 1905 262 1973 276
rect 1905 230 1927 262
rect 1959 230 1973 262
rect 1905 176 1973 230
rect 1905 144 1927 176
rect 1959 144 1973 176
rect 1905 128 1973 144
<< pdiff >>
rect 91 594 159 612
rect 91 562 105 594
rect 137 562 159 594
rect 91 526 159 562
rect 91 494 105 526
rect 137 494 159 526
rect 91 458 159 494
rect 91 426 105 458
rect 137 426 159 458
rect 91 412 159 426
rect 185 594 255 612
rect 185 562 207 594
rect 239 585 255 594
rect 700 628 760 642
rect 700 596 714 628
rect 746 596 760 628
rect 700 585 760 596
rect 825 585 880 631
rect 239 562 269 585
rect 185 526 269 562
rect 185 494 207 526
rect 239 494 269 526
rect 185 458 269 494
rect 185 426 207 458
rect 239 426 269 458
rect 185 412 269 426
rect 216 385 269 412
rect 295 385 461 585
rect 487 569 563 585
rect 487 537 509 569
rect 541 537 563 569
rect 487 501 563 537
rect 487 469 509 501
rect 541 469 563 501
rect 487 433 563 469
rect 487 401 509 433
rect 541 401 563 433
rect 487 385 563 401
rect 589 385 653 585
rect 679 385 779 585
rect 805 431 880 585
rect 906 574 1083 631
rect 906 542 928 574
rect 960 542 1029 574
rect 1061 542 1083 574
rect 906 478 1083 542
rect 906 446 928 478
rect 960 446 1029 478
rect 1061 446 1083 478
rect 906 431 1083 446
rect 1109 431 1163 631
rect 1189 615 1257 631
rect 1189 583 1211 615
rect 1243 583 1257 615
rect 1189 431 1257 583
rect 1299 622 1367 636
rect 1299 590 1313 622
rect 1345 590 1367 622
rect 1299 553 1367 590
rect 1299 521 1313 553
rect 1345 521 1367 553
rect 1299 483 1367 521
rect 1299 451 1313 483
rect 1345 451 1367 483
rect 1299 436 1367 451
rect 1393 621 1482 636
rect 1393 589 1419 621
rect 1451 589 1482 621
rect 1393 552 1482 589
rect 1393 520 1419 552
rect 1451 520 1482 552
rect 1393 482 1482 520
rect 1393 450 1419 482
rect 1451 450 1482 482
rect 1393 436 1482 450
rect 1508 574 1576 636
rect 1818 631 1883 636
rect 1508 542 1530 574
rect 1562 542 1576 574
rect 1508 482 1576 542
rect 1508 450 1530 482
rect 1562 450 1576 482
rect 1508 436 1576 450
rect 1658 574 1726 631
rect 1658 542 1672 574
rect 1704 542 1726 574
rect 1658 483 1726 542
rect 1658 451 1672 483
rect 1704 451 1726 483
rect 805 385 860 431
rect 1658 431 1726 451
rect 1752 619 1883 631
rect 1752 587 1829 619
rect 1861 587 1883 619
rect 1752 551 1883 587
rect 1752 519 1829 551
rect 1861 519 1883 551
rect 1752 431 1883 519
rect 1832 412 1883 431
rect 1909 605 1977 636
rect 1909 573 1931 605
rect 1963 573 1977 605
rect 1909 412 1977 573
<< ndiffc >>
rect 85 200 117 232
rect 85 132 117 164
rect 207 132 239 164
rect 420 190 452 222
rect 712 132 744 164
rect 925 132 957 164
rect 1119 150 1151 182
rect 1233 183 1265 215
rect 1399 242 1431 274
rect 1501 174 1533 206
rect 1707 230 1739 262
rect 1707 162 1739 194
rect 1233 92 1265 124
rect 1817 230 1849 262
rect 1817 162 1849 194
rect 1927 230 1959 262
rect 1927 144 1959 176
<< pdiffc >>
rect 105 562 137 594
rect 105 494 137 526
rect 105 426 137 458
rect 207 562 239 594
rect 714 596 746 628
rect 207 494 239 526
rect 207 426 239 458
rect 509 537 541 569
rect 509 469 541 501
rect 509 401 541 433
rect 928 542 960 574
rect 1029 542 1061 574
rect 928 446 960 478
rect 1029 446 1061 478
rect 1211 583 1243 615
rect 1313 590 1345 622
rect 1313 521 1345 553
rect 1313 451 1345 483
rect 1419 589 1451 621
rect 1419 520 1451 552
rect 1419 450 1451 482
rect 1530 542 1562 574
rect 1530 450 1562 482
rect 1672 542 1704 574
rect 1672 451 1704 483
rect 1829 587 1861 619
rect 1829 519 1861 551
rect 1931 573 1963 605
<< psubdiff >>
rect 0 16 2016 30
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 608 16
rect 640 -16 704 16
rect 736 -16 800 16
rect 832 -16 896 16
rect 928 -16 992 16
rect 1024 -16 1088 16
rect 1120 -16 1184 16
rect 1216 -16 1280 16
rect 1312 -16 1376 16
rect 1408 -16 1472 16
rect 1504 -16 1568 16
rect 1600 -16 1664 16
rect 1696 -16 1760 16
rect 1792 -16 1856 16
rect 1888 -16 1952 16
rect 1984 -16 2016 16
rect 0 -30 2016 -16
<< nsubdiff >>
rect 0 772 2016 786
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 608 772
rect 640 740 704 772
rect 736 740 800 772
rect 832 740 896 772
rect 928 740 992 772
rect 1024 740 1088 772
rect 1120 740 1184 772
rect 1216 740 1280 772
rect 1312 740 1376 772
rect 1408 740 1472 772
rect 1504 740 1568 772
rect 1600 740 1664 772
rect 1696 740 1760 772
rect 1792 740 1856 772
rect 1888 740 1952 772
rect 1984 740 2016 772
rect 0 726 2016 740
<< psubdiffcont >>
rect 32 -16 64 16
rect 128 -16 160 16
rect 224 -16 256 16
rect 320 -16 352 16
rect 416 -16 448 16
rect 512 -16 544 16
rect 608 -16 640 16
rect 704 -16 736 16
rect 800 -16 832 16
rect 896 -16 928 16
rect 992 -16 1024 16
rect 1088 -16 1120 16
rect 1184 -16 1216 16
rect 1280 -16 1312 16
rect 1376 -16 1408 16
rect 1472 -16 1504 16
rect 1568 -16 1600 16
rect 1664 -16 1696 16
rect 1760 -16 1792 16
rect 1856 -16 1888 16
rect 1952 -16 1984 16
<< nsubdiffcont >>
rect 32 740 64 772
rect 128 740 160 772
rect 224 740 256 772
rect 320 740 352 772
rect 416 740 448 772
rect 512 740 544 772
rect 608 740 640 772
rect 704 740 736 772
rect 800 740 832 772
rect 896 740 928 772
rect 992 740 1024 772
rect 1088 740 1120 772
rect 1184 740 1216 772
rect 1280 740 1312 772
rect 1376 740 1408 772
rect 1472 740 1504 772
rect 1568 740 1600 772
rect 1664 740 1696 772
rect 1760 740 1792 772
rect 1856 740 1888 772
rect 1952 740 1984 772
<< poly >>
rect 159 657 906 685
rect 159 612 185 657
rect 269 585 295 621
rect 461 585 487 657
rect 880 631 906 657
rect 1083 631 1109 667
rect 1163 631 1189 667
rect 1367 636 1393 672
rect 1482 636 1508 672
rect 563 585 589 621
rect 653 585 679 621
rect 779 585 805 621
rect 159 353 185 412
rect 1726 631 1752 667
rect 1883 636 1909 672
rect 880 412 906 431
rect 269 353 295 385
rect 461 370 487 385
rect 137 336 205 353
rect 137 304 157 336
rect 189 304 205 336
rect 137 287 205 304
rect 248 336 314 353
rect 248 304 265 336
rect 297 304 314 336
rect 248 287 314 304
rect 350 333 416 350
rect 350 301 367 333
rect 399 301 416 333
rect 139 246 165 287
rect 282 246 308 287
rect 350 284 416 301
rect 356 246 382 284
rect 461 261 500 370
rect 563 334 589 385
rect 653 353 679 385
rect 779 353 805 385
rect 880 382 1004 412
rect 1083 399 1109 431
rect 644 336 710 353
rect 536 317 602 334
rect 536 285 553 317
rect 585 285 602 317
rect 536 268 602 285
rect 644 304 661 336
rect 693 304 710 336
rect 644 287 710 304
rect 752 336 818 353
rect 752 304 769 336
rect 801 304 818 336
rect 752 287 818 304
rect 860 317 926 334
rect 474 246 500 261
rect 644 246 670 287
rect 784 246 810 287
rect 860 285 877 317
rect 909 285 926 317
rect 860 268 926 285
rect 974 291 1004 382
rect 1046 382 1109 399
rect 1046 350 1063 382
rect 1095 350 1109 382
rect 1046 333 1109 350
rect 1163 399 1189 431
rect 1163 382 1280 399
rect 1163 350 1231 382
rect 1263 350 1280 382
rect 1163 291 1280 350
rect 1367 342 1393 436
rect 1482 362 1508 436
rect 1570 382 1636 399
rect 1570 362 1587 382
rect 860 246 886 268
rect 974 261 1023 291
rect 997 246 1023 261
rect 1071 261 1280 291
rect 1351 312 1393 342
rect 1453 350 1587 362
rect 1619 350 1636 382
rect 1453 332 1636 350
rect 1726 380 1752 431
rect 1883 380 1909 412
rect 1726 363 1791 380
rect 1351 288 1377 312
rect 1453 288 1479 332
rect 1726 331 1742 363
rect 1774 331 1791 363
rect 1726 314 1791 331
rect 1833 363 1909 380
rect 1833 331 1850 363
rect 1882 331 1909 363
rect 1833 314 1909 331
rect 1071 246 1097 261
rect 1765 276 1791 314
rect 1879 276 1905 314
rect 139 82 165 118
rect 282 82 308 118
rect 356 82 382 118
rect 474 82 500 118
rect 644 82 670 118
rect 784 82 810 118
rect 860 82 886 118
rect 997 82 1023 118
rect 1071 82 1097 118
rect 1351 88 1377 160
rect 1453 124 1479 160
rect 1765 88 1791 148
rect 1879 92 1905 128
rect 1351 62 1791 88
<< polycont >>
rect 157 304 189 336
rect 265 304 297 336
rect 367 301 399 333
rect 553 285 585 317
rect 661 304 693 336
rect 769 304 801 336
rect 877 285 909 317
rect 1063 350 1095 382
rect 1231 350 1263 382
rect 1587 350 1619 382
rect 1742 331 1774 363
rect 1850 331 1882 363
<< metal1 >>
rect 0 772 2016 800
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 608 772
rect 640 740 704 772
rect 736 740 800 772
rect 832 740 896 772
rect 928 740 992 772
rect 1024 740 1088 772
rect 1120 740 1184 772
rect 1216 740 1280 772
rect 1312 740 1376 772
rect 1408 740 1472 772
rect 1504 740 1568 772
rect 1600 740 1664 772
rect 1696 740 1760 772
rect 1792 740 1856 772
rect 1888 740 1952 772
rect 1984 740 2016 772
rect 0 712 2016 740
rect 66 594 149 597
rect 66 562 105 594
rect 137 562 149 594
rect 66 526 149 562
rect 66 494 105 526
rect 137 494 149 526
rect 66 458 149 494
rect 66 426 105 458
rect 137 426 149 458
rect 66 424 149 426
rect 197 594 249 712
rect 704 628 756 712
rect 704 596 714 628
rect 746 596 756 628
rect 704 594 756 596
rect 803 625 1154 659
rect 197 562 207 594
rect 239 562 249 594
rect 197 526 249 562
rect 197 494 207 526
rect 239 494 249 526
rect 197 458 249 494
rect 197 426 207 458
rect 239 426 249 458
rect 197 424 249 426
rect 452 569 554 581
rect 452 537 509 569
rect 541 545 554 569
rect 803 545 848 625
rect 541 537 848 545
rect 452 511 848 537
rect 905 574 1077 589
rect 905 542 928 574
rect 960 542 1029 574
rect 1061 542 1077 574
rect 452 501 554 511
rect 452 469 509 501
rect 541 469 554 501
rect 905 478 1077 542
rect 1114 545 1154 625
rect 1190 615 1256 712
rect 1190 583 1211 615
rect 1243 583 1256 615
rect 1190 581 1256 583
rect 1302 622 1356 640
rect 1302 590 1313 622
rect 1345 590 1356 622
rect 1302 553 1356 590
rect 1302 545 1313 553
rect 1114 521 1313 545
rect 1345 521 1356 553
rect 1114 511 1356 521
rect 452 433 554 469
rect 66 240 100 424
rect 452 401 509 433
rect 541 401 554 433
rect 452 390 554 401
rect 141 336 208 384
rect 141 304 157 336
rect 189 304 208 336
rect 141 287 208 304
rect 248 336 314 384
rect 248 304 265 336
rect 297 304 314 336
rect 248 287 314 304
rect 350 333 416 350
rect 350 301 367 333
rect 399 301 416 333
rect 350 284 416 301
rect 350 240 383 284
rect 452 240 484 390
rect 644 336 708 474
rect 66 232 383 240
rect 66 200 85 232
rect 117 204 383 232
rect 117 200 128 204
rect 66 164 128 200
rect 66 132 85 164
rect 117 132 128 164
rect 66 118 128 132
rect 197 164 249 168
rect 197 132 207 164
rect 239 132 249 164
rect 197 44 249 132
rect 350 129 383 204
rect 419 222 484 240
rect 419 190 420 222
rect 452 190 484 222
rect 419 174 484 190
rect 536 317 602 334
rect 536 285 553 317
rect 585 285 602 317
rect 644 304 661 336
rect 693 304 708 336
rect 644 287 708 304
rect 744 336 818 474
rect 905 446 928 478
rect 960 446 1029 478
rect 1061 474 1077 478
rect 1302 483 1356 511
rect 1061 446 1177 474
rect 905 440 1177 446
rect 744 304 769 336
rect 801 304 818 336
rect 960 382 1107 394
rect 960 350 1063 382
rect 1095 350 1107 382
rect 744 287 818 304
rect 860 317 922 334
rect 536 242 602 285
rect 860 285 877 317
rect 909 285 922 317
rect 860 242 922 285
rect 960 333 1107 350
rect 960 242 994 333
rect 1143 276 1177 440
rect 1302 451 1313 483
rect 1345 451 1356 483
rect 1302 434 1356 451
rect 1214 382 1280 400
rect 1214 350 1231 382
rect 1263 350 1280 382
rect 1214 312 1280 350
rect 536 210 994 242
rect 1030 242 1275 276
rect 536 129 570 210
rect 1030 174 1064 242
rect 1223 215 1275 242
rect 350 95 570 129
rect 699 164 754 167
rect 699 132 712 164
rect 744 132 754 164
rect 699 44 754 132
rect 910 164 1064 174
rect 910 132 925 164
rect 957 132 1064 164
rect 910 119 1064 132
rect 1109 182 1161 202
rect 1109 150 1119 182
rect 1151 150 1161 182
rect 1109 44 1161 150
rect 1223 183 1233 215
rect 1265 183 1275 215
rect 1223 124 1275 183
rect 1316 196 1356 434
rect 1402 625 1782 659
rect 1402 621 1460 625
rect 1402 589 1419 621
rect 1451 589 1460 621
rect 1402 552 1460 589
rect 1402 520 1419 552
rect 1451 520 1460 552
rect 1402 482 1460 520
rect 1402 450 1419 482
rect 1451 450 1460 482
rect 1402 301 1460 450
rect 1393 274 1460 301
rect 1393 242 1399 274
rect 1431 267 1460 274
rect 1502 574 1572 584
rect 1502 542 1530 574
rect 1562 542 1572 574
rect 1502 482 1572 542
rect 1502 450 1530 482
rect 1562 450 1572 482
rect 1502 444 1572 450
rect 1639 574 1714 584
rect 1639 542 1672 574
rect 1704 542 1714 574
rect 1639 483 1714 542
rect 1639 451 1672 483
rect 1704 451 1714 483
rect 1502 297 1534 444
rect 1639 434 1714 451
rect 1750 480 1782 625
rect 1819 619 1871 712
rect 1819 587 1829 619
rect 1861 587 1871 619
rect 1819 551 1871 587
rect 1928 605 1981 615
rect 1928 573 1931 605
rect 1963 573 1981 605
rect 1928 556 1981 573
rect 1819 519 1829 551
rect 1861 519 1871 551
rect 1819 517 1871 519
rect 1750 446 1892 480
rect 1639 399 1671 434
rect 1570 382 1671 399
rect 1570 350 1587 382
rect 1619 350 1671 382
rect 1570 333 1671 350
rect 1431 242 1442 267
rect 1502 265 1603 297
rect 1393 232 1442 242
rect 1490 206 1535 216
rect 1490 196 1501 206
rect 1316 174 1501 196
rect 1533 174 1535 206
rect 1316 164 1535 174
rect 1223 92 1233 124
rect 1265 120 1275 124
rect 1571 120 1603 265
rect 1639 277 1671 333
rect 1707 363 1791 397
rect 1707 331 1742 363
rect 1774 331 1791 363
rect 1707 313 1791 331
rect 1839 363 1892 446
rect 1839 331 1850 363
rect 1882 331 1892 363
rect 1839 314 1892 331
rect 1639 262 1749 277
rect 1933 272 1981 556
rect 1639 230 1707 262
rect 1739 230 1749 262
rect 1639 194 1749 230
rect 1639 162 1707 194
rect 1739 162 1749 194
rect 1639 151 1749 162
rect 1807 262 1859 265
rect 1807 230 1817 262
rect 1849 230 1859 262
rect 1807 194 1859 230
rect 1807 162 1817 194
rect 1849 162 1859 194
rect 1265 92 1603 120
rect 1223 88 1603 92
rect 1807 44 1859 162
rect 1895 262 1981 272
rect 1895 230 1927 262
rect 1959 230 1981 262
rect 1895 176 1981 230
rect 1895 144 1927 176
rect 1959 144 1981 176
rect 1895 124 1981 144
rect 0 16 2016 44
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 608 16
rect 640 -16 704 16
rect 736 -16 800 16
rect 832 -16 896 16
rect 928 -16 992 16
rect 1024 -16 1088 16
rect 1120 -16 1184 16
rect 1216 -16 1280 16
rect 1312 -16 1376 16
rect 1408 -16 1472 16
rect 1504 -16 1568 16
rect 1600 -16 1664 16
rect 1696 -16 1760 16
rect 1792 -16 1856 16
rect 1888 -16 1952 16
rect 1984 -16 2016 16
rect 0 -44 2016 -16
<< labels >>
flabel metal1 s 1895 124 1981 272 0 FreeSans 400 0 0 0 X
port 2 nsew
flabel metal1 s 644 287 708 474 0 FreeSans 400 0 0 0 A1
port 3 nsew
flabel metal1 s 744 287 818 474 0 FreeSans 400 0 0 0 A2
port 4 nsew
flabel metal1 s 141 287 208 384 0 FreeSans 400 0 0 0 S0
port 5 nsew
flabel metal1 s 0 712 2016 800 0 FreeSans 400 0 0 0 VDD
port 6 nsew
flabel metal1 s 0 -44 2016 44 0 FreeSans 400 0 0 0 VSS
port 7 nsew
flabel metal1 s 1707 313 1791 397 0 FreeSans 400 0 0 0 S1
port 8 nsew
flabel metal1 s 248 287 314 384 0 FreeSans 400 0 0 0 A0
port 9 nsew
flabel metal1 s 1214 312 1280 400 0 FreeSans 400 0 0 0 A3
port 10 nsew
<< properties >>
string FIXED_BBOX 0 0 2016 756
string GDS_END 173986
string GDS_FILE ../gds/controller.gds
string GDS_START 161988
<< end >>
