magic
tech ihp-sg13g2
timestamp 1747537721
<< nwell >>
rect -24 175 216 417
<< pwell >>
rect 16 28 171 149
rect -13 -28 205 28
<< nmos >>
rect 63 97 76 136
rect 111 48 124 136
<< pmos >>
rect 63 247 76 277
rect 111 225 124 330
<< ndiff >>
rect 29 125 63 136
rect 29 109 36 125
rect 52 109 63 125
rect 29 97 63 109
rect 76 97 111 136
rect 83 70 111 97
rect 29 51 111 70
rect 29 35 57 51
rect 73 48 111 51
rect 124 119 158 136
rect 124 103 135 119
rect 151 103 158 119
rect 124 71 158 103
rect 124 55 135 71
rect 151 55 158 71
rect 124 48 158 55
rect 73 35 101 48
rect 29 18 101 35
<< pdiff >>
rect 29 338 101 360
rect 29 322 54 338
rect 70 330 101 338
rect 70 322 111 330
rect 29 304 111 322
rect 85 277 111 304
rect 29 270 63 277
rect 29 254 36 270
rect 52 254 63 270
rect 29 247 63 254
rect 76 247 111 277
rect 88 225 111 247
rect 124 282 158 330
rect 124 266 135 282
rect 151 266 158 282
rect 124 248 158 266
rect 124 232 135 248
rect 151 232 158 248
rect 124 225 158 232
<< ndiffc >>
rect 36 109 52 125
rect 57 35 73 51
rect 135 103 151 119
rect 135 55 151 71
<< pdiffc >>
rect 54 322 70 338
rect 36 254 52 270
rect 135 266 151 282
rect 135 232 151 248
<< psubdiff >>
rect 29 15 101 18
rect 0 8 192 15
rect 0 -8 16 8
rect 32 -8 64 8
rect 80 -8 112 8
rect 128 -8 160 8
rect 176 -8 192 8
rect 0 -15 192 -8
<< nsubdiff >>
rect 0 386 192 393
rect 0 370 16 386
rect 32 370 64 386
rect 80 370 112 386
rect 128 370 160 386
rect 176 370 192 386
rect 0 363 192 370
rect 29 360 101 363
<< psubdiffcont >>
rect 16 -8 32 8
rect 64 -8 80 8
rect 112 -8 128 8
rect 160 -8 176 8
<< nsubdiffcont >>
rect 16 370 32 386
rect 64 370 80 386
rect 112 370 128 386
rect 160 370 176 386
<< poly >>
rect 111 330 124 349
rect 63 277 76 296
rect 63 239 76 247
rect 29 232 76 239
rect 29 216 36 232
rect 52 226 76 232
rect 52 216 67 226
rect 29 209 67 216
rect 54 157 67 209
rect 111 208 124 225
rect 85 201 124 208
rect 85 185 92 201
rect 108 193 124 201
rect 108 185 115 193
rect 85 181 115 185
rect 85 180 114 181
rect 85 179 113 180
rect 85 178 112 179
rect 133 173 160 174
rect 132 172 160 173
rect 131 171 160 172
rect 130 167 160 171
rect 130 157 137 167
rect 54 144 76 157
rect 63 136 76 144
rect 111 151 137 157
rect 153 151 160 167
rect 111 144 160 151
rect 111 136 124 144
rect 63 78 76 97
rect 111 29 124 48
<< polycont >>
rect 36 216 52 232
rect 92 185 108 201
rect 137 151 153 167
<< metal1 >>
rect 0 386 192 400
rect 0 370 16 386
rect 32 370 64 386
rect 80 370 112 386
rect 128 370 160 386
rect 176 370 192 386
rect 0 356 192 370
rect 45 338 78 356
rect 45 322 54 338
rect 70 322 78 338
rect 45 316 78 322
rect 130 282 158 287
rect 31 270 57 276
rect 31 254 36 270
rect 52 254 57 270
rect 31 232 57 254
rect 31 216 36 232
rect 52 216 57 232
rect 31 211 57 216
rect 130 266 135 282
rect 151 266 158 282
rect 130 248 158 266
rect 130 232 135 248
rect 151 232 158 248
rect 87 201 111 206
rect 87 185 92 201
rect 108 185 111 201
rect 87 129 111 185
rect 130 167 158 232
rect 130 151 137 167
rect 153 151 158 167
rect 130 146 158 151
rect 31 125 111 129
rect 31 109 36 125
rect 52 109 111 125
rect 31 103 111 109
rect 129 119 158 123
rect 129 103 135 119
rect 151 103 158 119
rect 129 77 158 103
rect 109 71 158 77
rect 46 51 81 60
rect 46 35 57 51
rect 73 35 81 51
rect 109 55 135 71
rect 151 55 158 71
rect 109 48 158 55
rect 46 22 81 35
rect 0 8 192 22
rect 0 -8 16 8
rect 32 -8 64 8
rect 80 -8 112 8
rect 128 -8 160 8
rect 176 -8 192 8
rect 0 -22 192 -8
<< labels >>
flabel metal1 s 129 48 158 123 0 FreeSans 200 0 0 0 L_LO
port 2 nsew
flabel metal1 s 0 356 192 400 0 FreeSans 200 0 0 0 VDD
port 3 nsew
flabel metal1 s 0 -22 192 22 0 FreeSans 200 0 0 0 VSS
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 192 378
string GDS_END 261516
string GDS_FILE ../gds/controller.gds
string GDS_START 257776
<< end >>
