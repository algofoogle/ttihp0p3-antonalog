magic
tech ihp-sg13g2
timestamp 1747489030
<< pwell >>
rect -1401 -512 1941 392
<< psubdiff >>
rect -1370 354 1910 361
rect -1370 338 -1324 354
rect 1864 338 1910 354
rect -1370 331 1910 338
rect -1370 315 -1340 331
rect -1370 -435 -1363 315
rect -1347 -435 -1340 315
rect -1370 -451 -1340 -435
rect 1880 315 1910 331
rect 1880 -435 1887 315
rect 1903 -435 1910 315
rect 1880 -451 1910 -435
rect -1370 -458 1910 -451
rect -1370 -474 -1324 -458
rect 1864 -474 1910 -458
rect -1370 -481 1910 -474
<< psubdiffcont >>
rect -1324 338 1864 354
rect -1363 -435 -1347 315
rect 1887 -435 1903 315
rect -1324 -474 1864 -458
<< metal1 >>
rect -1363 338 -1324 354
rect 1864 338 1903 354
rect -1363 315 -1311 338
rect -1347 -360 -1311 315
rect 1887 315 1903 338
rect -1292 240 -1066 283
rect -1040 240 -814 283
rect -788 240 -562 283
rect -536 240 -436 313
rect -662 183 -562 240
rect -410 183 -310 283
rect -284 240 -58 283
rect -32 240 194 283
rect 220 240 320 313
rect -662 140 -310 183
rect 94 183 194 240
rect 346 183 446 283
rect 472 240 698 283
rect 724 240 950 283
rect 976 240 1076 313
rect 94 140 446 183
rect 850 183 950 240
rect 1102 183 1202 283
rect 1228 240 1454 283
rect 1480 240 1706 313
rect 1732 240 1832 313
rect 850 140 1202 183
rect -1040 -303 -688 -260
rect -1040 -360 -940 -303
rect -1347 -435 -1192 -360
rect -1166 -403 -940 -360
rect -914 -433 -814 -360
rect -788 -403 -688 -303
rect -284 -303 68 -260
rect -284 -360 -184 -303
rect -662 -403 -436 -360
rect -410 -403 -184 -360
rect -158 -433 -58 -360
rect -32 -403 68 -303
rect 472 -303 824 -260
rect 472 -360 572 -303
rect 94 -403 320 -360
rect 346 -403 572 -360
rect 598 -433 698 -360
rect 724 -403 824 -303
rect 1228 -303 1580 -260
rect 1228 -360 1328 -303
rect 850 -403 1076 -360
rect 1102 -403 1328 -360
rect 1354 -433 1454 -360
rect 1480 -403 1580 -303
rect 1606 -403 1832 -360
rect -1363 -458 -1192 -435
rect 1887 -458 1903 -435
rect -1363 -474 -1324 -458
rect 1864 -474 1903 -458
use rhigh  res
array 0 24 126 0 0 686
timestamp 1746838591
transform 1 0 -1292 0 1 -360
box 0 -43 100 643
<< labels >>
flabel metal1 -1292 240 -1066 283 0 FreeSans 160 0 0 0 wg0
flabel metal1 -1166 -403 -940 -360 0 FreeSans 160 0 0 0 wJ0
flabel metal1 -1040 240 -814 283 0 FreeSans 160 0 0 0 wi0
flabel metal1 -899 -418 -869 -388 0 FreeSans 160 0 0 0 IN[0]
port 0 nsew
flabel metal1 -788 240 -562 283 0 FreeSans 160 0 0 0 wJ1
flabel metal1 -662 -403 -436 -360 0 FreeSans 160 0 0 0 wi1
flabel metal1 -521 268 -491 298 0 FreeSans 160 0 0 0 IN[1]
port 1 nsew
flabel metal1 -410 -403 -184 -360 0 FreeSans 160 0 0 0 wJ2
flabel metal1 -284 240 -58 283 0 FreeSans 160 0 0 0 wi2
flabel metal1 -143 -418 -113 -388 0 FreeSans 160 0 0 0 IN[2]
port 2 nsew
flabel metal1 -32 240 194 283 0 FreeSans 160 0 0 0 wJ3
flabel metal1 94 -403 320 -360 0 FreeSans 160 0 0 0 wi3
flabel metal1 235 268 265 298 0 FreeSans 160 0 0 0 IN[3]
port 3 nsew
flabel metal1 346 -403 572 -360 0 FreeSans 160 0 0 0 wJ4
flabel metal1 472 240 698 283 0 FreeSans 160 0 0 0 wi4
flabel metal1 613 -418 643 -388 0 FreeSans 160 0 0 0 IN[4]
port 4 nsew
flabel metal1 724 240 950 283 0 FreeSans 160 0 0 0 wJ5
flabel metal1 850 -403 1076 -360 0 FreeSans 160 0 0 0 wi5
flabel metal1 991 268 1021 298 0 FreeSans 160 0 0 0 IN[5]
port 5 nsew
flabel metal1 1102 -403 1328 -360 0 FreeSans 160 0 0 0 wJ6
flabel metal1 1228 240 1454 283 0 FreeSans 160 0 0 0 wi6
flabel metal1 1369 -418 1399 -388 0 FreeSans 160 0 0 0 IN[6]
port 6 nsew
flabel metal1 1606 -403 1832 -360 0 FreeSans 160 0 0 0 wi7
flabel metal1 1747 268 1777 298 0 FreeSans 160 0 0 0 IN[7]
port 7 nsew
flabel metal1 1495 268 1525 298 0 FreeSans 160 0 0 0 OUT
port 8 nsew
flabel metal1 -1285 -435 -1255 -405 0 FreeSans 160 0 0 0 GND
port 9 nsew
<< end >>
