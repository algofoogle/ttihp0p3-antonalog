magic
tech ihp-sg13g2
magscale 1 2
timestamp 1746812698
<< error_s >>
rect 8245 28980 8287 28989
rect 9013 28980 9055 28989
rect 25141 28980 25183 28989
rect 25381 28980 25423 28989
rect 37700 28980 37758 28981
rect 8245 28940 8246 28980
rect 9013 28940 9014 28980
rect 25141 28940 25142 28980
rect 25381 28940 25382 28980
rect 37700 28940 37709 28980
rect 8245 28931 8287 28940
rect 9013 28931 9055 28940
rect 25141 28931 25183 28940
rect 25381 28931 25423 28940
rect 37700 28939 37758 28940
rect 9301 28896 9343 28905
rect 11108 28896 11166 28897
rect 11972 28896 12030 28897
rect 19556 28896 19614 28897
rect 21860 28896 21918 28897
rect 9301 28856 9302 28896
rect 11108 28856 11117 28896
rect 11972 28856 11981 28896
rect 19556 28856 19565 28896
rect 21860 28856 21869 28896
rect 9301 28847 9343 28856
rect 11108 28855 11166 28856
rect 11972 28855 12030 28856
rect 19556 28855 19614 28856
rect 21860 28855 21918 28856
rect 9205 28812 9247 28821
rect 9380 28812 9438 28813
rect 9596 28812 9638 28821
rect 9764 28812 9822 28813
rect 10352 28812 10394 28821
rect 10532 28812 10590 28813
rect 11797 28812 11839 28821
rect 12356 28812 12414 28813
rect 14852 28812 14910 28813
rect 17348 28812 17406 28813
rect 21476 28812 21534 28813
rect 22820 28812 22878 28813
rect 24935 28812 24977 28821
rect 25525 28812 25567 28821
rect 25717 28812 25759 28821
rect 26948 28812 27006 28813
rect 29732 28812 29790 28813
rect 33764 28812 33822 28813
rect 34148 28812 34206 28813
rect 34724 28812 34782 28813
rect 37525 28812 37567 28821
rect 37861 28812 37903 28821
rect 38005 28812 38047 28821
rect 9205 28772 9206 28812
rect 9380 28772 9389 28812
rect 9596 28772 9597 28812
rect 9764 28772 9773 28812
rect 10352 28772 10353 28812
rect 10532 28772 10541 28812
rect 11797 28772 11798 28812
rect 12356 28772 12365 28812
rect 14852 28772 14861 28812
rect 17348 28772 17357 28812
rect 21476 28772 21485 28812
rect 22820 28772 22829 28812
rect 24935 28772 24936 28812
rect 25237 28803 25279 28812
rect 9205 28763 9247 28772
rect 9380 28771 9438 28772
rect 9596 28763 9638 28772
rect 9764 28771 9822 28772
rect 10352 28763 10394 28772
rect 10532 28771 10590 28772
rect 11797 28763 11839 28772
rect 12356 28771 12414 28772
rect 14852 28771 14910 28772
rect 17348 28771 17406 28772
rect 21476 28771 21534 28772
rect 22820 28771 22878 28772
rect 24935 28763 24977 28772
rect 25237 28763 25238 28803
rect 25525 28772 25526 28812
rect 25717 28772 25718 28812
rect 26948 28772 26957 28812
rect 29732 28772 29741 28812
rect 33764 28772 33773 28812
rect 34148 28772 34157 28812
rect 34724 28772 34733 28812
rect 37525 28772 37526 28812
rect 37861 28772 37862 28812
rect 38005 28772 38006 28812
rect 38188 28803 38234 28812
rect 25525 28763 25567 28772
rect 25717 28763 25759 28772
rect 26948 28771 27006 28772
rect 29732 28771 29790 28772
rect 33764 28771 33822 28772
rect 34148 28771 34206 28772
rect 34724 28771 34782 28772
rect 37525 28763 37567 28772
rect 37861 28763 37903 28772
rect 38005 28763 38047 28772
rect 38188 28763 38189 28803
rect 25237 28754 25279 28763
rect 38188 28754 38234 28763
rect 14485 28728 14527 28737
rect 16981 28728 17023 28737
rect 22453 28728 22495 28737
rect 26389 28728 26431 28737
rect 26581 28728 26623 28737
rect 29365 28728 29407 28737
rect 34357 28728 34399 28737
rect 38341 28728 38383 28737
rect 14485 28688 14486 28728
rect 14861 28688 14870 28728
rect 16981 28688 16982 28728
rect 17933 28688 17942 28728
rect 21581 28688 21590 28728
rect 22453 28688 22454 28728
rect 23117 28688 23126 28728
rect 26389 28688 26390 28728
rect 26581 28688 26582 28728
rect 29365 28688 29366 28728
rect 29933 28688 29942 28728
rect 34357 28688 34358 28728
rect 34733 28688 34742 28728
rect 38341 28688 38342 28728
rect 14485 28679 14527 28688
rect 16981 28679 17023 28688
rect 22453 28679 22495 28688
rect 26389 28679 26431 28688
rect 26581 28679 26623 28688
rect 29365 28679 29407 28688
rect 34357 28679 34399 28688
rect 38341 28679 38383 28688
rect 8629 28644 8671 28653
rect 9764 28644 9822 28645
rect 10165 28644 10207 28653
rect 10933 28644 10975 28653
rect 22261 28644 22303 28653
rect 24757 28644 24799 28653
rect 8629 28604 8630 28644
rect 9764 28604 9773 28644
rect 10165 28604 10166 28644
rect 10933 28604 10934 28644
rect 22261 28604 22262 28644
rect 24757 28604 24758 28644
rect 8629 28595 8671 28604
rect 9764 28603 9822 28604
rect 10165 28595 10207 28604
rect 10933 28595 10975 28604
rect 22261 28595 22303 28604
rect 24757 28595 24799 28604
rect 10532 28560 10590 28561
rect 14293 28560 14335 28569
rect 16789 28560 16831 28569
rect 19285 28560 19327 28569
rect 24932 28560 24990 28561
rect 28885 28560 28927 28569
rect 31669 28560 31711 28569
rect 31861 28560 31903 28569
rect 36661 28560 36703 28569
rect 36853 28560 36895 28569
rect 10532 28520 10541 28560
rect 14293 28520 14294 28560
rect 16789 28520 16790 28560
rect 19285 28520 19286 28560
rect 24932 28520 24941 28560
rect 28885 28520 28886 28560
rect 31669 28520 31670 28560
rect 31861 28520 31862 28560
rect 36661 28520 36662 28560
rect 36853 28520 36854 28560
rect 10532 28519 10590 28520
rect 14293 28511 14335 28520
rect 16789 28511 16831 28520
rect 19285 28511 19327 28520
rect 24932 28519 24990 28520
rect 28885 28511 28927 28520
rect 31669 28511 31711 28520
rect 31861 28511 31903 28520
rect 36661 28511 36703 28520
rect 36853 28511 36895 28520
rect 9493 28224 9535 28233
rect 10052 28224 10110 28225
rect 14084 28224 14142 28225
rect 15332 28224 15390 28225
rect 17252 28224 17310 28225
rect 19477 28224 19519 28233
rect 22357 28224 22399 28233
rect 26581 28224 26623 28233
rect 30325 28224 30367 28233
rect 33781 28224 33823 28233
rect 35701 28224 35743 28233
rect 9493 28184 9494 28224
rect 10052 28184 10061 28224
rect 14084 28184 14093 28224
rect 15332 28184 15341 28224
rect 17252 28184 17261 28224
rect 19477 28184 19478 28224
rect 22357 28184 22358 28224
rect 26581 28184 26582 28224
rect 30325 28184 30326 28224
rect 33781 28184 33782 28224
rect 35701 28184 35702 28224
rect 9493 28175 9535 28184
rect 10052 28183 10110 28184
rect 14084 28183 14142 28184
rect 15332 28183 15390 28184
rect 17252 28183 17310 28184
rect 19477 28175 19519 28184
rect 22357 28175 22399 28184
rect 26581 28175 26623 28184
rect 30325 28175 30367 28184
rect 33781 28175 33823 28184
rect 35701 28175 35743 28184
rect 8533 28140 8575 28149
rect 13909 28140 13951 28149
rect 18517 28140 18559 28149
rect 20149 28140 20191 28149
rect 20821 28140 20863 28149
rect 23029 28140 23071 28149
rect 8533 28100 8534 28140
rect 13909 28100 13910 28140
rect 18517 28100 18518 28140
rect 20149 28100 20150 28140
rect 20821 28100 20822 28140
rect 23029 28100 23030 28140
rect 8533 28091 8575 28100
rect 13909 28091 13951 28100
rect 18517 28091 18559 28100
rect 20149 28091 20191 28100
rect 20821 28091 20863 28100
rect 23029 28091 23071 28100
rect 10628 28056 10686 28057
rect 15157 28056 15199 28065
rect 20917 28056 20959 28065
rect 28004 28056 28062 28057
rect 10628 28016 10637 28056
rect 10925 28016 10934 28056
rect 15157 28016 15158 28056
rect 20917 28016 20918 28056
rect 25709 28016 25718 28056
rect 28004 28016 28013 28056
rect 37517 28016 37526 28056
rect 10628 28015 10686 28016
rect 14377 28005 14419 28014
rect 15157 28007 15199 28016
rect 20917 28007 20959 28016
rect 28004 28015 28062 28016
rect 9493 27972 9535 27981
rect 9685 27972 9727 27981
rect 9877 27972 9919 27981
rect 10052 27972 10110 27973
rect 12164 27972 12222 27973
rect 12548 27972 12606 27973
rect 12949 27972 12991 27981
rect 13037 27972 13095 27973
rect 13285 27972 13327 27981
rect 9493 27932 9494 27972
rect 9685 27932 9686 27972
rect 9877 27932 9878 27972
rect 10052 27932 10061 27972
rect 12164 27932 12173 27972
rect 12548 27932 12557 27972
rect 12949 27932 12950 27972
rect 13037 27932 13046 27972
rect 13285 27932 13286 27972
rect 14377 27965 14378 28005
rect 14468 27972 14526 27973
rect 15541 27972 15583 27981
rect 15629 27972 15687 27973
rect 16021 27972 16063 27981
rect 16109 27972 16167 27973
rect 16309 27972 16351 27981
rect 17549 27972 17607 27973
rect 17845 27972 17887 27981
rect 18325 27972 18367 27981
rect 18805 27972 18847 27981
rect 19189 27972 19231 27981
rect 19303 27972 19361 27973
rect 19430 27972 19488 27973
rect 19652 27972 19710 27973
rect 20341 27972 20383 27981
rect 20590 27972 20648 27973
rect 20746 27972 20788 27981
rect 21044 27972 21102 27973
rect 21205 27972 21247 27981
rect 22148 27972 22206 27973
rect 23221 27972 23263 27981
rect 24452 27972 24510 27973
rect 26869 27972 26911 27981
rect 27253 27972 27295 27981
rect 27733 27972 27775 27981
rect 28693 27972 28735 27981
rect 28928 27972 28970 27981
rect 29060 27972 29118 27973
rect 29173 27972 29215 27981
rect 30133 27972 30175 27981
rect 30997 27972 31039 27981
rect 31861 27972 31903 27981
rect 32725 27972 32767 27981
rect 33589 27972 33631 27981
rect 34453 27972 34495 27981
rect 35317 27972 35359 27981
rect 37604 27972 37662 27973
rect 38293 27972 38335 27981
rect 14377 27956 14419 27965
rect 14468 27932 14477 27972
rect 15541 27932 15542 27972
rect 15629 27932 15638 27972
rect 16021 27932 16022 27972
rect 16109 27932 16118 27972
rect 16309 27932 16310 27972
rect 17549 27932 17558 27972
rect 17845 27932 17846 27972
rect 18325 27932 18326 27972
rect 18805 27932 18806 27972
rect 19189 27932 19190 27972
rect 19303 27932 19312 27972
rect 19430 27932 19439 27972
rect 19652 27932 19661 27972
rect 20341 27932 20342 27972
rect 20590 27932 20599 27972
rect 20746 27932 20747 27972
rect 21044 27932 21053 27972
rect 21205 27932 21206 27972
rect 22148 27932 22157 27972
rect 23221 27932 23222 27972
rect 24452 27932 24461 27972
rect 26869 27932 26870 27972
rect 26965 27963 27007 27972
rect 9493 27923 9535 27932
rect 9685 27923 9727 27932
rect 9877 27923 9919 27932
rect 10052 27931 10110 27932
rect 12164 27931 12222 27932
rect 12548 27931 12606 27932
rect 12949 27923 12991 27932
rect 13037 27931 13095 27932
rect 13285 27923 13327 27932
rect 14468 27931 14526 27932
rect 15541 27923 15583 27932
rect 15629 27931 15687 27932
rect 16021 27923 16063 27932
rect 16109 27931 16167 27932
rect 16309 27923 16351 27932
rect 17549 27931 17607 27932
rect 17845 27923 17887 27932
rect 18325 27923 18367 27932
rect 18805 27923 18847 27932
rect 19189 27923 19231 27932
rect 19303 27931 19361 27932
rect 19430 27931 19488 27932
rect 19652 27931 19710 27932
rect 20341 27923 20383 27932
rect 20590 27931 20648 27932
rect 20746 27923 20788 27932
rect 21044 27931 21102 27932
rect 21205 27923 21247 27932
rect 22148 27931 22206 27932
rect 23221 27923 23263 27932
rect 24452 27931 24510 27932
rect 26869 27923 26911 27932
rect 26965 27923 26966 27963
rect 27253 27932 27254 27972
rect 27733 27932 27734 27972
rect 28693 27932 28694 27972
rect 28928 27932 28929 27972
rect 29060 27932 29069 27972
rect 29173 27932 29174 27972
rect 30133 27932 30134 27972
rect 30997 27932 30998 27972
rect 31861 27932 31862 27972
rect 32725 27932 32726 27972
rect 33589 27932 33590 27972
rect 34453 27932 34454 27972
rect 35317 27932 35318 27972
rect 37604 27932 37613 27972
rect 38293 27932 38294 27972
rect 27253 27923 27295 27932
rect 27733 27923 27775 27932
rect 28693 27923 28735 27932
rect 28928 27923 28970 27932
rect 29060 27931 29118 27932
rect 29173 27923 29215 27932
rect 30133 27923 30175 27932
rect 30997 27923 31039 27932
rect 31861 27923 31903 27932
rect 32725 27923 32767 27932
rect 33589 27923 33631 27932
rect 34453 27923 34495 27932
rect 35317 27923 35359 27932
rect 37604 27931 37662 27932
rect 38293 27923 38335 27932
rect 26965 27914 27007 27923
rect 12743 27888 12785 27897
rect 15335 27888 15377 27897
rect 15815 27888 15857 27897
rect 17255 27888 17297 27897
rect 19971 27888 20013 27897
rect 22436 27888 22494 27889
rect 23893 27888 23935 27897
rect 24068 27888 24126 27889
rect 29252 27888 29310 27889
rect 32900 27888 32958 27889
rect 37988 27888 38046 27889
rect 12743 27848 12744 27888
rect 15335 27848 15336 27888
rect 15815 27848 15816 27888
rect 17255 27848 17256 27888
rect 19971 27848 19972 27888
rect 22436 27848 22445 27888
rect 23893 27848 23894 27888
rect 24068 27848 24077 27888
rect 29252 27848 29261 27888
rect 32900 27848 32909 27888
rect 37988 27848 37997 27888
rect 12743 27839 12785 27848
rect 15335 27839 15377 27848
rect 15815 27839 15857 27848
rect 17255 27839 17297 27848
rect 19971 27839 20013 27848
rect 22436 27847 22494 27848
rect 23893 27839 23935 27848
rect 24068 27847 24126 27848
rect 29252 27847 29310 27848
rect 32900 27847 32958 27848
rect 37988 27847 38046 27848
rect 8917 27804 8959 27813
rect 9301 27804 9343 27813
rect 10261 27804 10303 27813
rect 12836 27804 12894 27805
rect 14917 27804 14959 27813
rect 15541 27804 15583 27813
rect 15908 27804 15966 27805
rect 16981 27804 17023 27813
rect 17461 27804 17503 27813
rect 17732 27804 17790 27805
rect 18037 27804 18079 27813
rect 18212 27804 18270 27805
rect 18692 27804 18750 27805
rect 18997 27804 19039 27813
rect 19748 27804 19806 27805
rect 19861 27804 19903 27813
rect 20389 27804 20431 27813
rect 21877 27804 21919 27813
rect 26389 27804 26431 27813
rect 27541 27804 27583 27813
rect 27812 27804 27870 27805
rect 29461 27804 29503 27813
rect 31189 27804 31231 27813
rect 32053 27804 32095 27813
rect 34645 27804 34687 27813
rect 35701 27804 35743 27813
rect 38180 27804 38238 27805
rect 38485 27804 38527 27813
rect 8917 27764 8918 27804
rect 9301 27764 9302 27804
rect 10261 27764 10262 27804
rect 12836 27764 12845 27804
rect 14917 27764 14918 27804
rect 15541 27764 15542 27804
rect 15908 27764 15917 27804
rect 16981 27764 16982 27804
rect 17461 27764 17462 27804
rect 17732 27764 17741 27804
rect 18037 27764 18038 27804
rect 18212 27764 18221 27804
rect 18692 27764 18701 27804
rect 18997 27764 18998 27804
rect 19748 27764 19757 27804
rect 19861 27764 19862 27804
rect 20389 27764 20390 27804
rect 21877 27764 21878 27804
rect 26389 27764 26390 27804
rect 27541 27764 27542 27804
rect 27812 27764 27821 27804
rect 29461 27764 29462 27804
rect 31189 27764 31190 27804
rect 32053 27764 32054 27804
rect 34645 27764 34646 27804
rect 35701 27764 35702 27804
rect 38180 27764 38189 27804
rect 38485 27764 38486 27804
rect 8917 27755 8959 27764
rect 9301 27755 9343 27764
rect 10261 27755 10303 27764
rect 12836 27763 12894 27764
rect 14612 27762 14670 27763
rect 14612 27722 14621 27762
rect 14917 27755 14959 27764
rect 15541 27755 15583 27764
rect 15908 27763 15966 27764
rect 16981 27755 17023 27764
rect 17461 27755 17503 27764
rect 17732 27763 17790 27764
rect 18037 27755 18079 27764
rect 18212 27763 18270 27764
rect 18692 27763 18750 27764
rect 18997 27755 19039 27764
rect 19748 27763 19806 27764
rect 19861 27755 19903 27764
rect 20389 27755 20431 27764
rect 21877 27755 21919 27764
rect 26389 27755 26431 27764
rect 27541 27755 27583 27764
rect 27812 27763 27870 27764
rect 29461 27755 29503 27764
rect 31189 27755 31231 27764
rect 32053 27755 32095 27764
rect 34645 27755 34687 27764
rect 35701 27755 35743 27764
rect 38180 27763 38238 27764
rect 38485 27755 38527 27764
rect 14612 27721 14670 27722
rect 25412 27510 25470 27511
rect 10069 27468 10111 27477
rect 12421 27468 12463 27477
rect 16213 27468 16255 27477
rect 18709 27468 18751 27477
rect 19573 27468 19615 27477
rect 20132 27468 20190 27469
rect 20900 27468 20958 27469
rect 21013 27468 21055 27477
rect 23749 27468 23791 27477
rect 25412 27470 25421 27510
rect 25412 27469 25470 27470
rect 26293 27468 26335 27477
rect 27908 27468 27966 27469
rect 32581 27468 32623 27477
rect 32900 27468 32958 27469
rect 34453 27468 34495 27477
rect 35221 27468 35263 27477
rect 38677 27468 38719 27477
rect 10069 27428 10070 27468
rect 12421 27428 12422 27468
rect 16213 27428 16214 27468
rect 18709 27428 18710 27468
rect 19573 27428 19574 27468
rect 20132 27428 20141 27468
rect 20900 27428 20909 27468
rect 21013 27428 21014 27468
rect 23749 27428 23750 27468
rect 10069 27419 10111 27428
rect 12421 27419 12463 27428
rect 16213 27419 16255 27428
rect 18709 27419 18751 27428
rect 19573 27419 19615 27428
rect 20132 27427 20190 27428
rect 20900 27427 20958 27428
rect 21013 27419 21055 27428
rect 23749 27419 23791 27428
rect 25537 27426 25579 27435
rect 26293 27428 26294 27468
rect 27908 27428 27917 27468
rect 32581 27428 32582 27468
rect 32900 27428 32909 27468
rect 34453 27428 34454 27468
rect 35221 27428 35222 27468
rect 38677 27428 38678 27468
rect 10405 27384 10447 27393
rect 11413 27384 11455 27393
rect 12085 27384 12127 27393
rect 25537 27386 25538 27426
rect 26293 27419 26335 27428
rect 27908 27427 27966 27428
rect 32581 27419 32623 27428
rect 32900 27427 32958 27428
rect 34453 27419 34495 27428
rect 35221 27419 35263 27428
rect 38677 27419 38719 27428
rect 13892 27384 13950 27385
rect 16388 27384 16446 27385
rect 21284 27384 21342 27385
rect 10405 27344 10406 27384
rect 11413 27344 11414 27384
rect 12085 27344 12086 27384
rect 13892 27344 13901 27384
rect 16388 27344 16397 27384
rect 21284 27344 21293 27384
rect 25537 27377 25579 27386
rect 29444 27384 29502 27385
rect 33829 27384 33871 27393
rect 10405 27335 10447 27344
rect 11413 27335 11455 27344
rect 12085 27335 12127 27344
rect 13892 27343 13950 27344
rect 16388 27343 16446 27344
rect 21284 27343 21342 27344
rect 25457 27342 25499 27351
rect 29444 27344 29453 27384
rect 33829 27344 33830 27384
rect 29444 27343 29502 27344
rect 9493 27300 9535 27309
rect 9668 27300 9726 27301
rect 10741 27300 10783 27309
rect 11701 27300 11743 27309
rect 11972 27300 12030 27301
rect 12565 27300 12607 27309
rect 14276 27300 14334 27301
rect 16772 27300 16830 27301
rect 18901 27300 18943 27309
rect 19861 27300 19903 27309
rect 20069 27300 20127 27301
rect 20250 27300 20292 27309
rect 20354 27300 20412 27301
rect 20612 27300 20670 27301
rect 20802 27300 20860 27301
rect 21123 27300 21165 27309
rect 21668 27300 21726 27301
rect 23893 27300 23935 27309
rect 24068 27300 24126 27301
rect 24757 27300 24799 27309
rect 25457 27302 25458 27342
rect 33829 27335 33871 27344
rect 9493 27260 9494 27300
rect 9668 27260 9677 27300
rect 10252 27291 10298 27300
rect 9493 27251 9535 27260
rect 9668 27259 9726 27260
rect 10252 27251 10253 27291
rect 10741 27260 10742 27300
rect 11701 27260 11702 27300
rect 11972 27260 11981 27300
rect 12565 27260 12566 27300
rect 14276 27260 14285 27300
rect 16772 27260 16781 27300
rect 18901 27260 18902 27300
rect 19861 27260 19862 27300
rect 20069 27260 20078 27300
rect 20250 27260 20251 27300
rect 20354 27260 20363 27300
rect 20485 27289 20527 27298
rect 10741 27251 10783 27260
rect 11701 27251 11743 27260
rect 11972 27259 12030 27260
rect 12565 27251 12607 27260
rect 14276 27259 14334 27260
rect 16772 27259 16830 27260
rect 13748 27258 13806 27259
rect 10252 27242 10298 27251
rect 8245 27216 8287 27225
rect 13748 27218 13757 27258
rect 18901 27251 18943 27260
rect 19861 27251 19903 27260
rect 20069 27259 20127 27260
rect 20250 27251 20292 27260
rect 20354 27259 20412 27260
rect 20485 27249 20486 27289
rect 20612 27260 20621 27300
rect 20802 27260 20811 27300
rect 21123 27260 21124 27300
rect 21668 27260 21677 27300
rect 23893 27260 23894 27300
rect 24068 27260 24077 27300
rect 24757 27260 24758 27300
rect 25457 27293 25499 27302
rect 25748 27300 25806 27301
rect 25904 27300 25946 27309
rect 26101 27300 26143 27309
rect 26965 27300 27007 27309
rect 27157 27300 27199 27309
rect 27445 27300 27487 27309
rect 28069 27300 28111 27309
rect 28213 27300 28255 27309
rect 28772 27300 28830 27301
rect 29828 27300 29886 27301
rect 31957 27300 31999 27309
rect 32132 27300 32190 27301
rect 32245 27300 32287 27309
rect 33205 27300 33247 27309
rect 34165 27300 34207 27309
rect 34741 27300 34783 27309
rect 35125 27300 35167 27309
rect 36181 27300 36223 27309
rect 36740 27300 36798 27301
rect 25748 27260 25757 27300
rect 25904 27260 25905 27300
rect 26101 27260 26102 27300
rect 26965 27260 26966 27300
rect 27157 27260 27158 27300
rect 27445 27260 27446 27300
rect 28069 27260 28070 27300
rect 28213 27260 28214 27300
rect 28772 27260 28781 27300
rect 29828 27260 29837 27300
rect 31957 27260 31958 27300
rect 32132 27260 32141 27300
rect 32245 27260 32246 27300
rect 32428 27291 32474 27300
rect 20612 27259 20670 27260
rect 20802 27259 20860 27260
rect 21123 27251 21165 27260
rect 21668 27259 21726 27260
rect 23893 27251 23935 27260
rect 24068 27259 24126 27260
rect 24757 27251 24799 27260
rect 25748 27259 25806 27260
rect 25904 27251 25946 27260
rect 26101 27251 26143 27260
rect 26965 27251 27007 27260
rect 27157 27251 27199 27260
rect 27445 27251 27487 27260
rect 28069 27251 28111 27260
rect 28213 27251 28255 27260
rect 28772 27259 28830 27260
rect 29828 27259 29886 27260
rect 31957 27251 31999 27260
rect 32132 27259 32190 27260
rect 32245 27251 32287 27260
rect 32428 27251 32429 27291
rect 33205 27260 33206 27300
rect 33676 27291 33722 27300
rect 33205 27251 33247 27260
rect 33676 27251 33677 27291
rect 34165 27260 34166 27300
rect 34293 27276 34335 27285
rect 34165 27251 34207 27260
rect 20485 27240 20527 27249
rect 32428 27242 32474 27251
rect 33676 27242 33722 27251
rect 34293 27236 34294 27276
rect 34741 27260 34742 27300
rect 35125 27260 35126 27300
rect 36181 27260 36182 27300
rect 36740 27260 36749 27300
rect 34741 27251 34783 27260
rect 35125 27251 35167 27260
rect 36181 27251 36223 27260
rect 36740 27259 36798 27260
rect 34293 27227 34335 27236
rect 13748 27217 13806 27218
rect 13556 27216 13614 27217
rect 25621 27216 25663 27225
rect 33115 27216 33157 27225
rect 36373 27216 36415 27225
rect 8245 27176 8246 27216
rect 13556 27176 13565 27216
rect 14189 27176 14198 27216
rect 22253 27176 22262 27216
rect 25621 27176 25622 27216
rect 33115 27176 33116 27216
rect 36373 27176 36374 27216
rect 36557 27176 36566 27216
rect 8245 27167 8287 27176
rect 13556 27175 13614 27176
rect 25621 27167 25663 27176
rect 33115 27167 33157 27176
rect 36373 27167 36415 27176
rect 8005 27132 8047 27141
rect 8917 27132 8959 27141
rect 9301 27132 9343 27141
rect 9668 27132 9726 27133
rect 23605 27132 23647 27141
rect 24949 27132 24991 27141
rect 26005 27132 26047 27141
rect 27781 27132 27823 27141
rect 31765 27132 31807 27141
rect 32245 27132 32287 27141
rect 35509 27132 35551 27141
rect 8005 27092 8006 27132
rect 8917 27092 8918 27132
rect 9301 27092 9302 27132
rect 9668 27092 9677 27132
rect 23605 27092 23606 27132
rect 24949 27092 24950 27132
rect 26005 27092 26006 27132
rect 27781 27092 27782 27132
rect 31765 27092 31766 27132
rect 32245 27092 32246 27132
rect 35509 27092 35510 27132
rect 8005 27083 8047 27092
rect 8917 27083 8959 27092
rect 9301 27083 9343 27092
rect 9668 27091 9726 27092
rect 23605 27083 23647 27092
rect 24949 27083 24991 27092
rect 26005 27083 26047 27092
rect 27781 27083 27823 27092
rect 31765 27083 31807 27092
rect 32245 27083 32287 27092
rect 35509 27083 35551 27092
rect 13237 27048 13279 27057
rect 29173 27048 29215 27057
rect 13237 27008 13238 27048
rect 29173 27008 29174 27048
rect 13237 26999 13279 27008
rect 29173 26999 29215 27008
rect 12949 26712 12991 26721
rect 15236 26712 15294 26713
rect 16261 26712 16303 26721
rect 28484 26712 28542 26713
rect 34261 26712 34303 26721
rect 35509 26712 35551 26721
rect 12949 26672 12950 26712
rect 15236 26672 15245 26712
rect 16261 26672 16262 26712
rect 28484 26672 28493 26712
rect 34261 26672 34262 26712
rect 35509 26672 35510 26712
rect 12949 26663 12991 26672
rect 15236 26671 15294 26672
rect 16261 26663 16303 26672
rect 28484 26671 28542 26672
rect 34261 26663 34303 26672
rect 35509 26663 35551 26672
rect 9013 26628 9055 26637
rect 9781 26628 9823 26637
rect 16597 26628 16639 26637
rect 18181 26628 18223 26637
rect 18997 26628 19039 26637
rect 21589 26628 21631 26637
rect 22165 26628 22207 26637
rect 26101 26628 26143 26637
rect 32629 26628 32671 26637
rect 33781 26628 33823 26637
rect 38389 26628 38431 26637
rect 9013 26588 9014 26628
rect 9781 26588 9782 26628
rect 15013 26619 15055 26628
rect 9013 26579 9055 26588
rect 9781 26579 9823 26588
rect 15013 26579 15014 26619
rect 16597 26588 16598 26628
rect 18181 26588 18182 26628
rect 18997 26588 18998 26628
rect 21589 26588 21590 26628
rect 22165 26588 22166 26628
rect 26101 26588 26102 26628
rect 32629 26588 32630 26628
rect 33077 26619 33119 26628
rect 16597 26579 16639 26588
rect 18181 26579 18223 26588
rect 18997 26579 19039 26588
rect 21589 26579 21631 26588
rect 22165 26579 22207 26588
rect 26101 26579 26143 26588
rect 32629 26579 32671 26588
rect 33077 26579 33078 26619
rect 33781 26588 33782 26628
rect 38389 26588 38390 26628
rect 33781 26579 33823 26588
rect 38389 26579 38431 26588
rect 15013 26570 15055 26579
rect 33077 26570 33119 26579
rect 8053 26544 8095 26553
rect 8629 26544 8671 26553
rect 10052 26544 10110 26545
rect 10453 26544 10495 26553
rect 16021 26544 16063 26553
rect 16981 26544 17023 26553
rect 21253 26544 21295 26553
rect 22069 26544 22111 26553
rect 23797 26544 23839 26553
rect 32725 26544 32767 26553
rect 34741 26544 34783 26553
rect 8053 26504 8054 26544
rect 8629 26504 8630 26544
rect 10052 26504 10061 26544
rect 10453 26504 10454 26544
rect 10637 26504 10646 26544
rect 16021 26504 16022 26544
rect 16981 26504 16982 26544
rect 21253 26504 21254 26544
rect 22069 26504 22070 26544
rect 23797 26504 23798 26544
rect 24941 26504 24950 26544
rect 29165 26504 29174 26544
rect 32725 26504 32726 26544
rect 34741 26504 34742 26544
rect 8053 26495 8095 26504
rect 8629 26495 8671 26504
rect 10052 26503 10110 26504
rect 10453 26495 10495 26504
rect 16021 26495 16063 26504
rect 16981 26495 17023 26504
rect 21253 26495 21295 26504
rect 22069 26495 22111 26504
rect 23797 26495 23839 26504
rect 32725 26495 32767 26504
rect 34741 26495 34783 26504
rect 19706 26471 19748 26480
rect 9205 26460 9247 26469
rect 9397 26460 9439 26469
rect 9920 26460 9962 26469
rect 10150 26460 10208 26461
rect 10820 26460 10878 26461
rect 13621 26460 13663 26469
rect 13909 26460 13951 26469
rect 14293 26460 14335 26469
rect 14677 26460 14719 26469
rect 15044 26460 15102 26461
rect 15737 26460 15795 26461
rect 17348 26460 17406 26461
rect 17749 26460 17791 26469
rect 18037 26460 18079 26469
rect 18260 26460 18318 26461
rect 18805 26460 18847 26469
rect 18920 26460 18962 26469
rect 19093 26460 19135 26469
rect 19313 26460 19371 26461
rect 19460 26460 19518 26461
rect 19585 26460 19627 26469
rect 9205 26420 9206 26460
rect 9397 26420 9398 26460
rect 9920 26420 9921 26460
rect 10150 26420 10159 26460
rect 10820 26420 10829 26460
rect 13333 26451 13375 26460
rect 9205 26411 9247 26420
rect 9397 26411 9439 26420
rect 9920 26411 9962 26420
rect 10150 26419 10208 26420
rect 10820 26419 10878 26420
rect 13333 26411 13334 26451
rect 13621 26420 13622 26460
rect 13909 26420 13910 26460
rect 14293 26420 14294 26460
rect 14677 26420 14678 26460
rect 15044 26420 15053 26460
rect 15737 26420 15746 26460
rect 17348 26420 17357 26460
rect 17749 26420 17750 26460
rect 18037 26420 18038 26460
rect 18260 26420 18269 26460
rect 18805 26420 18806 26460
rect 18920 26420 18921 26460
rect 19093 26420 19094 26460
rect 19313 26420 19322 26460
rect 19460 26420 19469 26460
rect 19585 26420 19586 26460
rect 19706 26431 19707 26471
rect 19844 26460 19902 26461
rect 20146 26460 20188 26469
rect 20263 26460 20321 26461
rect 20389 26460 20431 26469
rect 20609 26460 20667 26461
rect 21059 26460 21117 26461
rect 21925 26460 21967 26469
rect 22240 26460 22282 26469
rect 22388 26460 22446 26461
rect 23221 26460 23263 26469
rect 23396 26460 23438 26469
rect 23605 26460 23647 26469
rect 24164 26460 24222 26461
rect 26389 26460 26431 26469
rect 27253 26460 27295 26469
rect 27541 26460 27583 26469
rect 27956 26460 28014 26461
rect 28781 26460 28839 26461
rect 29348 26460 29406 26461
rect 32149 26460 32191 26469
rect 32389 26460 32431 26469
rect 32846 26460 32888 26469
rect 33092 26460 33150 26461
rect 33493 26460 33535 26469
rect 33668 26460 33726 26461
rect 33781 26460 33823 26469
rect 33956 26460 34014 26461
rect 34400 26460 34442 26469
rect 34532 26460 34590 26461
rect 34645 26460 34687 26469
rect 34916 26460 34974 26461
rect 36181 26460 36223 26469
rect 37045 26460 37087 26469
rect 37909 26460 37951 26469
rect 38197 26460 38239 26469
rect 19706 26422 19748 26431
rect 19844 26420 19853 26460
rect 20146 26420 20147 26460
rect 20263 26420 20272 26460
rect 20389 26420 20390 26460
rect 20609 26420 20618 26460
rect 21059 26420 21068 26460
rect 21925 26420 21926 26460
rect 22240 26420 22241 26460
rect 22388 26420 22397 26460
rect 23221 26420 23222 26460
rect 23396 26420 23397 26460
rect 23605 26420 23606 26460
rect 24164 26420 24173 26460
rect 26389 26420 26390 26460
rect 27253 26420 27254 26460
rect 27541 26420 27542 26460
rect 27956 26420 27965 26460
rect 28781 26420 28790 26460
rect 29348 26420 29357 26460
rect 32149 26420 32150 26460
rect 32389 26420 32390 26460
rect 13621 26411 13663 26420
rect 13909 26411 13951 26420
rect 14293 26411 14335 26420
rect 14677 26411 14719 26420
rect 15044 26419 15102 26420
rect 15737 26419 15795 26420
rect 17348 26419 17406 26420
rect 17749 26411 17791 26420
rect 18037 26411 18079 26420
rect 18260 26419 18318 26420
rect 18805 26411 18847 26420
rect 18920 26411 18962 26420
rect 19093 26411 19135 26420
rect 19313 26419 19371 26420
rect 19460 26419 19518 26420
rect 19585 26411 19627 26420
rect 19844 26419 19902 26420
rect 20146 26411 20188 26420
rect 20263 26419 20321 26420
rect 20389 26411 20431 26420
rect 20609 26419 20667 26420
rect 21059 26419 21117 26420
rect 21925 26411 21967 26420
rect 22240 26411 22282 26420
rect 22388 26419 22446 26420
rect 23221 26411 23263 26420
rect 23396 26411 23438 26420
rect 23605 26411 23647 26420
rect 24164 26419 24222 26420
rect 26389 26411 26431 26420
rect 27253 26411 27295 26420
rect 27541 26411 27583 26420
rect 27956 26419 28014 26420
rect 28781 26419 28839 26420
rect 29348 26419 29406 26420
rect 32149 26411 32191 26420
rect 32389 26411 32431 26420
rect 32561 26418 32603 26427
rect 32846 26420 32847 26460
rect 33092 26420 33101 26460
rect 33493 26420 33494 26460
rect 33668 26420 33677 26460
rect 33781 26420 33782 26460
rect 33956 26420 33965 26460
rect 34400 26420 34401 26460
rect 34532 26420 34541 26460
rect 34645 26420 34646 26460
rect 34916 26420 34925 26460
rect 36181 26420 36182 26460
rect 37045 26420 37046 26460
rect 37909 26420 37910 26460
rect 38197 26420 38198 26460
rect 13333 26402 13375 26411
rect 8293 26376 8335 26385
rect 13237 26376 13279 26385
rect 15572 26376 15630 26377
rect 16741 26376 16783 26385
rect 19844 26376 19902 26377
rect 28487 26376 28529 26385
rect 32561 26378 32562 26418
rect 32846 26411 32888 26420
rect 33092 26419 33150 26420
rect 33493 26411 33535 26420
rect 33668 26419 33726 26420
rect 33781 26411 33823 26420
rect 33956 26419 34014 26420
rect 34400 26411 34442 26420
rect 34532 26419 34590 26420
rect 34645 26411 34687 26420
rect 34916 26419 34974 26420
rect 36181 26411 36223 26420
rect 37045 26411 37087 26420
rect 37909 26411 37951 26420
rect 38197 26411 38239 26420
rect 28964 26376 29022 26377
rect 8293 26336 8294 26376
rect 13237 26336 13238 26376
rect 15572 26336 15581 26376
rect 16741 26336 16742 26376
rect 19844 26336 19853 26376
rect 28487 26336 28488 26376
rect 28964 26336 28973 26376
rect 32561 26369 32603 26378
rect 34069 26376 34111 26385
rect 34272 26376 34314 26385
rect 35232 26376 35274 26385
rect 36356 26376 36414 26377
rect 34069 26336 34070 26376
rect 34272 26336 34273 26376
rect 35232 26336 35233 26376
rect 36356 26336 36365 26376
rect 8293 26327 8335 26336
rect 13237 26327 13279 26336
rect 15572 26335 15630 26336
rect 16741 26327 16783 26336
rect 19844 26335 19902 26336
rect 28487 26327 28529 26336
rect 28964 26335 29022 26336
rect 34069 26327 34111 26336
rect 34272 26327 34314 26336
rect 35232 26327 35274 26336
rect 36356 26335 36414 26336
rect 8389 26292 8431 26301
rect 9380 26292 9438 26293
rect 10244 26292 10302 26293
rect 12757 26292 12799 26301
rect 14389 26292 14431 26301
rect 15236 26292 15294 26293
rect 18469 26292 18511 26301
rect 20437 26292 20479 26301
rect 20773 26292 20815 26301
rect 22549 26292 22591 26301
rect 23588 26292 23646 26293
rect 27061 26292 27103 26301
rect 27733 26292 27775 26301
rect 28165 26292 28207 26301
rect 28693 26292 28735 26301
rect 31285 26292 31327 26301
rect 31477 26292 31519 26301
rect 33284 26292 33342 26293
rect 35012 26292 35070 26293
rect 35125 26292 35167 26301
rect 37237 26292 37279 26301
rect 38084 26292 38142 26293
rect 8389 26252 8390 26292
rect 9380 26252 9389 26292
rect 10244 26252 10253 26292
rect 12757 26252 12758 26292
rect 14389 26252 14390 26292
rect 15236 26252 15245 26292
rect 18469 26252 18470 26292
rect 20437 26252 20438 26292
rect 20773 26252 20774 26292
rect 22549 26252 22550 26292
rect 23588 26252 23597 26292
rect 27061 26252 27062 26292
rect 27733 26252 27734 26292
rect 28165 26252 28166 26292
rect 28693 26252 28694 26292
rect 31285 26252 31286 26292
rect 31477 26252 31478 26292
rect 33284 26252 33293 26292
rect 35012 26252 35021 26292
rect 35125 26252 35126 26292
rect 37237 26252 37238 26292
rect 38084 26252 38093 26292
rect 8389 26243 8431 26252
rect 9380 26251 9438 26252
rect 10244 26251 10302 26252
rect 12757 26243 12799 26252
rect 14389 26243 14431 26252
rect 15236 26251 15294 26252
rect 18469 26243 18511 26252
rect 20437 26243 20479 26252
rect 20773 26243 20815 26252
rect 22549 26243 22591 26252
rect 23588 26251 23646 26252
rect 27061 26243 27103 26252
rect 27733 26243 27775 26252
rect 28165 26243 28207 26252
rect 28693 26243 28735 26252
rect 31285 26243 31327 26252
rect 31477 26243 31519 26252
rect 33284 26251 33342 26252
rect 35012 26251 35070 26252
rect 35125 26243 35167 26252
rect 37237 26243 37279 26252
rect 38084 26251 38142 26252
rect 9109 25956 9151 25965
rect 32612 25956 32670 25957
rect 33973 25956 34015 25965
rect 38677 25956 38719 25965
rect 9109 25916 9110 25956
rect 32612 25916 32621 25956
rect 33973 25916 33974 25956
rect 38677 25916 38678 25956
rect 9109 25907 9151 25916
rect 32612 25915 32670 25916
rect 33973 25907 34015 25916
rect 38677 25907 38719 25916
rect 9284 25872 9342 25873
rect 13508 25872 13566 25873
rect 35015 25872 35057 25881
rect 35221 25872 35263 25881
rect 9284 25832 9293 25872
rect 13508 25832 13517 25872
rect 35015 25832 35016 25872
rect 35221 25832 35222 25872
rect 9284 25831 9342 25832
rect 13508 25831 13566 25832
rect 35015 25823 35057 25832
rect 35221 25823 35263 25832
rect 9668 25788 9726 25789
rect 11797 25788 11839 25797
rect 32053 25788 32095 25797
rect 32288 25788 32330 25797
rect 32533 25788 32575 25797
rect 33301 25788 33343 25797
rect 33418 25788 33476 25789
rect 33589 25788 33631 25797
rect 33770 25788 33812 25797
rect 34309 25788 34351 25797
rect 34539 25788 34581 25797
rect 34724 25788 34782 25789
rect 34837 25788 34879 25797
rect 35509 25788 35551 25797
rect 36740 25788 36798 25789
rect 9668 25748 9677 25788
rect 11797 25748 11798 25788
rect 32053 25748 32054 25788
rect 32288 25748 32289 25788
rect 32533 25748 32534 25788
rect 32812 25779 32858 25788
rect 9668 25747 9726 25748
rect 11797 25739 11839 25748
rect 32053 25739 32095 25748
rect 32288 25739 32330 25748
rect 32533 25739 32575 25748
rect 32812 25739 32813 25779
rect 33301 25748 33302 25788
rect 33418 25748 33427 25788
rect 33589 25748 33590 25788
rect 33770 25748 33771 25788
rect 34069 25779 34111 25788
rect 33301 25739 33343 25748
rect 33418 25747 33476 25748
rect 33589 25739 33631 25748
rect 33770 25739 33812 25748
rect 34069 25739 34070 25779
rect 34309 25748 34310 25788
rect 34539 25748 34540 25788
rect 34724 25748 34733 25788
rect 34837 25748 34838 25788
rect 35317 25779 35359 25788
rect 34309 25739 34351 25748
rect 34539 25739 34581 25748
rect 34724 25747 34782 25748
rect 34837 25739 34879 25748
rect 35317 25739 35318 25779
rect 35509 25748 35510 25788
rect 36740 25748 36749 25788
rect 35509 25739 35551 25748
rect 36740 25747 36798 25748
rect 32812 25730 32858 25739
rect 34069 25730 34111 25739
rect 35317 25730 35359 25739
rect 8725 25704 8767 25713
rect 32197 25704 32239 25713
rect 32420 25704 32478 25705
rect 32965 25704 33007 25713
rect 36373 25704 36415 25713
rect 8725 25664 8726 25704
rect 32197 25664 32198 25704
rect 32420 25664 32429 25704
rect 32965 25664 32966 25704
rect 36373 25664 36374 25704
rect 37133 25664 37142 25704
rect 8725 25655 8767 25664
rect 32197 25655 32239 25664
rect 32420 25663 32478 25664
rect 32965 25655 33007 25664
rect 36373 25655 36415 25664
rect 8341 25620 8383 25629
rect 11605 25620 11647 25629
rect 12949 25620 12991 25629
rect 13333 25620 13375 25629
rect 33493 25620 33535 25629
rect 34213 25620 34255 25629
rect 34837 25620 34879 25629
rect 8341 25580 8342 25620
rect 11605 25580 11606 25620
rect 12949 25580 12950 25620
rect 13333 25580 13334 25620
rect 33493 25580 33494 25620
rect 34213 25580 34214 25620
rect 34837 25580 34838 25620
rect 8341 25571 8383 25580
rect 11605 25571 11647 25580
rect 12949 25571 12991 25580
rect 13333 25571 13375 25580
rect 33493 25571 33535 25580
rect 34213 25571 34255 25580
rect 34837 25571 34879 25580
rect 8485 25536 8527 25545
rect 12469 25536 12511 25545
rect 13909 25536 13951 25545
rect 33764 25536 33822 25537
rect 35012 25536 35070 25537
rect 36181 25536 36223 25545
rect 8485 25496 8486 25536
rect 12469 25496 12470 25536
rect 13909 25496 13910 25536
rect 33764 25496 33773 25536
rect 35012 25496 35021 25536
rect 36181 25496 36182 25536
rect 8485 25487 8527 25496
rect 12469 25487 12511 25496
rect 13909 25487 13951 25496
rect 33764 25495 33822 25496
rect 35012 25495 35070 25496
rect 36181 25487 36223 25496
rect 8437 25200 8479 25209
rect 11989 25200 12031 25209
rect 13573 25200 13615 25209
rect 32869 25200 32911 25209
rect 35509 25200 35551 25209
rect 8437 25160 8438 25200
rect 11989 25160 11990 25200
rect 13573 25160 13574 25200
rect 32869 25160 32870 25200
rect 35509 25160 35510 25200
rect 8437 25151 8479 25160
rect 11989 25151 12031 25160
rect 13573 25151 13615 25160
rect 32869 25151 32911 25160
rect 35509 25151 35551 25160
rect 34645 25116 34687 25125
rect 34645 25076 34646 25116
rect 34645 25067 34687 25076
rect 36373 25032 36415 25041
rect 8909 24992 8918 25032
rect 36373 24992 36374 25032
rect 37613 24992 37622 25032
rect 36373 24983 36415 24992
rect 9956 24948 10014 24949
rect 11509 24948 11551 24957
rect 11797 24948 11839 24957
rect 12661 24948 12703 24957
rect 12949 24948 12991 24957
rect 13333 24948 13375 24957
rect 14039 24948 14068 24949
rect 32101 24948 32159 24949
rect 32245 24948 32287 24957
rect 32480 24948 32522 24957
rect 32725 24948 32767 24957
rect 33013 24948 33055 24957
rect 33248 24948 33290 24957
rect 33493 24948 33535 24957
rect 33860 24948 33918 24949
rect 34176 24948 34218 24957
rect 34340 24948 34398 24949
rect 34645 24948 34687 24957
rect 35029 24948 35071 24957
rect 35173 24948 35215 24957
rect 36181 24948 36223 24957
rect 36740 24948 36798 24949
rect 9956 24908 9965 24948
rect 11509 24908 11510 24948
rect 11797 24908 11798 24948
rect 12373 24939 12415 24948
rect 9956 24907 10014 24908
rect 11509 24899 11551 24908
rect 11797 24899 11839 24908
rect 12373 24899 12374 24939
rect 12661 24908 12662 24948
rect 12949 24908 12950 24948
rect 13333 24908 13334 24948
rect 14039 24908 14048 24948
rect 32101 24908 32110 24948
rect 32245 24908 32246 24948
rect 32480 24908 32481 24948
rect 32620 24939 32666 24948
rect 12661 24899 12703 24908
rect 12949 24899 12991 24908
rect 13333 24899 13375 24908
rect 14039 24907 14068 24908
rect 32101 24907 32159 24908
rect 32245 24899 32287 24908
rect 32480 24899 32522 24908
rect 32620 24899 32621 24939
rect 32725 24908 32726 24948
rect 33013 24908 33014 24948
rect 33248 24908 33249 24948
rect 33388 24939 33434 24948
rect 32725 24899 32767 24908
rect 33013 24899 33055 24908
rect 33248 24899 33290 24908
rect 33388 24899 33389 24939
rect 33493 24908 33494 24948
rect 33860 24908 33869 24948
rect 34176 24908 34177 24948
rect 34340 24908 34349 24948
rect 34645 24908 34646 24948
rect 35029 24908 35030 24948
rect 35173 24908 35174 24948
rect 36181 24908 36182 24948
rect 36740 24908 36749 24948
rect 33493 24899 33535 24908
rect 33860 24907 33918 24908
rect 34176 24899 34218 24908
rect 34340 24907 34398 24908
rect 34645 24899 34687 24908
rect 35029 24899 35071 24908
rect 35173 24899 35215 24908
rect 36181 24899 36223 24908
rect 36740 24907 36798 24908
rect 12373 24890 12415 24899
rect 32620 24890 32666 24899
rect 33388 24890 33434 24899
rect 8036 24864 8094 24865
rect 10340 24864 10398 24865
rect 10820 24864 10878 24865
rect 12277 24864 12319 24873
rect 13844 24864 13902 24865
rect 34820 24864 34878 24865
rect 8036 24824 8045 24864
rect 10340 24824 10349 24864
rect 10820 24824 10829 24864
rect 12277 24824 12278 24864
rect 13844 24824 13853 24864
rect 34820 24824 34829 24864
rect 8036 24823 8094 24824
rect 10340 24823 10398 24824
rect 10820 24823 10878 24824
rect 12277 24815 12319 24824
rect 13844 24823 13902 24824
rect 34820 24823 34878 24824
rect 11653 24780 11695 24789
rect 32437 24780 32479 24789
rect 33205 24780 33247 24789
rect 33956 24780 34014 24781
rect 34069 24780 34111 24789
rect 35125 24780 35167 24789
rect 38677 24780 38719 24789
rect 11653 24740 11654 24780
rect 32437 24740 32438 24780
rect 33205 24740 33206 24780
rect 33956 24740 33965 24780
rect 34069 24740 34070 24780
rect 35125 24740 35126 24780
rect 38677 24740 38678 24780
rect 11653 24731 11695 24740
rect 32437 24731 32479 24740
rect 33205 24731 33247 24740
rect 33956 24739 34014 24740
rect 34069 24731 34111 24740
rect 35125 24731 35167 24740
rect 38677 24731 38719 24740
rect 9092 24444 9150 24445
rect 10964 24444 11022 24445
rect 11396 24444 11454 24445
rect 11509 24444 11551 24453
rect 12181 24444 12223 24453
rect 12469 24444 12511 24453
rect 13028 24444 13086 24445
rect 35893 24444 35935 24453
rect 9092 24404 9101 24444
rect 10964 24404 10973 24444
rect 11396 24404 11405 24444
rect 11509 24404 11510 24444
rect 12181 24404 12182 24444
rect 12469 24404 12470 24444
rect 13028 24404 13037 24444
rect 35893 24404 35894 24444
rect 9092 24403 9150 24404
rect 10964 24403 11022 24404
rect 11396 24403 11454 24404
rect 11509 24395 11551 24404
rect 12181 24395 12223 24404
rect 12469 24395 12511 24404
rect 13028 24403 13086 24404
rect 35893 24395 35935 24404
rect 9572 24360 9630 24361
rect 9685 24360 9727 24369
rect 10645 24360 10687 24369
rect 12068 24360 12126 24361
rect 12935 24360 12977 24369
rect 13508 24360 13566 24361
rect 32533 24360 32575 24369
rect 34357 24360 34399 24369
rect 9572 24320 9581 24360
rect 9685 24320 9686 24360
rect 10645 24320 10646 24360
rect 12068 24320 12077 24360
rect 12935 24320 12936 24360
rect 13508 24320 13517 24360
rect 32533 24320 32534 24360
rect 33196 24351 33242 24360
rect 9572 24319 9630 24320
rect 9685 24311 9727 24320
rect 10645 24311 10687 24320
rect 12068 24319 12126 24320
rect 12935 24311 12977 24320
rect 13508 24319 13566 24320
rect 32533 24311 32575 24320
rect 33196 24311 33197 24351
rect 34357 24320 34358 24360
rect 34357 24311 34399 24320
rect 33196 24302 33242 24311
rect 8245 24276 8287 24285
rect 8420 24276 8478 24277
rect 8629 24276 8671 24285
rect 8804 24276 8862 24277
rect 8996 24276 9054 24277
rect 9315 24276 9357 24285
rect 9482 24276 9524 24285
rect 9973 24276 10015 24285
rect 11129 24276 11187 24277
rect 11306 24276 11348 24285
rect 11975 24276 12017 24285
rect 12565 24276 12607 24285
rect 12794 24276 12852 24277
rect 13141 24276 13183 24285
rect 32228 24276 32286 24277
rect 32900 24276 32958 24277
rect 33284 24276 33342 24277
rect 33461 24276 33519 24277
rect 33860 24276 33918 24277
rect 34052 24276 34110 24277
rect 34165 24276 34207 24285
rect 34604 24276 34662 24277
rect 34837 24276 34879 24285
rect 35446 24276 35504 24277
rect 35605 24276 35647 24285
rect 36757 24276 36799 24285
rect 36949 24276 36991 24285
rect 37796 24276 37854 24277
rect 38485 24276 38527 24285
rect 8245 24236 8246 24276
rect 8420 24236 8429 24276
rect 8629 24236 8630 24276
rect 8804 24236 8813 24276
rect 8996 24236 9005 24276
rect 9315 24236 9316 24276
rect 9482 24236 9483 24276
rect 9781 24267 9823 24276
rect 8245 24227 8287 24236
rect 8420 24235 8478 24236
rect 8629 24227 8671 24236
rect 8804 24235 8862 24236
rect 8996 24235 9054 24236
rect 9315 24227 9357 24236
rect 9482 24227 9524 24236
rect 9781 24227 9782 24267
rect 9973 24236 9974 24276
rect 11129 24236 11138 24276
rect 11306 24236 11307 24276
rect 11605 24267 11647 24276
rect 9973 24227 10015 24236
rect 11129 24235 11187 24236
rect 11306 24227 11348 24236
rect 11605 24227 11606 24267
rect 11975 24236 11976 24276
rect 12277 24267 12319 24276
rect 11975 24227 12017 24236
rect 12277 24227 12278 24267
rect 12565 24236 12566 24276
rect 12794 24236 12803 24276
rect 13141 24236 13142 24276
rect 13237 24267 13279 24276
rect 12565 24227 12607 24236
rect 12794 24235 12852 24236
rect 13141 24227 13183 24236
rect 13237 24227 13238 24267
rect 32228 24236 32237 24276
rect 32900 24236 32909 24276
rect 33013 24267 33055 24276
rect 32228 24235 32286 24236
rect 32900 24235 32958 24236
rect 33013 24227 33014 24267
rect 33284 24236 33293 24276
rect 33461 24236 33470 24276
rect 33860 24236 33869 24276
rect 34052 24236 34061 24276
rect 34165 24236 34166 24276
rect 34470 24261 34512 24270
rect 33284 24235 33342 24236
rect 33461 24235 33519 24236
rect 33860 24235 33918 24236
rect 34052 24235 34110 24236
rect 34165 24227 34207 24236
rect 9781 24218 9823 24227
rect 11605 24218 11647 24227
rect 12277 24218 12319 24227
rect 13237 24218 13279 24227
rect 33013 24218 33055 24227
rect 34470 24221 34471 24261
rect 34604 24236 34613 24276
rect 34837 24236 34838 24276
rect 35446 24236 35455 24276
rect 35605 24236 35606 24276
rect 35739 24244 35797 24245
rect 34604 24235 34662 24236
rect 34837 24227 34879 24236
rect 35446 24235 35504 24236
rect 35605 24227 35647 24236
rect 34470 24212 34512 24221
rect 35739 24204 35748 24244
rect 36757 24236 36758 24276
rect 36949 24236 36950 24276
rect 37796 24236 37805 24276
rect 38485 24236 38486 24276
rect 36757 24227 36799 24236
rect 36949 24227 36991 24236
rect 37796 24235 37854 24236
rect 38485 24227 38527 24236
rect 35739 24203 35797 24204
rect 12469 24192 12511 24201
rect 12684 24192 12726 24201
rect 32053 24192 32095 24201
rect 32629 24192 32671 24201
rect 34724 24192 34782 24193
rect 34933 24192 34975 24201
rect 35252 24192 35310 24193
rect 12469 24152 12470 24192
rect 12684 24152 12685 24192
rect 32053 24152 32054 24192
rect 32629 24152 32630 24192
rect 34724 24152 34733 24192
rect 34933 24152 34934 24192
rect 35252 24152 35261 24192
rect 12469 24143 12511 24152
rect 12684 24143 12726 24152
rect 32053 24143 32095 24152
rect 32629 24143 32671 24152
rect 34724 24151 34782 24152
rect 34933 24143 34975 24152
rect 35252 24151 35310 24152
rect 8420 24108 8478 24109
rect 8804 24108 8862 24109
rect 8420 24068 8429 24108
rect 8804 24068 8813 24108
rect 8420 24067 8478 24068
rect 8804 24067 8862 24068
rect 9301 24024 9343 24033
rect 32900 24024 32958 24025
rect 36085 24024 36127 24033
rect 37621 24024 37663 24033
rect 9301 23984 9302 24024
rect 32900 23984 32909 24024
rect 36085 23984 36086 24024
rect 37621 23984 37622 24024
rect 9301 23975 9343 23984
rect 32900 23983 32958 23984
rect 36085 23975 36127 23984
rect 37621 23975 37663 23984
rect 13412 23688 13470 23689
rect 33301 23688 33343 23697
rect 34549 23688 34591 23697
rect 35125 23688 35167 23697
rect 13412 23648 13421 23688
rect 33301 23648 33302 23688
rect 34549 23648 34550 23688
rect 35125 23648 35126 23688
rect 13412 23647 13470 23648
rect 33301 23639 33343 23648
rect 34549 23639 34591 23648
rect 35125 23639 35167 23648
rect 36757 23604 36799 23613
rect 36757 23564 36758 23604
rect 36757 23555 36799 23564
rect 9781 23520 9823 23529
rect 11156 23520 11214 23521
rect 11509 23520 11551 23529
rect 12757 23520 12799 23529
rect 13237 23520 13279 23529
rect 32900 23520 32958 23521
rect 35227 23520 35269 23529
rect 38660 23520 38718 23521
rect 9781 23480 9782 23520
rect 10012 23511 10058 23520
rect 9781 23471 9823 23480
rect 10012 23471 10013 23511
rect 11156 23480 11165 23520
rect 11509 23480 11510 23520
rect 11740 23511 11786 23520
rect 11156 23479 11214 23480
rect 11509 23471 11551 23480
rect 11740 23471 11741 23511
rect 12757 23480 12758 23520
rect 13237 23480 13238 23520
rect 12757 23471 12799 23480
rect 13237 23471 13279 23480
rect 13861 23478 13903 23487
rect 32900 23480 32909 23520
rect 35227 23480 35228 23520
rect 37805 23480 37814 23520
rect 38660 23480 38669 23520
rect 32900 23479 32958 23480
rect 33908 23478 33966 23479
rect 10012 23462 10058 23471
rect 11740 23462 11786 23471
rect 13707 23469 13765 23470
rect 9109 23436 9151 23445
rect 9284 23436 9342 23437
rect 9600 23436 9642 23445
rect 9877 23436 9919 23445
rect 10106 23436 10164 23437
rect 10693 23436 10751 23437
rect 10837 23436 10879 23445
rect 11321 23436 11379 23437
rect 11605 23436 11647 23445
rect 11834 23436 11892 23437
rect 12181 23436 12223 23445
rect 12373 23436 12415 23445
rect 12896 23436 12938 23445
rect 13028 23436 13086 23437
rect 13141 23436 13183 23445
rect 9109 23396 9110 23436
rect 9284 23396 9293 23436
rect 9600 23396 9601 23436
rect 9877 23396 9878 23436
rect 10106 23396 10115 23436
rect 10693 23396 10702 23436
rect 10837 23396 10838 23436
rect 11321 23396 11330 23436
rect 11605 23396 11606 23436
rect 11834 23396 11843 23436
rect 12181 23396 12182 23436
rect 12373 23396 12374 23436
rect 12896 23396 12897 23436
rect 13028 23396 13037 23436
rect 13141 23396 13142 23436
rect 13707 23429 13716 23469
rect 13861 23438 13862 23478
rect 13861 23429 13903 23438
rect 13988 23436 14046 23437
rect 32043 23436 32085 23445
rect 32228 23436 32286 23437
rect 32341 23436 32383 23445
rect 32780 23436 32838 23437
rect 33013 23436 33055 23445
rect 33344 23436 33386 23445
rect 33440 23436 33498 23437
rect 33589 23436 33631 23445
rect 33778 23436 33820 23445
rect 33908 23438 33917 23478
rect 35227 23471 35269 23480
rect 38660 23479 38718 23480
rect 33908 23437 33966 23438
rect 34022 23436 34080 23437
rect 34244 23436 34302 23437
rect 34549 23436 34591 23445
rect 34837 23436 34879 23445
rect 35317 23436 35359 23445
rect 36089 23436 36147 23437
rect 38276 23436 38334 23437
rect 13707 23428 13765 23429
rect 13988 23396 13997 23436
rect 32043 23396 32044 23436
rect 32228 23396 32237 23436
rect 32341 23396 32342 23436
rect 32780 23396 32789 23436
rect 33013 23396 33014 23436
rect 33344 23396 33345 23436
rect 33440 23396 33449 23436
rect 33589 23396 33590 23436
rect 33778 23396 33779 23436
rect 34022 23396 34031 23436
rect 34244 23396 34253 23436
rect 34549 23396 34550 23436
rect 34837 23396 34838 23436
rect 35317 23396 35318 23436
rect 36089 23396 36098 23436
rect 38276 23396 38285 23436
rect 9109 23387 9151 23396
rect 9284 23395 9342 23396
rect 9600 23387 9642 23396
rect 9877 23387 9919 23396
rect 10106 23395 10164 23396
rect 10693 23395 10751 23396
rect 10837 23387 10879 23396
rect 11321 23395 11379 23396
rect 11605 23387 11647 23396
rect 11834 23395 11892 23396
rect 12181 23387 12223 23396
rect 12373 23387 12415 23396
rect 12896 23387 12938 23396
rect 13028 23395 13086 23396
rect 13141 23387 13183 23396
rect 13988 23395 14046 23396
rect 32043 23387 32085 23396
rect 32228 23395 32286 23396
rect 32341 23387 32383 23396
rect 32780 23395 32838 23396
rect 33013 23387 33055 23396
rect 33344 23387 33386 23396
rect 33440 23395 33498 23396
rect 33589 23387 33631 23396
rect 33778 23387 33820 23396
rect 34022 23395 34080 23396
rect 34244 23395 34302 23396
rect 34549 23387 34591 23396
rect 34837 23387 34879 23396
rect 35317 23387 35359 23396
rect 36089 23395 36147 23396
rect 38276 23395 38334 23396
rect 8132 23352 8190 23353
rect 9493 23352 9535 23361
rect 12277 23352 12319 23361
rect 13418 23352 13460 23361
rect 32132 23352 32190 23353
rect 35924 23352 35982 23353
rect 8132 23312 8141 23352
rect 9493 23312 9494 23352
rect 12277 23312 12278 23352
rect 13418 23312 13419 23352
rect 32132 23312 32141 23352
rect 35924 23312 35933 23352
rect 8132 23311 8190 23312
rect 9493 23303 9535 23312
rect 12277 23303 12319 23312
rect 13418 23303 13460 23312
rect 32132 23311 32190 23312
rect 35924 23311 35982 23312
rect 9380 23268 9438 23269
rect 10532 23268 10590 23269
rect 12517 23268 12559 23277
rect 13621 23268 13663 23277
rect 33092 23268 33150 23269
rect 34069 23268 34111 23277
rect 36373 23268 36415 23277
rect 9380 23228 9389 23268
rect 10532 23228 10541 23268
rect 12517 23228 12518 23268
rect 13621 23228 13622 23268
rect 33092 23228 33101 23268
rect 34069 23228 34070 23268
rect 36373 23228 36374 23268
rect 9380 23227 9438 23228
rect 10532 23227 10590 23228
rect 12517 23219 12559 23228
rect 13621 23219 13663 23228
rect 33092 23227 33150 23228
rect 34069 23219 34111 23228
rect 36373 23219 36415 23228
rect 8708 22932 8766 22933
rect 10933 22932 10975 22941
rect 12740 22932 12798 22933
rect 13316 22932 13374 22933
rect 13717 22932 13759 22941
rect 32965 22932 33007 22941
rect 33781 22932 33823 22941
rect 34652 22932 34710 22933
rect 34981 22932 35023 22941
rect 36037 22932 36079 22941
rect 8708 22892 8717 22932
rect 10933 22892 10934 22932
rect 12740 22892 12749 22932
rect 13316 22892 13325 22932
rect 13717 22892 13718 22932
rect 32965 22892 32966 22932
rect 33781 22892 33782 22932
rect 34652 22892 34661 22932
rect 34981 22892 34982 22932
rect 36037 22892 36038 22932
rect 8708 22891 8766 22892
rect 10933 22883 10975 22892
rect 12740 22891 12798 22892
rect 13316 22891 13374 22892
rect 13717 22883 13759 22892
rect 32965 22883 33007 22892
rect 33781 22883 33823 22892
rect 34652 22891 34710 22892
rect 34981 22883 35023 22892
rect 36037 22883 36079 22892
rect 10247 22848 10289 22857
rect 11040 22848 11082 22857
rect 12164 22848 12222 22849
rect 13429 22848 13471 22857
rect 33685 22848 33727 22857
rect 35399 22848 35441 22857
rect 36356 22848 36414 22849
rect 10247 22808 10248 22848
rect 11040 22808 11041 22848
rect 12164 22808 12173 22848
rect 13429 22808 13430 22848
rect 33685 22808 33686 22848
rect 35399 22808 35400 22848
rect 36356 22808 36365 22848
rect 10247 22799 10289 22808
rect 11040 22799 11082 22808
rect 12164 22807 12222 22808
rect 13429 22799 13471 22808
rect 33685 22799 33727 22808
rect 35399 22799 35441 22808
rect 36356 22807 36414 22808
rect 8533 22764 8575 22773
rect 8720 22764 8778 22765
rect 8917 22764 8959 22773
rect 9022 22764 9064 22773
rect 9244 22764 9286 22773
rect 9445 22764 9487 22773
rect 10453 22764 10495 22773
rect 10724 22764 10782 22765
rect 10837 22764 10879 22773
rect 11840 22764 11882 22773
rect 12085 22764 12127 22773
rect 12901 22764 12943 22773
rect 13045 22764 13087 22773
rect 13223 22764 13265 22773
rect 13813 22764 13855 22773
rect 14030 22764 14068 22773
rect 32000 22764 32042 22773
rect 32245 22764 32287 22773
rect 32532 22764 32574 22773
rect 32708 22764 32766 22765
rect 32821 22764 32863 22773
rect 33109 22764 33151 22773
rect 33877 22764 33919 22773
rect 34532 22764 34590 22765
rect 35605 22764 35647 22773
rect 36740 22764 36798 22765
rect 8533 22724 8534 22764
rect 8720 22724 8729 22764
rect 8917 22724 8918 22764
rect 9022 22724 9023 22764
rect 9244 22724 9245 22764
rect 9445 22724 9446 22764
rect 10453 22724 10454 22764
rect 10549 22755 10591 22764
rect 8533 22715 8575 22724
rect 8720 22723 8778 22724
rect 8917 22715 8959 22724
rect 9022 22715 9064 22724
rect 9244 22715 9286 22724
rect 9445 22715 9487 22724
rect 10453 22715 10495 22724
rect 10549 22715 10550 22755
rect 10724 22724 10733 22764
rect 10837 22724 10838 22764
rect 11404 22755 11450 22764
rect 10724 22723 10782 22724
rect 10837 22715 10879 22724
rect 11404 22715 11405 22755
rect 11840 22724 11841 22764
rect 12085 22724 12086 22764
rect 12901 22724 12902 22764
rect 13045 22724 13046 22764
rect 13223 22724 13224 22764
rect 13525 22755 13567 22764
rect 11840 22715 11882 22724
rect 12085 22715 12127 22724
rect 12901 22715 12943 22724
rect 13045 22715 13087 22724
rect 13223 22715 13265 22724
rect 13525 22715 13526 22755
rect 13813 22724 13814 22764
rect 14030 22724 14031 22764
rect 32000 22724 32001 22764
rect 32245 22724 32246 22764
rect 32532 22724 32533 22764
rect 32708 22724 32717 22764
rect 32821 22724 32822 22764
rect 33109 22724 33110 22764
rect 33580 22755 33626 22764
rect 13813 22715 13855 22724
rect 14030 22715 14068 22724
rect 32000 22715 32042 22724
rect 32245 22715 32287 22724
rect 32532 22715 32574 22724
rect 32708 22723 32766 22724
rect 32821 22715 32863 22724
rect 33109 22715 33151 22724
rect 33580 22715 33581 22755
rect 33877 22724 33878 22764
rect 34449 22755 34491 22764
rect 33877 22715 33919 22724
rect 34449 22715 34450 22755
rect 34532 22724 34541 22764
rect 34828 22755 34874 22764
rect 34532 22723 34590 22724
rect 34828 22715 34829 22755
rect 35605 22724 35606 22764
rect 35701 22755 35743 22764
rect 35884 22755 35930 22764
rect 35605 22715 35647 22724
rect 35701 22715 35702 22755
rect 35884 22715 35885 22755
rect 36740 22724 36749 22764
rect 36740 22723 36798 22724
rect 10549 22706 10591 22715
rect 11404 22706 11450 22715
rect 13525 22706 13567 22715
rect 33580 22706 33626 22715
rect 34449 22706 34491 22715
rect 34828 22706 34874 22715
rect 35701 22706 35743 22715
rect 35884 22706 35930 22715
rect 8245 22680 8287 22689
rect 11557 22680 11599 22689
rect 11972 22680 12030 22681
rect 12373 22680 12415 22689
rect 13932 22680 13974 22689
rect 32132 22680 32190 22681
rect 32341 22680 32383 22689
rect 8245 22640 8246 22680
rect 9148 22671 9194 22680
rect 8245 22631 8287 22640
rect 9148 22631 9149 22671
rect 11557 22640 11558 22680
rect 11972 22640 11981 22680
rect 12373 22640 12374 22680
rect 13932 22640 13933 22680
rect 32132 22640 32141 22680
rect 32341 22640 32342 22680
rect 37805 22640 37814 22680
rect 11557 22631 11599 22640
rect 11972 22639 12030 22640
rect 12373 22631 12415 22640
rect 13932 22631 13974 22640
rect 32132 22639 32190 22640
rect 32341 22631 32383 22640
rect 9148 22622 9194 22631
rect 12613 22596 12655 22605
rect 32821 22596 32863 22605
rect 12613 22556 12614 22596
rect 32821 22556 32822 22596
rect 12613 22547 12655 22556
rect 32821 22547 32863 22556
rect 8005 22512 8047 22521
rect 10069 22512 10111 22521
rect 10244 22512 10302 22513
rect 33397 22512 33439 22521
rect 34148 22512 34206 22513
rect 35396 22512 35454 22513
rect 38677 22512 38719 22521
rect 8005 22472 8006 22512
rect 10069 22472 10070 22512
rect 10244 22472 10253 22512
rect 33397 22472 33398 22512
rect 34148 22472 34157 22512
rect 35396 22472 35405 22512
rect 38677 22472 38678 22512
rect 8005 22463 8047 22472
rect 10069 22463 10111 22472
rect 10244 22471 10302 22472
rect 33397 22463 33439 22472
rect 34148 22471 34206 22472
rect 35396 22471 35454 22472
rect 38677 22463 38719 22472
rect 8005 22176 8047 22185
rect 8629 22176 8671 22185
rect 10933 22176 10975 22185
rect 12356 22176 12414 22177
rect 33205 22176 33247 22185
rect 33781 22176 33823 22185
rect 35108 22176 35166 22177
rect 37237 22176 37279 22185
rect 8005 22136 8006 22176
rect 8629 22136 8630 22176
rect 10933 22136 10934 22176
rect 12356 22136 12365 22176
rect 33205 22136 33206 22176
rect 33781 22136 33782 22176
rect 35108 22136 35117 22176
rect 37237 22136 37238 22176
rect 8005 22127 8047 22136
rect 8629 22127 8671 22136
rect 10933 22127 10975 22136
rect 12356 22135 12414 22136
rect 33205 22127 33247 22136
rect 33781 22127 33823 22136
rect 35108 22135 35166 22136
rect 37237 22127 37279 22136
rect 8245 22008 8287 22017
rect 11317 22008 11359 22017
rect 12565 22008 12607 22017
rect 32132 22008 32190 22009
rect 32708 22008 32766 22009
rect 36356 22008 36414 22009
rect 8245 21968 8246 22008
rect 11317 21968 11318 22008
rect 11740 21999 11786 22008
rect 8245 21959 8287 21968
rect 11317 21959 11359 21968
rect 11740 21959 11741 21999
rect 12565 21968 12566 22008
rect 32132 21968 32141 22008
rect 32708 21968 32717 22008
rect 36356 21968 36365 22008
rect 12565 21959 12607 21968
rect 32132 21967 32190 21968
rect 32708 21967 32766 21968
rect 36356 21967 36414 21968
rect 11740 21950 11786 21959
rect 8533 21924 8575 21933
rect 8725 21924 8767 21933
rect 8917 21924 8959 21933
rect 9109 21929 9151 21938
rect 8533 21884 8534 21924
rect 8725 21884 8726 21924
rect 8917 21884 8918 21924
rect 9109 21889 9110 21929
rect 9301 21924 9343 21933
rect 9493 21924 9535 21933
rect 9967 21924 10025 21925
rect 10484 21924 10542 21925
rect 10628 21924 10686 21925
rect 11605 21924 11647 21933
rect 11834 21924 11892 21925
rect 12181 21924 12223 21933
rect 12356 21924 12414 21925
rect 12661 21924 12703 21933
rect 12780 21924 12822 21933
rect 12890 21924 12948 21925
rect 13045 21924 13087 21933
rect 13220 21924 13278 21925
rect 13430 21924 13472 21933
rect 13619 21924 13661 21933
rect 13813 21924 13855 21933
rect 14005 21924 14047 21933
rect 32516 21924 32574 21925
rect 33013 21924 33055 21933
rect 33493 21924 33535 21933
rect 33668 21924 33726 21925
rect 33781 21924 33823 21933
rect 34052 21924 34110 21925
rect 34368 21924 34410 21933
rect 34549 21924 34591 21933
rect 34683 21924 34741 21925
rect 35317 21924 35359 21933
rect 35780 21924 35838 21925
rect 35893 21924 35935 21933
rect 37045 21924 37087 21933
rect 37909 21924 37951 21933
rect 38293 21924 38335 21933
rect 38581 21924 38623 21933
rect 8533 21875 8575 21884
rect 8725 21875 8767 21884
rect 8917 21875 8959 21884
rect 9109 21880 9151 21889
rect 9301 21884 9302 21924
rect 9493 21884 9494 21924
rect 9967 21884 9976 21924
rect 10484 21884 10493 21924
rect 10628 21884 10637 21924
rect 11605 21884 11606 21924
rect 11834 21884 11843 21924
rect 12181 21884 12182 21924
rect 12356 21884 12365 21924
rect 12661 21884 12662 21924
rect 12780 21884 12781 21924
rect 12890 21884 12899 21924
rect 13045 21884 13046 21924
rect 13220 21884 13229 21924
rect 13430 21884 13431 21924
rect 13619 21884 13620 21924
rect 13813 21884 13814 21924
rect 14005 21884 14006 21924
rect 32516 21884 32525 21924
rect 33013 21884 33014 21924
rect 33493 21884 33494 21924
rect 33668 21884 33677 21924
rect 33781 21884 33782 21924
rect 34052 21884 34061 21924
rect 34368 21884 34369 21924
rect 34549 21884 34550 21924
rect 34683 21884 34692 21924
rect 35020 21915 35066 21924
rect 9301 21875 9343 21884
rect 9493 21875 9535 21884
rect 9967 21883 10025 21884
rect 10484 21883 10542 21884
rect 10628 21883 10686 21884
rect 11605 21875 11647 21884
rect 11834 21883 11892 21884
rect 12181 21875 12223 21884
rect 12356 21883 12414 21884
rect 12661 21875 12703 21884
rect 12780 21875 12822 21884
rect 12890 21883 12948 21884
rect 13045 21875 13087 21884
rect 13220 21883 13278 21884
rect 13430 21875 13472 21884
rect 13619 21875 13661 21884
rect 13813 21875 13855 21884
rect 14005 21875 14047 21884
rect 32516 21883 32574 21884
rect 33013 21875 33055 21884
rect 33493 21875 33535 21884
rect 33668 21883 33726 21884
rect 33781 21875 33823 21884
rect 34052 21883 34110 21884
rect 34368 21875 34410 21884
rect 34549 21875 34591 21884
rect 34683 21883 34741 21884
rect 35020 21875 35021 21915
rect 35317 21884 35318 21924
rect 35780 21884 35789 21924
rect 35893 21884 35894 21924
rect 37045 21884 37046 21924
rect 37909 21884 37910 21924
rect 38293 21884 38294 21924
rect 38581 21884 38582 21924
rect 35317 21875 35359 21884
rect 35780 21883 35838 21884
rect 35893 21875 35935 21884
rect 37045 21875 37087 21884
rect 37909 21875 37951 21884
rect 38293 21875 38335 21884
rect 38581 21875 38623 21884
rect 35020 21866 35066 21875
rect 9013 21840 9055 21849
rect 9674 21840 9716 21849
rect 10944 21840 10986 21849
rect 11509 21840 11551 21849
rect 13525 21840 13567 21849
rect 35125 21840 35167 21849
rect 38084 21840 38142 21841
rect 9013 21800 9014 21840
rect 9674 21800 9675 21840
rect 10944 21800 10945 21840
rect 11509 21800 11510 21840
rect 13525 21800 13526 21840
rect 35125 21800 35126 21840
rect 38084 21800 38093 21840
rect 9013 21791 9055 21800
rect 9674 21791 9716 21800
rect 10944 21791 10986 21800
rect 11509 21791 11551 21800
rect 13525 21791 13567 21800
rect 35125 21791 35167 21800
rect 38084 21799 38142 21800
rect 9397 21756 9439 21765
rect 9764 21756 9822 21757
rect 9877 21756 9919 21765
rect 10292 21756 10350 21757
rect 10724 21756 10782 21757
rect 11077 21756 11119 21765
rect 13141 21756 13183 21765
rect 13813 21756 13855 21765
rect 32228 21756 32286 21757
rect 32900 21756 32958 21757
rect 33188 21756 33246 21757
rect 34148 21756 34206 21757
rect 34261 21756 34303 21765
rect 34837 21756 34879 21765
rect 36181 21756 36223 21765
rect 38372 21756 38430 21757
rect 9397 21716 9398 21756
rect 9764 21716 9773 21756
rect 9877 21716 9878 21756
rect 10292 21716 10301 21756
rect 10724 21716 10733 21756
rect 11077 21716 11078 21756
rect 13141 21716 13142 21756
rect 13813 21716 13814 21756
rect 32228 21716 32237 21756
rect 32900 21716 32909 21756
rect 33188 21716 33197 21756
rect 34148 21716 34157 21756
rect 34261 21716 34262 21756
rect 34837 21716 34838 21756
rect 36181 21716 36182 21756
rect 38372 21716 38381 21756
rect 9397 21707 9439 21716
rect 9764 21715 9822 21716
rect 9877 21707 9919 21716
rect 10292 21715 10350 21716
rect 10724 21715 10782 21716
rect 11077 21707 11119 21716
rect 13141 21707 13183 21716
rect 13813 21707 13855 21716
rect 32228 21715 32286 21716
rect 32900 21715 32958 21716
rect 33188 21715 33246 21716
rect 34148 21715 34206 21716
rect 34261 21707 34303 21716
rect 34837 21707 34879 21716
rect 36181 21707 36223 21716
rect 38372 21715 38430 21716
rect 10069 21420 10111 21429
rect 10628 21420 10686 21421
rect 12757 21420 12799 21429
rect 13604 21420 13662 21421
rect 13717 21420 13759 21429
rect 32372 21420 32430 21421
rect 36373 21420 36415 21429
rect 10069 21380 10070 21420
rect 10628 21380 10637 21420
rect 12757 21380 12758 21420
rect 13604 21380 13613 21420
rect 13717 21380 13718 21420
rect 32372 21380 32381 21420
rect 36373 21380 36374 21420
rect 10069 21371 10111 21380
rect 10628 21379 10686 21380
rect 12757 21371 12799 21380
rect 13604 21379 13662 21380
rect 13717 21371 13759 21380
rect 32372 21379 32430 21380
rect 36373 21371 36415 21380
rect 11461 21336 11503 21345
rect 12074 21336 12116 21345
rect 12277 21336 12319 21345
rect 32149 21336 32191 21345
rect 33301 21336 33343 21345
rect 35221 21336 35263 21345
rect 36181 21336 36223 21345
rect 38660 21336 38718 21337
rect 11461 21296 11462 21336
rect 12074 21296 12075 21336
rect 12277 21296 12278 21336
rect 32149 21296 32150 21336
rect 33301 21296 33302 21336
rect 35221 21296 35222 21336
rect 36181 21296 36182 21336
rect 38660 21296 38669 21336
rect 11461 21287 11503 21296
rect 12074 21287 12116 21296
rect 12277 21287 12319 21296
rect 32149 21287 32191 21296
rect 33301 21287 33343 21296
rect 35221 21287 35263 21296
rect 36181 21287 36223 21296
rect 38660 21295 38718 21296
rect 9109 21252 9151 21261
rect 9536 21252 9578 21261
rect 9781 21252 9823 21261
rect 10165 21252 10207 21261
rect 10394 21252 10452 21253
rect 10789 21252 10831 21261
rect 10933 21252 10975 21261
rect 12554 21252 12596 21261
rect 13141 21252 13183 21261
rect 13370 21252 13428 21253
rect 13514 21252 13556 21261
rect 14005 21252 14047 21261
rect 32516 21252 32574 21253
rect 33397 21252 33439 21261
rect 33626 21252 33684 21253
rect 34103 21252 34161 21253
rect 34538 21252 34580 21261
rect 34645 21252 34687 21261
rect 35012 21252 35070 21253
rect 35313 21252 35355 21261
rect 35557 21252 35599 21261
rect 38276 21252 38334 21253
rect 9109 21212 9110 21252
rect 9536 21212 9537 21252
rect 9781 21212 9782 21252
rect 10165 21212 10166 21252
rect 10394 21212 10403 21252
rect 10789 21212 10790 21252
rect 10933 21212 10934 21252
rect 12373 21243 12415 21252
rect 9109 21203 9151 21212
rect 9536 21203 9578 21212
rect 9781 21203 9823 21212
rect 10165 21203 10207 21212
rect 10394 21211 10452 21212
rect 10789 21203 10831 21212
rect 10933 21203 10975 21212
rect 12373 21203 12374 21243
rect 12554 21212 12555 21252
rect 12853 21243 12895 21252
rect 12554 21203 12596 21212
rect 12853 21203 12854 21243
rect 13141 21212 13142 21252
rect 13370 21212 13379 21252
rect 13514 21212 13515 21252
rect 13813 21243 13855 21252
rect 13141 21203 13183 21212
rect 13370 21211 13428 21212
rect 13514 21203 13556 21212
rect 13813 21203 13814 21243
rect 14005 21212 14006 21252
rect 32516 21212 32525 21252
rect 32629 21243 32671 21252
rect 14005 21203 14047 21212
rect 32516 21211 32574 21212
rect 32629 21203 32630 21243
rect 33397 21212 33398 21252
rect 33626 21212 33635 21252
rect 34103 21212 34112 21252
rect 34538 21212 34539 21252
rect 34645 21212 34646 21252
rect 35012 21212 35021 21252
rect 35313 21212 35314 21252
rect 35557 21212 35558 21252
rect 38276 21212 38285 21252
rect 33397 21203 33439 21212
rect 33626 21211 33684 21212
rect 34103 21211 34161 21212
rect 34538 21203 34580 21212
rect 34645 21203 34687 21212
rect 35012 21211 35070 21212
rect 35313 21203 35355 21212
rect 35557 21203 35599 21212
rect 38276 21211 38334 21212
rect 12373 21194 12415 21203
rect 12853 21194 12895 21203
rect 13813 21194 13855 21203
rect 32629 21194 32671 21203
rect 9668 21168 9726 21169
rect 9877 21168 9919 21177
rect 11317 21168 11359 21177
rect 11701 21168 11743 21177
rect 13045 21168 13087 21177
rect 32245 21168 32287 21177
rect 33516 21168 33558 21177
rect 33908 21168 33966 21169
rect 9668 21128 9677 21168
rect 9877 21128 9878 21168
rect 10300 21159 10346 21168
rect 9668 21127 9726 21128
rect 9877 21119 9919 21128
rect 10300 21119 10301 21159
rect 11317 21128 11318 21168
rect 11701 21128 11702 21168
rect 13045 21128 13046 21168
rect 13276 21159 13322 21168
rect 11317 21119 11359 21128
rect 11701 21119 11743 21128
rect 13045 21119 13087 21128
rect 13276 21119 13277 21159
rect 32245 21128 32246 21168
rect 33516 21128 33517 21168
rect 33908 21128 33917 21168
rect 32245 21119 32287 21128
rect 33516 21119 33558 21128
rect 33908 21127 33966 21128
rect 10300 21110 10346 21119
rect 13276 21110 13322 21119
rect 8324 21000 8382 21001
rect 11077 21000 11119 21009
rect 12068 21000 12126 21001
rect 12548 21000 12606 21001
rect 32917 21000 32959 21009
rect 34645 21000 34687 21009
rect 8324 20960 8333 21000
rect 11077 20960 11078 21000
rect 12068 20960 12077 21000
rect 12548 20960 12557 21000
rect 32917 20960 32918 21000
rect 34645 20960 34646 21000
rect 8324 20959 8382 20960
rect 11077 20951 11119 20960
rect 12068 20959 12126 20960
rect 12548 20959 12606 20960
rect 32917 20951 32959 20960
rect 34645 20951 34687 20960
rect 9572 20664 9630 20665
rect 11125 20664 11167 20673
rect 11780 20664 11838 20665
rect 13316 20664 13374 20665
rect 38677 20664 38719 20673
rect 9572 20624 9581 20664
rect 11125 20624 11126 20664
rect 11780 20624 11789 20664
rect 13316 20624 13325 20664
rect 38677 20624 38678 20664
rect 9572 20623 9630 20624
rect 11125 20615 11167 20624
rect 11780 20623 11838 20624
rect 13316 20623 13374 20624
rect 38677 20615 38719 20624
rect 9013 20580 9055 20589
rect 9013 20540 9014 20580
rect 9013 20531 9055 20540
rect 8245 20496 8287 20505
rect 12853 20496 12895 20505
rect 13068 20496 13110 20505
rect 33973 20496 34015 20505
rect 34453 20496 34495 20505
rect 34668 20496 34710 20505
rect 8245 20456 8246 20496
rect 12853 20456 12854 20496
rect 13068 20456 13069 20496
rect 33973 20456 33974 20496
rect 34453 20456 34454 20496
rect 34668 20456 34669 20496
rect 37997 20456 38006 20496
rect 8245 20447 8287 20456
rect 12853 20447 12895 20456
rect 13068 20447 13110 20456
rect 33973 20447 34015 20456
rect 34453 20447 34495 20456
rect 34668 20447 34710 20456
rect 9205 20412 9247 20421
rect 9397 20412 9439 20421
rect 9578 20412 9620 20421
rect 9869 20412 9927 20413
rect 10340 20412 10398 20413
rect 10453 20412 10495 20421
rect 10820 20412 10878 20413
rect 11139 20412 11181 20421
rect 11413 20412 11455 20421
rect 11532 20412 11574 20421
rect 11642 20412 11700 20413
rect 11783 20412 11825 20421
rect 12077 20412 12135 20413
rect 12469 20412 12511 20421
rect 12661 20412 12703 20421
rect 12949 20412 12991 20421
rect 13178 20412 13236 20413
rect 13322 20412 13364 20421
rect 13613 20412 13671 20413
rect 13760 20412 13802 20421
rect 13892 20412 13950 20413
rect 14005 20412 14047 20421
rect 32053 20412 32095 20421
rect 32228 20412 32286 20413
rect 32725 20412 32767 20421
rect 33013 20412 33055 20421
rect 33397 20412 33439 20421
rect 34052 20412 34110 20413
rect 34549 20412 34591 20421
rect 34778 20412 34836 20413
rect 35025 20412 35067 20421
rect 35221 20412 35263 20421
rect 35509 20412 35551 20421
rect 36740 20412 36798 20413
rect 9205 20372 9206 20412
rect 9397 20372 9398 20412
rect 9578 20372 9579 20412
rect 9869 20372 9878 20412
rect 10340 20372 10349 20412
rect 10453 20372 10454 20412
rect 10820 20372 10829 20412
rect 11139 20372 11140 20412
rect 11413 20372 11414 20412
rect 11532 20372 11533 20412
rect 11642 20372 11651 20412
rect 11783 20372 11784 20412
rect 12077 20372 12086 20412
rect 12469 20372 12470 20412
rect 12661 20372 12662 20412
rect 12949 20372 12950 20412
rect 13178 20372 13187 20412
rect 13322 20372 13323 20412
rect 13613 20372 13622 20412
rect 13760 20372 13761 20412
rect 13892 20372 13901 20412
rect 14005 20372 14006 20412
rect 32053 20372 32054 20412
rect 32228 20372 32237 20412
rect 32725 20372 32726 20412
rect 33013 20372 33014 20412
rect 33397 20372 33398 20412
rect 34052 20372 34061 20412
rect 34549 20372 34550 20412
rect 34778 20372 34787 20412
rect 35025 20372 35026 20412
rect 35221 20372 35222 20412
rect 35509 20372 35510 20412
rect 36740 20372 36749 20412
rect 9205 20363 9247 20372
rect 9397 20363 9439 20372
rect 9578 20363 9620 20372
rect 9869 20371 9927 20372
rect 10340 20371 10398 20372
rect 10453 20363 10495 20372
rect 10820 20371 10878 20372
rect 11139 20363 11181 20372
rect 11413 20363 11455 20372
rect 11532 20363 11574 20372
rect 11642 20371 11700 20372
rect 11783 20363 11825 20372
rect 12077 20371 12135 20372
rect 12469 20363 12511 20372
rect 12661 20363 12703 20372
rect 12949 20363 12991 20372
rect 13178 20371 13236 20372
rect 13322 20363 13364 20372
rect 13613 20371 13671 20372
rect 13760 20363 13802 20372
rect 13892 20371 13950 20372
rect 14005 20363 14047 20372
rect 32053 20363 32095 20372
rect 32228 20371 32286 20372
rect 32725 20363 32767 20372
rect 33013 20363 33055 20372
rect 33397 20363 33439 20372
rect 34052 20371 34110 20372
rect 34549 20363 34591 20372
rect 34778 20371 34836 20372
rect 35025 20363 35067 20372
rect 35221 20363 35263 20372
rect 35509 20363 35551 20372
rect 36740 20371 36798 20372
rect 10659 20328 10701 20337
rect 32149 20328 32191 20337
rect 36356 20328 36414 20329
rect 10659 20288 10660 20328
rect 32149 20288 32150 20328
rect 36356 20288 36365 20328
rect 10659 20279 10701 20288
rect 32149 20279 32191 20288
rect 36356 20287 36414 20288
rect 8005 20244 8047 20253
rect 9205 20244 9247 20253
rect 9781 20244 9823 20253
rect 10549 20244 10591 20253
rect 10916 20244 10974 20245
rect 11317 20244 11359 20253
rect 11989 20244 12031 20253
rect 12644 20244 12702 20245
rect 13525 20244 13567 20253
rect 32516 20244 32574 20245
rect 33205 20244 33247 20253
rect 33476 20244 33534 20245
rect 35029 20244 35071 20253
rect 36181 20244 36223 20253
rect 8005 20204 8006 20244
rect 9205 20204 9206 20244
rect 9781 20204 9782 20244
rect 10549 20204 10550 20244
rect 10916 20204 10925 20244
rect 11317 20204 11318 20244
rect 11989 20204 11990 20244
rect 12644 20204 12653 20244
rect 13525 20204 13526 20244
rect 32516 20204 32525 20244
rect 33205 20204 33206 20244
rect 33476 20204 33485 20244
rect 33684 20235 33726 20244
rect 8005 20195 8047 20204
rect 9205 20195 9247 20204
rect 9781 20195 9823 20204
rect 10549 20195 10591 20204
rect 10916 20203 10974 20204
rect 11317 20195 11359 20204
rect 11989 20195 12031 20204
rect 12644 20203 12702 20204
rect 13525 20195 13567 20204
rect 32516 20203 32574 20204
rect 33205 20195 33247 20204
rect 33476 20203 33534 20204
rect 33684 20195 33685 20235
rect 35029 20204 35030 20244
rect 36181 20204 36182 20244
rect 35029 20195 35071 20204
rect 36181 20195 36223 20204
rect 33684 20186 33726 20195
rect 8149 19908 8191 19917
rect 12661 19908 12703 19917
rect 13892 19908 13950 19909
rect 33092 19908 33150 19909
rect 8149 19868 8150 19908
rect 12661 19868 12662 19908
rect 13892 19868 13901 19908
rect 33092 19868 33101 19908
rect 8149 19859 8191 19868
rect 12661 19859 12703 19868
rect 13892 19867 13950 19868
rect 33092 19867 33150 19868
rect 37813 19824 37855 19833
rect 37813 19784 37814 19824
rect 37813 19775 37855 19784
rect 10052 19740 10110 19741
rect 11317 19740 11359 19749
rect 11605 19740 11647 19749
rect 11834 19740 11892 19741
rect 12373 19740 12415 19749
rect 12500 19740 12558 19741
rect 13141 19740 13183 19749
rect 13316 19740 13374 19741
rect 13541 19740 13599 19741
rect 13700 19740 13758 19741
rect 13825 19740 13867 19749
rect 32149 19740 32191 19749
rect 32264 19740 32306 19749
rect 32437 19740 32479 19749
rect 32629 19740 32671 19749
rect 32804 19740 32862 19741
rect 32996 19740 33054 19741
rect 33312 19740 33354 19749
rect 33589 19740 33631 19749
rect 33781 19740 33823 19749
rect 34261 19740 34303 19749
rect 34436 19740 34494 19741
rect 34549 19740 34591 19749
rect 36644 19740 36702 19741
rect 37028 19740 37086 19741
rect 37223 19740 37265 19749
rect 37333 19740 37375 19749
rect 37525 19740 37567 19749
rect 37717 19740 37759 19749
rect 38005 19740 38047 19749
rect 10052 19700 10061 19740
rect 11317 19700 11318 19740
rect 11605 19700 11606 19740
rect 11834 19700 11843 19740
rect 12373 19700 12374 19740
rect 12500 19700 12509 19740
rect 13141 19700 13142 19740
rect 13316 19700 13325 19740
rect 13541 19700 13550 19740
rect 13700 19700 13709 19740
rect 13825 19700 13826 19740
rect 13984 19729 14042 19730
rect 10052 19699 10110 19700
rect 11317 19691 11359 19700
rect 11605 19691 11647 19700
rect 11834 19699 11892 19700
rect 12373 19691 12415 19700
rect 12500 19699 12558 19700
rect 13141 19691 13183 19700
rect 13316 19699 13374 19700
rect 13541 19699 13599 19700
rect 13700 19699 13758 19700
rect 13825 19691 13867 19700
rect 13984 19689 13993 19729
rect 32149 19700 32150 19740
rect 32264 19700 32265 19740
rect 32437 19700 32438 19740
rect 32629 19700 32630 19740
rect 32804 19700 32813 19740
rect 32996 19700 33005 19740
rect 33312 19700 33313 19740
rect 33589 19700 33590 19740
rect 33781 19700 33782 19740
rect 34261 19700 34262 19740
rect 34436 19700 34445 19740
rect 34549 19700 34550 19740
rect 36644 19700 36653 19740
rect 37028 19700 37037 19740
rect 37223 19700 37224 19740
rect 37333 19700 37334 19740
rect 37525 19700 37526 19740
rect 37717 19700 37718 19740
rect 38005 19700 38006 19740
rect 38188 19731 38234 19740
rect 32149 19691 32191 19700
rect 32264 19691 32306 19700
rect 32437 19691 32479 19700
rect 32629 19691 32671 19700
rect 32804 19699 32862 19700
rect 32996 19699 33054 19700
rect 33312 19691 33354 19700
rect 33589 19691 33631 19700
rect 33781 19691 33823 19700
rect 34261 19691 34303 19700
rect 34436 19699 34494 19700
rect 34549 19691 34591 19700
rect 36644 19699 36702 19700
rect 37028 19699 37086 19700
rect 37223 19691 37265 19700
rect 37333 19691 37375 19700
rect 37525 19691 37567 19700
rect 37717 19691 37759 19700
rect 38005 19691 38047 19700
rect 38188 19691 38189 19731
rect 13984 19688 14042 19689
rect 38188 19682 38234 19691
rect 10436 19656 10494 19657
rect 11509 19656 11551 19665
rect 33476 19656 33534 19657
rect 35108 19656 35166 19657
rect 38341 19656 38383 19665
rect 9389 19616 9398 19656
rect 10436 19616 10445 19656
rect 11509 19616 11510 19656
rect 11740 19647 11786 19656
rect 10436 19615 10494 19616
rect 11509 19607 11551 19616
rect 11740 19607 11741 19647
rect 33476 19616 33485 19656
rect 35108 19616 35117 19656
rect 38341 19616 38342 19656
rect 33476 19615 33534 19616
rect 35108 19615 35166 19616
rect 38341 19607 38383 19616
rect 11740 19598 11786 19607
rect 13316 19572 13374 19573
rect 32149 19572 32191 19581
rect 34357 19572 34399 19581
rect 37237 19572 37279 19581
rect 13316 19532 13325 19572
rect 32149 19532 32150 19572
rect 34357 19532 34358 19572
rect 37237 19532 37238 19572
rect 13316 19531 13374 19532
rect 32149 19523 32191 19532
rect 34357 19523 34399 19532
rect 37237 19523 37279 19532
rect 8533 19488 8575 19497
rect 10645 19488 10687 19497
rect 32804 19488 32862 19489
rect 33301 19488 33343 19497
rect 34741 19488 34783 19497
rect 8533 19448 8534 19488
rect 10645 19448 10646 19488
rect 32804 19448 32813 19488
rect 33301 19448 33302 19488
rect 34741 19448 34742 19488
rect 8533 19439 8575 19448
rect 10645 19439 10687 19448
rect 32804 19447 32862 19448
rect 33301 19439 33343 19448
rect 34741 19439 34783 19448
rect 13717 19152 13759 19161
rect 33572 19152 33630 19153
rect 35125 19152 35167 19161
rect 13717 19112 13718 19152
rect 33572 19112 33581 19152
rect 35125 19112 35126 19152
rect 13717 19103 13759 19112
rect 33572 19111 33630 19112
rect 35125 19103 35167 19112
rect 9397 19068 9439 19077
rect 9781 19068 9823 19077
rect 11125 19068 11167 19077
rect 11605 19068 11647 19077
rect 32180 19068 32238 19069
rect 9397 19028 9398 19068
rect 9781 19028 9782 19068
rect 11125 19028 11126 19068
rect 11605 19028 11606 19068
rect 32180 19028 32189 19068
rect 9397 19019 9439 19028
rect 9781 19019 9823 19028
rect 11125 19019 11167 19028
rect 11605 19019 11647 19028
rect 32180 19027 32238 19028
rect 10165 18984 10207 18993
rect 33013 18984 33055 18993
rect 35108 18984 35166 18985
rect 35492 18984 35550 18985
rect 10165 18944 10166 18984
rect 33013 18944 33014 18984
rect 35108 18944 35117 18984
rect 35492 18944 35501 18984
rect 10165 18935 10207 18944
rect 33013 18935 33055 18944
rect 35108 18943 35166 18944
rect 35492 18943 35550 18944
rect 13600 18911 13658 18912
rect 13726 18911 13784 18912
rect 9685 18900 9727 18909
rect 9860 18900 9918 18901
rect 9973 18900 10015 18909
rect 10261 18900 10303 18909
rect 10380 18900 10422 18909
rect 10490 18900 10548 18901
rect 10820 18900 10878 18901
rect 10933 18900 10975 18909
rect 11797 18900 11839 18909
rect 12181 18900 12223 18909
rect 12300 18900 12342 18909
rect 12410 18900 12468 18901
rect 12663 18900 12705 18909
rect 12853 18900 12895 18909
rect 13157 18900 13215 18901
rect 13316 18900 13374 18901
rect 13460 18900 13518 18901
rect 9685 18860 9686 18900
rect 9860 18860 9869 18900
rect 9973 18860 9974 18900
rect 10261 18860 10262 18900
rect 10380 18860 10381 18900
rect 10490 18860 10499 18900
rect 10820 18860 10829 18900
rect 10933 18860 10934 18900
rect 11797 18860 11798 18900
rect 12181 18860 12182 18900
rect 12300 18860 12301 18900
rect 12410 18860 12419 18900
rect 12663 18860 12664 18900
rect 12853 18860 12854 18900
rect 13157 18860 13166 18900
rect 13316 18860 13325 18900
rect 13460 18860 13469 18900
rect 13600 18871 13609 18911
rect 13726 18871 13735 18911
rect 32053 18900 32095 18909
rect 32389 18900 32431 18909
rect 32533 18900 32575 18909
rect 33109 18900 33151 18909
rect 33228 18900 33270 18909
rect 33340 18900 33382 18909
rect 33973 18900 34015 18909
rect 34244 18900 34302 18901
rect 34933 18900 34975 18909
rect 37028 18900 37086 18901
rect 37601 18900 37659 18901
rect 38081 18900 38139 18901
rect 13600 18870 13658 18871
rect 13726 18870 13784 18871
rect 32053 18860 32054 18900
rect 32389 18860 32390 18900
rect 32533 18860 32534 18900
rect 33109 18860 33110 18900
rect 33228 18860 33229 18900
rect 33340 18860 33341 18900
rect 33973 18860 33974 18900
rect 34244 18860 34253 18900
rect 34933 18860 34934 18900
rect 37028 18860 37037 18900
rect 37601 18860 37610 18900
rect 38081 18860 38090 18900
rect 9685 18851 9727 18860
rect 9860 18859 9918 18860
rect 9973 18851 10015 18860
rect 10261 18851 10303 18860
rect 10380 18851 10422 18860
rect 10490 18859 10548 18860
rect 10820 18859 10878 18860
rect 10933 18851 10975 18860
rect 11797 18851 11839 18860
rect 12181 18851 12223 18860
rect 12300 18851 12342 18860
rect 12410 18859 12468 18860
rect 12663 18851 12705 18860
rect 12853 18851 12895 18860
rect 13157 18859 13215 18860
rect 13316 18859 13374 18860
rect 13460 18859 13518 18860
rect 32053 18851 32095 18860
rect 32389 18851 32431 18860
rect 32533 18851 32575 18860
rect 33109 18851 33151 18860
rect 33228 18851 33270 18860
rect 33340 18851 33382 18860
rect 33973 18851 34015 18860
rect 34244 18859 34302 18860
rect 34933 18851 34975 18860
rect 37028 18859 37086 18860
rect 37601 18859 37659 18860
rect 38081 18859 38139 18860
rect 12085 18816 12127 18825
rect 37412 18816 37470 18817
rect 12085 18776 12086 18816
rect 37412 18776 37421 18816
rect 12085 18767 12127 18776
rect 37412 18775 37470 18776
rect 10837 18732 10879 18741
rect 12853 18732 12895 18741
rect 33781 18732 33823 18741
rect 37765 18732 37807 18741
rect 38245 18732 38287 18741
rect 10837 18692 10838 18732
rect 12853 18692 12854 18732
rect 33781 18692 33782 18732
rect 37765 18692 37766 18732
rect 38245 18692 38246 18732
rect 10837 18683 10879 18692
rect 12853 18683 12895 18692
rect 33781 18683 33823 18692
rect 37765 18683 37807 18692
rect 38245 18683 38287 18692
rect 9572 18396 9630 18397
rect 10724 18396 10782 18397
rect 11684 18396 11742 18397
rect 11876 18396 11934 18397
rect 12356 18396 12414 18397
rect 32533 18396 32575 18405
rect 33566 18396 33624 18397
rect 34549 18396 34591 18405
rect 34933 18396 34975 18405
rect 36949 18396 36991 18405
rect 37124 18396 37182 18397
rect 37429 18396 37471 18405
rect 9572 18356 9581 18396
rect 10724 18356 10733 18396
rect 11684 18356 11693 18396
rect 11876 18356 11885 18396
rect 12356 18356 12365 18396
rect 32533 18356 32534 18396
rect 33566 18356 33575 18396
rect 34549 18356 34550 18396
rect 34933 18356 34934 18396
rect 36949 18356 36950 18396
rect 37124 18356 37133 18396
rect 37429 18356 37430 18396
rect 9572 18355 9630 18356
rect 10724 18355 10782 18356
rect 11684 18355 11742 18356
rect 11876 18355 11934 18356
rect 12356 18355 12414 18356
rect 32533 18347 32575 18356
rect 33566 18355 33624 18356
rect 34549 18347 34591 18356
rect 34933 18347 34975 18356
rect 36949 18347 36991 18356
rect 37124 18355 37182 18356
rect 37429 18347 37471 18356
rect 10436 18312 10494 18313
rect 11204 18312 11262 18313
rect 34100 18312 34158 18313
rect 10436 18272 10445 18312
rect 11204 18272 11213 18312
rect 12652 18303 12698 18312
rect 13420 18303 13466 18312
rect 10436 18271 10494 18272
rect 11204 18271 11262 18272
rect 12652 18263 12653 18303
rect 13420 18263 13421 18303
rect 34100 18272 34109 18312
rect 34100 18271 34158 18272
rect 12652 18254 12698 18263
rect 13420 18254 13466 18263
rect 9685 18228 9727 18237
rect 10645 18228 10687 18237
rect 10880 18228 10922 18237
rect 11125 18228 11167 18237
rect 11605 18228 11647 18237
rect 11989 18228 12031 18237
rect 12356 18228 12414 18229
rect 12740 18228 12798 18229
rect 12874 18228 12932 18229
rect 13135 18228 13193 18229
rect 13280 18228 13338 18229
rect 13508 18228 13566 18229
rect 13684 18228 13742 18229
rect 32053 18228 32095 18237
rect 32170 18228 32228 18229
rect 32341 18228 32383 18237
rect 32629 18228 32671 18237
rect 32858 18228 32916 18229
rect 33109 18228 33151 18237
rect 33223 18228 33281 18229
rect 33350 18228 33408 18229
rect 33668 18228 33726 18229
rect 34453 18228 34495 18237
rect 34574 18228 34616 18237
rect 34976 18228 35018 18237
rect 35090 18228 35148 18229
rect 35221 18228 35263 18237
rect 36085 18228 36127 18237
rect 36277 18228 36319 18237
rect 37237 18228 37279 18237
rect 37621 18228 37663 18237
rect 9685 18188 9686 18228
rect 10645 18188 10646 18228
rect 10880 18188 10881 18228
rect 11125 18188 11126 18228
rect 11605 18188 11606 18228
rect 11989 18188 11990 18228
rect 12356 18188 12365 18228
rect 12469 18219 12511 18228
rect 9685 18179 9727 18188
rect 10645 18179 10687 18188
rect 10880 18179 10922 18188
rect 11125 18179 11167 18188
rect 11605 18179 11647 18188
rect 11989 18179 12031 18188
rect 12356 18187 12414 18188
rect 12469 18179 12470 18219
rect 12740 18188 12749 18228
rect 12874 18188 12883 18228
rect 13135 18188 13144 18228
rect 13280 18188 13289 18228
rect 13508 18188 13517 18228
rect 13684 18188 13693 18228
rect 13892 18227 13950 18228
rect 12740 18187 12798 18188
rect 12874 18187 12932 18188
rect 13135 18187 13193 18188
rect 13280 18187 13338 18188
rect 13508 18187 13566 18188
rect 13684 18187 13742 18188
rect 13892 18187 13901 18227
rect 32053 18188 32054 18228
rect 32170 18188 32179 18228
rect 32341 18188 32342 18228
rect 32629 18188 32630 18228
rect 32858 18188 32867 18228
rect 33109 18188 33110 18228
rect 33223 18188 33232 18228
rect 33350 18188 33359 18228
rect 33668 18188 33677 18228
rect 33781 18219 33823 18228
rect 13892 18186 13950 18187
rect 32053 18179 32095 18188
rect 32170 18187 32228 18188
rect 32341 18179 32383 18188
rect 32629 18179 32671 18188
rect 32858 18187 32916 18188
rect 33109 18179 33151 18188
rect 33223 18187 33281 18188
rect 33350 18187 33408 18188
rect 33668 18187 33726 18188
rect 33781 18179 33782 18219
rect 34453 18188 34454 18228
rect 34574 18188 34575 18228
rect 34976 18188 34977 18228
rect 35090 18188 35099 18228
rect 35221 18188 35222 18228
rect 36085 18188 36086 18228
rect 36277 18188 36278 18228
rect 37237 18188 37238 18228
rect 37621 18188 37622 18228
rect 34453 18179 34495 18188
rect 34574 18179 34616 18188
rect 34976 18179 35018 18188
rect 35090 18187 35148 18188
rect 35221 18179 35263 18188
rect 36085 18179 36127 18188
rect 36277 18179 36319 18188
rect 37237 18179 37279 18188
rect 37621 18179 37663 18188
rect 12469 18170 12511 18179
rect 33781 18170 33823 18179
rect 11012 18144 11070 18145
rect 11012 18104 11021 18144
rect 32764 18135 32810 18144
rect 11012 18103 11070 18104
rect 32764 18095 32765 18135
rect 32764 18086 32810 18095
rect 11413 18060 11455 18069
rect 12181 18060 12223 18069
rect 32149 18060 32191 18069
rect 34244 18060 34302 18061
rect 38005 18060 38047 18069
rect 38389 18060 38431 18069
rect 11413 18020 11414 18060
rect 12181 18020 12182 18060
rect 32149 18020 32150 18060
rect 34244 18020 34253 18060
rect 38005 18020 38006 18060
rect 38389 18020 38390 18060
rect 11413 18011 11455 18020
rect 12181 18011 12223 18020
rect 32149 18011 32191 18020
rect 34244 18019 34302 18020
rect 38005 18011 38047 18020
rect 38389 18011 38431 18020
rect 9877 17976 9919 17985
rect 13124 17976 13182 17977
rect 33397 17976 33439 17985
rect 35413 17976 35455 17985
rect 37717 17976 37759 17985
rect 9877 17936 9878 17976
rect 13124 17936 13133 17976
rect 33397 17936 33398 17976
rect 35413 17936 35414 17976
rect 37717 17936 37718 17976
rect 9877 17927 9919 17936
rect 13124 17935 13182 17936
rect 33397 17927 33439 17936
rect 35413 17927 35455 17936
rect 37717 17927 37759 17936
rect 8917 17640 8959 17649
rect 11029 17640 11071 17649
rect 32804 17640 32862 17641
rect 34837 17640 34879 17649
rect 38197 17640 38239 17649
rect 8917 17600 8918 17640
rect 11029 17600 11030 17640
rect 32804 17600 32813 17640
rect 34837 17600 34838 17640
rect 38197 17600 38198 17640
rect 8917 17591 8959 17600
rect 11029 17591 11071 17600
rect 32804 17599 32862 17600
rect 34837 17591 34879 17600
rect 38197 17591 38239 17600
rect 32437 17556 32479 17565
rect 37717 17556 37759 17565
rect 32437 17516 32438 17556
rect 37717 17516 37718 17556
rect 32437 17507 32479 17516
rect 37717 17507 37759 17516
rect 33157 17472 33199 17481
rect 33572 17472 33630 17473
rect 33781 17472 33823 17481
rect 35588 17472 35646 17473
rect 37508 17472 37566 17473
rect 11452 17463 11498 17472
rect 11452 17423 11453 17463
rect 33157 17432 33158 17472
rect 33572 17432 33581 17472
rect 33781 17432 33782 17472
rect 35588 17432 35597 17472
rect 37325 17432 37334 17472
rect 37508 17432 37517 17472
rect 32804 17430 32862 17431
rect 11452 17414 11498 17423
rect 32437 17421 32479 17430
rect 8821 17388 8863 17397
rect 9236 17388 9294 17389
rect 9589 17388 9631 17397
rect 10148 17388 10206 17389
rect 10261 17388 10303 17397
rect 10837 17388 10879 17397
rect 11317 17388 11359 17397
rect 11546 17388 11604 17389
rect 32139 17388 32181 17397
rect 32324 17388 32382 17389
rect 8821 17348 8822 17388
rect 9014 17361 9072 17362
rect 8821 17339 8863 17348
rect 9014 17321 9023 17361
rect 9236 17348 9245 17388
rect 9589 17348 9590 17388
rect 10148 17348 10157 17388
rect 10261 17348 10262 17388
rect 10837 17348 10838 17388
rect 11317 17348 11318 17388
rect 11546 17348 11555 17388
rect 32139 17348 32140 17388
rect 32324 17348 32333 17388
rect 32437 17381 32438 17421
rect 32629 17388 32671 17397
rect 32804 17390 32813 17430
rect 33157 17423 33199 17432
rect 33572 17431 33630 17432
rect 33781 17423 33823 17432
rect 35588 17431 35646 17432
rect 37508 17431 37566 17432
rect 32804 17389 32862 17390
rect 32993 17388 33051 17389
rect 33452 17388 33510 17389
rect 33685 17388 33727 17397
rect 34357 17388 34399 17397
rect 34837 17388 34879 17397
rect 35029 17388 35071 17397
rect 37124 17388 37182 17389
rect 38101 17388 38143 17397
rect 38293 17388 38335 17397
rect 38474 17388 38516 17397
rect 38677 17388 38719 17397
rect 32437 17372 32479 17381
rect 32629 17348 32630 17388
rect 32993 17348 33002 17388
rect 33452 17348 33461 17388
rect 33685 17348 33686 17388
rect 34060 17379 34106 17388
rect 9236 17347 9294 17348
rect 9589 17339 9631 17348
rect 10148 17347 10206 17348
rect 10261 17339 10303 17348
rect 10837 17339 10879 17348
rect 11317 17339 11359 17348
rect 11546 17347 11604 17348
rect 32139 17339 32181 17348
rect 32324 17347 32382 17348
rect 32629 17339 32671 17348
rect 32993 17347 33051 17348
rect 33452 17347 33510 17348
rect 33685 17339 33727 17348
rect 34060 17339 34061 17379
rect 34357 17348 34358 17388
rect 34837 17348 34838 17388
rect 35029 17348 35030 17388
rect 37124 17348 37133 17388
rect 38101 17348 38102 17388
rect 38293 17348 38294 17388
rect 38474 17348 38475 17388
rect 38677 17348 38678 17388
rect 34357 17339 34399 17348
rect 34837 17339 34879 17348
rect 35029 17339 35071 17348
rect 37124 17347 37182 17348
rect 38101 17339 38143 17348
rect 38293 17339 38335 17348
rect 38474 17339 38516 17348
rect 38677 17339 38719 17348
rect 34060 17330 34106 17339
rect 9014 17320 9072 17321
rect 11221 17304 11263 17313
rect 11221 17264 11222 17304
rect 11221 17255 11263 17264
rect 11684 17263 11690 17305
rect 34165 17304 34207 17313
rect 34165 17264 34166 17304
rect 34165 17255 34207 17264
rect 9685 17220 9727 17229
rect 10549 17220 10591 17229
rect 10724 17220 10782 17221
rect 35221 17220 35263 17229
rect 38485 17220 38527 17229
rect 9685 17180 9686 17220
rect 10549 17180 10550 17220
rect 10724 17180 10733 17220
rect 35221 17180 35222 17220
rect 38485 17180 38486 17220
rect 9685 17171 9727 17180
rect 10549 17171 10591 17180
rect 10724 17179 10782 17180
rect 35221 17171 35263 17180
rect 38485 17171 38527 17180
rect 9397 16884 9439 16893
rect 9758 16884 9816 16885
rect 10820 16884 10878 16885
rect 11300 16884 11358 16885
rect 11509 16884 11551 16893
rect 32629 16884 32671 16893
rect 34453 16884 34495 16893
rect 34820 16884 34878 16885
rect 37220 16884 37278 16885
rect 9397 16844 9398 16884
rect 9758 16844 9767 16884
rect 10820 16844 10829 16884
rect 11300 16844 11309 16884
rect 11509 16844 11510 16884
rect 32629 16844 32630 16884
rect 34453 16844 34454 16884
rect 34820 16844 34829 16884
rect 37220 16844 37229 16884
rect 9397 16835 9439 16844
rect 9758 16843 9816 16844
rect 10820 16843 10878 16844
rect 11300 16843 11358 16844
rect 11509 16835 11551 16844
rect 32629 16835 32671 16844
rect 34453 16835 34495 16844
rect 34820 16843 34878 16844
rect 37220 16843 37278 16844
rect 11012 16800 11070 16801
rect 11012 16760 11021 16800
rect 11012 16759 11070 16760
rect 8996 16716 9054 16717
rect 9109 16716 9151 16725
rect 9860 16716 9918 16717
rect 10496 16716 10538 16725
rect 10741 16716 10783 16725
rect 11221 16716 11263 16725
rect 32885 16716 32943 16717
rect 32996 16716 33054 16717
rect 33445 16716 33487 16725
rect 33589 16716 33631 16725
rect 34165 16716 34207 16725
rect 34292 16716 34350 16717
rect 34406 16716 34464 16717
rect 34933 16716 34975 16725
rect 35317 16716 35359 16725
rect 36181 16716 36223 16725
rect 36373 16716 36415 16725
rect 37525 16716 37567 16725
rect 8996 16676 9005 16716
rect 9109 16676 9110 16716
rect 9860 16676 9869 16716
rect 9973 16707 10015 16716
rect 8996 16675 9054 16676
rect 9109 16667 9151 16676
rect 9860 16675 9918 16676
rect 9973 16667 9974 16707
rect 10496 16676 10497 16716
rect 10741 16676 10742 16716
rect 11221 16676 11222 16716
rect 10496 16667 10538 16676
rect 10741 16667 10783 16676
rect 11221 16667 11263 16676
rect 11605 16674 11647 16683
rect 32885 16676 32894 16716
rect 32996 16676 33005 16716
rect 33445 16676 33446 16716
rect 33589 16676 33590 16716
rect 34165 16676 34166 16716
rect 34292 16676 34301 16716
rect 34406 16676 34415 16716
rect 34933 16676 34934 16716
rect 35317 16676 35318 16716
rect 36181 16676 36182 16716
rect 36373 16676 36374 16716
rect 37525 16676 37526 16716
rect 37996 16707 38042 16716
rect 32885 16675 32943 16676
rect 32996 16675 33054 16676
rect 32782 16674 32840 16675
rect 9973 16658 10015 16667
rect 11605 16634 11606 16674
rect 32782 16634 32791 16674
rect 33445 16667 33487 16676
rect 33589 16667 33631 16676
rect 34165 16667 34207 16676
rect 34292 16675 34350 16676
rect 34406 16675 34464 16676
rect 34933 16667 34975 16676
rect 35317 16667 35359 16676
rect 36181 16667 36223 16676
rect 36373 16667 36415 16676
rect 37525 16667 37567 16676
rect 37996 16667 37997 16707
rect 37996 16658 38042 16667
rect 10628 16632 10686 16633
rect 10628 16592 10637 16632
rect 11605 16625 11647 16634
rect 32782 16633 32840 16634
rect 37435 16632 37477 16641
rect 38149 16632 38191 16641
rect 37435 16592 37436 16632
rect 38149 16592 38150 16632
rect 10628 16591 10686 16592
rect 37435 16583 37477 16592
rect 38149 16583 38191 16592
rect 33236 16548 33294 16549
rect 33781 16548 33823 16557
rect 38485 16548 38527 16557
rect 33236 16508 33245 16548
rect 33781 16508 33782 16548
rect 38485 16508 38486 16548
rect 33236 16507 33294 16508
rect 33781 16499 33823 16508
rect 38485 16499 38527 16508
rect 10261 16464 10303 16473
rect 32245 16464 32287 16473
rect 35509 16464 35551 16473
rect 37045 16464 37087 16473
rect 10261 16424 10262 16464
rect 32245 16424 32246 16464
rect 35509 16424 35510 16464
rect 37045 16424 37046 16464
rect 10261 16415 10303 16424
rect 32245 16415 32287 16424
rect 35509 16415 35551 16424
rect 37045 16415 37087 16424
rect 9349 16128 9391 16137
rect 11588 16128 11646 16129
rect 32341 16128 32383 16137
rect 32629 16128 32671 16137
rect 35029 16128 35071 16137
rect 38101 16128 38143 16137
rect 9349 16088 9350 16128
rect 11588 16088 11597 16128
rect 32341 16088 32342 16128
rect 32629 16088 32630 16128
rect 35029 16088 35030 16128
rect 38101 16088 38102 16128
rect 9349 16079 9391 16088
rect 11588 16087 11646 16088
rect 32341 16079 32383 16088
rect 32629 16079 32671 16088
rect 35029 16079 35071 16088
rect 38101 16079 38143 16088
rect 33301 16044 33343 16053
rect 38389 16044 38431 16053
rect 11381 16035 11423 16044
rect 11381 15995 11382 16035
rect 33301 16004 33302 16044
rect 38389 16004 38390 16044
rect 33301 15995 33343 16004
rect 38389 15995 38431 16004
rect 11381 15986 11423 15995
rect 32458 15960 32500 15969
rect 32821 15960 32863 15969
rect 33036 15960 33078 15969
rect 34148 15960 34206 15961
rect 35876 15960 35934 15961
rect 32458 15920 32459 15960
rect 32821 15920 32822 15960
rect 33036 15920 33037 15960
rect 34148 15920 34157 15960
rect 35876 15920 35885 15960
rect 37613 15920 37622 15960
rect 32458 15911 32500 15920
rect 32576 15909 32618 15918
rect 32821 15911 32863 15920
rect 33036 15911 33078 15920
rect 34148 15919 34206 15920
rect 35876 15919 35934 15920
rect 8725 15876 8767 15885
rect 9013 15876 9055 15885
rect 9493 15876 9535 15885
rect 9685 15876 9727 15885
rect 10645 15876 10687 15885
rect 10733 15876 10791 15877
rect 11396 15876 11454 15877
rect 32245 15876 32287 15885
rect 8725 15836 8726 15876
rect 9013 15836 9014 15876
rect 9493 15836 9494 15876
rect 9685 15836 9686 15876
rect 10645 15836 10646 15876
rect 10733 15836 10742 15876
rect 11396 15836 11405 15876
rect 32245 15836 32246 15876
rect 32576 15869 32577 15909
rect 32917 15876 32959 15885
rect 33151 15876 33193 15885
rect 33322 15876 33364 15885
rect 33589 15876 33631 15885
rect 33781 15876 33823 15885
rect 34016 15876 34058 15885
rect 34261 15876 34303 15885
rect 34741 15876 34783 15885
rect 34829 15876 34887 15877
rect 35029 15876 35071 15885
rect 35210 15876 35268 15877
rect 37412 15876 37470 15877
rect 38005 15876 38047 15885
rect 38197 15876 38239 15885
rect 32576 15860 32618 15869
rect 32917 15836 32918 15876
rect 33151 15836 33152 15876
rect 33322 15836 33323 15876
rect 33589 15836 33590 15876
rect 33781 15836 33782 15876
rect 34016 15836 34017 15876
rect 34261 15836 34262 15876
rect 34741 15836 34742 15876
rect 34829 15836 34838 15876
rect 35029 15836 35030 15876
rect 35210 15836 35219 15876
rect 37412 15836 37421 15876
rect 38005 15836 38006 15876
rect 38197 15836 38198 15876
rect 8725 15827 8767 15836
rect 9013 15827 9055 15836
rect 9493 15827 9535 15836
rect 9685 15827 9727 15836
rect 10645 15827 10687 15836
rect 10733 15835 10791 15836
rect 11396 15835 11454 15836
rect 32245 15827 32287 15836
rect 32917 15827 32959 15836
rect 33151 15827 33193 15836
rect 33322 15827 33364 15836
rect 33589 15827 33631 15836
rect 33781 15827 33823 15836
rect 34016 15827 34058 15836
rect 34261 15827 34303 15836
rect 34741 15827 34783 15836
rect 34829 15835 34887 15836
rect 35029 15827 35071 15836
rect 35210 15835 35268 15836
rect 37412 15835 37470 15836
rect 38005 15827 38047 15836
rect 38197 15827 38239 15836
rect 10439 15792 10481 15801
rect 34340 15792 34398 15793
rect 34535 15792 34577 15801
rect 35492 15792 35550 15793
rect 37796 15792 37854 15793
rect 10439 15752 10440 15792
rect 34340 15752 34349 15792
rect 34535 15752 34536 15792
rect 35492 15752 35501 15792
rect 37796 15752 37805 15792
rect 10439 15743 10481 15752
rect 34340 15751 34398 15752
rect 34535 15743 34577 15752
rect 35492 15751 35550 15752
rect 37796 15751 37854 15752
rect 9493 15708 9535 15717
rect 10532 15708 10590 15709
rect 34628 15708 34686 15709
rect 9493 15668 9494 15708
rect 10532 15668 10541 15708
rect 34628 15668 34637 15708
rect 9493 15659 9535 15668
rect 10532 15667 10590 15668
rect 34628 15667 34686 15668
rect 8948 15372 9006 15373
rect 9493 15372 9535 15381
rect 11029 15372 11071 15381
rect 11396 15372 11454 15373
rect 37045 15372 37087 15381
rect 38245 15372 38287 15381
rect 8948 15332 8957 15372
rect 9493 15332 9494 15372
rect 11029 15332 11030 15372
rect 11396 15332 11405 15372
rect 37045 15332 37046 15372
rect 38245 15332 38246 15372
rect 8948 15331 9006 15332
rect 9493 15323 9535 15332
rect 11029 15323 11071 15332
rect 11396 15331 11454 15332
rect 37045 15323 37087 15332
rect 38245 15323 38287 15332
rect 36613 15288 36655 15297
rect 36613 15248 36614 15288
rect 36613 15239 36655 15248
rect 8437 15204 8479 15213
rect 8612 15204 8670 15205
rect 9113 15204 9171 15205
rect 9284 15204 9342 15205
rect 9589 15204 9631 15213
rect 9956 15204 10014 15205
rect 10069 15204 10111 15213
rect 10549 15204 10591 15213
rect 10837 15204 10879 15213
rect 33572 15204 33630 15205
rect 34436 15204 34494 15205
rect 34549 15204 34591 15213
rect 35012 15204 35070 15205
rect 35317 15204 35359 15213
rect 35588 15204 35646 15205
rect 36277 15204 36319 15213
rect 36425 15204 36483 15205
rect 36949 15204 36991 15213
rect 37140 15204 37182 15213
rect 37514 15204 37572 15205
rect 8437 15164 8438 15204
rect 8612 15164 8621 15204
rect 9113 15164 9122 15204
rect 9284 15164 9293 15204
rect 9589 15164 9590 15204
rect 9956 15164 9965 15204
rect 10069 15164 10070 15204
rect 10549 15164 10550 15204
rect 10837 15164 10838 15204
rect 33572 15164 33581 15204
rect 34436 15164 34445 15204
rect 34549 15164 34550 15204
rect 35012 15164 35021 15204
rect 35317 15164 35318 15204
rect 35588 15164 35597 15204
rect 36277 15164 36278 15204
rect 36425 15164 36434 15204
rect 36949 15164 36950 15204
rect 37140 15164 37141 15204
rect 8437 15155 8479 15164
rect 8612 15163 8670 15164
rect 9113 15163 9171 15164
rect 9284 15163 9342 15164
rect 9589 15155 9631 15164
rect 9956 15163 10014 15164
rect 10069 15155 10111 15164
rect 10549 15155 10591 15164
rect 10837 15155 10879 15164
rect 33572 15163 33630 15164
rect 34436 15163 34494 15164
rect 34549 15155 34591 15164
rect 35012 15163 35070 15164
rect 35317 15155 35359 15164
rect 35588 15163 35646 15164
rect 36277 15155 36319 15164
rect 36425 15163 36483 15164
rect 36949 15155 36991 15164
rect 37140 15155 37182 15164
rect 37333 15162 37375 15171
rect 37514 15164 37523 15204
rect 37514 15163 37572 15164
rect 11611 15120 11653 15129
rect 37333 15122 37334 15162
rect 32036 15120 32094 15121
rect 33956 15120 34014 15121
rect 11611 15080 11612 15120
rect 32036 15080 32045 15120
rect 33581 15080 33590 15120
rect 33956 15080 33965 15120
rect 37333 15113 37375 15122
rect 38485 15120 38527 15129
rect 38485 15080 38486 15120
rect 11611 15071 11653 15080
rect 32036 15079 32094 15080
rect 33956 15079 34014 15080
rect 38485 15071 38527 15080
rect 10244 15036 10302 15037
rect 35317 15036 35359 15045
rect 37717 15036 37759 15045
rect 10244 14996 10253 15036
rect 35317 14996 35318 15036
rect 37717 14996 37718 15036
rect 10244 14995 10302 14996
rect 35317 14987 35359 14996
rect 37717 14987 37759 14996
rect 8612 14952 8670 14953
rect 34724 14952 34782 14953
rect 37333 14952 37375 14961
rect 8612 14912 8621 14952
rect 34724 14912 34733 14952
rect 37333 14912 37334 14952
rect 8612 14911 8670 14912
rect 34724 14911 34782 14912
rect 37333 14903 37375 14912
rect 33205 14616 33247 14625
rect 35221 14616 35263 14625
rect 33205 14576 33206 14616
rect 35221 14576 35222 14616
rect 33205 14567 33247 14576
rect 35221 14567 35263 14576
rect 38197 14532 38239 14541
rect 38197 14492 38198 14532
rect 38197 14483 38239 14492
rect 9476 14448 9534 14449
rect 9685 14448 9727 14457
rect 13141 14448 13183 14457
rect 33812 14448 33870 14449
rect 34309 14448 34351 14457
rect 37124 14448 37182 14449
rect 9476 14408 9485 14448
rect 9685 14408 9686 14448
rect 13141 14408 13142 14448
rect 13372 14439 13418 14448
rect 9476 14407 9534 14408
rect 9685 14399 9727 14408
rect 13141 14399 13183 14408
rect 13372 14399 13373 14439
rect 33812 14408 33821 14448
rect 34309 14408 34310 14448
rect 37124 14408 37133 14448
rect 33812 14407 33870 14408
rect 34309 14399 34351 14408
rect 37124 14407 37182 14408
rect 13372 14390 13418 14399
rect 12644 14375 12702 14376
rect 8951 14364 9009 14365
rect 9344 14364 9386 14373
rect 9589 14364 9631 14373
rect 10436 14364 10494 14365
rect 10549 14364 10591 14373
rect 11701 14364 11743 14373
rect 11828 14364 11886 14365
rect 12197 14364 12255 14365
rect 12378 14364 12420 14373
rect 12482 14364 12540 14365
rect 8951 14324 8960 14364
rect 9344 14324 9345 14364
rect 9589 14324 9590 14364
rect 10436 14324 10445 14364
rect 10549 14324 10550 14364
rect 11701 14324 11702 14364
rect 11828 14324 11837 14364
rect 12197 14324 12206 14364
rect 12378 14324 12379 14364
rect 12482 14324 12491 14364
rect 12644 14335 12653 14375
rect 12766 14364 12824 14365
rect 13237 14364 13279 14373
rect 13477 14364 13519 14373
rect 13616 14364 13658 14373
rect 13796 14364 13854 14365
rect 14048 14364 14066 14373
rect 32533 14364 32575 14373
rect 32708 14364 32766 14365
rect 33205 14364 33247 14373
rect 33322 14364 33380 14365
rect 33493 14364 33535 14373
rect 33977 14364 34035 14365
rect 34145 14364 34203 14365
rect 36740 14364 36798 14365
rect 37268 14364 37326 14365
rect 37813 14364 37855 14373
rect 38005 14364 38047 14373
rect 38581 14364 38623 14373
rect 12644 14334 12702 14335
rect 12766 14324 12775 14364
rect 13237 14324 13238 14364
rect 13477 14324 13478 14364
rect 13616 14324 13617 14364
rect 13796 14324 13805 14364
rect 14048 14324 14049 14364
rect 32533 14324 32534 14364
rect 32708 14324 32717 14364
rect 33205 14324 33206 14364
rect 33322 14324 33331 14364
rect 33493 14324 33494 14364
rect 33977 14324 33986 14364
rect 34145 14324 34154 14364
rect 36740 14324 36749 14364
rect 37268 14324 37277 14364
rect 37813 14324 37814 14364
rect 38005 14324 38006 14364
rect 38581 14324 38582 14364
rect 8951 14323 9009 14324
rect 9344 14315 9386 14324
rect 9589 14315 9631 14324
rect 10436 14323 10494 14324
rect 10549 14315 10591 14324
rect 11701 14315 11743 14324
rect 11828 14323 11886 14324
rect 12197 14323 12255 14324
rect 12378 14315 12420 14324
rect 12482 14323 12540 14324
rect 12766 14323 12824 14324
rect 13237 14315 13279 14324
rect 13477 14315 13519 14324
rect 13616 14315 13658 14324
rect 13796 14323 13854 14324
rect 14048 14315 14066 14324
rect 32533 14315 32575 14324
rect 32708 14323 32766 14324
rect 33205 14315 33247 14324
rect 33322 14323 33380 14324
rect 33493 14315 33535 14324
rect 33977 14323 34035 14324
rect 34145 14323 34203 14324
rect 36740 14323 36798 14324
rect 37268 14323 37326 14324
rect 37813 14315 37855 14324
rect 38005 14315 38047 14324
rect 38581 14315 38623 14324
rect 33024 14280 33066 14289
rect 34820 14280 34878 14281
rect 33024 14240 33025 14280
rect 34820 14240 34829 14280
rect 33024 14231 33066 14240
rect 34820 14239 34878 14240
rect 8756 14196 8814 14197
rect 10837 14196 10879 14205
rect 11989 14196 12031 14205
rect 12260 14196 12318 14197
rect 13717 14196 13759 14205
rect 32804 14196 32862 14197
rect 32917 14196 32959 14205
rect 37477 14196 37519 14205
rect 37988 14196 38046 14197
rect 8756 14156 8765 14196
rect 10837 14156 10838 14196
rect 11989 14156 11990 14196
rect 12260 14156 12269 14196
rect 13717 14156 13718 14196
rect 32804 14156 32813 14196
rect 32917 14156 32918 14196
rect 37477 14156 37478 14196
rect 37988 14156 37997 14196
rect 8756 14155 8814 14156
rect 10837 14147 10879 14156
rect 11989 14147 12031 14156
rect 12260 14155 12318 14156
rect 13717 14147 13759 14156
rect 32804 14155 32862 14156
rect 32917 14147 32959 14156
rect 37477 14147 37519 14156
rect 37988 14155 38046 14156
rect 8629 13860 8671 13869
rect 9397 13860 9439 13869
rect 9781 13860 9823 13869
rect 11684 13860 11742 13861
rect 11972 13860 12030 13861
rect 13333 13860 13375 13869
rect 13717 13860 13759 13869
rect 37141 13860 37183 13869
rect 8629 13820 8630 13860
rect 9397 13820 9398 13860
rect 9781 13820 9782 13860
rect 11684 13820 11693 13860
rect 11972 13820 11981 13860
rect 13333 13820 13334 13860
rect 13717 13820 13718 13860
rect 37141 13820 37142 13860
rect 8629 13811 8671 13820
rect 9397 13811 9439 13820
rect 9781 13811 9823 13820
rect 11684 13819 11742 13820
rect 11972 13819 12030 13820
rect 13333 13811 13375 13820
rect 13717 13811 13759 13820
rect 37141 13811 37183 13820
rect 9891 13776 9933 13785
rect 10340 13776 10398 13777
rect 37525 13776 37567 13785
rect 9891 13736 9892 13776
rect 10340 13736 10349 13776
rect 37525 13736 37526 13776
rect 9891 13727 9933 13736
rect 10340 13735 10398 13736
rect 37525 13727 37567 13736
rect 8341 13692 8383 13701
rect 8468 13692 8526 13693
rect 8996 13692 9054 13693
rect 9109 13692 9151 13701
rect 9572 13692 9630 13693
rect 9685 13692 9727 13701
rect 10016 13692 10058 13701
rect 10261 13692 10303 13701
rect 11360 13692 11402 13701
rect 11492 13692 11550 13693
rect 11605 13692 11647 13701
rect 12181 13692 12223 13701
rect 12469 13692 12511 13701
rect 12661 13692 12703 13701
rect 12853 13692 12895 13701
rect 13237 13692 13279 13701
rect 13412 13692 13470 13693
rect 13624 13692 13682 13693
rect 13796 13692 13854 13693
rect 32804 13692 32862 13693
rect 33397 13692 33439 13701
rect 33589 13692 33631 13701
rect 34148 13692 34206 13693
rect 37045 13692 37087 13701
rect 37218 13692 37260 13701
rect 37429 13692 37471 13701
rect 37621 13692 37663 13701
rect 8341 13652 8342 13692
rect 8468 13652 8477 13692
rect 8996 13652 9005 13692
rect 9109 13652 9110 13692
rect 9572 13652 9581 13692
rect 9685 13652 9686 13692
rect 10016 13652 10017 13692
rect 10261 13652 10262 13692
rect 11360 13652 11361 13692
rect 11492 13652 11501 13692
rect 11605 13652 11606 13692
rect 12181 13652 12182 13692
rect 12469 13652 12470 13692
rect 12661 13652 12662 13692
rect 12853 13652 12854 13692
rect 13237 13652 13238 13692
rect 13412 13652 13421 13692
rect 13624 13652 13633 13692
rect 13796 13652 13805 13692
rect 32804 13652 32813 13692
rect 33397 13652 33398 13692
rect 33589 13652 33590 13692
rect 34148 13652 34157 13692
rect 37045 13652 37046 13692
rect 37218 13652 37219 13692
rect 37429 13652 37430 13692
rect 37621 13652 37622 13692
rect 8341 13643 8383 13652
rect 8468 13651 8526 13652
rect 8996 13651 9054 13652
rect 9109 13643 9151 13652
rect 9572 13651 9630 13652
rect 9685 13643 9727 13652
rect 10016 13643 10058 13652
rect 10261 13643 10303 13652
rect 11360 13643 11402 13652
rect 11492 13651 11550 13652
rect 11605 13643 11647 13652
rect 12181 13643 12223 13652
rect 12469 13643 12511 13652
rect 12661 13643 12703 13652
rect 12853 13643 12895 13652
rect 13237 13643 13279 13652
rect 13412 13651 13470 13652
rect 13624 13651 13682 13652
rect 13796 13651 13854 13652
rect 32804 13651 32862 13652
rect 33397 13643 33439 13652
rect 33589 13643 33631 13652
rect 34148 13651 34206 13652
rect 37045 13643 37087 13652
rect 37218 13643 37260 13652
rect 37429 13643 37471 13652
rect 37621 13643 37663 13652
rect 10148 13608 10206 13609
rect 33188 13608 33246 13609
rect 33781 13608 33823 13617
rect 35701 13608 35743 13617
rect 10148 13568 10157 13608
rect 33188 13568 33197 13608
rect 33781 13568 33782 13608
rect 35701 13568 35702 13608
rect 10148 13567 10206 13568
rect 33188 13567 33246 13568
rect 33781 13559 33823 13568
rect 35701 13559 35743 13568
rect 33397 13524 33439 13533
rect 36277 13524 36319 13533
rect 36661 13524 36703 13533
rect 37909 13524 37951 13533
rect 38293 13524 38335 13533
rect 33397 13484 33398 13524
rect 36277 13484 36278 13524
rect 36661 13484 36662 13524
rect 37909 13484 37910 13524
rect 38293 13484 38294 13524
rect 33397 13475 33439 13484
rect 36277 13475 36319 13484
rect 36661 13475 36703 13484
rect 37909 13475 37951 13484
rect 38293 13475 38335 13484
rect 12661 13440 12703 13449
rect 36085 13440 36127 13449
rect 12661 13400 12662 13440
rect 36085 13400 36086 13440
rect 12661 13391 12703 13400
rect 36085 13391 36127 13400
rect 8821 13104 8863 13113
rect 9685 13104 9727 13113
rect 12181 13104 12223 13113
rect 13045 13104 13087 13113
rect 14005 13104 14047 13113
rect 34549 13104 34591 13113
rect 35989 13104 36031 13113
rect 36548 13104 36606 13105
rect 37717 13104 37759 13113
rect 38101 13104 38143 13113
rect 8821 13064 8822 13104
rect 9685 13064 9686 13104
rect 12181 13064 12182 13104
rect 13045 13064 13046 13104
rect 14005 13064 14006 13104
rect 34549 13064 34550 13104
rect 35989 13064 35990 13104
rect 36548 13064 36557 13104
rect 37717 13064 37718 13104
rect 38101 13064 38102 13104
rect 8821 13055 8863 13064
rect 9685 13055 9727 13064
rect 12181 13055 12223 13064
rect 13045 13055 13087 13064
rect 14005 13055 14047 13064
rect 34549 13055 34591 13064
rect 35989 13055 36031 13064
rect 36548 13063 36606 13064
rect 37717 13055 37759 13064
rect 38101 13055 38143 13064
rect 10741 13020 10783 13029
rect 13525 13020 13567 13029
rect 36757 13020 36799 13029
rect 38389 13020 38431 13029
rect 10741 12980 10742 13020
rect 13525 12980 13526 13020
rect 36757 12980 36758 13020
rect 38389 12980 38390 13020
rect 10741 12971 10783 12980
rect 13525 12971 13567 12980
rect 36757 12971 36799 12980
rect 38389 12971 38431 12980
rect 9397 12936 9439 12945
rect 32996 12936 33054 12937
rect 34651 12936 34693 12945
rect 9397 12896 9398 12936
rect 32996 12896 33005 12936
rect 34651 12896 34652 12936
rect 9397 12887 9439 12896
rect 32996 12895 33054 12896
rect 11897 12885 11939 12894
rect 34651 12887 34693 12896
rect 8341 12852 8383 12861
rect 8516 12852 8574 12853
rect 8716 12852 8774 12853
rect 8916 12852 8958 12861
rect 9061 12852 9103 12861
rect 9188 12852 9246 12853
rect 9301 12852 9343 12861
rect 9589 12852 9631 12861
rect 9781 12852 9823 12861
rect 10069 12852 10111 12861
rect 10549 12852 10591 12861
rect 10933 12852 10975 12861
rect 11317 12852 11359 12861
rect 11780 12852 11838 12853
rect 8341 12812 8342 12852
rect 8516 12812 8525 12852
rect 8716 12812 8725 12852
rect 8916 12812 8917 12852
rect 9061 12812 9062 12852
rect 9188 12812 9197 12852
rect 9301 12812 9302 12852
rect 9589 12812 9590 12852
rect 9781 12812 9782 12852
rect 10069 12812 10070 12852
rect 10549 12812 10550 12852
rect 10933 12812 10934 12852
rect 11317 12812 11318 12852
rect 11780 12812 11789 12852
rect 11897 12845 11898 12885
rect 12373 12852 12415 12861
rect 12565 12852 12607 12861
rect 12740 12852 12798 12853
rect 13333 12852 13375 12861
rect 13700 12852 13758 12853
rect 32533 12852 32575 12861
rect 33397 12852 33439 12861
rect 33877 12852 33919 12861
rect 34261 12852 34303 12861
rect 34741 12852 34783 12861
rect 35365 12852 35407 12861
rect 35509 12852 35551 12861
rect 35989 12852 36031 12861
rect 36181 12852 36223 12861
rect 36373 12852 36415 12861
rect 36542 12852 36584 12861
rect 36757 12852 36799 12861
rect 36949 12852 36991 12861
rect 37141 12852 37183 12861
rect 37333 12852 37375 12861
rect 37621 12852 37663 12861
rect 37813 12852 37855 12861
rect 38005 12852 38047 12861
rect 38197 12852 38239 12861
rect 11897 12836 11939 12845
rect 12373 12812 12374 12852
rect 12565 12812 12566 12852
rect 12740 12812 12749 12852
rect 13333 12812 13334 12852
rect 13700 12812 13709 12852
rect 32533 12812 32534 12852
rect 33397 12812 33398 12852
rect 33877 12812 33878 12852
rect 34261 12812 34262 12852
rect 34741 12812 34742 12852
rect 35365 12812 35366 12852
rect 35509 12812 35510 12852
rect 35989 12812 35990 12852
rect 36181 12812 36182 12852
rect 36373 12812 36374 12852
rect 36542 12812 36543 12852
rect 36757 12812 36758 12852
rect 36949 12812 36950 12852
rect 37141 12812 37142 12852
rect 37333 12812 37334 12852
rect 37621 12812 37622 12852
rect 37813 12812 37814 12852
rect 38005 12812 38006 12852
rect 38197 12812 38198 12852
rect 8341 12803 8383 12812
rect 8516 12811 8574 12812
rect 8716 12811 8774 12812
rect 8916 12803 8958 12812
rect 9061 12803 9103 12812
rect 9188 12811 9246 12812
rect 9301 12803 9343 12812
rect 9589 12803 9631 12812
rect 9781 12803 9823 12812
rect 10069 12803 10111 12812
rect 10549 12803 10591 12812
rect 10933 12803 10975 12812
rect 11317 12803 11359 12812
rect 11780 12811 11838 12812
rect 12373 12803 12415 12812
rect 12565 12803 12607 12812
rect 12740 12811 12798 12812
rect 13333 12803 13375 12812
rect 13700 12811 13758 12812
rect 32533 12803 32575 12812
rect 33397 12803 33439 12812
rect 33877 12803 33919 12812
rect 34261 12803 34303 12812
rect 34741 12803 34783 12812
rect 35365 12803 35407 12812
rect 35509 12803 35551 12812
rect 35989 12803 36031 12812
rect 36181 12803 36223 12812
rect 36373 12803 36415 12812
rect 36542 12803 36584 12812
rect 36757 12803 36799 12812
rect 36949 12803 36991 12812
rect 37141 12803 37183 12812
rect 37333 12803 37375 12812
rect 37621 12803 37663 12812
rect 37813 12803 37855 12812
rect 38005 12803 38047 12812
rect 38197 12803 38239 12812
rect 9685 12768 9727 12777
rect 12469 12768 12511 12777
rect 12853 12768 12895 12777
rect 13059 12768 13101 12777
rect 13813 12768 13855 12777
rect 14019 12768 14061 12777
rect 37237 12768 37279 12777
rect 9685 12728 9686 12768
rect 12469 12728 12470 12768
rect 12853 12728 12854 12768
rect 13059 12728 13060 12768
rect 13813 12728 13814 12768
rect 14019 12728 14020 12768
rect 37237 12728 37238 12768
rect 9685 12719 9727 12728
rect 12469 12719 12511 12728
rect 12853 12719 12895 12728
rect 13059 12719 13101 12728
rect 13813 12719 13855 12728
rect 14019 12719 14061 12728
rect 37237 12719 37279 12728
rect 8437 12684 8479 12693
rect 9956 12684 10014 12685
rect 10261 12684 10303 12693
rect 10436 12684 10494 12685
rect 11413 12684 11455 12693
rect 13220 12684 13278 12685
rect 32341 12684 32383 12693
rect 33764 12684 33822 12685
rect 35204 12684 35262 12685
rect 8437 12644 8438 12684
rect 9956 12644 9965 12684
rect 10261 12644 10262 12684
rect 10436 12644 10445 12684
rect 11413 12644 11414 12684
rect 11692 12675 11738 12684
rect 8437 12635 8479 12644
rect 9956 12643 10014 12644
rect 10261 12635 10303 12644
rect 10436 12643 10494 12644
rect 11413 12635 11455 12644
rect 11692 12635 11693 12675
rect 13220 12644 13229 12684
rect 32341 12644 32342 12684
rect 33764 12644 33773 12684
rect 35204 12644 35213 12684
rect 13220 12643 13278 12644
rect 32341 12635 32383 12644
rect 33764 12643 33822 12644
rect 35204 12643 35262 12644
rect 11692 12626 11738 12635
rect 11204 12390 11262 12391
rect 9205 12348 9247 12357
rect 10165 12348 10207 12357
rect 11204 12350 11213 12390
rect 11204 12349 11262 12350
rect 12548 12348 12606 12349
rect 13316 12348 13374 12349
rect 32804 12348 32862 12349
rect 34069 12348 34111 12357
rect 34532 12348 34590 12349
rect 36757 12348 36799 12357
rect 37045 12348 37087 12357
rect 37525 12348 37567 12357
rect 9205 12308 9206 12348
rect 10165 12308 10166 12348
rect 12548 12308 12557 12348
rect 13316 12308 13325 12348
rect 32804 12308 32813 12348
rect 34069 12308 34070 12348
rect 34532 12308 34541 12348
rect 36757 12308 36758 12348
rect 37045 12308 37046 12348
rect 37525 12308 37526 12348
rect 9205 12299 9247 12308
rect 10165 12299 10207 12308
rect 12548 12307 12606 12308
rect 13316 12307 13374 12308
rect 32804 12307 32862 12308
rect 34069 12299 34111 12308
rect 34532 12307 34590 12308
rect 36757 12299 36799 12308
rect 37045 12299 37087 12308
rect 37525 12299 37567 12308
rect 8341 12264 8383 12273
rect 8341 12224 8342 12264
rect 8341 12215 8383 12224
rect 37230 12199 37272 12208
rect 8245 12180 8287 12189
rect 8437 12180 8479 12189
rect 8804 12180 8862 12181
rect 8917 12180 8959 12189
rect 9877 12180 9919 12189
rect 10004 12180 10062 12181
rect 10532 12180 10590 12181
rect 10645 12180 10687 12189
rect 11242 12180 11284 12189
rect 11540 12180 11598 12181
rect 12236 12180 12294 12181
rect 12469 12180 12511 12189
rect 12992 12180 13034 12189
rect 13237 12180 13279 12189
rect 32039 12180 32081 12189
rect 32149 12180 32191 12189
rect 32492 12180 32550 12181
rect 32725 12180 32767 12189
rect 33013 12180 33055 12189
rect 33301 12180 33343 12189
rect 33668 12180 33726 12181
rect 33781 12180 33823 12189
rect 34837 12180 34879 12189
rect 35989 12180 36031 12189
rect 36661 12180 36703 12189
rect 36836 12180 36894 12181
rect 37045 12180 37087 12189
rect 8245 12140 8246 12180
rect 8437 12140 8438 12180
rect 8804 12140 8813 12180
rect 8917 12140 8918 12180
rect 9877 12140 9878 12180
rect 10004 12140 10013 12180
rect 10532 12140 10541 12180
rect 10645 12140 10646 12180
rect 11242 12140 11243 12180
rect 11540 12140 11549 12180
rect 12236 12140 12245 12180
rect 12469 12140 12470 12180
rect 12992 12140 12993 12180
rect 13237 12140 13238 12180
rect 32039 12140 32040 12180
rect 32149 12140 32150 12180
rect 32492 12140 32501 12180
rect 32725 12140 32726 12180
rect 33013 12140 33014 12180
rect 33301 12140 33302 12180
rect 33668 12140 33677 12180
rect 33781 12140 33782 12180
rect 34837 12140 34838 12180
rect 35989 12140 35990 12180
rect 36661 12140 36662 12180
rect 36836 12140 36845 12180
rect 37045 12140 37046 12180
rect 37230 12159 37231 12199
rect 37621 12180 37663 12189
rect 37230 12150 37272 12159
rect 8245 12131 8287 12140
rect 8437 12131 8479 12140
rect 8804 12139 8862 12140
rect 8917 12131 8959 12140
rect 9877 12131 9919 12140
rect 10004 12139 10062 12140
rect 10532 12139 10590 12140
rect 10645 12131 10687 12140
rect 11242 12131 11284 12140
rect 11540 12139 11598 12140
rect 12236 12139 12294 12140
rect 12469 12131 12511 12140
rect 12992 12131 13034 12140
rect 13237 12131 13279 12140
rect 32039 12131 32081 12140
rect 32149 12131 32191 12140
rect 32492 12139 32550 12140
rect 32338 12138 32396 12139
rect 11413 12096 11455 12105
rect 32338 12098 32347 12138
rect 32725 12131 32767 12140
rect 33013 12131 33055 12140
rect 33301 12131 33343 12140
rect 33668 12139 33726 12140
rect 33781 12131 33823 12140
rect 34837 12131 34879 12140
rect 35989 12131 36031 12140
rect 36661 12131 36703 12140
rect 36836 12139 36894 12140
rect 37045 12131 37087 12140
rect 37429 12138 37471 12147
rect 37621 12140 37622 12180
rect 32338 12097 32396 12098
rect 12356 12096 12414 12097
rect 13124 12096 13182 12097
rect 32612 12096 32670 12097
rect 34747 12096 34789 12105
rect 37429 12098 37430 12138
rect 37621 12131 37663 12140
rect 11413 12056 11414 12096
rect 12356 12056 12365 12096
rect 13124 12056 13133 12096
rect 32612 12056 32621 12096
rect 34747 12056 34748 12096
rect 37429 12089 37471 12098
rect 11413 12047 11455 12056
rect 12356 12055 12414 12056
rect 13124 12055 13182 12056
rect 32612 12055 32670 12056
rect 34747 12047 34789 12056
rect 11317 12012 11359 12021
rect 32245 12012 32287 12021
rect 36277 12012 36319 12021
rect 37813 12012 37855 12021
rect 38197 12012 38239 12021
rect 11317 11972 11318 12012
rect 32245 11972 32246 12012
rect 36277 11972 36278 12012
rect 37813 11972 37814 12012
rect 38197 11972 38198 12012
rect 11317 11963 11359 11972
rect 32245 11963 32287 11972
rect 36277 11963 36319 11972
rect 37813 11963 37855 11972
rect 38197 11963 38239 11972
rect 10820 11928 10878 11929
rect 33013 11928 33055 11937
rect 35588 11928 35646 11929
rect 10820 11888 10829 11928
rect 33013 11888 33014 11928
rect 35588 11888 35597 11928
rect 10820 11887 10878 11888
rect 33013 11879 33055 11888
rect 35588 11887 35646 11888
rect 9061 11592 9103 11601
rect 10741 11592 10783 11601
rect 12644 11592 12702 11593
rect 13813 11592 13855 11601
rect 32437 11592 32479 11601
rect 35204 11592 35262 11593
rect 9061 11552 9062 11592
rect 10741 11552 10742 11592
rect 12644 11552 12653 11592
rect 13813 11552 13814 11592
rect 32437 11552 32438 11592
rect 35204 11552 35213 11592
rect 9061 11543 9103 11552
rect 10741 11543 10783 11552
rect 12644 11551 12702 11552
rect 13813 11543 13855 11552
rect 32437 11543 32479 11552
rect 35204 11551 35262 11552
rect 9668 11508 9726 11509
rect 35893 11508 35935 11517
rect 37813 11508 37855 11517
rect 38197 11508 38239 11517
rect 9668 11468 9677 11508
rect 35893 11468 35894 11508
rect 37813 11468 37814 11508
rect 38197 11468 38198 11508
rect 9668 11467 9726 11468
rect 35893 11459 35935 11468
rect 37813 11459 37855 11468
rect 38197 11459 38239 11468
rect 10052 11424 10110 11425
rect 11012 11424 11070 11425
rect 11221 11424 11263 11433
rect 32539 11424 32581 11433
rect 33403 11424 33445 11433
rect 10052 11384 10061 11424
rect 11012 11384 11021 11424
rect 11221 11384 11222 11424
rect 32539 11384 32540 11424
rect 33403 11384 33404 11424
rect 10052 11383 10110 11384
rect 11012 11383 11070 11384
rect 11221 11375 11263 11384
rect 32539 11375 32581 11384
rect 33403 11375 33445 11384
rect 8053 11340 8095 11349
rect 8245 11340 8287 11349
rect 8437 11340 8479 11349
rect 8821 11340 8863 11349
rect 9380 11340 9438 11341
rect 9493 11340 9535 11349
rect 9925 11340 9967 11349
rect 10165 11340 10207 11349
rect 10436 11340 10494 11341
rect 10549 11340 10591 11349
rect 10892 11340 10950 11341
rect 11125 11340 11167 11349
rect 11413 11340 11455 11349
rect 11797 11340 11839 11349
rect 12356 11340 12414 11341
rect 12469 11340 12511 11349
rect 12949 11340 12991 11349
rect 13237 11340 13279 11349
rect 13861 11340 13903 11349
rect 14005 11340 14047 11349
rect 32629 11340 32671 11349
rect 33493 11340 33535 11349
rect 34261 11340 34303 11349
rect 34549 11340 34591 11349
rect 34724 11340 34782 11341
rect 35029 11340 35071 11349
rect 35413 11340 35455 11349
rect 35501 11340 35559 11341
rect 36757 11340 36799 11349
rect 8053 11300 8054 11340
rect 8245 11300 8246 11340
rect 8437 11300 8438 11340
rect 8821 11300 8822 11340
rect 9380 11300 9389 11340
rect 9493 11300 9494 11340
rect 9925 11300 9926 11340
rect 10165 11300 10166 11340
rect 10436 11300 10445 11340
rect 10549 11300 10550 11340
rect 10892 11300 10901 11340
rect 11125 11300 11126 11340
rect 11413 11300 11414 11340
rect 11797 11300 11798 11340
rect 12356 11300 12365 11340
rect 12469 11300 12470 11340
rect 12949 11300 12950 11340
rect 13237 11300 13238 11340
rect 13861 11300 13862 11340
rect 14005 11300 14006 11340
rect 32629 11300 32630 11340
rect 33493 11300 33494 11340
rect 34261 11300 34262 11340
rect 34549 11300 34550 11340
rect 34724 11300 34733 11340
rect 35029 11300 35030 11340
rect 35413 11300 35414 11340
rect 35501 11300 35510 11340
rect 36757 11300 36758 11340
rect 8053 11291 8095 11300
rect 8245 11291 8287 11300
rect 8437 11291 8479 11300
rect 8821 11291 8863 11300
rect 9380 11299 9438 11300
rect 9493 11291 9535 11300
rect 9925 11291 9967 11300
rect 10165 11291 10207 11300
rect 10436 11299 10494 11300
rect 10549 11291 10591 11300
rect 10892 11299 10950 11300
rect 11125 11291 11167 11300
rect 11413 11291 11455 11300
rect 11797 11291 11839 11300
rect 12356 11299 12414 11300
rect 12469 11291 12511 11300
rect 12949 11291 12991 11300
rect 13237 11291 13279 11300
rect 13861 11291 13903 11300
rect 14005 11291 14047 11300
rect 32629 11291 32671 11300
rect 33493 11291 33535 11300
rect 34261 11291 34303 11300
rect 34549 11291 34591 11300
rect 34724 11299 34782 11300
rect 35029 11291 35071 11300
rect 35413 11291 35455 11300
rect 35501 11299 35559 11300
rect 36757 11291 36799 11300
rect 10244 11256 10302 11257
rect 10755 11256 10797 11265
rect 13573 11256 13615 11265
rect 34933 11256 34975 11265
rect 35207 11256 35249 11265
rect 10244 11216 10253 11256
rect 10755 11216 10756 11256
rect 13573 11216 13574 11256
rect 34933 11216 34934 11256
rect 35207 11216 35208 11256
rect 10244 11215 10302 11216
rect 10755 11207 10797 11216
rect 13573 11207 13615 11216
rect 34933 11207 34975 11216
rect 35207 11207 35249 11216
rect 8228 11172 8286 11173
rect 11893 11172 11935 11181
rect 33188 11172 33246 11173
rect 34052 11172 34110 11173
rect 35413 11172 35455 11181
rect 36085 11172 36127 11181
rect 8228 11132 8237 11172
rect 11893 11132 11894 11172
rect 33188 11132 33197 11172
rect 34052 11132 34061 11172
rect 35413 11132 35414 11172
rect 36085 11132 36086 11172
rect 8228 11131 8286 11132
rect 11893 11123 11935 11132
rect 33188 11131 33246 11132
rect 34052 11131 34110 11132
rect 35413 11123 35455 11132
rect 36085 11123 36127 11132
rect 8341 10836 8383 10845
rect 9205 10836 9247 10845
rect 11605 10836 11647 10845
rect 12164 10836 12222 10837
rect 33236 10836 33294 10837
rect 34837 10836 34879 10845
rect 8341 10796 8342 10836
rect 9205 10796 9206 10836
rect 11605 10796 11606 10836
rect 12164 10796 12173 10836
rect 33236 10796 33245 10836
rect 34837 10796 34838 10836
rect 8341 10787 8383 10796
rect 9205 10787 9247 10796
rect 11605 10787 11647 10796
rect 12164 10795 12222 10796
rect 33236 10795 33294 10796
rect 34837 10787 34879 10796
rect 9781 10752 9823 10761
rect 13717 10752 13759 10761
rect 32615 10752 32657 10761
rect 32708 10752 32766 10753
rect 33685 10752 33727 10761
rect 34357 10752 34399 10761
rect 9781 10712 9782 10752
rect 13717 10712 13718 10752
rect 32615 10712 32616 10752
rect 32708 10712 32717 10752
rect 33685 10712 33686 10752
rect 34357 10712 34358 10752
rect 9781 10703 9823 10712
rect 13717 10703 13759 10712
rect 32615 10703 32657 10712
rect 32708 10711 32766 10712
rect 33685 10703 33727 10712
rect 34357 10703 34399 10712
rect 8341 10668 8383 10677
rect 8533 10668 8575 10677
rect 8725 10668 8767 10677
rect 9109 10668 9151 10677
rect 9685 10668 9727 10677
rect 9881 10668 9923 10677
rect 10069 10668 10111 10677
rect 10357 10668 10399 10677
rect 10496 10668 10538 10677
rect 10741 10668 10783 10677
rect 11029 10668 11071 10677
rect 11146 10668 11204 10669
rect 11317 10668 11359 10677
rect 11509 10668 11551 10677
rect 11701 10668 11743 10677
rect 12085 10668 12127 10677
rect 12512 10668 12554 10677
rect 12757 10668 12799 10677
rect 13045 10668 13087 10677
rect 13220 10668 13278 10669
rect 13621 10668 13663 10677
rect 13813 10668 13855 10677
rect 32005 10668 32047 10677
rect 32149 10668 32191 10677
rect 32821 10668 32863 10677
rect 33401 10668 33459 10669
rect 33572 10668 33614 10677
rect 33776 10668 33834 10669
rect 33973 10668 34015 10677
rect 34148 10668 34206 10669
rect 34453 10668 34495 10677
rect 34682 10668 34740 10669
rect 36740 10668 36798 10669
rect 8341 10628 8342 10668
rect 8533 10628 8534 10668
rect 8725 10628 8726 10668
rect 9109 10628 9110 10668
rect 9685 10628 9686 10668
rect 9881 10628 9882 10668
rect 10069 10628 10070 10668
rect 10357 10628 10358 10668
rect 10496 10628 10497 10668
rect 10741 10628 10742 10668
rect 11029 10628 11030 10668
rect 11146 10628 11155 10668
rect 11317 10628 11318 10668
rect 11509 10628 11510 10668
rect 11701 10628 11702 10668
rect 8341 10619 8383 10628
rect 8533 10619 8575 10628
rect 8725 10619 8767 10628
rect 9109 10619 9151 10628
rect 9685 10619 9727 10628
rect 9881 10619 9923 10628
rect 10069 10619 10111 10628
rect 10357 10619 10399 10628
rect 10496 10619 10538 10628
rect 10741 10619 10783 10628
rect 11029 10619 11071 10628
rect 11146 10627 11204 10628
rect 11317 10619 11359 10628
rect 11509 10619 11551 10628
rect 11701 10619 11743 10628
rect 11845 10626 11887 10635
rect 12085 10628 12086 10668
rect 12512 10628 12513 10668
rect 12757 10628 12758 10668
rect 13045 10628 13046 10668
rect 13220 10628 13229 10668
rect 13621 10628 13622 10668
rect 13813 10628 13814 10668
rect 32005 10628 32006 10668
rect 32149 10628 32150 10668
rect 32821 10628 32822 10668
rect 32917 10659 32959 10668
rect 10622 10584 10664 10593
rect 10837 10584 10879 10593
rect 11845 10586 11846 10626
rect 12085 10619 12127 10628
rect 12512 10619 12554 10628
rect 12757 10619 12799 10628
rect 13045 10619 13087 10628
rect 13220 10627 13278 10628
rect 13621 10619 13663 10628
rect 13813 10619 13855 10628
rect 32005 10619 32047 10628
rect 32149 10619 32191 10628
rect 32821 10619 32863 10628
rect 32917 10619 32918 10659
rect 33401 10628 33410 10668
rect 33572 10628 33573 10668
rect 33776 10628 33785 10668
rect 33973 10628 33974 10668
rect 34148 10628 34157 10668
rect 34453 10628 34454 10668
rect 34682 10628 34691 10668
rect 36740 10628 36749 10668
rect 33401 10627 33459 10628
rect 33572 10619 33614 10628
rect 33776 10627 33834 10628
rect 33973 10619 34015 10628
rect 34148 10627 34206 10628
rect 34453 10619 34495 10628
rect 34682 10627 34740 10628
rect 36740 10627 36798 10628
rect 32917 10610 32959 10619
rect 10622 10544 10623 10584
rect 10837 10544 10838 10584
rect 11845 10577 11887 10586
rect 11972 10584 12030 10585
rect 12644 10584 12702 10585
rect 12853 10584 12895 10593
rect 37124 10584 37182 10585
rect 11972 10544 11981 10584
rect 12644 10544 12653 10584
rect 12853 10544 12854 10584
rect 34588 10575 34634 10584
rect 10622 10535 10664 10544
rect 10837 10535 10879 10544
rect 11972 10543 12030 10544
rect 12644 10543 12702 10544
rect 12853 10535 12895 10544
rect 34588 10535 34589 10575
rect 35885 10544 35894 10584
rect 37124 10544 37133 10584
rect 37124 10543 37182 10544
rect 34588 10526 34634 10535
rect 13273 10500 13315 10509
rect 34148 10500 34206 10501
rect 13273 10460 13274 10500
rect 34148 10460 34157 10500
rect 13273 10451 13315 10460
rect 34148 10459 34206 10460
rect 10069 10416 10111 10425
rect 11029 10416 11071 10425
rect 10069 10376 10070 10416
rect 11029 10376 11030 10416
rect 10069 10367 10111 10376
rect 11029 10367 11071 10376
rect 8437 10080 8479 10089
rect 10724 10080 10782 10081
rect 13765 10080 13807 10089
rect 35605 10080 35647 10089
rect 8437 10040 8438 10080
rect 10724 10040 10733 10080
rect 13765 10040 13766 10080
rect 35605 10040 35606 10080
rect 8437 10031 8479 10040
rect 10724 10039 10782 10040
rect 13765 10031 13807 10040
rect 35605 10031 35647 10040
rect 8053 9996 8095 10005
rect 35797 9996 35839 10005
rect 8053 9956 8054 9996
rect 35797 9956 35798 9996
rect 8053 9947 8095 9956
rect 35797 9947 35839 9956
rect 10340 9912 10398 9913
rect 12187 9912 12229 9921
rect 32539 9912 32581 9921
rect 33349 9912 33391 9921
rect 9389 9872 9398 9912
rect 10340 9872 10349 9912
rect 12187 9872 12188 9912
rect 32539 9872 32540 9912
rect 33349 9872 33350 9912
rect 10340 9871 10398 9872
rect 12187 9863 12229 9872
rect 32539 9863 32581 9872
rect 33349 9863 33391 9872
rect 9956 9828 10014 9829
rect 10730 9828 10772 9837
rect 11021 9828 11079 9829
rect 11221 9828 11263 9837
rect 11605 9828 11647 9837
rect 12277 9828 12319 9837
rect 12853 9828 12895 9837
rect 13076 9828 13134 9829
rect 13429 9828 13471 9837
rect 14005 9828 14047 9837
rect 32629 9828 32671 9837
rect 33205 9828 33247 9837
rect 34165 9828 34207 9837
rect 34549 9828 34591 9837
rect 34637 9828 34695 9829
rect 34933 9828 34975 9837
rect 36469 9828 36511 9837
rect 9956 9788 9965 9828
rect 10730 9788 10731 9828
rect 11021 9788 11030 9828
rect 11221 9788 11222 9828
rect 11605 9788 11606 9828
rect 12277 9788 12278 9828
rect 12853 9788 12854 9828
rect 13076 9788 13085 9828
rect 13429 9788 13430 9828
rect 14005 9788 14006 9828
rect 32629 9788 32630 9828
rect 33205 9788 33206 9828
rect 34165 9788 34166 9828
rect 34549 9788 34550 9828
rect 34637 9788 34646 9828
rect 34933 9788 34934 9828
rect 36469 9788 36470 9828
rect 9956 9787 10014 9788
rect 10730 9779 10772 9788
rect 11021 9787 11079 9788
rect 11221 9779 11263 9788
rect 11605 9779 11647 9788
rect 12277 9779 12319 9788
rect 12853 9779 12895 9788
rect 13076 9787 13134 9788
rect 13429 9779 13471 9788
rect 14005 9779 14047 9788
rect 32629 9779 32671 9788
rect 33205 9779 33247 9788
rect 34165 9779 34207 9788
rect 34549 9779 34591 9788
rect 34637 9787 34695 9788
rect 34933 9779 34975 9788
rect 36469 9779 36511 9788
rect 34343 9744 34385 9753
rect 34436 9744 34494 9745
rect 34343 9704 34344 9744
rect 34436 9704 34445 9744
rect 34343 9695 34385 9704
rect 34436 9703 34494 9704
rect 10933 9660 10975 9669
rect 11701 9660 11743 9669
rect 11972 9660 12030 9661
rect 12709 9660 12751 9669
rect 13525 9660 13567 9669
rect 32053 9660 32095 9669
rect 32324 9660 32382 9661
rect 33493 9660 33535 9669
rect 10933 9620 10934 9660
rect 11701 9620 11702 9660
rect 11972 9620 11981 9660
rect 12709 9620 12710 9660
rect 13525 9620 13526 9660
rect 32053 9620 32054 9660
rect 32324 9620 32333 9660
rect 33493 9620 33494 9660
rect 10933 9611 10975 9620
rect 11701 9611 11743 9620
rect 11972 9619 12030 9620
rect 12709 9611 12751 9620
rect 13525 9611 13567 9620
rect 32053 9611 32095 9620
rect 32324 9619 32382 9620
rect 33493 9611 33535 9620
rect 8869 9324 8911 9333
rect 10436 9324 10494 9325
rect 10741 9324 10783 9333
rect 11204 9324 11262 9325
rect 13220 9324 13278 9325
rect 13700 9324 13758 9325
rect 14005 9324 14047 9333
rect 35509 9324 35551 9333
rect 8869 9284 8870 9324
rect 10436 9284 10445 9324
rect 10741 9284 10742 9324
rect 11204 9284 11213 9324
rect 13220 9284 13229 9324
rect 13700 9284 13709 9324
rect 14005 9284 14006 9324
rect 35509 9284 35510 9324
rect 8869 9275 8911 9284
rect 10436 9283 10494 9284
rect 10741 9275 10783 9284
rect 11204 9283 11262 9284
rect 13220 9283 13278 9284
rect 13700 9283 13758 9284
rect 14005 9275 14047 9284
rect 35509 9275 35551 9284
rect 10165 9240 10207 9249
rect 32533 9240 32575 9249
rect 33188 9240 33246 9241
rect 10165 9200 10166 9240
rect 32533 9200 32534 9240
rect 33188 9200 33197 9240
rect 10165 9191 10207 9200
rect 32533 9191 32575 9200
rect 33188 9199 33246 9200
rect 10069 9156 10111 9165
rect 10244 9156 10302 9157
rect 10549 9156 10591 9165
rect 11509 9156 11551 9165
rect 12238 9156 12296 9157
rect 12394 9156 12436 9165
rect 12686 9156 12728 9165
rect 13333 9156 13375 9165
rect 13813 9156 13855 9165
rect 32053 9156 32095 9165
rect 32245 9156 32287 9165
rect 32432 9156 32474 9165
rect 32617 9156 32659 9165
rect 32821 9156 32863 9165
rect 33013 9156 33055 9165
rect 33572 9156 33630 9157
rect 8716 9147 8762 9156
rect 8716 9107 8717 9147
rect 10069 9116 10070 9156
rect 10244 9116 10253 9156
rect 10549 9116 10550 9156
rect 11509 9116 11510 9156
rect 12238 9116 12247 9156
rect 12394 9116 12395 9156
rect 12686 9116 12687 9156
rect 13333 9116 13334 9156
rect 13813 9116 13814 9156
rect 32053 9116 32054 9156
rect 32245 9116 32246 9156
rect 32432 9116 32433 9156
rect 32617 9116 32618 9156
rect 32821 9116 32822 9156
rect 33013 9116 33014 9156
rect 33572 9116 33581 9156
rect 10069 9107 10111 9116
rect 10244 9115 10302 9116
rect 10549 9107 10591 9116
rect 11509 9107 11551 9116
rect 12238 9115 12296 9116
rect 12394 9107 12436 9116
rect 12686 9107 12728 9116
rect 13333 9107 13375 9116
rect 13813 9107 13855 9116
rect 32053 9107 32095 9116
rect 32245 9107 32287 9116
rect 32432 9107 32474 9116
rect 32617 9107 32659 9116
rect 32821 9107 32863 9116
rect 33013 9107 33055 9116
rect 33572 9115 33630 9116
rect 8716 9098 8762 9107
rect 11419 9072 11461 9081
rect 12565 9072 12607 9081
rect 11419 9032 11420 9072
rect 12565 9032 12566 9072
rect 11419 9023 11461 9032
rect 12565 9023 12607 9032
rect 9397 8988 9439 8997
rect 12469 8988 12511 8997
rect 32612 8988 32670 8989
rect 35701 8988 35743 8997
rect 9397 8948 9398 8988
rect 12469 8948 12470 8988
rect 32612 8948 32621 8988
rect 35701 8948 35702 8988
rect 9397 8939 9439 8948
rect 12469 8939 12511 8948
rect 32612 8947 32670 8948
rect 35701 8939 35743 8948
rect 13525 8904 13567 8913
rect 32821 8904 32863 8913
rect 35125 8904 35167 8913
rect 13525 8864 13526 8904
rect 32821 8864 32822 8904
rect 35125 8864 35126 8904
rect 13525 8855 13567 8864
rect 32821 8855 32863 8864
rect 35125 8855 35167 8864
rect 13429 8568 13471 8577
rect 13429 8528 13430 8568
rect 13429 8519 13471 8528
rect 11605 8484 11647 8493
rect 11605 8444 11606 8484
rect 12053 8475 12095 8484
rect 11605 8435 11647 8444
rect 12053 8435 12054 8475
rect 12053 8426 12095 8435
rect 9524 8400 9582 8401
rect 33877 8400 33919 8409
rect 9524 8360 9533 8400
rect 33877 8360 33878 8400
rect 9524 8359 9582 8360
rect 32468 8358 32526 8359
rect 9719 8316 9777 8317
rect 9973 8316 10015 8325
rect 10637 8316 10695 8317
rect 10837 8316 10879 8325
rect 11221 8316 11263 8325
rect 12068 8316 12126 8317
rect 12469 8316 12511 8325
rect 13510 8316 13552 8325
rect 32468 8318 32477 8358
rect 33877 8351 33919 8360
rect 32468 8317 32526 8318
rect 13616 8316 13674 8317
rect 32629 8316 32671 8325
rect 32821 8316 32863 8325
rect 33536 8316 33578 8325
rect 33668 8316 33726 8317
rect 33781 8316 33823 8325
rect 34628 8316 34686 8317
rect 34944 8316 34986 8325
rect 9719 8276 9728 8316
rect 9973 8276 9974 8316
rect 10637 8276 10646 8316
rect 10837 8276 10838 8316
rect 11221 8276 11222 8316
rect 12068 8276 12077 8316
rect 12469 8276 12470 8316
rect 13510 8276 13511 8316
rect 13616 8276 13625 8316
rect 32629 8276 32630 8316
rect 32821 8276 32822 8316
rect 33536 8276 33537 8316
rect 33668 8276 33677 8316
rect 33781 8276 33782 8316
rect 34628 8276 34637 8316
rect 34944 8276 34945 8316
rect 9719 8275 9777 8276
rect 9973 8267 10015 8276
rect 10637 8275 10695 8276
rect 10837 8267 10879 8276
rect 11221 8267 11263 8276
rect 12068 8275 12126 8276
rect 12469 8267 12511 8276
rect 13510 8267 13552 8276
rect 13616 8275 13674 8276
rect 32629 8267 32671 8276
rect 32821 8267 32863 8276
rect 33536 8267 33578 8276
rect 33668 8275 33726 8276
rect 33781 8267 33823 8276
rect 34628 8275 34686 8276
rect 34944 8267 34986 8276
rect 10343 8232 10385 8241
rect 12277 8232 12319 8241
rect 32725 8232 32767 8241
rect 34837 8232 34879 8241
rect 10343 8192 10344 8232
rect 12277 8192 12278 8232
rect 32725 8192 32726 8232
rect 34837 8192 34838 8232
rect 10343 8183 10385 8192
rect 12277 8183 12319 8192
rect 32725 8183 32767 8192
rect 34837 8183 34879 8192
rect 9860 8148 9918 8149
rect 10165 8148 10207 8157
rect 10436 8148 10494 8149
rect 10549 8148 10591 8157
rect 11317 8148 11359 8157
rect 13141 8148 13183 8157
rect 32276 8148 32334 8149
rect 34724 8148 34782 8149
rect 9860 8108 9869 8148
rect 10165 8108 10166 8148
rect 10436 8108 10445 8148
rect 10549 8108 10550 8148
rect 11317 8108 11318 8148
rect 13141 8108 13142 8148
rect 32276 8108 32285 8148
rect 34724 8108 34733 8148
rect 9860 8107 9918 8108
rect 10165 8099 10207 8108
rect 10436 8107 10494 8108
rect 10549 8099 10591 8108
rect 11317 8099 11359 8108
rect 13141 8099 13183 8108
rect 32276 8107 32334 8108
rect 34724 8107 34782 8108
rect 12469 7812 12511 7821
rect 13621 7812 13663 7821
rect 12469 7772 12470 7812
rect 13621 7772 13622 7812
rect 12469 7763 12511 7772
rect 13621 7763 13663 7772
rect 10148 7728 10206 7729
rect 10148 7688 10157 7728
rect 10148 7687 10206 7688
rect 9781 7644 9823 7653
rect 9998 7644 10040 7653
rect 10532 7644 10590 7645
rect 12983 7644 13041 7645
rect 13333 7644 13375 7653
rect 13472 7644 13514 7653
rect 13813 7644 13855 7653
rect 13928 7644 13970 7653
rect 9781 7604 9782 7644
rect 9998 7604 9999 7644
rect 10532 7604 10541 7644
rect 12983 7604 12992 7644
rect 13333 7604 13334 7644
rect 13472 7604 13473 7644
rect 13813 7604 13814 7644
rect 13928 7604 13929 7644
rect 9781 7595 9823 7604
rect 9998 7595 10040 7604
rect 10532 7603 10590 7604
rect 12983 7603 13041 7604
rect 13333 7595 13375 7604
rect 13472 7595 13514 7604
rect 13813 7595 13855 7604
rect 13928 7595 13970 7604
rect 9685 7560 9727 7569
rect 12788 7560 12846 7561
rect 9685 7520 9686 7560
rect 9916 7551 9962 7560
rect 9685 7511 9727 7520
rect 9916 7511 9917 7551
rect 11597 7520 11606 7560
rect 12788 7520 12797 7560
rect 12788 7519 12846 7520
rect 9916 7502 9962 7511
rect 12085 7392 12127 7401
rect 13813 7392 13855 7401
rect 12085 7352 12086 7392
rect 13813 7352 13814 7392
rect 12085 7343 12127 7352
rect 13813 7343 13855 7352
rect 13141 7056 13183 7065
rect 13141 7016 13142 7056
rect 13141 7007 13183 7016
rect 12277 6972 12319 6981
rect 12277 6932 12278 6972
rect 12277 6923 12319 6932
rect 9863 6804 9905 6813
rect 10157 6804 10215 6805
rect 10340 6804 10398 6805
rect 11029 6804 11071 6813
rect 11300 6804 11358 6805
rect 11964 6804 12006 6813
rect 12076 6804 12134 6805
rect 12469 6804 12511 6813
rect 13508 6804 13566 6805
rect 13621 6804 13663 6813
rect 14005 6804 14047 6813
rect 9863 6764 9864 6804
rect 10157 6764 10166 6804
rect 10340 6764 10349 6804
rect 11029 6764 11030 6804
rect 11300 6764 11309 6804
rect 11964 6764 11965 6804
rect 12076 6764 12085 6804
rect 12469 6764 12470 6804
rect 13508 6764 13517 6804
rect 13621 6764 13622 6804
rect 14005 6764 14006 6804
rect 9863 6755 9905 6764
rect 10157 6763 10215 6764
rect 10340 6763 10398 6764
rect 11029 6755 11071 6764
rect 11300 6763 11358 6764
rect 11964 6755 12006 6764
rect 12076 6763 12134 6764
rect 12469 6755 12511 6764
rect 13508 6763 13566 6764
rect 13621 6755 13663 6764
rect 14005 6755 14047 6764
rect 9956 6720 10014 6721
rect 11509 6720 11551 6729
rect 11619 6720 11661 6729
rect 13796 6720 13854 6721
rect 9956 6680 9965 6720
rect 11509 6680 11510 6720
rect 11619 6680 11620 6720
rect 13796 6680 13805 6720
rect 9956 6679 10014 6680
rect 11509 6671 11551 6680
rect 11619 6671 11661 6680
rect 13796 6679 13854 6680
rect 10069 6636 10111 6645
rect 11396 6636 11454 6637
rect 11989 6636 12031 6645
rect 13525 6636 13567 6645
rect 10069 6596 10070 6636
rect 11396 6596 11405 6636
rect 11989 6596 11990 6636
rect 13525 6596 13526 6636
rect 10069 6587 10111 6596
rect 11396 6595 11454 6596
rect 11989 6587 12031 6596
rect 13525 6587 13567 6596
rect 14773 6300 14815 6309
rect 17749 6300 17791 6309
rect 18788 6300 18846 6301
rect 19652 6300 19710 6301
rect 19957 6300 19999 6309
rect 22933 6300 22975 6309
rect 25813 6300 25855 6309
rect 26084 6300 26142 6301
rect 28837 6300 28879 6309
rect 29269 6300 29311 6309
rect 29653 6300 29695 6309
rect 14773 6260 14774 6300
rect 17749 6260 17750 6300
rect 18788 6260 18797 6300
rect 19652 6260 19661 6300
rect 19957 6260 19958 6300
rect 22933 6260 22934 6300
rect 25813 6260 25814 6300
rect 26084 6260 26093 6300
rect 28837 6260 28838 6300
rect 29269 6260 29270 6300
rect 29653 6260 29654 6300
rect 14773 6251 14815 6260
rect 17749 6251 17791 6260
rect 18788 6259 18846 6260
rect 19652 6259 19710 6260
rect 19957 6251 19999 6260
rect 22933 6251 22975 6260
rect 25813 6251 25855 6260
rect 26084 6259 26142 6260
rect 28837 6251 28879 6260
rect 29269 6251 29311 6260
rect 29653 6251 29695 6260
rect 12452 6216 12510 6217
rect 20228 6216 20286 6217
rect 20612 6216 20670 6217
rect 26307 6216 26349 6225
rect 29379 6216 29421 6225
rect 12452 6176 12461 6216
rect 20228 6176 20237 6216
rect 20612 6176 20621 6216
rect 26307 6176 26308 6216
rect 29379 6176 29380 6216
rect 12452 6175 12510 6176
rect 20228 6175 20286 6176
rect 20612 6175 20670 6176
rect 26307 6167 26349 6176
rect 29379 6167 29421 6176
rect 12836 6132 12894 6133
rect 15812 6132 15870 6133
rect 18613 6132 18655 6141
rect 19093 6132 19135 6141
rect 19765 6132 19807 6141
rect 20139 6132 20181 6141
rect 20324 6132 20382 6133
rect 20437 6132 20479 6141
rect 20996 6132 21054 6133
rect 23876 6132 23934 6133
rect 25988 6132 26046 6133
rect 28309 6132 28351 6141
rect 28505 6132 28547 6141
rect 28693 6132 28735 6141
rect 29060 6132 29118 6133
rect 29173 6132 29215 6141
rect 29557 6132 29599 6141
rect 29749 6132 29791 6141
rect 12836 6092 12845 6132
rect 14956 6123 15002 6132
rect 12836 6091 12894 6092
rect 14956 6083 14957 6123
rect 15812 6092 15821 6132
rect 18613 6092 18614 6132
rect 19093 6092 19094 6132
rect 19765 6092 19766 6132
rect 20139 6092 20140 6132
rect 20324 6092 20333 6132
rect 20437 6092 20438 6132
rect 20996 6092 21005 6132
rect 23876 6092 23885 6132
rect 25988 6092 25997 6132
rect 27532 6123 27578 6132
rect 15812 6091 15870 6092
rect 18613 6083 18655 6092
rect 19093 6083 19135 6092
rect 19765 6083 19807 6092
rect 20139 6083 20181 6092
rect 20324 6091 20382 6092
rect 20437 6083 20479 6092
rect 20996 6091 21054 6092
rect 23876 6091 23934 6092
rect 25988 6091 26046 6092
rect 27532 6083 27533 6123
rect 28309 6092 28310 6132
rect 28505 6092 28506 6132
rect 28693 6092 28694 6132
rect 29060 6092 29069 6132
rect 29173 6092 29174 6132
rect 29557 6092 29558 6132
rect 29749 6092 29750 6132
rect 28309 6083 28351 6092
rect 28505 6083 28547 6092
rect 28693 6083 28735 6092
rect 29060 6091 29118 6092
rect 29173 6083 29215 6092
rect 29557 6083 29599 6092
rect 29749 6083 29791 6092
rect 14956 6074 15002 6083
rect 27532 6074 27578 6083
rect 15109 6048 15151 6057
rect 15445 6048 15487 6057
rect 19003 6048 19045 6057
rect 22549 6048 22591 6057
rect 23509 6048 23551 6057
rect 25429 6048 25471 6057
rect 27685 6048 27727 6057
rect 13613 6008 13622 6048
rect 15109 6008 15110 6048
rect 15445 6008 15446 6048
rect 16397 6008 16406 6048
rect 19003 6008 19004 6048
rect 21773 6008 21782 6048
rect 22549 6008 22550 6048
rect 23509 6008 23510 6048
rect 24557 6008 24566 6048
rect 25429 6008 25430 6048
rect 27685 6008 27686 6048
rect 15109 5999 15151 6008
rect 15445 5999 15487 6008
rect 19003 5999 19045 6008
rect 22549 5999 22591 6008
rect 23509 5999 23551 6008
rect 25429 5999 25471 6008
rect 27685 5999 27727 6008
rect 14773 5964 14815 5973
rect 17941 5964 17983 5973
rect 14773 5924 14774 5964
rect 17941 5924 17942 5964
rect 14773 5915 14815 5924
rect 17941 5915 17983 5924
rect 14389 5880 14431 5889
rect 17365 5880 17407 5889
rect 17749 5880 17791 5889
rect 26293 5880 26335 5889
rect 28405 5880 28447 5889
rect 14389 5840 14390 5880
rect 17365 5840 17366 5880
rect 17749 5840 17750 5880
rect 26293 5840 26294 5880
rect 28405 5840 28406 5880
rect 14389 5831 14431 5840
rect 17365 5831 17407 5840
rect 17749 5831 17791 5840
rect 26293 5831 26335 5840
rect 28405 5831 28447 5840
rect 15253 5544 15295 5553
rect 20629 5544 20671 5553
rect 23509 5544 23551 5553
rect 15253 5504 15254 5544
rect 20629 5504 20630 5544
rect 23509 5504 23510 5544
rect 15253 5495 15295 5504
rect 20629 5495 20671 5504
rect 23509 5495 23551 5504
rect 13621 5460 13663 5469
rect 15877 5460 15919 5469
rect 19189 5460 19231 5469
rect 21109 5460 21151 5469
rect 21877 5460 21919 5469
rect 24565 5460 24607 5469
rect 13621 5420 13622 5460
rect 15877 5420 15878 5460
rect 19189 5420 19190 5460
rect 21109 5420 21110 5460
rect 21877 5420 21878 5460
rect 24565 5420 24566 5460
rect 13621 5411 13663 5420
rect 15877 5411 15919 5420
rect 19189 5411 19231 5420
rect 21109 5411 21151 5420
rect 21877 5411 21919 5420
rect 24565 5411 24607 5420
rect 15660 5376 15702 5385
rect 17204 5376 17262 5377
rect 17989 5376 18031 5385
rect 22580 5376 22638 5377
rect 15660 5336 15661 5376
rect 17204 5336 17213 5376
rect 17989 5336 17990 5376
rect 22580 5336 22589 5376
rect 15660 5327 15702 5336
rect 17204 5335 17262 5336
rect 17989 5327 18031 5336
rect 22580 5335 22638 5336
rect 14948 5292 15006 5293
rect 15541 5292 15583 5301
rect 15770 5292 15828 5293
rect 16021 5292 16063 5301
rect 17399 5292 17457 5293
rect 17780 5292 17838 5293
rect 19093 5292 19135 5301
rect 19285 5292 19327 5301
rect 20629 5292 20671 5301
rect 20821 5292 20863 5301
rect 21205 5292 21247 5301
rect 21493 5292 21535 5301
rect 22775 5292 22833 5293
rect 23204 5292 23262 5293
rect 23523 5292 23565 5301
rect 14948 5252 14957 5292
rect 15541 5252 15542 5292
rect 15770 5252 15779 5292
rect 16021 5252 16022 5292
rect 17399 5252 17408 5292
rect 17780 5252 17789 5292
rect 19093 5252 19094 5292
rect 19285 5252 19286 5292
rect 20629 5252 20630 5292
rect 20821 5252 20822 5292
rect 21205 5252 21206 5292
rect 21493 5252 21494 5292
rect 22775 5252 22784 5292
rect 23204 5252 23213 5292
rect 23523 5252 23524 5292
rect 14948 5251 15006 5252
rect 15541 5243 15583 5252
rect 15770 5251 15828 5252
rect 16021 5243 16063 5252
rect 17399 5251 17457 5252
rect 17780 5251 17838 5252
rect 19093 5243 19135 5252
rect 19285 5243 19327 5252
rect 20629 5243 20671 5252
rect 20821 5243 20863 5252
rect 21205 5243 21247 5252
rect 21493 5243 21535 5252
rect 22775 5251 22833 5252
rect 23204 5251 23262 5252
rect 23523 5243 23565 5252
rect 15267 5208 15309 5217
rect 15445 5208 15487 5217
rect 23317 5208 23359 5217
rect 15267 5168 15268 5208
rect 15445 5168 15446 5208
rect 23317 5168 23318 5208
rect 15267 5159 15309 5168
rect 15445 5159 15487 5168
rect 23317 5159 23359 5168
rect 15044 5124 15102 5125
rect 21109 5124 21151 5133
rect 21380 5124 21438 5125
rect 21685 5124 21727 5133
rect 15044 5084 15053 5124
rect 21109 5084 21110 5124
rect 21380 5084 21389 5124
rect 21685 5084 21686 5124
rect 15044 5083 15102 5084
rect 21109 5075 21151 5084
rect 21380 5083 21438 5084
rect 21685 5075 21727 5084
<< metal1 >>
rect 2687 27560 3127 27569
rect 2687 27120 2688 27560
rect 3126 27120 3824 27560
rect 2687 27111 3127 27120
rect 3705 26378 3785 26387
rect 3705 26298 3706 26378
rect 3784 26298 3785 26378
rect 3705 26289 3785 26298
rect 5265 25482 5345 25491
rect 5265 25402 5266 25482
rect 5344 25402 5345 25482
rect 5265 25393 5345 25402
rect 3703 24596 3783 24605
rect 3703 24516 3704 24596
rect 3782 24516 3783 24596
rect 3703 24507 3783 24516
rect 5265 23708 5345 23717
rect 5265 23628 5266 23708
rect 5344 23628 5345 23708
rect 5265 23619 5345 23628
rect 3695 22820 3775 22829
rect 3695 22740 3696 22820
rect 3774 22740 3775 22820
rect 3695 22731 3775 22740
rect 5249 21940 5329 21949
rect 5249 21860 5250 21940
rect 5328 21860 5329 21940
rect 5249 21851 5329 21860
rect 3695 21020 3775 21029
rect 3695 20940 3696 21020
rect 3774 20940 3775 21020
rect 3695 20931 3775 20940
rect 5227 20646 5407 20655
rect 5227 20466 5228 20646
rect 5406 20466 5407 20646
rect 5227 20457 5407 20466
rect 2657 20324 3097 20333
rect 2657 19884 2658 20324
rect 3096 19924 3662 20324
rect 5249 20150 5329 20159
rect 5249 20070 5250 20150
rect 5328 20070 5329 20150
rect 5249 20061 5329 20070
rect 3096 19884 5642 19924
rect 2657 19875 3097 19884
rect 3222 19680 5642 19884
rect 3218 19628 5642 19680
rect 3218 19174 5712 19628
rect 3218 18784 3936 19174
rect 3719 18054 3799 18063
rect 3719 17974 3720 18054
rect 3798 17974 3799 18054
rect 3719 17965 3799 17974
rect 5275 17158 5355 17167
rect 5275 17078 5276 17158
rect 5354 17078 5355 17158
rect 5275 17069 5355 17078
rect 3713 16276 3793 16285
rect 3713 16196 3714 16276
rect 3792 16196 3793 16276
rect 3713 16187 3793 16196
rect 5285 15388 5383 15389
rect 5285 15310 5294 15388
rect 5374 15310 5383 15388
rect 5285 15309 5383 15310
rect 3719 14484 3799 14493
rect 3719 14404 3720 14484
rect 3798 14404 3799 14484
rect 3719 14395 3799 14404
rect 5265 13612 5345 13621
rect 5265 13532 5266 13612
rect 5344 13532 5345 13612
rect 5265 13523 5345 13532
rect 3709 12720 3789 12729
rect 3709 12640 3710 12720
rect 3788 12640 3789 12720
rect 3709 12631 3789 12640
rect 5219 12338 5399 12347
rect 5219 12158 5220 12338
rect 5398 12158 5399 12338
rect 5219 12149 5399 12158
rect 5269 11834 5349 11843
rect 2621 11752 3061 11761
rect 5269 11754 5270 11834
rect 5348 11754 5349 11834
rect 2621 11312 2622 11752
rect 3060 11746 3152 11752
rect 3060 11584 3680 11746
rect 5269 11745 5349 11754
rect 3060 11320 5664 11584
rect 3060 11318 5696 11320
rect 3060 11312 3152 11318
rect 2621 11303 3061 11312
rect 3428 11006 5696 11318
rect 3462 10842 5696 11006
rect 3462 10452 3900 10842
rect 3723 9720 3803 9729
rect 3723 9640 3724 9720
rect 3802 9640 3803 9720
rect 3723 9631 3803 9640
rect 5281 8842 5361 8851
rect 5281 8762 5282 8842
rect 5360 8762 5361 8842
rect 5281 8753 5361 8762
rect 3729 7948 3809 7957
rect 3729 7868 3730 7948
rect 3808 7868 3809 7948
rect 3729 7859 3809 7868
rect 5285 7054 5365 7063
rect 5285 6974 5286 7054
rect 5364 6974 5365 7054
rect 5285 6965 5365 6974
rect 3729 6176 3809 6185
rect 3729 6096 3730 6176
rect 3808 6096 3809 6176
rect 3729 6087 3809 6096
rect 5271 5286 5351 5295
rect 5271 5206 5272 5286
rect 5350 5206 5351 5286
rect 5271 5197 5351 5206
rect 3713 4398 3793 4407
rect 3713 4318 3714 4398
rect 3792 4318 3793 4398
rect 3713 4309 3793 4318
rect 5223 4010 5403 4019
rect 5223 3830 5224 4010
rect 5402 3830 5403 4010
rect 5223 3821 5403 3830
rect 5271 3504 5351 3513
rect 5271 3424 5272 3504
rect 5350 3424 5351 3504
rect 5271 3415 5351 3424
rect 2581 3334 3021 3343
rect 2581 2894 2582 3334
rect 3020 3328 3112 3334
rect 3020 3312 3226 3328
rect 3020 3299 3370 3312
rect 3020 2949 5639 3299
rect 3020 2906 3370 2949
rect 3020 2900 3226 2906
rect 3020 2894 3112 2900
rect 2581 2885 3021 2894
<< via1 >>
rect 2688 27120 3126 27560
rect 3706 26298 3784 26378
rect 5266 25402 5344 25482
rect 3704 24516 3782 24596
rect 5266 23628 5344 23708
rect 3696 22740 3774 22820
rect 5250 21860 5328 21940
rect 3696 20940 3774 21020
rect 5228 20466 5406 20646
rect 2658 19884 3096 20324
rect 5250 20070 5328 20150
rect 3720 17974 3798 18054
rect 5276 17078 5354 17158
rect 3714 16196 3792 16276
rect 5294 15310 5374 15388
rect 3720 14404 3798 14484
rect 5266 13532 5344 13612
rect 3710 12640 3788 12720
rect 5220 12158 5398 12338
rect 5270 11754 5348 11834
rect 2622 11312 3060 11752
rect 3724 9640 3802 9720
rect 5282 8762 5360 8842
rect 3730 7868 3808 7948
rect 5286 6974 5364 7054
rect 3730 6096 3808 6176
rect 5272 5206 5350 5286
rect 3714 4318 3792 4398
rect 5224 3830 5402 4010
rect 5272 3424 5350 3504
rect 2582 2894 3020 3334
<< metal2 >>
rect 2686 27560 3126 27569
rect 2679 27120 2686 27560
rect 3126 27120 3135 27560
rect 2686 27111 3126 27120
rect 3697 26298 3706 26378
rect 3784 26298 7298 26378
rect 5257 25402 5266 25482
rect 5344 25402 7106 25482
rect 3695 24516 3704 24596
rect 3782 24516 6900 24596
rect 5257 23628 5266 23708
rect 5344 23628 6650 23708
rect 3687 22740 3696 22820
rect 3774 22740 6422 22820
rect 5241 21860 5250 21940
rect 5328 21860 6188 21940
rect 3007 21600 3016 21780
rect 3196 21600 3205 21780
rect 3016 20646 3196 21600
rect 6108 21440 6188 21860
rect 6342 21860 6422 22740
rect 6570 22280 6650 23628
rect 6820 22700 6900 24516
rect 7026 23120 7106 25402
rect 7218 23540 7298 26298
rect 7218 23460 7726 23540
rect 7026 23040 7682 23120
rect 6820 22620 7698 22700
rect 6570 22200 7690 22280
rect 6342 21780 7674 21860
rect 6108 21360 7682 21440
rect 3687 20940 3696 21020
rect 3774 20940 7690 21020
rect 3016 20466 5228 20646
rect 5406 20466 5415 20646
rect 7116 20520 7690 20600
rect 2656 20324 3096 20333
rect 2649 19884 2656 20324
rect 3096 19884 3105 20324
rect 7116 20150 7196 20520
rect 5241 20070 5250 20150
rect 5328 20070 7196 20150
rect 2656 19875 3096 19884
rect 3711 17974 3720 18054
rect 3798 17974 7262 18054
rect 5267 17078 5276 17158
rect 5354 17078 7020 17158
rect 6940 16400 7020 17078
rect 7182 16820 7262 17974
rect 7182 16740 7686 16820
rect 6940 16320 7586 16400
rect 3705 16196 3714 16276
rect 3792 16196 6784 16276
rect 6704 15980 6784 16196
rect 6704 15900 7592 15980
rect 5294 15480 7680 15560
rect 5294 15388 5374 15480
rect 5294 15301 5374 15310
rect 5860 15060 7672 15140
rect 5860 14484 5940 15060
rect 3711 14404 3720 14484
rect 3798 14404 5940 14484
rect 6276 14640 7596 14720
rect 6276 13612 6356 14640
rect 5257 13532 5266 13612
rect 5344 13532 6356 13612
rect 6676 14220 7596 14300
rect 6676 12720 6756 14220
rect 3701 12640 3710 12720
rect 3788 12640 6756 12720
rect 7064 13800 7600 13880
rect 2707 12158 2716 12338
rect 2896 12158 5220 12338
rect 5398 12158 5407 12338
rect 7064 11834 7144 13800
rect 2620 11752 3060 11761
rect 5261 11754 5270 11834
rect 5348 11754 7144 11834
rect 2613 11312 2620 11752
rect 3060 11312 3069 11752
rect 2620 11303 3060 11312
rect 5326 10020 7680 10100
rect 5326 9720 5406 10020
rect 3715 9640 3724 9720
rect 3802 9640 5406 9720
rect 5598 9600 7590 9680
rect 5598 8842 5678 9600
rect 5273 8762 5282 8842
rect 5360 8762 5678 8842
rect 5814 9180 7586 9260
rect 5814 7948 5894 9180
rect 3721 7868 3730 7948
rect 3808 7868 5894 7948
rect 6030 8760 7580 8840
rect 6030 7054 6110 8760
rect 5277 6974 5286 7054
rect 5364 6974 6110 7054
rect 6240 8340 7596 8420
rect 6240 6176 6320 8340
rect 3721 6096 3730 6176
rect 3808 6096 6320 6176
rect 6440 7920 7586 8000
rect 6440 5286 6520 7920
rect 5263 5206 5272 5286
rect 5350 5206 6520 5286
rect 6646 7500 7590 7580
rect 6646 4398 6726 7500
rect 3705 4318 3714 4398
rect 3792 4318 6726 4398
rect 6888 7080 7616 7160
rect 1634 4010 1814 4019
rect 1814 3830 5224 4010
rect 5402 3830 5411 4010
rect 1634 3821 1814 3830
rect 6888 3504 6968 7080
rect 5263 3424 5272 3504
rect 5350 3424 6968 3504
rect 2580 3334 3020 3343
rect 2573 2894 2580 3334
rect 3020 2894 3029 3334
rect 2580 2885 3020 2894
<< via2 >>
rect 2686 27120 2688 27560
rect 2688 27120 3126 27560
rect 3016 21600 3196 21780
rect 2656 19884 2658 20324
rect 2658 19884 3096 20324
rect 2716 12158 2896 12338
rect 2620 11312 2622 11752
rect 2622 11312 3060 11752
rect 1634 3830 1814 4010
rect 2580 2894 2582 3334
rect 2582 2894 3020 3334
<< metal3 >>
rect 10502 30465 10621 30479
rect 10502 30373 10515 30465
rect 10607 30373 10621 30465
rect 10502 30019 10621 30373
rect 11270 30465 11389 30479
rect 11270 30373 11283 30465
rect 11375 30373 11389 30465
rect 11270 30019 11389 30373
rect 12038 30465 12157 30479
rect 12038 30373 12051 30465
rect 12143 30373 12157 30465
rect 12038 30019 12157 30373
rect 12806 30465 12925 30479
rect 12806 30373 12819 30465
rect 12911 30373 12925 30465
rect 12806 30019 12925 30373
rect 13574 30465 13693 30479
rect 13574 30373 13587 30465
rect 13679 30373 13693 30465
rect 13574 30019 13693 30373
rect 14342 30465 14461 30479
rect 14342 30373 14355 30465
rect 14447 30373 14461 30465
rect 14342 30019 14461 30373
rect 15110 30465 15229 30479
rect 15110 30373 15123 30465
rect 15215 30373 15229 30465
rect 15110 30019 15229 30373
rect 15878 30465 15997 30479
rect 15878 30373 15891 30465
rect 15983 30373 15997 30465
rect 15878 30019 15997 30373
rect 16646 30465 16765 30479
rect 16646 30373 16659 30465
rect 16751 30373 16765 30465
rect 16646 30019 16765 30373
rect 17414 30465 17533 30479
rect 17414 30373 17427 30465
rect 17519 30373 17533 30465
rect 17414 30019 17533 30373
rect 18182 30465 18301 30479
rect 18182 30373 18195 30465
rect 18287 30373 18301 30465
rect 18182 30019 18301 30373
rect 18950 30465 19069 30479
rect 18950 30373 18963 30465
rect 19055 30373 19069 30465
rect 18950 30019 19069 30373
rect 19718 30465 19837 30479
rect 19718 30373 19731 30465
rect 19823 30373 19837 30465
rect 19718 30019 19837 30373
rect 20486 30465 20605 30479
rect 20486 30373 20499 30465
rect 20591 30373 20605 30465
rect 20486 30019 20605 30373
rect 21254 30465 21373 30479
rect 21254 30373 21267 30465
rect 21359 30373 21373 30465
rect 21254 30019 21373 30373
rect 22022 30465 22141 30479
rect 22022 30373 22035 30465
rect 22127 30373 22141 30465
rect 22022 30019 22141 30373
rect 22790 30465 22909 30479
rect 22790 30373 22803 30465
rect 22895 30373 22909 30465
rect 22790 30019 22909 30373
rect 23558 30465 23677 30479
rect 23558 30373 23571 30465
rect 23663 30373 23677 30465
rect 23558 30019 23677 30373
rect 30471 30362 30480 30458
rect 30576 30362 30585 30458
rect 31239 30362 31248 30458
rect 31344 30362 31353 30458
rect 32007 30362 32016 30458
rect 32112 30362 32121 30458
rect 32775 30362 32784 30458
rect 32880 30362 32889 30458
rect 33543 30362 33552 30458
rect 33648 30362 33657 30458
rect 34311 30362 34320 30458
rect 34416 30362 34425 30458
rect 35079 30362 35088 30458
rect 35184 30362 35193 30458
rect 35847 30362 35856 30458
rect 35952 30362 35961 30458
rect 36615 30362 36624 30458
rect 36720 30362 36729 30458
rect 37383 30362 37392 30458
rect 37488 30362 37497 30458
rect 38151 30362 38160 30458
rect 38256 30362 38265 30458
rect 30480 30010 30576 30362
rect 31248 30010 31344 30362
rect 32016 30010 32112 30362
rect 32784 30010 32880 30362
rect 33552 30010 33648 30362
rect 34320 30010 34416 30362
rect 35088 30010 35184 30362
rect 35856 30010 35952 30362
rect 36624 30010 36720 30362
rect 37392 30010 37488 30362
rect 38160 30010 38256 30362
rect 2677 27120 2686 27560
rect 3126 27120 3135 27560
rect 3007 24596 3016 24776
rect 3196 24596 3205 24776
rect 3016 21780 3196 24596
rect 3016 21591 3196 21600
rect 2181 21396 2190 21576
rect 2370 21396 2379 21576
rect 2190 19098 2370 21396
rect 2647 19884 2656 20324
rect 3096 19884 3105 20324
rect 2190 18918 2896 19098
rect 1625 18196 1634 18376
rect 1814 18196 1823 18376
rect 1634 4010 1814 18196
rect 2716 12338 2896 18918
rect 2716 12149 2896 12158
rect 2611 11312 2620 11752
rect 3060 11312 3069 11752
rect 1625 3830 1634 4010
rect 1814 3830 1823 4010
rect 2571 2894 2580 3334
rect 3020 2894 3029 3334
<< via3 >>
rect 10515 30373 10607 30465
rect 11283 30373 11375 30465
rect 12051 30373 12143 30465
rect 12819 30373 12911 30465
rect 13587 30373 13679 30465
rect 14355 30373 14447 30465
rect 15123 30373 15215 30465
rect 15891 30373 15983 30465
rect 16659 30373 16751 30465
rect 17427 30373 17519 30465
rect 18195 30373 18287 30465
rect 18963 30373 19055 30465
rect 19731 30373 19823 30465
rect 20499 30373 20591 30465
rect 21267 30373 21359 30465
rect 22035 30373 22127 30465
rect 22803 30373 22895 30465
rect 23571 30373 23663 30465
rect 30480 30362 30576 30458
rect 31248 30362 31344 30458
rect 32016 30362 32112 30458
rect 32784 30362 32880 30458
rect 33552 30362 33648 30458
rect 34320 30362 34416 30458
rect 35088 30362 35184 30458
rect 35856 30362 35952 30458
rect 36624 30362 36720 30458
rect 37392 30362 37488 30458
rect 38160 30362 38256 30458
rect 2686 27120 3126 27560
rect 3016 24596 3196 24776
rect 2190 21396 2370 21576
rect 2656 19884 3096 20324
rect 1634 18196 1814 18376
rect 2620 11312 3060 11752
rect 2580 2894 3020 3334
<< metal4 >>
rect 10515 30465 10607 30474
rect 11283 30465 11375 30474
rect 12051 30465 12143 30474
rect 12819 30465 12911 30474
rect 13587 30465 13679 30474
rect 14355 30465 14447 30474
rect 15123 30465 15215 30474
rect 15891 30465 15983 30474
rect 16659 30465 16751 30474
rect 17427 30465 17519 30474
rect 18195 30465 18287 30474
rect 18963 30465 19055 30474
rect 19731 30465 19823 30474
rect 20499 30465 20591 30474
rect 21267 30465 21359 30474
rect 22035 30465 22127 30474
rect 22803 30465 22895 30474
rect 23571 30465 23663 30474
rect 10508 30375 10515 30462
rect 10607 30375 10613 30462
rect 11276 30375 11283 30462
rect 11375 30375 11381 30462
rect 12044 30375 12051 30462
rect 12143 30375 12149 30462
rect 12812 30375 12819 30462
rect 12911 30375 12917 30462
rect 13580 30375 13587 30462
rect 13679 30375 13685 30462
rect 14348 30375 14355 30462
rect 14447 30375 14453 30462
rect 15116 30375 15123 30462
rect 15215 30375 15221 30462
rect 15884 30375 15891 30462
rect 15983 30375 15989 30462
rect 16652 30375 16659 30462
rect 16751 30375 16757 30462
rect 17420 30375 17427 30462
rect 17519 30375 17525 30462
rect 18188 30375 18195 30462
rect 18287 30375 18293 30462
rect 18956 30375 18963 30462
rect 19055 30375 19061 30462
rect 19724 30375 19731 30462
rect 19823 30375 19829 30462
rect 20492 30375 20499 30462
rect 20591 30375 20597 30462
rect 21260 30375 21267 30462
rect 21359 30375 21365 30462
rect 22028 30375 22035 30462
rect 22127 30375 22133 30462
rect 22796 30375 22803 30462
rect 22895 30375 22901 30462
rect 23564 30375 23571 30462
rect 23663 30375 23669 30462
rect 30480 30458 30576 30467
rect 31248 30458 31344 30467
rect 32016 30458 32112 30467
rect 32784 30458 32880 30467
rect 33552 30458 33648 30467
rect 34320 30458 34416 30467
rect 35088 30458 35184 30467
rect 35856 30458 35952 30467
rect 36624 30458 36720 30467
rect 37392 30458 37488 30467
rect 38160 30458 38256 30467
rect 10515 30364 10607 30373
rect 11283 30364 11375 30373
rect 12051 30364 12143 30373
rect 12819 30364 12911 30373
rect 13587 30364 13679 30373
rect 14355 30364 14447 30373
rect 15123 30364 15215 30373
rect 15891 30364 15983 30373
rect 16659 30364 16751 30373
rect 17427 30364 17519 30373
rect 18195 30364 18287 30373
rect 18963 30364 19055 30373
rect 19731 30364 19823 30373
rect 20499 30364 20591 30373
rect 21267 30364 21359 30373
rect 22035 30364 22127 30373
rect 22803 30364 22895 30373
rect 23571 30364 23663 30373
rect 30471 30362 30480 30458
rect 30576 30362 30585 30458
rect 31239 30362 31248 30458
rect 31344 30362 31353 30458
rect 32007 30362 32016 30458
rect 32112 30362 32121 30458
rect 32775 30362 32784 30458
rect 32880 30362 32889 30458
rect 33543 30362 33552 30458
rect 33648 30362 33657 30458
rect 34311 30362 34320 30458
rect 34416 30362 34425 30458
rect 35079 30362 35088 30458
rect 35184 30362 35193 30458
rect 35847 30362 35856 30458
rect 35952 30362 35961 30458
rect 36615 30362 36624 30458
rect 36720 30362 36729 30458
rect 37383 30362 37392 30458
rect 37488 30362 37497 30458
rect 38151 30362 38160 30458
rect 38256 30362 38265 30458
rect 30480 30353 30576 30362
rect 31248 30353 31344 30362
rect 32016 30353 32112 30362
rect 32784 30353 32880 30362
rect 33552 30353 33648 30362
rect 34320 30353 34416 30362
rect 35088 30353 35184 30362
rect 35856 30353 35952 30362
rect 36624 30353 36720 30362
rect 37392 30353 37488 30362
rect 38160 30353 38256 30362
rect 2686 27560 3126 27569
rect 2686 27111 3126 27120
rect 416 24776 596 24785
rect 3016 24776 3196 24785
rect 596 24596 3016 24776
rect 416 24587 596 24596
rect 3016 24587 3196 24596
rect 418 21576 598 21585
rect 2190 21576 2370 21585
rect 598 21396 2190 21576
rect 418 21387 598 21396
rect 2190 21387 2370 21396
rect 2656 20324 3096 20333
rect 2656 19875 3096 19884
rect 392 18376 572 18385
rect 1634 18376 1814 18385
rect 572 18196 1634 18376
rect 392 18187 572 18196
rect 1634 18187 1814 18196
rect 2620 11752 3060 11761
rect 2620 11303 3060 11312
rect 2580 3334 3020 3343
rect 2580 2885 3020 2894
rect 7113 1659 7718 1668
rect 7718 1584 38332 1659
rect 7718 1144 11718 1584
rect 12158 1144 19492 1584
rect 19932 1578 38332 1584
rect 19932 1144 27266 1578
rect 7718 1138 27266 1144
rect 27706 1570 38332 1578
rect 27706 1138 35040 1570
rect 7718 1130 35040 1138
rect 35480 1130 38332 1570
rect 7718 1054 38332 1130
rect 7113 1045 7718 1054
<< via4 >>
rect 10517 30375 10604 30462
rect 11285 30375 11372 30462
rect 12053 30375 12140 30462
rect 12821 30375 12908 30462
rect 13589 30375 13676 30462
rect 14357 30375 14444 30462
rect 15125 30375 15212 30462
rect 15893 30375 15980 30462
rect 16661 30375 16748 30462
rect 17429 30375 17516 30462
rect 18197 30375 18284 30462
rect 18965 30375 19052 30462
rect 19733 30375 19820 30462
rect 20501 30375 20588 30462
rect 21269 30375 21356 30462
rect 22037 30375 22124 30462
rect 22805 30375 22892 30462
rect 23573 30375 23660 30462
rect 30480 30362 30576 30458
rect 31248 30362 31344 30458
rect 32016 30362 32112 30458
rect 32784 30362 32880 30458
rect 33552 30362 33648 30458
rect 34320 30362 34416 30458
rect 35088 30362 35184 30458
rect 35856 30362 35952 30458
rect 36624 30362 36720 30458
rect 37392 30362 37488 30458
rect 38160 30362 38256 30458
rect 2686 27120 3126 27560
rect 416 24596 596 24776
rect 418 21396 598 21576
rect 2656 19884 3096 20324
rect 392 18196 572 18376
rect 2620 11312 3060 11752
rect 2580 2894 3020 3334
rect 7113 1054 7718 1659
rect 11718 1144 12158 1584
rect 19492 1144 19932 1584
rect 27266 1138 27706 1578
rect 35040 1130 35480 1570
<< metal5 >>
rect 958 30596 1732 30678
rect 791 30592 1732 30596
rect 5922 30592 5982 30996
rect 6690 30592 6750 30996
rect 7458 30592 7518 30996
rect 8226 30592 8286 30996
rect 8994 30592 9054 30996
rect 9762 30592 9822 30996
rect 791 30532 9822 30592
rect 791 30456 1732 30532
rect 10530 30522 10590 30996
rect 11298 30522 11358 30996
rect 12066 30522 12126 30996
rect 12834 30522 12894 30996
rect 13602 30522 13662 30996
rect 14370 30522 14430 30996
rect 15138 30522 15198 30996
rect 15906 30522 15966 30996
rect 16674 30522 16734 30996
rect 17442 30522 17502 30996
rect 18210 30522 18270 30996
rect 18978 30522 19038 30996
rect 19746 30522 19806 30996
rect 20514 30522 20574 30996
rect 21282 30522 21342 30996
rect 22050 30522 22110 30996
rect 22818 30522 22878 30996
rect 23586 30522 23646 30996
rect 24354 30796 24414 30996
rect 25122 30796 25182 30996
rect 25890 30796 25950 30996
rect 26658 30796 26718 30996
rect 27426 30796 27486 30996
rect 28194 30796 28254 30996
rect 28962 30796 29022 30996
rect 29730 30796 29790 30996
rect 30498 30522 30558 30996
rect 31266 30522 31326 30996
rect 32034 30522 32094 30996
rect 32802 30522 32862 30996
rect 33570 30522 33630 30996
rect 34338 30522 34398 30996
rect 35106 30522 35166 30996
rect 35874 30522 35934 30996
rect 36642 30522 36702 30996
rect 37410 30522 37470 30996
rect 38178 30522 38238 30996
rect 800 30446 1732 30456
rect 10517 30462 10604 30522
rect 800 27560 1240 30446
rect 10517 30366 10604 30375
rect 11285 30462 11372 30522
rect 11285 30366 11372 30375
rect 12053 30462 12140 30522
rect 12053 30366 12140 30375
rect 12821 30462 12908 30522
rect 12821 30366 12908 30375
rect 13589 30462 13676 30522
rect 13589 30366 13676 30375
rect 14357 30462 14444 30522
rect 14357 30366 14444 30375
rect 15125 30462 15212 30522
rect 15125 30366 15212 30375
rect 15893 30462 15980 30522
rect 15893 30366 15980 30375
rect 16661 30462 16748 30522
rect 16661 30366 16748 30375
rect 17429 30462 17516 30522
rect 17429 30366 17516 30375
rect 18197 30462 18284 30522
rect 18197 30366 18284 30375
rect 18965 30462 19052 30522
rect 18965 30366 19052 30375
rect 19733 30462 19820 30522
rect 19733 30366 19820 30375
rect 20501 30462 20588 30522
rect 20501 30366 20588 30375
rect 21269 30462 21356 30522
rect 21269 30366 21356 30375
rect 22037 30462 22124 30522
rect 22037 30366 22124 30375
rect 22805 30462 22892 30522
rect 22805 30366 22892 30375
rect 23573 30462 23660 30522
rect 23573 30366 23660 30375
rect 30480 30458 30576 30522
rect 30480 30353 30576 30362
rect 31248 30458 31344 30522
rect 31248 30353 31344 30362
rect 32016 30458 32112 30522
rect 32016 30353 32112 30362
rect 32784 30458 32880 30522
rect 32784 30353 32880 30362
rect 33552 30458 33648 30522
rect 33552 30353 33648 30362
rect 34320 30458 34416 30522
rect 34320 30353 34416 30362
rect 35088 30458 35184 30522
rect 35088 30353 35184 30362
rect 35856 30458 35952 30522
rect 35856 30353 35952 30362
rect 36624 30458 36720 30522
rect 36624 30353 36720 30362
rect 37392 30458 37488 30522
rect 37392 30353 37488 30362
rect 38160 30458 38256 30522
rect 38160 30353 38256 30362
rect 800 27120 2686 27560
rect 3126 27120 3135 27560
rect 0 24596 416 24776
rect 596 24596 605 24776
rect 0 21396 418 21576
rect 598 21396 607 21576
rect 800 20324 1240 27120
rect 800 19884 2656 20324
rect 3096 19884 3105 20324
rect 0 18196 392 18376
rect 572 18196 581 18376
rect 0 14996 200 15176
rect 800 11752 1240 19884
rect 800 11312 2620 11752
rect 3060 11312 3069 11752
rect 800 3334 1240 11312
rect 800 2894 2580 3334
rect 3020 2894 3029 3334
rect 800 1576 1240 2894
rect 6420 1576 7113 1659
rect 800 1136 7113 1576
rect 800 0 1240 1136
rect 6420 1054 7113 1136
rect 7718 1054 7727 1659
rect 10448 796 10968 2534
rect 11718 1584 12158 2488
rect 11718 1135 12158 1144
rect 18214 796 18734 2540
rect 19492 1584 19932 2372
rect 19492 1135 19932 1144
rect 25998 796 26518 2556
rect 27266 1578 27706 2372
rect 27266 1129 27706 1138
rect 33750 796 34270 2482
rect 35040 1570 35480 2372
rect 35040 1121 35480 1130
rect 39800 796 40240 30596
rect 7168 356 40240 796
rect 7254 276 40240 356
rect 39800 0 40240 276
use r2r_dac  blue_dac
timestamp 1746810912
transform 0 1 3516 -1 0 10920
box -142 -18 7922 2062
use controller  controller_0
timestamp 1746801438
transform 1 0 7402 0 1 1156
box 0 700 31805 29000
use r2r_dac  green_dac
timestamp 1746810912
transform 0 1 3512 -1 0 19246
box -142 -18 7922 2062
use r2r_dac  red_dac
timestamp 1746810912
transform 0 1 3492 -1 0 27566
box -142 -18 7922 2062
<< labels >>
flabel metal5 s 37410 30796 37470 30996 4 FreeSans 320 0 0 0 clk
port 2 nsew
flabel metal5 s 38178 30796 38238 30996 4 FreeSans 320 0 0 0 ena
port 3 nsew
flabel metal5 s 36642 30796 36702 30996 4 FreeSans 320 0 0 0 rst_n
port 4 nsew
flabel metal5 s 35874 30796 35934 30996 4 FreeSans 320 0 0 0 ui_in[0]
port 5 nsew
flabel metal5 s 35106 30796 35166 30996 4 FreeSans 320 0 0 0 ui_in[1]
port 6 nsew
flabel metal5 s 34338 30796 34398 30996 4 FreeSans 320 0 0 0 ui_in[2]
port 7 nsew
flabel metal5 s 33570 30796 33630 30996 4 FreeSans 320 0 0 0 ui_in[3]
port 8 nsew
flabel metal5 s 32802 30796 32862 30996 4 FreeSans 320 0 0 0 ui_in[4]
port 9 nsew
flabel metal5 s 32034 30796 32094 30996 4 FreeSans 320 0 0 0 ui_in[5]
port 10 nsew
flabel metal5 s 31266 30796 31326 30996 4 FreeSans 320 0 0 0 ui_in[6]
port 11 nsew
flabel metal5 s 30498 30796 30558 30996 4 FreeSans 320 0 0 0 ui_in[7]
port 12 nsew
flabel metal5 s 29730 30796 29790 30996 4 FreeSans 320 0 0 0 uio_in[0]
port 13 nsew
flabel metal5 s 28962 30796 29022 30996 4 FreeSans 320 0 0 0 uio_in[1]
port 14 nsew
flabel metal5 s 28194 30796 28254 30996 4 FreeSans 320 0 0 0 uio_in[2]
port 15 nsew
flabel metal5 s 27426 30796 27486 30996 4 FreeSans 320 0 0 0 uio_in[3]
port 16 nsew
flabel metal5 s 26658 30796 26718 30996 4 FreeSans 320 0 0 0 uio_in[4]
port 17 nsew
flabel metal5 s 25890 30796 25950 30996 4 FreeSans 320 0 0 0 uio_in[5]
port 18 nsew
flabel metal5 s 25122 30796 25182 30996 4 FreeSans 320 0 0 0 uio_in[6]
port 19 nsew
flabel metal5 s 24354 30796 24414 30996 4 FreeSans 320 0 0 0 uio_in[7]
port 20 nsew
flabel metal5 s 11298 30796 11358 30996 4 FreeSans 320 0 0 0 uio_oe[0]
port 21 nsew
flabel metal5 s 10530 30796 10590 30996 4 FreeSans 320 0 0 0 uio_oe[1]
port 22 nsew
flabel metal5 s 9762 30796 9822 30996 4 FreeSans 320 0 0 0 uio_oe[2]
port 23 nsew
flabel metal5 s 8994 30796 9054 30996 4 FreeSans 320 0 0 0 uio_oe[3]
port 24 nsew
flabel metal5 s 8226 30796 8286 30996 4 FreeSans 320 0 0 0 uio_oe[4]
port 25 nsew
flabel metal5 s 7458 30796 7518 30996 4 FreeSans 320 0 0 0 uio_oe[5]
port 26 nsew
flabel metal5 s 6690 30796 6750 30996 4 FreeSans 320 0 0 0 uio_oe[6]
port 27 nsew
flabel metal5 s 5922 30796 5982 30996 4 FreeSans 320 0 0 0 uio_oe[7]
port 28 nsew
flabel metal5 s 17442 30796 17502 30996 4 FreeSans 320 0 0 0 uio_out[0]
port 29 nsew
flabel metal5 s 16674 30796 16734 30996 4 FreeSans 320 0 0 0 uio_out[1]
port 30 nsew
flabel metal5 s 15906 30796 15966 30996 4 FreeSans 320 0 0 0 uio_out[2]
port 31 nsew
flabel metal5 s 15138 30796 15198 30996 4 FreeSans 320 0 0 0 uio_out[3]
port 32 nsew
flabel metal5 s 14370 30796 14430 30996 4 FreeSans 320 0 0 0 uio_out[4]
port 33 nsew
flabel metal5 s 13602 30796 13662 30996 4 FreeSans 320 0 0 0 uio_out[5]
port 34 nsew
flabel metal5 s 12834 30796 12894 30996 4 FreeSans 320 0 0 0 uio_out[6]
port 35 nsew
flabel metal5 s 12066 30796 12126 30996 4 FreeSans 320 0 0 0 uio_out[7]
port 36 nsew
flabel metal5 s 23586 30796 23646 30996 4 FreeSans 320 0 0 0 uo_out[0]
port 37 nsew
flabel metal5 s 22818 30796 22878 30996 4 FreeSans 320 0 0 0 uo_out[1]
port 38 nsew
flabel metal5 s 22050 30796 22110 30996 4 FreeSans 320 0 0 0 uo_out[2]
port 39 nsew
flabel metal5 s 21282 30796 21342 30996 4 FreeSans 320 0 0 0 uo_out[3]
port 40 nsew
flabel metal5 s 20514 30796 20574 30996 4 FreeSans 320 0 0 0 uo_out[4]
port 41 nsew
flabel metal5 s 19746 30796 19806 30996 4 FreeSans 320 0 0 0 uo_out[5]
port 42 nsew
flabel metal5 s 18978 30796 19038 30996 4 FreeSans 320 0 0 0 uo_out[6]
port 43 nsew
flabel metal5 s 18210 30796 18270 30996 4 FreeSans 320 0 0 0 uo_out[7]
port 44 nsew
flabel metal5 s 0 24596 200 24776 0 FreeSans 320 0 0 0 ua[0]
port 45 nsew
flabel metal5 s 0 21396 200 21576 0 FreeSans 320 0 0 0 ua[1]
port 46 nsew
flabel metal5 s 0 18196 200 18376 0 FreeSans 320 0 0 0 ua[2]
port 47 nsew
flabel metal5 s 0 14996 200 15176 0 FreeSans 320 0 0 0 ua[3]
port 48 nsew
flabel metal5 s 800 0 1240 30596 0 FreeSans 320 0 0 0 VGND
port 49 nsew
flabel metal5 s 39800 0 40240 30596 0 FreeSans 320 0 0 0 VPWR
port 50 nsew
<< properties >>
string FIXED_BBOX 0 0 40416 30996
<< end >>
