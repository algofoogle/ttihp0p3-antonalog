magic
tech ihp-sg13g2
magscale 1 2
timestamp 1747537721
<< nwell >>
rect -48 350 432 834
<< pwell >>
rect 50 56 366 292
rect -26 -56 410 56
<< nmos >>
rect 144 118 170 266
rect 246 118 272 266
<< pmos >>
rect 144 412 170 636
rect 212 412 238 636
<< ndiff >>
rect 76 252 144 266
rect 76 220 90 252
rect 122 220 144 252
rect 76 164 144 220
rect 76 132 90 164
rect 122 132 144 164
rect 76 118 144 132
rect 170 252 246 266
rect 170 220 192 252
rect 224 220 246 252
rect 170 164 246 220
rect 170 132 192 164
rect 224 132 246 164
rect 170 118 246 132
rect 272 252 340 266
rect 272 220 294 252
rect 326 220 340 252
rect 272 164 340 220
rect 272 132 294 164
rect 326 132 340 164
rect 272 118 340 132
<< pdiff >>
rect 72 622 144 636
rect 72 590 90 622
rect 122 590 144 622
rect 72 553 144 590
rect 72 521 90 553
rect 122 521 144 553
rect 72 483 144 521
rect 72 451 90 483
rect 122 451 144 483
rect 72 412 144 451
rect 170 412 212 636
rect 238 622 306 636
rect 238 590 260 622
rect 292 590 306 622
rect 238 553 306 590
rect 238 521 260 553
rect 292 521 306 553
rect 238 483 306 521
rect 238 451 260 483
rect 292 451 306 483
rect 238 412 306 451
<< ndiffc >>
rect 90 220 122 252
rect 90 132 122 164
rect 192 220 224 252
rect 192 132 224 164
rect 294 220 326 252
rect 294 132 326 164
<< pdiffc >>
rect 90 590 122 622
rect 90 521 122 553
rect 90 451 122 483
rect 260 590 292 622
rect 260 521 292 553
rect 260 451 292 483
<< psubdiff >>
rect 0 16 384 30
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 384 16
rect 0 -30 384 -16
<< nsubdiff >>
rect 0 772 384 786
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 384 772
rect 0 726 384 740
<< psubdiffcont >>
rect 32 -16 64 16
rect 128 -16 160 16
rect 224 -16 256 16
rect 320 -16 352 16
<< nsubdiffcont >>
rect 32 740 64 772
rect 128 740 160 772
rect 224 740 256 772
rect 320 740 352 772
<< poly >>
rect 144 636 170 672
rect 212 636 238 672
rect 144 397 170 412
rect 128 370 170 397
rect 70 353 170 370
rect 70 321 87 353
rect 119 321 170 353
rect 70 304 170 321
rect 212 397 238 412
rect 212 370 248 397
rect 212 353 308 370
rect 212 321 259 353
rect 291 321 308 353
rect 212 304 308 321
rect 144 266 170 304
rect 246 266 272 304
rect 144 82 170 118
rect 246 82 272 118
<< polycont >>
rect 87 321 119 353
rect 259 321 291 353
<< metal1 >>
rect 0 772 384 800
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 384 772
rect 0 712 384 740
rect 80 622 132 712
rect 80 590 90 622
rect 122 590 132 622
rect 80 553 132 590
rect 80 521 90 553
rect 122 521 132 553
rect 80 483 132 521
rect 248 622 308 625
rect 248 590 260 622
rect 292 590 308 622
rect 248 553 308 590
rect 248 521 260 553
rect 292 521 308 553
rect 248 487 308 521
rect 80 451 90 483
rect 122 451 132 483
rect 80 448 132 451
rect 174 483 308 487
rect 174 451 260 483
rect 292 451 308 483
rect 174 447 308 451
rect 70 353 136 400
rect 70 321 87 353
rect 119 321 136 353
rect 70 304 136 321
rect 174 270 208 447
rect 244 353 308 400
rect 244 321 259 353
rect 291 321 308 353
rect 244 304 308 321
rect 80 252 132 257
rect 80 220 90 252
rect 122 220 132 252
rect 80 164 132 220
rect 80 132 90 164
rect 122 132 132 164
rect 80 44 132 132
rect 174 252 227 270
rect 174 220 192 252
rect 224 220 227 252
rect 174 164 227 220
rect 174 132 192 164
rect 224 132 227 164
rect 174 121 227 132
rect 284 252 336 257
rect 284 220 294 252
rect 326 220 336 252
rect 284 164 336 220
rect 284 132 294 164
rect 326 132 336 164
rect 284 44 336 132
rect 0 16 384 44
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 384 16
rect 0 -44 384 -16
<< labels >>
flabel metal1 s 70 304 136 400 0 FreeSans 400 0 0 0 A
port 2 nsew
flabel metal1 s 0 712 384 800 0 FreeSans 400 0 0 0 VDD
port 3 nsew
flabel metal1 s 248 447 308 625 0 FreeSans 400 0 0 0 Y
port 4 nsew
flabel metal1 s 0 -44 384 44 0 FreeSans 400 0 0 0 VSS
port 5 nsew
flabel metal1 s 244 304 308 400 0 FreeSans 400 0 0 0 B
port 6 nsew
<< properties >>
string FIXED_BBOX 0 0 384 756
string GDS_END 11110
string GDS_FILE ../gds/controller.gds
string GDS_START 7312
<< end >>
