magic
tech ihp-sg13g2
magscale 1 2
timestamp 1747056038
<< nwell >>
rect -54 350 720 834
<< pwell >>
rect 24 56 652 314
rect -26 -56 698 56
<< nmos >>
rect 118 160 144 288
rect 226 144 252 288
rect 328 144 354 288
rect 430 144 456 288
rect 532 144 558 288
<< pmos >>
rect 118 412 144 612
rect 226 412 252 636
rect 328 412 354 636
rect 430 412 456 636
rect 532 412 558 636
<< ndiff >>
rect 50 274 118 288
rect 50 242 64 274
rect 96 242 118 274
rect 50 160 118 242
rect 144 274 226 288
rect 144 242 172 274
rect 204 242 226 274
rect 144 190 226 242
rect 144 160 172 190
rect 158 158 172 160
rect 204 158 226 190
rect 158 144 226 158
rect 252 262 328 288
rect 252 230 274 262
rect 306 230 328 262
rect 252 190 328 230
rect 252 158 274 190
rect 306 158 328 190
rect 252 144 328 158
rect 354 190 430 288
rect 354 158 376 190
rect 408 158 430 190
rect 354 144 430 158
rect 456 262 532 288
rect 456 230 478 262
rect 510 230 532 262
rect 456 190 532 230
rect 456 158 478 190
rect 510 158 532 190
rect 456 144 532 158
rect 558 262 626 288
rect 558 230 580 262
rect 612 230 626 262
rect 558 190 626 230
rect 558 158 580 190
rect 612 158 626 190
rect 558 144 626 158
<< pdiff >>
rect 158 622 226 636
rect 158 612 172 622
rect 50 598 118 612
rect 50 566 64 598
rect 96 566 118 598
rect 50 528 118 566
rect 50 496 64 528
rect 96 496 118 528
rect 50 458 118 496
rect 50 426 64 458
rect 96 426 118 458
rect 50 412 118 426
rect 144 590 172 612
rect 204 590 226 622
rect 144 543 226 590
rect 144 511 172 543
rect 204 511 226 543
rect 144 458 226 511
rect 144 426 172 458
rect 204 426 226 458
rect 144 412 226 426
rect 252 622 328 636
rect 252 590 274 622
rect 306 590 328 622
rect 252 543 328 590
rect 252 511 274 543
rect 306 511 328 543
rect 252 412 328 511
rect 354 527 430 636
rect 354 495 376 527
rect 408 495 430 527
rect 354 458 430 495
rect 354 426 376 458
rect 408 426 430 458
rect 354 412 430 426
rect 456 622 532 636
rect 456 590 478 622
rect 510 590 532 622
rect 456 543 532 590
rect 456 511 478 543
rect 510 511 532 543
rect 456 458 532 511
rect 456 426 478 458
rect 510 426 532 458
rect 456 412 532 426
rect 558 622 626 636
rect 558 590 580 622
rect 612 590 626 622
rect 558 543 626 590
rect 558 511 580 543
rect 612 511 626 543
rect 558 458 626 511
rect 558 426 580 458
rect 612 426 626 458
rect 558 412 626 426
<< ndiffc >>
rect 64 242 96 274
rect 172 242 204 274
rect 172 158 204 190
rect 274 230 306 262
rect 274 158 306 190
rect 376 158 408 190
rect 478 230 510 262
rect 478 158 510 190
rect 580 230 612 262
rect 580 158 612 190
<< pdiffc >>
rect 64 566 96 598
rect 64 496 96 528
rect 64 426 96 458
rect 172 590 204 622
rect 172 511 204 543
rect 172 426 204 458
rect 274 590 306 622
rect 274 511 306 543
rect 376 495 408 527
rect 376 426 408 458
rect 478 590 510 622
rect 478 511 510 543
rect 478 426 510 458
rect 580 590 612 622
rect 580 511 612 543
rect 580 426 612 458
<< psubdiff >>
rect 0 16 672 30
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 608 16
rect 640 -16 672 16
rect 0 -30 672 -16
<< nsubdiff >>
rect 0 772 672 786
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 608 772
rect 640 740 672 772
rect 0 726 672 740
<< psubdiffcont >>
rect 32 -16 64 16
rect 128 -16 160 16
rect 224 -16 256 16
rect 320 -16 352 16
rect 416 -16 448 16
rect 512 -16 544 16
rect 608 -16 640 16
<< nsubdiffcont >>
rect 32 740 64 772
rect 128 740 160 772
rect 224 740 256 772
rect 320 740 352 772
rect 416 740 448 772
rect 512 740 544 772
rect 608 740 640 772
<< poly >>
rect 118 612 144 648
rect 226 636 252 672
rect 328 636 354 672
rect 430 636 456 672
rect 532 636 558 672
rect 118 288 144 412
rect 226 387 252 412
rect 180 373 252 387
rect 180 341 194 373
rect 226 341 252 373
rect 180 327 252 341
rect 226 288 252 327
rect 328 379 354 412
rect 430 379 456 412
rect 328 365 496 379
rect 328 333 450 365
rect 482 333 496 365
rect 328 319 496 333
rect 328 288 354 319
rect 430 288 456 319
rect 532 288 558 412
rect 118 140 144 160
rect 70 126 144 140
rect 70 94 84 126
rect 116 94 144 126
rect 70 80 144 94
rect 226 71 252 144
rect 328 108 354 144
rect 430 108 456 144
rect 532 71 558 144
rect 226 45 558 71
rect 226 44 252 45
rect 532 44 558 45
<< polycont >>
rect 194 341 226 373
rect 450 333 482 365
rect 84 94 116 126
<< metal1 >>
rect 0 772 672 800
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 608 772
rect 640 740 672 772
rect 0 712 672 740
rect 162 622 214 712
rect 54 598 106 608
rect 54 566 64 598
rect 96 566 106 598
rect 54 528 106 566
rect 54 496 64 528
rect 96 496 106 528
rect 54 458 106 496
rect 54 426 64 458
rect 96 426 106 458
rect 54 373 106 426
rect 162 590 172 622
rect 204 590 214 622
rect 162 543 214 590
rect 162 511 172 543
rect 204 511 214 543
rect 162 458 214 511
rect 264 622 520 652
rect 264 590 274 622
rect 306 616 478 622
rect 306 590 316 616
rect 264 543 316 590
rect 468 590 478 616
rect 510 590 520 622
rect 264 511 274 543
rect 306 511 316 543
rect 264 495 316 511
rect 366 527 418 580
rect 366 495 376 527
rect 408 495 418 527
rect 162 426 172 458
rect 204 426 214 458
rect 366 458 418 495
rect 366 440 376 458
rect 162 416 214 426
rect 272 426 376 440
rect 408 426 418 458
rect 272 400 418 426
rect 468 543 520 590
rect 468 511 478 543
rect 510 511 520 543
rect 468 458 520 511
rect 468 426 478 458
rect 510 426 520 458
rect 468 416 520 426
rect 570 622 622 712
rect 570 590 580 622
rect 612 590 622 622
rect 570 543 622 590
rect 570 511 580 543
rect 612 511 622 543
rect 570 458 622 511
rect 570 426 580 458
rect 612 426 622 458
rect 570 416 622 426
rect 54 341 194 373
rect 226 341 236 373
rect 54 274 106 341
rect 54 242 64 274
rect 96 242 106 274
rect 54 232 106 242
rect 162 274 214 284
rect 162 242 172 274
rect 204 242 214 274
rect 272 272 316 400
rect 434 333 450 365
rect 482 333 592 365
rect 434 308 592 333
rect 74 126 126 192
rect 74 94 84 126
rect 116 94 126 126
rect 74 80 126 94
rect 162 190 214 242
rect 162 158 172 190
rect 204 158 214 190
rect 162 44 214 158
rect 264 262 520 272
rect 264 230 274 262
rect 306 232 478 262
rect 306 230 316 232
rect 264 190 316 230
rect 468 230 478 232
rect 510 230 520 262
rect 264 158 274 190
rect 306 158 316 190
rect 264 144 316 158
rect 366 190 418 196
rect 366 158 376 190
rect 408 158 418 190
rect 366 44 418 158
rect 468 190 520 230
rect 468 158 478 190
rect 510 158 520 190
rect 468 144 520 158
rect 570 262 622 272
rect 570 230 580 262
rect 612 230 622 262
rect 570 190 622 230
rect 570 158 580 190
rect 612 158 622 190
rect 570 44 622 158
rect 0 16 672 44
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 608 16
rect 640 -16 672 16
rect 0 -44 672 -16
<< labels >>
flabel metal1 s 434 308 592 365 0 FreeSans 400 0 0 0 A
port 2 nsew
flabel metal1 s 74 80 126 192 0 FreeSans 400 0 0 0 B_N
port 3 nsew
flabel metal1 s 0 712 672 800 0 FreeSans 400 0 0 0 VDD
port 4 nsew
flabel metal1 s 264 232 520 272 0 FreeSans 400 0 0 0 Y
port 5 nsew
flabel metal1 s 0 -44 672 44 0 FreeSans 400 0 0 0 VSS
port 6 nsew
<< properties >>
string FIXED_BBOX 0 0 672 756
string GDS_END 225190
string GDS_FILE ../gds/controller.gds
string GDS_START 220062
<< end >>
