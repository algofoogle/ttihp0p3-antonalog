magic
tech ihp-sg13g2
timestamp 1747537721
<< nwell >>
rect -24 175 264 417
<< pwell >>
rect 103 116 210 135
rect -2 28 210 116
rect -13 -28 253 28
<< nmos >>
rect 45 48 58 103
rect 96 48 109 103
rect 150 48 163 122
<< pmos >>
rect 45 246 58 330
rect 96 246 109 330
rect 150 218 163 330
<< ndiff >>
rect 116 105 150 122
rect 116 103 123 105
rect 11 96 45 103
rect 11 80 18 96
rect 34 80 45 96
rect 11 48 45 80
rect 58 96 96 103
rect 58 80 69 96
rect 85 80 96 96
rect 58 48 96 80
rect 109 89 123 103
rect 139 89 150 105
rect 109 71 150 89
rect 109 55 122 71
rect 138 55 150 71
rect 109 48 150 55
rect 163 115 197 122
rect 163 99 174 115
rect 190 99 197 115
rect 163 71 197 99
rect 163 55 174 71
rect 190 55 197 71
rect 163 48 197 55
<< pdiff >>
rect 11 323 45 330
rect 11 307 18 323
rect 34 307 45 323
rect 11 269 45 307
rect 11 253 18 269
rect 34 253 45 269
rect 11 246 45 253
rect 58 246 96 330
rect 109 323 150 330
rect 109 307 122 323
rect 138 307 150 323
rect 109 283 150 307
rect 109 267 122 283
rect 138 267 150 283
rect 109 249 150 267
rect 109 246 123 249
rect 116 233 123 246
rect 139 233 150 249
rect 116 218 150 233
rect 163 323 199 330
rect 163 307 175 323
rect 191 307 199 323
rect 163 283 199 307
rect 163 267 175 283
rect 191 267 199 283
rect 163 241 199 267
rect 163 225 175 241
rect 191 225 199 241
rect 163 218 199 225
<< ndiffc >>
rect 18 80 34 96
rect 69 80 85 96
rect 123 89 139 105
rect 122 55 138 71
rect 174 99 190 115
rect 174 55 190 71
<< pdiffc >>
rect 18 307 34 323
rect 18 253 34 269
rect 122 307 138 323
rect 122 267 138 283
rect 123 233 139 249
rect 175 307 191 323
rect 175 267 191 283
rect 175 225 191 241
<< psubdiff >>
rect 0 8 240 15
rect 0 -8 16 8
rect 32 -8 64 8
rect 80 -8 112 8
rect 128 -8 160 8
rect 176 -8 208 8
rect 224 -8 240 8
rect 0 -15 240 -8
<< nsubdiff >>
rect 0 386 240 393
rect 0 370 16 386
rect 32 370 64 386
rect 80 370 112 386
rect 128 370 160 386
rect 176 370 208 386
rect 224 370 240 386
rect 0 363 240 370
<< psubdiffcont >>
rect 16 -8 32 8
rect 64 -8 80 8
rect 112 -8 128 8
rect 160 -8 176 8
rect 208 -8 224 8
<< nsubdiffcont >>
rect 16 370 32 386
rect 64 370 80 386
rect 112 370 128 386
rect 160 370 176 386
rect 208 370 224 386
<< poly >>
rect 45 330 58 352
rect 96 330 109 352
rect 150 330 163 353
rect 45 239 58 246
rect 45 232 78 239
rect 45 216 54 232
rect 70 216 78 232
rect 45 209 78 216
rect 45 103 58 209
rect 96 191 109 246
rect 84 184 114 191
rect 84 168 91 184
rect 107 168 114 184
rect 84 161 114 168
rect 96 103 109 161
rect 150 160 163 218
rect 135 153 167 160
rect 135 137 143 153
rect 159 137 167 153
rect 135 129 167 137
rect 150 122 163 129
rect 45 22 58 48
rect 96 22 109 48
rect 150 22 163 48
<< polycont >>
rect 54 216 70 232
rect 91 168 107 184
rect 143 137 159 153
<< metal1 >>
rect 0 386 240 400
rect 0 370 16 386
rect 32 370 64 386
rect 80 370 112 386
rect 128 370 160 386
rect 176 370 208 386
rect 224 370 240 386
rect 0 356 240 370
rect 118 323 144 356
rect 13 307 18 323
rect 34 307 39 323
rect 13 269 39 307
rect 13 253 18 269
rect 34 253 39 269
rect 117 307 122 323
rect 138 307 144 323
rect 117 283 144 307
rect 117 267 122 283
rect 138 267 144 283
rect 13 139 31 253
rect 65 235 90 265
rect 49 232 90 235
rect 49 216 54 232
rect 70 216 90 232
rect 117 249 144 267
rect 117 233 123 249
rect 139 233 144 249
rect 117 225 144 233
rect 170 307 175 323
rect 191 307 196 323
rect 170 283 196 307
rect 170 267 175 283
rect 191 267 196 283
rect 170 241 196 267
rect 170 225 175 241
rect 191 225 196 241
rect 49 213 90 216
rect 71 184 113 194
rect 71 168 91 184
rect 107 168 113 184
rect 71 157 113 168
rect 135 153 161 158
rect 135 139 143 153
rect 13 137 143 139
rect 159 137 161 153
rect 13 131 161 137
rect 13 123 152 131
rect 13 116 90 123
rect 64 96 90 116
rect 179 115 195 225
rect 13 80 18 96
rect 34 80 39 96
rect 64 80 69 96
rect 85 80 90 96
rect 118 89 123 105
rect 139 89 144 105
rect 13 22 39 80
rect 118 71 144 89
rect 118 55 122 71
rect 138 55 144 71
rect 169 99 174 115
rect 190 99 195 115
rect 169 71 195 99
rect 169 55 174 71
rect 190 55 195 71
rect 118 22 144 55
rect 0 8 240 22
rect 0 -8 16 8
rect 32 -8 64 8
rect 80 -8 112 8
rect 128 -8 160 8
rect 176 -8 208 8
rect 224 -8 240 8
rect 0 -22 240 -8
<< labels >>
flabel metal1 s 71 157 113 194 0 FreeSans 200 0 0 0 A
port 2 nsew
flabel metal1 s 0 -22 240 22 0 FreeSans 200 0 0 0 VSS
port 3 nsew
flabel metal1 s 65 213 90 265 0 FreeSans 200 0 0 0 B
port 4 nsew
flabel metal1 s 179 115 195 225 0 FreeSans 200 0 0 0 X
port 5 nsew
flabel metal1 s 0 356 240 400 0 FreeSans 200 0 0 0 VDD
port 6 nsew
<< properties >>
string FIXED_BBOX 0 0 240 378
string GDS_END 65488
string GDS_FILE ../gds/controller.gds
string GDS_START 61194
<< end >>
