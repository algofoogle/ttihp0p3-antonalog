magic
tech ihp-sg13g2
timestamp 1747537721
<< nwell >>
rect -24 175 216 417
<< pwell >>
rect 13 28 172 146
rect -13 -28 205 28
<< nmos >>
rect 60 59 73 133
rect 111 59 124 133
<< pmos >>
rect 59 206 72 318
rect 111 206 124 318
<< ndiff >>
rect 26 125 60 133
rect 26 109 33 125
rect 49 109 60 125
rect 26 83 60 109
rect 26 67 33 83
rect 49 67 60 83
rect 26 59 60 67
rect 73 125 111 133
rect 73 109 84 125
rect 100 109 111 125
rect 73 83 111 109
rect 73 67 84 83
rect 100 67 111 83
rect 73 59 111 67
rect 124 125 159 133
rect 124 109 136 125
rect 152 109 159 125
rect 124 83 159 109
rect 124 67 136 83
rect 152 67 159 83
rect 124 59 159 67
<< pdiff >>
rect 25 309 59 318
rect 25 293 32 309
rect 48 293 59 309
rect 25 275 59 293
rect 25 259 32 275
rect 48 259 59 275
rect 25 239 59 259
rect 25 223 32 239
rect 48 223 59 239
rect 25 206 59 223
rect 72 309 111 318
rect 72 293 84 309
rect 100 293 111 309
rect 72 270 111 293
rect 72 254 84 270
rect 100 254 111 270
rect 72 230 111 254
rect 72 214 84 230
rect 100 214 111 230
rect 72 206 111 214
rect 124 309 158 318
rect 124 293 135 309
rect 151 293 158 309
rect 124 270 158 293
rect 124 254 135 270
rect 151 254 158 270
rect 124 230 158 254
rect 124 214 135 230
rect 151 214 158 230
rect 124 206 158 214
<< ndiffc >>
rect 33 109 49 125
rect 33 67 49 83
rect 84 109 100 125
rect 84 67 100 83
rect 136 109 152 125
rect 136 67 152 83
<< pdiffc >>
rect 32 293 48 309
rect 32 259 48 275
rect 32 223 48 239
rect 84 293 100 309
rect 84 254 100 270
rect 84 214 100 230
rect 135 293 151 309
rect 135 254 151 270
rect 135 214 151 230
<< psubdiff >>
rect 0 8 192 15
rect 0 -8 16 8
rect 32 -8 64 8
rect 80 -8 112 8
rect 128 -8 160 8
rect 176 -8 192 8
rect 0 -15 192 -8
<< nsubdiff >>
rect 0 386 192 393
rect 0 370 16 386
rect 32 370 64 386
rect 80 370 112 386
rect 128 370 160 386
rect 176 370 192 386
rect 0 363 192 370
<< psubdiffcont >>
rect 16 -8 32 8
rect 64 -8 80 8
rect 112 -8 128 8
rect 160 -8 176 8
<< nsubdiffcont >>
rect 16 370 32 386
rect 64 370 80 386
rect 112 370 128 386
rect 160 370 176 386
<< poly >>
rect 59 318 72 336
rect 111 318 124 336
rect 59 198 72 206
rect 111 198 124 206
rect 59 185 78 198
rect 30 176 78 185
rect 30 160 39 176
rect 55 167 78 176
rect 105 167 124 198
rect 55 160 124 167
rect 30 152 124 160
rect 60 133 73 152
rect 111 133 124 152
rect 60 41 73 59
rect 111 41 124 59
<< polycont >>
rect 39 160 55 176
<< metal1 >>
rect 0 386 192 400
rect 0 370 16 386
rect 32 370 64 386
rect 80 370 112 386
rect 128 370 160 386
rect 176 370 192 386
rect 0 356 192 370
rect 27 309 53 356
rect 27 293 32 309
rect 48 293 53 309
rect 27 275 53 293
rect 27 259 32 275
rect 48 259 53 275
rect 27 239 53 259
rect 27 223 32 239
rect 48 223 53 239
rect 27 218 53 223
rect 82 309 102 318
rect 82 293 84 309
rect 100 293 102 309
rect 82 270 102 293
rect 82 254 84 270
rect 100 254 102 270
rect 82 230 102 254
rect 82 214 84 230
rect 100 214 102 230
rect 18 176 63 200
rect 18 160 39 176
rect 55 160 63 176
rect 18 152 63 160
rect 28 125 54 130
rect 28 109 33 125
rect 49 109 54 125
rect 28 83 54 109
rect 28 67 33 83
rect 49 67 54 83
rect 28 22 54 67
rect 82 125 102 214
rect 132 309 153 356
rect 132 293 135 309
rect 151 293 153 309
rect 132 270 153 293
rect 132 254 135 270
rect 151 254 153 270
rect 132 230 153 254
rect 132 214 135 230
rect 151 214 153 230
rect 132 209 153 214
rect 82 109 84 125
rect 100 109 102 125
rect 82 83 102 109
rect 82 67 84 83
rect 100 67 102 83
rect 82 57 102 67
rect 134 125 154 130
rect 134 109 136 125
rect 152 109 154 125
rect 134 83 154 109
rect 134 67 136 83
rect 152 67 154 83
rect 134 22 154 67
rect 0 8 192 22
rect 0 -8 16 8
rect 32 -8 64 8
rect 80 -8 112 8
rect 128 -8 160 8
rect 176 -8 192 8
rect 0 -22 192 -8
<< labels >>
flabel metal1 s 0 -22 192 22 0 FreeSans 200 0 0 0 VSS
port 2 nsew
flabel metal1 s 0 356 192 400 0 FreeSans 200 0 0 0 VDD
port 3 nsew
flabel metal1 s 82 57 102 318 0 FreeSans 200 0 0 0 Y
port 4 nsew
flabel metal1 s 18 152 63 200 0 FreeSans 200 0 0 0 A
port 5 nsew
<< properties >>
string FIXED_BBOX 0 0 192 378
string GDS_END 93350
string GDS_FILE ../gds/controller.gds
string GDS_START 89662
<< end >>
