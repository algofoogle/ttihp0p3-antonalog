magic
tech ihp-sg13g2
magscale 1 2
timestamp 1746816402
<< nwell >>
rect -48 350 720 834
<< pwell >>
rect 68 56 640 296
rect -26 -56 698 56
<< nmos >>
rect 162 160 188 270
rect 291 122 317 270
rect 411 122 437 270
rect 496 122 522 270
<< pmos >>
rect 184 412 210 580
rect 292 412 318 636
rect 394 412 420 636
rect 496 412 522 636
<< ndiff >>
rect 94 231 162 270
rect 94 199 108 231
rect 140 199 162 231
rect 94 160 162 199
rect 188 182 291 270
rect 188 160 227 182
rect 202 150 227 160
rect 259 150 291 182
rect 202 122 291 150
rect 317 122 411 270
rect 437 122 496 270
rect 522 252 614 270
rect 522 220 565 252
rect 597 220 614 252
rect 522 171 614 220
rect 522 139 544 171
rect 576 139 614 171
rect 522 122 614 139
<< pdiff >>
rect 224 621 292 636
rect 224 589 238 621
rect 270 589 292 621
rect 224 580 292 589
rect 116 566 184 580
rect 116 534 130 566
rect 162 534 184 566
rect 116 483 184 534
rect 116 451 130 483
rect 162 451 184 483
rect 116 412 184 451
rect 210 551 292 580
rect 210 519 238 551
rect 270 519 292 551
rect 210 467 292 519
rect 210 435 238 467
rect 270 435 292 467
rect 210 412 292 435
rect 318 621 394 636
rect 318 589 340 621
rect 372 589 394 621
rect 318 553 394 589
rect 318 521 340 553
rect 372 521 394 553
rect 318 483 394 521
rect 318 451 340 483
rect 372 451 394 483
rect 318 412 394 451
rect 420 621 496 636
rect 420 589 442 621
rect 474 589 496 621
rect 420 551 496 589
rect 420 519 442 551
rect 474 519 496 551
rect 420 412 496 519
rect 522 621 590 636
rect 522 589 544 621
rect 576 589 590 621
rect 522 540 590 589
rect 522 508 544 540
rect 576 508 590 540
rect 522 461 590 508
rect 522 429 544 461
rect 576 429 590 461
rect 522 412 590 429
<< ndiffc >>
rect 108 199 140 231
rect 227 150 259 182
rect 565 220 597 252
rect 544 139 576 171
<< pdiffc >>
rect 238 589 270 621
rect 130 534 162 566
rect 130 451 162 483
rect 238 519 270 551
rect 238 435 270 467
rect 340 589 372 621
rect 340 521 372 553
rect 340 451 372 483
rect 442 589 474 621
rect 442 519 474 551
rect 544 589 576 621
rect 544 508 576 540
rect 544 429 576 461
<< psubdiff >>
rect 0 16 672 30
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 608 16
rect 640 -16 672 16
rect 0 -30 672 -16
<< nsubdiff >>
rect 0 772 672 786
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 608 772
rect 640 740 672 772
rect 0 726 672 740
<< psubdiffcont >>
rect 32 -16 64 16
rect 128 -16 160 16
rect 224 -16 256 16
rect 320 -16 352 16
rect 416 -16 448 16
rect 512 -16 544 16
rect 608 -16 640 16
<< nsubdiffcont >>
rect 32 740 64 772
rect 128 740 160 772
rect 224 740 256 772
rect 320 740 352 772
rect 416 740 448 772
rect 512 740 544 772
rect 608 740 640 772
<< poly >>
rect 292 636 318 672
rect 394 636 420 672
rect 496 636 522 672
rect 184 580 210 616
rect 184 374 210 412
rect 292 374 318 412
rect 394 380 420 412
rect 151 360 211 374
rect 151 328 165 360
rect 197 328 211 360
rect 151 314 211 328
rect 270 360 330 374
rect 270 328 284 360
rect 316 328 330 360
rect 270 314 330 328
rect 393 363 453 380
rect 496 371 522 412
rect 393 331 407 363
rect 439 331 453 363
rect 393 317 453 331
rect 494 357 555 371
rect 494 325 509 357
rect 541 325 555 357
rect 162 270 188 314
rect 291 270 317 314
rect 411 270 437 317
rect 494 311 555 325
rect 496 270 522 311
rect 162 124 188 160
rect 291 86 317 122
rect 411 86 437 122
rect 496 86 522 122
<< polycont >>
rect 165 328 197 360
rect 284 328 316 360
rect 407 331 439 363
rect 509 325 541 357
<< metal1 >>
rect 0 772 672 800
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 608 772
rect 640 740 672 772
rect 0 712 672 740
rect 228 621 280 712
rect 228 589 238 621
rect 270 589 280 621
rect 88 566 172 572
rect 88 534 130 566
rect 162 534 172 566
rect 88 483 172 534
rect 88 451 130 483
rect 162 451 172 483
rect 88 447 172 451
rect 228 551 280 589
rect 228 519 238 551
rect 270 519 280 551
rect 228 467 280 519
rect 88 274 122 447
rect 228 435 238 467
rect 270 435 280 467
rect 330 621 382 626
rect 330 589 340 621
rect 372 589 382 621
rect 330 553 382 589
rect 330 521 340 553
rect 372 521 382 553
rect 330 483 382 521
rect 432 621 484 712
rect 432 589 442 621
rect 474 589 484 621
rect 432 551 484 589
rect 432 519 442 551
rect 474 519 484 551
rect 432 515 484 519
rect 528 621 626 640
rect 528 589 544 621
rect 576 589 626 621
rect 528 540 626 589
rect 330 451 340 483
rect 372 478 382 483
rect 528 508 544 540
rect 576 508 626 540
rect 528 478 626 508
rect 372 461 626 478
rect 372 451 544 461
rect 330 440 544 451
rect 228 434 280 435
rect 528 429 544 440
rect 576 429 626 461
rect 528 420 626 429
rect 158 360 234 397
rect 158 328 165 360
rect 197 328 234 360
rect 158 314 234 328
rect 270 360 336 397
rect 270 328 284 360
rect 316 328 336 360
rect 270 314 336 328
rect 380 363 450 400
rect 380 331 407 363
rect 439 331 450 363
rect 380 314 450 331
rect 486 357 556 374
rect 486 325 509 357
rect 541 325 556 357
rect 486 308 556 325
rect 486 274 518 308
rect 88 240 518 274
rect 592 272 626 420
rect 554 252 626 272
rect 88 231 142 240
rect 88 199 108 231
rect 140 199 142 231
rect 554 220 565 252
rect 597 220 626 252
rect 554 202 626 220
rect 88 176 142 199
rect 216 182 270 192
rect 216 150 227 182
rect 259 150 270 182
rect 216 44 270 150
rect 526 171 626 202
rect 526 139 544 171
rect 576 139 626 171
rect 526 124 626 139
rect 0 16 672 44
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 608 16
rect 640 -16 672 16
rect 0 -44 672 -16
<< labels >>
flabel metal1 s 158 314 234 397 0 FreeSans 400 0 0 0 A_N
port 2 nsew
flabel metal1 s 528 420 626 640 0 FreeSans 400 0 0 0 Y
port 3 nsew
flabel metal1 s 0 712 672 800 0 FreeSans 400 0 0 0 VDD
port 4 nsew
flabel metal1 s 0 -44 672 44 0 FreeSans 400 0 0 0 VSS
port 5 nsew
flabel metal1 s 380 314 450 400 0 FreeSans 400 0 0 0 B
port 6 nsew
flabel metal1 s 270 314 336 397 0 FreeSans 400 0 0 0 C
port 7 nsew
<< properties >>
string FIXED_BBOX 0 0 672 756
string GDS_END 128044
string GDS_FILE ../gds/controller.gds
string GDS_START 122214
<< end >>
