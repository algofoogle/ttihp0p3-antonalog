magic
tech ihp-sg13g2
timestamp 1747574105
<< pwell >>
rect -1423 412 1971 422
rect -1431 -542 1971 412
<< psubdiff >>
rect -1400 384 1940 391
rect -1400 368 -1324 384
rect 1864 368 1940 384
rect -1400 361 1940 368
rect -1400 315 -1370 361
rect -1400 -435 -1393 315
rect -1377 -435 -1370 315
rect -1400 -481 -1370 -435
rect 1910 315 1940 361
rect 1910 -435 1917 315
rect 1933 -435 1940 315
rect 1910 -481 1940 -435
rect -1400 -488 1940 -481
rect -1400 -504 -1324 -488
rect 1864 -504 1940 -488
rect -1400 -511 1940 -504
<< psubdiffcont >>
rect -1324 368 1864 384
rect -1393 -435 -1377 315
rect 1917 -435 1933 315
rect -1324 -504 1864 -488
<< metal1 >>
rect -1393 368 -1324 384
rect 1864 368 1933 384
rect -1393 315 -1311 368
rect -1377 -360 -1311 315
rect 1917 315 1933 368
rect -1292 240 -1066 283
rect -1040 240 -814 283
rect -788 240 -562 283
rect -536 240 -436 313
rect -662 183 -562 240
rect -410 183 -310 283
rect -284 240 -58 283
rect -32 240 194 283
rect 220 240 320 313
rect -662 140 -310 183
rect 94 183 194 240
rect 346 183 446 283
rect 472 240 698 283
rect 724 240 950 283
rect 976 240 1076 313
rect 94 140 446 183
rect 850 183 950 240
rect 1102 183 1202 283
rect 1228 240 1454 283
rect 1480 240 1706 313
rect 1732 240 1832 313
rect 850 140 1202 183
rect -1040 -303 -688 -260
rect -1040 -360 -940 -303
rect -1377 -435 -1192 -360
rect -1166 -403 -940 -360
rect -914 -433 -814 -360
rect -788 -403 -688 -303
rect -284 -303 68 -260
rect -284 -360 -184 -303
rect -662 -403 -436 -360
rect -410 -403 -184 -360
rect -158 -433 -58 -360
rect -32 -403 68 -303
rect 472 -303 824 -260
rect 472 -360 572 -303
rect 94 -403 320 -360
rect 346 -403 572 -360
rect 598 -433 698 -360
rect 724 -403 824 -303
rect 1228 -303 1580 -260
rect 1228 -360 1328 -303
rect 850 -403 1076 -360
rect 1102 -403 1328 -360
rect 1354 -433 1454 -360
rect 1480 -403 1580 -303
rect 1606 -403 1832 -360
rect -1393 -488 -1192 -435
rect 1917 -488 1933 -435
rect -1393 -504 -1324 -488
rect 1864 -504 1933 -488
use rhigh  res
array 0 24 126 0 0 686
timestamp 1746838591
transform 1 0 -1292 0 1 -360
box 0 -43 100 643
<< labels >>
flabel metal1 -1292 240 -1066 283 0 FreeSans 160 0 0 0 wg0
flabel metal1 -1166 -403 -940 -360 0 FreeSans 160 0 0 0 wJ0
flabel metal1 -1040 240 -814 283 0 FreeSans 160 0 0 0 wi0
flabel metal1 -899 -418 -869 -388 0 FreeSans 160 0 0 0 IN[0]
port 0 nsew
flabel metal1 -788 240 -562 283 0 FreeSans 160 0 0 0 wJ1
flabel metal1 -662 -403 -436 -360 0 FreeSans 160 0 0 0 wi1
flabel metal1 -521 268 -491 298 0 FreeSans 160 0 0 0 IN[1]
port 1 nsew
flabel metal1 -410 -403 -184 -360 0 FreeSans 160 0 0 0 wJ2
flabel metal1 -284 240 -58 283 0 FreeSans 160 0 0 0 wi2
flabel metal1 -143 -418 -113 -388 0 FreeSans 160 0 0 0 IN[2]
port 2 nsew
flabel metal1 -32 240 194 283 0 FreeSans 160 0 0 0 wJ3
flabel metal1 94 -403 320 -360 0 FreeSans 160 0 0 0 wi3
flabel metal1 235 268 265 298 0 FreeSans 160 0 0 0 IN[3]
port 3 nsew
flabel metal1 346 -403 572 -360 0 FreeSans 160 0 0 0 wJ4
flabel metal1 472 240 698 283 0 FreeSans 160 0 0 0 wi4
flabel metal1 613 -418 643 -388 0 FreeSans 160 0 0 0 IN[4]
port 4 nsew
flabel metal1 724 240 950 283 0 FreeSans 160 0 0 0 wJ5
flabel metal1 850 -403 1076 -360 0 FreeSans 160 0 0 0 wi5
flabel metal1 991 268 1021 298 0 FreeSans 160 0 0 0 IN[5]
port 5 nsew
flabel metal1 1102 -403 1328 -360 0 FreeSans 160 0 0 0 wJ6
flabel metal1 1228 240 1454 283 0 FreeSans 160 0 0 0 wi6
flabel metal1 1369 -418 1399 -388 0 FreeSans 160 0 0 0 IN[6]
port 6 nsew
flabel metal1 1606 -403 1832 -360 0 FreeSans 160 0 0 0 wi7
flabel metal1 1747 268 1777 298 0 FreeSans 160 0 0 0 IN[7]
port 7 nsew
flabel metal1 1495 268 1525 298 0 FreeSans 160 0 0 0 OUT
port 8 nsew
flabel metal1 -1285 -435 -1255 -405 0 FreeSans 160 0 0 0 GND
port 9 nsew
<< end >>
