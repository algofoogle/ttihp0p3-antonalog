magic
tech ihp-sg13g2
timestamp 1747537721
<< nwell >>
rect -24 175 360 417
<< pwell >>
rect 213 127 317 146
rect 23 28 317 127
rect -13 -28 349 28
<< nmos >>
rect 70 59 83 114
rect 121 59 134 114
rect 206 59 219 114
rect 257 59 270 133
<< pmos >>
rect 70 206 83 306
rect 109 206 122 306
rect 166 206 179 306
rect 251 206 264 318
<< ndiff >>
rect 226 114 257 133
rect 36 94 70 114
rect 36 78 43 94
rect 59 78 70 94
rect 36 59 70 78
rect 83 88 121 114
rect 83 72 94 88
rect 110 72 121 88
rect 83 59 121 72
rect 134 92 206 114
rect 134 76 145 92
rect 161 76 179 92
rect 195 76 206 92
rect 134 59 206 76
rect 219 88 257 114
rect 219 72 230 88
rect 246 72 257 88
rect 219 59 257 72
rect 270 125 304 133
rect 270 109 281 125
rect 297 109 304 125
rect 270 82 304 109
rect 270 66 281 82
rect 297 66 304 82
rect 270 59 304 66
<< pdiff >>
rect 214 306 251 318
rect 36 298 70 306
rect 36 282 43 298
rect 59 282 70 298
rect 36 241 70 282
rect 36 225 43 241
rect 59 225 70 241
rect 36 206 70 225
rect 83 206 109 306
rect 122 206 166 306
rect 179 299 251 306
rect 179 283 190 299
rect 206 283 224 299
rect 240 283 251 299
rect 179 265 251 283
rect 179 249 190 265
rect 206 249 224 265
rect 240 249 251 265
rect 179 206 251 249
rect 264 310 298 318
rect 264 294 275 310
rect 291 294 298 310
rect 264 270 298 294
rect 264 254 275 270
rect 291 254 298 270
rect 264 230 298 254
rect 264 214 275 230
rect 291 214 298 230
rect 264 206 298 214
<< ndiffc >>
rect 43 78 59 94
rect 94 72 110 88
rect 145 76 161 92
rect 179 76 195 92
rect 230 72 246 88
rect 281 109 297 125
rect 281 66 297 82
<< pdiffc >>
rect 43 282 59 298
rect 43 225 59 241
rect 190 283 206 299
rect 224 283 240 299
rect 190 249 206 265
rect 224 249 240 265
rect 275 294 291 310
rect 275 254 291 270
rect 275 214 291 230
<< psubdiff >>
rect 0 8 336 15
rect 0 -8 16 8
rect 32 -8 64 8
rect 80 -8 112 8
rect 128 -8 160 8
rect 176 -8 208 8
rect 224 -8 256 8
rect 272 -8 304 8
rect 320 -8 336 8
rect 0 -15 336 -8
<< nsubdiff >>
rect 0 386 336 393
rect 0 370 16 386
rect 32 370 64 386
rect 80 370 112 386
rect 128 370 160 386
rect 176 370 208 386
rect 224 370 256 386
rect 272 370 304 386
rect 320 370 336 386
rect 0 363 336 370
<< psubdiffcont >>
rect 16 -8 32 8
rect 64 -8 80 8
rect 112 -8 128 8
rect 160 -8 176 8
rect 208 -8 224 8
rect 256 -8 272 8
rect 304 -8 320 8
<< nsubdiffcont >>
rect 16 370 32 386
rect 64 370 80 386
rect 112 370 128 386
rect 160 370 176 386
rect 208 370 224 386
rect 256 370 272 386
rect 304 370 320 386
<< poly >>
rect 70 306 83 324
rect 109 306 122 324
rect 166 306 179 324
rect 251 318 264 336
rect 70 190 83 206
rect 49 181 83 190
rect 49 165 58 181
rect 74 165 83 181
rect 49 157 83 165
rect 109 190 122 206
rect 166 190 179 206
rect 109 181 142 190
rect 109 165 117 181
rect 133 165 142 181
rect 109 157 142 165
rect 166 181 219 190
rect 251 183 264 206
rect 166 165 182 181
rect 198 165 219 181
rect 166 157 219 165
rect 70 114 83 157
rect 121 114 134 157
rect 206 114 219 157
rect 239 176 270 183
rect 239 160 246 176
rect 262 160 270 176
rect 239 153 270 160
rect 257 133 270 153
rect 70 41 83 59
rect 121 41 134 59
rect 206 41 219 59
rect 257 41 270 59
<< polycont >>
rect 58 165 74 181
rect 117 165 133 181
rect 182 165 198 181
rect 246 160 262 176
<< metal1 >>
rect 0 386 336 400
rect 0 370 16 386
rect 32 370 64 386
rect 80 370 112 386
rect 128 370 160 386
rect 176 370 208 386
rect 224 370 256 386
rect 272 370 304 386
rect 320 370 336 386
rect 0 356 336 370
rect 185 299 245 356
rect 38 298 64 299
rect 38 282 43 298
rect 59 282 64 298
rect 38 241 64 282
rect 185 283 190 299
rect 206 283 224 299
rect 240 283 245 299
rect 185 265 245 283
rect 185 249 190 265
rect 206 249 224 265
rect 240 249 245 265
rect 185 247 245 249
rect 270 310 305 320
rect 270 294 275 310
rect 291 294 305 310
rect 270 270 305 294
rect 270 254 275 270
rect 291 254 305 270
rect 38 225 43 241
rect 59 229 64 241
rect 270 230 305 254
rect 59 225 251 229
rect 38 212 251 225
rect 29 181 83 193
rect 29 165 58 181
rect 74 165 83 181
rect 29 150 83 165
rect 109 181 156 193
rect 109 165 117 181
rect 133 165 156 181
rect 109 150 156 165
rect 174 181 207 193
rect 174 165 182 181
rect 198 165 207 181
rect 174 150 207 165
rect 234 185 251 212
rect 270 214 275 230
rect 291 214 305 230
rect 270 204 305 214
rect 234 176 271 185
rect 234 160 246 176
rect 262 160 271 176
rect 234 152 271 160
rect 234 132 251 152
rect 38 111 251 132
rect 289 130 305 204
rect 276 125 305 130
rect 38 94 64 111
rect 38 78 43 94
rect 59 78 64 94
rect 144 92 196 111
rect 38 76 64 78
rect 89 88 115 89
rect 89 72 94 88
rect 110 72 115 88
rect 89 22 115 72
rect 144 76 145 92
rect 161 76 179 92
rect 195 76 196 92
rect 276 109 281 125
rect 297 109 305 125
rect 144 67 196 76
rect 225 88 251 89
rect 225 72 230 88
rect 246 72 251 88
rect 225 22 251 72
rect 276 82 305 109
rect 276 66 281 82
rect 297 66 305 82
rect 276 60 305 66
rect 0 8 336 22
rect 0 -8 16 8
rect 32 -8 64 8
rect 80 -8 112 8
rect 128 -8 160 8
rect 176 -8 208 8
rect 224 -8 256 8
rect 272 -8 304 8
rect 320 -8 336 8
rect 0 -22 336 -8
<< labels >>
flabel metal1 s 0 356 336 400 0 FreeSans 200 0 0 0 VDD
port 2 nsew
flabel metal1 s 0 -22 336 22 0 FreeSans 200 0 0 0 VSS
port 3 nsew
flabel metal1 s 29 150 83 193 0 FreeSans 200 0 0 0 C
port 4 nsew
flabel metal1 s 109 150 156 193 0 FreeSans 200 0 0 0 B
port 5 nsew
flabel metal1 s 174 150 207 193 0 FreeSans 200 0 0 0 A
port 6 nsew
flabel metal1 s 270 204 305 320 0 FreeSans 200 0 0 0 X
port 7 nsew
<< properties >>
string FIXED_BBOX 0 0 336 378
string GDS_END 128346
string GDS_FILE ../gds/controller.gds
string GDS_START 122822
<< end >>
