magic
tech ihp-sg13g2
magscale 1 2
timestamp 1747056038
<< nwell >>
rect -48 350 624 834
<< pwell >>
rect 6 56 570 270
rect -26 -56 602 56
<< nmos >>
rect 101 96 127 244
rect 202 96 228 244
rect 372 96 398 244
rect 450 96 476 244
<< pmos >>
rect 101 436 127 660
rect 224 436 250 660
rect 326 436 352 660
rect 450 436 476 660
<< ndiff >>
rect 32 230 101 244
rect 32 198 46 230
rect 78 198 101 230
rect 32 142 101 198
rect 32 110 46 142
rect 78 110 101 142
rect 32 96 101 110
rect 127 96 202 244
rect 228 220 372 244
rect 228 188 250 220
rect 282 188 318 220
rect 350 188 372 220
rect 228 96 372 188
rect 398 96 450 244
rect 476 230 544 244
rect 476 198 498 230
rect 530 198 544 230
rect 476 142 544 198
rect 476 110 498 142
rect 530 110 544 142
rect 476 96 544 110
<< pdiff >>
rect 33 646 101 660
rect 33 614 47 646
rect 79 614 101 646
rect 33 567 101 614
rect 33 535 47 567
rect 79 535 101 567
rect 33 482 101 535
rect 33 450 47 482
rect 79 450 101 482
rect 33 436 101 450
rect 127 646 224 660
rect 127 614 170 646
rect 202 614 224 646
rect 127 567 224 614
rect 127 535 170 567
rect 202 535 224 567
rect 127 482 224 535
rect 127 450 170 482
rect 202 450 224 482
rect 127 436 224 450
rect 250 570 326 660
rect 250 538 272 570
rect 304 538 326 570
rect 250 482 326 538
rect 250 450 272 482
rect 304 450 326 482
rect 250 436 326 450
rect 352 646 450 660
rect 352 614 374 646
rect 406 614 450 646
rect 352 567 450 614
rect 352 535 374 567
rect 406 535 450 567
rect 352 436 450 535
rect 476 646 544 660
rect 476 614 498 646
rect 530 614 544 646
rect 476 567 544 614
rect 476 535 498 567
rect 530 535 544 567
rect 476 482 544 535
rect 476 450 498 482
rect 530 450 544 482
rect 476 436 544 450
<< ndiffc >>
rect 46 198 78 230
rect 46 110 78 142
rect 250 188 282 220
rect 318 188 350 220
rect 498 198 530 230
rect 498 110 530 142
<< pdiffc >>
rect 47 614 79 646
rect 47 535 79 567
rect 47 450 79 482
rect 170 614 202 646
rect 170 535 202 567
rect 170 450 202 482
rect 272 538 304 570
rect 272 450 304 482
rect 374 614 406 646
rect 374 535 406 567
rect 498 614 530 646
rect 498 535 530 567
rect 498 450 530 482
<< psubdiff >>
rect 0 16 576 30
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 576 16
rect 0 -30 576 -16
<< nsubdiff >>
rect 0 772 576 786
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 576 772
rect 0 726 576 740
<< psubdiffcont >>
rect 32 -16 64 16
rect 128 -16 160 16
rect 224 -16 256 16
rect 320 -16 352 16
rect 416 -16 448 16
rect 512 -16 544 16
<< nsubdiffcont >>
rect 32 740 64 772
rect 128 740 160 772
rect 224 740 256 772
rect 320 740 352 772
rect 416 740 448 772
rect 512 740 544 772
<< poly >>
rect 101 660 127 696
rect 224 660 250 696
rect 326 660 352 696
rect 450 660 476 696
rect 101 422 127 436
rect 34 408 127 422
rect 224 418 250 436
rect 34 376 48 408
rect 80 396 127 408
rect 190 404 250 418
rect 80 376 95 396
rect 34 362 95 376
rect 190 372 204 404
rect 236 372 250 404
rect 326 414 352 436
rect 450 414 476 436
rect 326 400 414 414
rect 326 380 368 400
rect 190 350 250 372
rect 140 326 250 350
rect 101 322 250 326
rect 286 368 368 380
rect 400 368 414 400
rect 286 354 414 368
rect 450 400 544 414
rect 450 368 498 400
rect 530 368 544 400
rect 450 354 544 368
rect 101 298 166 322
rect 101 244 127 298
rect 286 286 312 354
rect 202 258 312 286
rect 354 304 414 318
rect 354 272 368 304
rect 400 272 414 304
rect 354 258 414 272
rect 202 244 228 258
rect 372 244 398 258
rect 450 244 476 354
rect 101 60 127 96
rect 202 60 228 96
rect 372 60 398 96
rect 450 60 476 96
<< polycont >>
rect 48 376 80 408
rect 204 372 236 404
rect 368 368 400 400
rect 498 368 530 400
rect 368 272 400 304
<< metal1 >>
rect 0 772 576 800
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 512 772
rect 544 740 576 772
rect 0 712 576 740
rect 36 646 90 712
rect 36 614 47 646
rect 79 614 90 646
rect 36 567 90 614
rect 36 535 47 567
rect 79 535 90 567
rect 36 482 90 535
rect 36 450 47 482
rect 79 450 90 482
rect 160 646 416 666
rect 160 614 170 646
rect 202 617 374 646
rect 202 614 212 617
rect 160 567 212 614
rect 364 614 374 617
rect 406 614 416 646
rect 160 535 170 567
rect 202 535 212 567
rect 160 482 212 535
rect 160 450 170 482
rect 202 450 212 482
rect 262 570 320 580
rect 262 538 272 570
rect 304 538 320 570
rect 262 482 320 538
rect 364 567 416 614
rect 364 535 374 567
rect 406 535 416 567
rect 364 524 416 535
rect 488 646 540 712
rect 488 614 498 646
rect 530 614 540 646
rect 488 567 540 614
rect 488 535 498 567
rect 530 535 540 567
rect 262 450 272 482
rect 304 450 320 482
rect 34 408 94 414
rect 34 376 48 408
rect 80 376 94 408
rect 34 298 94 376
rect 192 404 248 414
rect 192 372 204 404
rect 236 372 248 404
rect 34 266 156 298
rect 192 266 248 372
rect 36 198 46 230
rect 78 198 88 230
rect 36 142 88 198
rect 36 110 46 142
rect 78 110 88 142
rect 124 142 156 266
rect 284 230 320 450
rect 356 400 416 488
rect 488 482 540 535
rect 488 450 498 482
rect 530 450 540 482
rect 356 368 368 400
rect 400 368 416 400
rect 356 340 416 368
rect 484 400 544 414
rect 484 368 498 400
rect 530 368 544 400
rect 358 272 368 304
rect 400 272 418 304
rect 250 220 350 230
rect 282 188 318 220
rect 250 178 350 188
rect 386 142 418 272
rect 484 266 544 368
rect 124 110 418 142
rect 488 198 498 230
rect 530 198 540 230
rect 488 142 540 198
rect 488 110 498 142
rect 530 110 540 142
rect 36 44 88 110
rect 488 44 540 110
rect 0 16 576 44
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 512 16
rect 544 -16 576 16
rect 0 -44 576 -16
<< labels >>
flabel metal1 s 284 178 320 580 0 FreeSans 400 0 0 0 Y
port 2 nsew
flabel metal1 s 484 266 544 414 0 FreeSans 400 0 0 0 A2
port 3 nsew
flabel metal1 s 0 712 576 800 0 FreeSans 400 0 0 0 VDD
port 4 nsew
flabel metal1 s 192 266 248 414 0 FreeSans 400 0 0 0 B1
port 5 nsew
flabel metal1 s 0 -44 576 44 0 FreeSans 400 0 0 0 VSS
port 6 nsew
flabel metal1 s 34 266 94 414 0 FreeSans 400 0 0 0 A1
port 7 nsew
flabel metal1 s 356 340 416 488 0 FreeSans 400 0 0 0 B2
port 8 nsew
<< properties >>
string FIXED_BBOX 0 0 576 756
string GDS_END 148628
string GDS_FILE ../gds/controller.gds
string GDS_START 143522
<< end >>
