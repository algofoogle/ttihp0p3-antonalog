magic
tech ihp-sg13g2
magscale 1 2
timestamp 1747056038
<< nwell >>
rect -48 350 528 834
<< pwell >>
rect 1 56 447 292
rect -26 -56 506 56
<< nmos >>
rect 95 156 121 266
rect 265 118 291 266
rect 327 118 353 266
<< pmos >>
rect 95 412 121 580
rect 203 412 229 636
rect 305 412 331 636
<< ndiff >>
rect 27 226 95 266
rect 27 194 41 226
rect 73 194 95 226
rect 27 156 95 194
rect 121 200 265 266
rect 121 168 143 200
rect 175 198 265 200
rect 175 168 211 198
rect 121 166 211 168
rect 243 166 265 198
rect 121 156 265 166
rect 135 118 265 156
rect 291 118 327 266
rect 353 252 421 266
rect 353 220 375 252
rect 407 220 421 252
rect 353 164 421 220
rect 353 132 375 164
rect 407 132 421 164
rect 353 118 421 132
<< pdiff >>
rect 135 618 203 636
rect 135 586 149 618
rect 181 586 203 618
rect 135 580 203 586
rect 27 566 95 580
rect 27 534 41 566
rect 73 534 95 566
rect 27 482 95 534
rect 27 450 41 482
rect 73 450 95 482
rect 27 412 95 450
rect 121 550 203 580
rect 121 518 149 550
rect 181 518 203 550
rect 121 412 203 518
rect 229 622 305 636
rect 229 590 251 622
rect 283 590 305 622
rect 229 550 305 590
rect 229 518 251 550
rect 283 518 305 550
rect 229 412 305 518
rect 331 622 399 636
rect 331 590 353 622
rect 385 590 399 622
rect 331 412 399 590
<< ndiffc >>
rect 41 194 73 226
rect 143 168 175 200
rect 211 166 243 198
rect 375 220 407 252
rect 375 132 407 164
<< pdiffc >>
rect 149 586 181 618
rect 41 534 73 566
rect 41 450 73 482
rect 149 518 181 550
rect 251 590 283 622
rect 251 518 283 550
rect 353 590 385 622
<< psubdiff >>
rect 0 16 480 30
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 480 16
rect 0 -30 480 -16
<< nsubdiff >>
rect 0 772 480 786
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 480 772
rect 0 726 480 740
<< psubdiffcont >>
rect 32 -16 64 16
rect 128 -16 160 16
rect 224 -16 256 16
rect 320 -16 352 16
rect 416 -16 448 16
<< nsubdiffcont >>
rect 32 740 64 772
rect 128 740 160 772
rect 224 740 256 772
rect 320 740 352 772
rect 416 740 448 772
<< poly >>
rect 203 636 229 672
rect 305 636 331 672
rect 95 580 121 616
rect 95 370 121 412
rect 21 352 155 370
rect 21 320 37 352
rect 69 320 105 352
rect 137 320 155 352
rect 21 304 155 320
rect 203 366 229 412
rect 305 385 331 412
rect 203 352 263 366
rect 305 354 387 385
rect 203 320 217 352
rect 249 320 263 352
rect 203 309 263 320
rect 327 352 387 354
rect 327 320 341 352
rect 373 320 387 352
rect 95 266 121 304
rect 203 280 291 309
rect 265 266 291 280
rect 327 304 387 320
rect 327 266 353 304
rect 95 120 121 156
rect 265 82 291 118
rect 327 82 353 118
<< polycont >>
rect 37 320 69 352
rect 105 320 137 352
rect 217 320 249 352
rect 341 320 373 352
<< metal1 >>
rect 0 772 480 800
rect 0 740 32 772
rect 64 740 128 772
rect 160 740 224 772
rect 256 740 320 772
rect 352 740 416 772
rect 448 740 480 772
rect 0 712 480 740
rect 146 618 183 712
rect 146 586 149 618
rect 181 586 183 618
rect 38 566 76 580
rect 38 534 41 566
rect 73 534 76 566
rect 38 482 76 534
rect 146 550 183 586
rect 146 518 149 550
rect 181 518 183 550
rect 146 508 183 518
rect 241 622 293 625
rect 241 590 251 622
rect 283 590 293 622
rect 241 550 293 590
rect 343 622 395 712
rect 343 590 353 622
rect 385 590 395 622
rect 343 587 395 590
rect 241 518 251 550
rect 283 536 293 550
rect 283 518 451 536
rect 241 502 451 518
rect 38 450 41 482
rect 73 466 76 482
rect 73 450 379 466
rect 38 434 379 450
rect 21 352 155 378
rect 21 320 37 352
rect 69 320 105 352
rect 137 320 155 352
rect 21 306 155 320
rect 203 352 267 389
rect 203 320 217 352
rect 249 320 267 352
rect 325 352 379 434
rect 325 340 341 352
rect 203 310 267 320
rect 303 320 341 340
rect 373 320 379 352
rect 303 304 379 320
rect 303 270 337 304
rect 31 238 337 270
rect 417 263 451 502
rect 373 252 451 263
rect 31 226 83 238
rect 31 194 41 226
rect 73 194 83 226
rect 373 220 375 252
rect 407 220 451 252
rect 31 184 83 194
rect 133 200 253 201
rect 133 168 143 200
rect 175 198 253 200
rect 175 168 211 198
rect 133 166 211 168
rect 243 166 253 198
rect 133 44 253 166
rect 373 164 451 220
rect 373 132 375 164
rect 407 132 451 164
rect 373 122 451 132
rect 0 16 480 44
rect 0 -16 32 16
rect 64 -16 128 16
rect 160 -16 224 16
rect 256 -16 320 16
rect 352 -16 416 16
rect 448 -16 480 16
rect 0 -44 480 -16
<< labels >>
flabel metal1 s 0 -44 480 44 0 FreeSans 400 0 0 0 VSS
port 2 nsew
flabel metal1 s 21 306 155 378 0 FreeSans 400 0 0 0 A_N
port 3 nsew
flabel metal1 s 373 122 451 263 0 FreeSans 400 0 0 0 Y
port 4 nsew
flabel metal1 s 203 310 267 389 0 FreeSans 400 0 0 0 B
port 5 nsew
flabel metal1 s 0 712 480 800 0 FreeSans 400 0 0 0 VDD
port 6 nsew
<< properties >>
string FIXED_BBOX 0 0 480 756
string GDS_END 116984
string GDS_FILE ../gds/controller.gds
string GDS_START 112496
<< end >>
