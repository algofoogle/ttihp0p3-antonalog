magic
tech ihp-sg13g2
magscale 1 2
timestamp 1747574207
<< metal1 >>
rect 2026 30244 3192 30322
rect 2026 30118 2268 30244
rect 2936 30118 3192 30244
rect 2026 29124 2148 30118
rect 3040 30040 3192 30118
rect 4340 30118 4950 30256
rect 4340 30040 4496 30118
rect 2420 29730 2768 30014
rect 3040 29910 4496 30040
rect 3040 29750 3276 29910
rect 3484 29834 3630 29910
rect 3944 29882 4496 29910
rect 4768 30040 4950 30118
rect 4768 29916 7132 30040
rect 4768 29882 6184 29916
rect 3944 29750 4314 29882
rect 2420 29124 2768 29500
rect 3040 29124 3262 29750
rect 3652 29596 3846 29680
rect 3534 29124 3846 29596
rect 4118 29652 4314 29750
rect 4982 29876 6184 29882
rect 4982 29756 5250 29876
rect 5918 29756 6184 29876
rect 6392 29840 6538 29916
rect 6852 29756 7132 29916
rect 4982 29652 5174 29756
rect 4118 29124 4496 29652
rect 4768 29262 5174 29652
rect 5446 29354 5724 29646
rect 5996 29262 6170 29756
rect 6560 29602 6754 29686
rect 4768 29124 5258 29262
rect 5926 29130 6170 29262
rect 6442 29130 6754 29602
rect 7026 29130 7132 29756
rect 5926 29124 7132 29130
rect 2026 29012 7132 29124
<< via1 >>
rect 4336 25816 4524 26118
rect 4336 25060 4442 25220
rect 2990 24304 3096 24464
rect 4336 23548 4442 23708
rect 2990 22792 3096 22952
rect 4336 22036 4442 22196
rect 2990 21280 3096 21440
rect 4336 20524 4442 20684
rect 2990 20020 3096 20432
rect 2990 19768 3096 19928
rect 4336 18256 4524 18558
rect 4336 17500 4442 17660
rect 2990 16744 3096 16904
rect 4336 15988 4442 16148
rect 2990 15232 3096 15392
rect 4336 14476 4442 14636
rect 2990 13720 3096 13880
rect 4336 12964 4442 13124
rect 2990 12460 3096 12872
rect 2990 12208 3096 12368
rect 4336 10696 4524 10998
rect 4336 9940 4442 10100
rect 2990 9184 3096 9344
rect 4336 8428 4442 8588
rect 2990 7672 3096 7832
rect 4336 6916 4442 7076
rect 2990 6160 3096 6320
rect 4336 5404 4442 5564
rect 2990 4900 3096 5312
rect 2990 4648 3096 4808
<< metal2 >>
rect 2026 30244 3192 30322
rect 2026 30118 2268 30244
rect 2936 30118 3192 30244
rect 2026 29124 2148 30118
rect 3040 30040 3192 30118
rect 4340 30118 4950 30256
rect 4340 30040 4496 30118
rect 2420 29730 2768 30014
rect 3040 29910 4496 30040
rect 3040 29750 3276 29910
rect 3484 29834 3630 29910
rect 3944 29882 4496 29910
rect 4768 30040 4950 30118
rect 4768 29916 7132 30040
rect 4768 29882 6184 29916
rect 3944 29750 4314 29882
rect 2420 29124 2768 29500
rect 3040 29124 3262 29750
rect 3652 29596 3846 29680
rect 3534 29124 3846 29596
rect 4118 29652 4314 29750
rect 4982 29876 6184 29882
rect 4982 29756 5250 29876
rect 5918 29756 6184 29876
rect 6392 29840 6538 29916
rect 6852 29756 7132 29916
rect 4982 29652 5174 29756
rect 4118 29124 4496 29652
rect 4768 29262 5174 29652
rect 5446 29354 5724 29646
rect 5996 29262 6170 29756
rect 6560 29602 6754 29686
rect 4768 29124 5258 29262
rect 5926 29130 6170 29262
rect 6442 29130 6754 29602
rect 7026 29130 7132 29756
rect 5926 29124 7132 29130
rect 2026 29012 7132 29124
rect 4316 26518 4544 26538
rect 4316 26216 4336 26518
rect 4524 26216 4544 26518
rect 4316 26118 4544 26216
rect 4316 25816 4336 26118
rect 4524 25816 4544 26118
rect 4316 25796 4544 25816
rect 4316 25220 4462 25240
rect 4316 25060 4336 25220
rect 4442 25140 4752 25220
rect 4442 25060 4462 25140
rect 4316 25040 4462 25060
rect 2970 24464 3116 24484
rect 2970 24304 2990 24464
rect 3096 24384 4752 24464
rect 3096 24304 3116 24384
rect 2970 24284 3116 24304
rect 4316 23708 4462 23728
rect 4316 23548 4336 23708
rect 4442 23628 4752 23708
rect 4442 23548 4462 23628
rect 4316 23528 4462 23548
rect 7176 23460 7458 23540
rect 7176 23040 7458 23120
rect 2970 22952 3116 22972
rect 2970 22792 2990 22952
rect 3096 22872 4752 22952
rect 3096 22792 3116 22872
rect 2970 22772 3116 22792
rect 7176 22620 7458 22700
rect 4316 22196 4462 22216
rect 7176 22200 7458 22280
rect 4316 22036 4336 22196
rect 4442 22116 4752 22196
rect 4442 22036 4462 22116
rect 4316 22016 4462 22036
rect 7176 21780 7458 21860
rect 2970 21440 3116 21460
rect 2970 21280 2990 21440
rect 3096 21360 4752 21440
rect 7176 21360 7458 21440
rect 3096 21280 3116 21360
rect 2970 21260 3116 21280
rect 7176 20940 7458 21020
rect 4316 20684 4462 20704
rect 4316 20524 4336 20684
rect 4442 20604 4752 20684
rect 4442 20524 4462 20604
rect 4316 20504 4462 20524
rect 7176 20520 7458 20600
rect 2570 20432 3116 20452
rect 2570 20020 2590 20432
rect 2776 20020 2990 20432
rect 3096 20020 3116 20432
rect 2570 20000 3116 20020
rect 2970 19928 3116 19948
rect 2970 19768 2990 19928
rect 3096 19848 4752 19928
rect 3096 19768 3116 19848
rect 2970 19748 3116 19768
rect 4316 18958 4544 18978
rect 4316 18656 4336 18958
rect 4524 18656 4544 18958
rect 4316 18558 4544 18656
rect 4316 18256 4336 18558
rect 4524 18256 4544 18558
rect 4316 18236 4544 18256
rect 4316 17660 4462 17680
rect 4316 17500 4336 17660
rect 4442 17580 4752 17660
rect 4442 17500 4462 17580
rect 4316 17480 4462 17500
rect 2970 16904 3116 16924
rect 2970 16744 2990 16904
rect 3096 16824 4752 16904
rect 3096 16744 3116 16824
rect 2970 16724 3116 16744
rect 7176 16740 7458 16820
rect 7176 16320 7458 16400
rect 4316 16148 4462 16168
rect 4316 15988 4336 16148
rect 4442 16068 4752 16148
rect 4442 15988 4462 16068
rect 4316 15968 4462 15988
rect 7176 15900 7458 15980
rect 7176 15480 7458 15560
rect 2970 15392 3116 15412
rect 2970 15232 2990 15392
rect 3096 15312 4752 15392
rect 3096 15232 3116 15312
rect 2970 15212 3116 15232
rect 7176 15060 7458 15140
rect 4316 14636 4462 14656
rect 7176 14640 7458 14720
rect 4316 14476 4336 14636
rect 4442 14556 4752 14636
rect 4442 14476 4462 14556
rect 4316 14456 4462 14476
rect 7176 14220 7458 14300
rect 2970 13880 3116 13900
rect 2970 13720 2990 13880
rect 3096 13800 4752 13880
rect 7176 13800 7458 13880
rect 3096 13720 3116 13800
rect 2970 13700 3116 13720
rect 4316 13124 4462 13144
rect 4316 12964 4336 13124
rect 4442 13044 4752 13124
rect 4442 12964 4462 13044
rect 4316 12944 4462 12964
rect 2570 12872 3116 12892
rect 2570 12460 2590 12872
rect 2776 12460 2990 12872
rect 3096 12460 3116 12872
rect 2570 12440 3116 12460
rect 2970 12368 3116 12388
rect 2970 12208 2990 12368
rect 3096 12288 4752 12368
rect 3096 12208 3116 12288
rect 2970 12188 3116 12208
rect 4316 11398 4544 11418
rect 4316 11096 4336 11398
rect 4524 11096 4544 11398
rect 4316 10998 4544 11096
rect 4316 10696 4336 10998
rect 4524 10696 4544 10998
rect 4316 10676 4544 10696
rect 4316 10100 4462 10120
rect 4316 9940 4336 10100
rect 4442 10020 4752 10100
rect 7176 10020 7458 10100
rect 4442 9940 4462 10020
rect 4316 9920 4462 9940
rect 7176 9600 7458 9680
rect 2970 9344 3116 9364
rect 2970 9184 2990 9344
rect 3096 9264 4752 9344
rect 3096 9184 3116 9264
rect 2970 9164 3116 9184
rect 7176 9180 7458 9260
rect 7176 8760 7458 8840
rect 4316 8588 4462 8608
rect 4316 8428 4336 8588
rect 4442 8508 4752 8588
rect 4442 8428 4462 8508
rect 4316 8408 4462 8428
rect 7176 8340 7458 8420
rect 7176 7920 7458 8000
rect 2970 7832 3116 7852
rect 2970 7672 2990 7832
rect 3096 7752 4752 7832
rect 3096 7672 3116 7752
rect 2970 7652 3116 7672
rect 7176 7500 7458 7580
rect 4316 7076 4462 7096
rect 7176 7080 7458 7160
rect 4316 6916 4336 7076
rect 4442 6996 4752 7076
rect 4442 6916 4462 6996
rect 4316 6896 4462 6916
rect 2970 6320 3116 6340
rect 2970 6160 2990 6320
rect 3096 6240 4752 6320
rect 3096 6160 3116 6240
rect 2970 6140 3116 6160
rect 4316 5564 4462 5584
rect 4316 5404 4336 5564
rect 4442 5484 4752 5564
rect 4442 5404 4462 5484
rect 4316 5384 4462 5404
rect 2570 5312 3116 5332
rect 2570 4900 2590 5312
rect 2776 4900 2990 5312
rect 3096 4900 3116 5312
rect 2570 4880 3116 4900
rect 2970 4808 3116 4828
rect 2970 4648 2990 4808
rect 3096 4728 4752 4808
rect 3096 4648 3116 4728
rect 2970 4628 3116 4648
<< via2 >>
rect 4336 26216 4524 26518
rect 2590 20020 2776 20432
rect 4336 18656 4524 18958
rect 2590 12460 2776 12872
rect 4336 11096 4524 11398
rect 2590 4900 2776 5312
<< metal3 >>
rect 10502 30465 10621 30479
rect 10502 30373 10515 30465
rect 10607 30373 10621 30465
rect 2026 30244 3192 30322
rect 2026 30118 2268 30244
rect 2936 30118 3192 30244
rect 2026 29124 2148 30118
rect 3040 30040 3192 30118
rect 4340 30118 4950 30256
rect 4340 30040 4496 30118
rect 2420 29730 2768 30014
rect 3040 29910 4496 30040
rect 3040 29750 3276 29910
rect 3484 29834 3630 29910
rect 3944 29882 4496 29910
rect 4768 30040 4950 30118
rect 4768 29916 7132 30040
rect 10502 30019 10621 30373
rect 11270 30465 11389 30479
rect 11270 30373 11283 30465
rect 11375 30373 11389 30465
rect 11270 30019 11389 30373
rect 12038 30465 12157 30479
rect 12038 30373 12051 30465
rect 12143 30373 12157 30465
rect 12038 30019 12157 30373
rect 12806 30465 12925 30479
rect 12806 30373 12819 30465
rect 12911 30373 12925 30465
rect 12806 30019 12925 30373
rect 13574 30465 13693 30479
rect 13574 30373 13587 30465
rect 13679 30373 13693 30465
rect 13574 30019 13693 30373
rect 14342 30465 14461 30479
rect 14342 30373 14355 30465
rect 14447 30373 14461 30465
rect 14342 30019 14461 30373
rect 15110 30465 15229 30479
rect 15110 30373 15123 30465
rect 15215 30373 15229 30465
rect 15110 30019 15229 30373
rect 15878 30465 15997 30479
rect 15878 30373 15891 30465
rect 15983 30373 15997 30465
rect 15878 30019 15997 30373
rect 16646 30465 16765 30479
rect 16646 30373 16659 30465
rect 16751 30373 16765 30465
rect 16646 30019 16765 30373
rect 17414 30465 17533 30479
rect 17414 30373 17427 30465
rect 17519 30373 17533 30465
rect 17414 30019 17533 30373
rect 18182 30465 18301 30479
rect 18182 30373 18195 30465
rect 18287 30373 18301 30465
rect 18182 30019 18301 30373
rect 18950 30465 19069 30479
rect 18950 30373 18963 30465
rect 19055 30373 19069 30465
rect 18950 30019 19069 30373
rect 19718 30465 19837 30479
rect 19718 30373 19731 30465
rect 19823 30373 19837 30465
rect 19718 30019 19837 30373
rect 20486 30465 20605 30479
rect 20486 30373 20499 30465
rect 20591 30373 20605 30465
rect 20486 30019 20605 30373
rect 21254 30465 21373 30479
rect 21254 30373 21267 30465
rect 21359 30373 21373 30465
rect 21254 30019 21373 30373
rect 22022 30465 22141 30479
rect 22022 30373 22035 30465
rect 22127 30373 22141 30465
rect 22022 30019 22141 30373
rect 22790 30465 22909 30479
rect 22790 30373 22803 30465
rect 22895 30373 22909 30465
rect 22790 30019 22909 30373
rect 23558 30465 23677 30479
rect 23558 30373 23571 30465
rect 23663 30373 23677 30465
rect 23558 30019 23677 30373
rect 30471 30362 30480 30458
rect 30576 30362 30585 30458
rect 31239 30362 31248 30458
rect 31344 30362 31353 30458
rect 32007 30362 32016 30458
rect 32112 30362 32121 30458
rect 32775 30362 32784 30458
rect 32880 30362 32889 30458
rect 33543 30362 33552 30458
rect 33648 30362 33657 30458
rect 34311 30362 34320 30458
rect 34416 30362 34425 30458
rect 35079 30362 35088 30458
rect 35184 30362 35193 30458
rect 35847 30362 35856 30458
rect 35952 30362 35961 30458
rect 36615 30362 36624 30458
rect 36720 30362 36729 30458
rect 37383 30362 37392 30458
rect 37488 30362 37497 30458
rect 38151 30362 38160 30458
rect 38256 30362 38265 30458
rect 30480 30010 30576 30362
rect 31248 30010 31344 30362
rect 32016 30010 32112 30362
rect 32784 30010 32880 30362
rect 33552 30010 33648 30362
rect 34320 30010 34416 30362
rect 35088 30010 35184 30362
rect 35856 30010 35952 30362
rect 36624 30010 36720 30362
rect 37392 30010 37488 30362
rect 38160 30010 38256 30362
rect 4768 29882 6184 29916
rect 3944 29750 4314 29882
rect 2420 29124 2768 29500
rect 3040 29124 3262 29750
rect 3652 29596 3846 29680
rect 3534 29124 3846 29596
rect 4118 29652 4314 29750
rect 4982 29876 6184 29882
rect 4982 29756 5250 29876
rect 5918 29756 6184 29876
rect 6392 29840 6538 29916
rect 6852 29756 7132 29916
rect 4982 29652 5174 29756
rect 4118 29124 4496 29652
rect 4768 29262 5174 29652
rect 5446 29354 5724 29646
rect 5996 29262 6170 29756
rect 6560 29602 6754 29686
rect 4768 29124 5258 29262
rect 5926 29130 6170 29262
rect 6442 29130 6754 29602
rect 7026 29130 7132 29756
rect 5926 29124 7132 29130
rect 2026 29012 7132 29124
rect 4316 26518 4544 26538
rect 4316 26216 4336 26518
rect 4524 26216 4544 26518
rect 4316 26196 4544 26216
rect 425 21976 605 21985
rect 605 21796 2776 21976
rect 425 21787 605 21796
rect 2596 20452 2776 21796
rect 2570 20432 2796 20452
rect 2570 20020 2590 20432
rect 2776 20020 2796 20432
rect 2570 20000 2796 20020
rect 4316 18958 4544 18978
rect 418 18628 427 18808
rect 607 18628 2778 18808
rect 4316 18656 4336 18958
rect 4524 18656 4544 18958
rect 4316 18636 4544 18656
rect 2598 12892 2778 18628
rect 2570 12872 2796 12892
rect 2570 12460 2590 12872
rect 2776 12460 2796 12872
rect 2570 12440 2796 12460
rect 4316 11398 4544 11418
rect 4316 11096 4336 11398
rect 4524 11096 4544 11398
rect 4316 11076 4544 11096
rect 2570 5312 2796 5332
rect 401 5196 581 5205
rect 2570 5196 2590 5312
rect 581 5016 2590 5196
rect 401 5007 581 5016
rect 2570 4900 2590 5016
rect 2776 4900 2796 5312
rect 2570 4880 2796 4900
<< via3 >>
rect 10515 30373 10607 30465
rect 11283 30373 11375 30465
rect 12051 30373 12143 30465
rect 12819 30373 12911 30465
rect 13587 30373 13679 30465
rect 14355 30373 14447 30465
rect 15123 30373 15215 30465
rect 15891 30373 15983 30465
rect 16659 30373 16751 30465
rect 17427 30373 17519 30465
rect 18195 30373 18287 30465
rect 18963 30373 19055 30465
rect 19731 30373 19823 30465
rect 20499 30373 20591 30465
rect 21267 30373 21359 30465
rect 22035 30373 22127 30465
rect 22803 30373 22895 30465
rect 23571 30373 23663 30465
rect 30480 30362 30576 30458
rect 31248 30362 31344 30458
rect 32016 30362 32112 30458
rect 32784 30362 32880 30458
rect 33552 30362 33648 30458
rect 34320 30362 34416 30458
rect 35088 30362 35184 30458
rect 35856 30362 35952 30458
rect 36624 30362 36720 30458
rect 37392 30362 37488 30458
rect 38160 30362 38256 30458
rect 4336 26216 4524 26518
rect 425 21796 605 21976
rect 427 18628 607 18808
rect 4336 18656 4524 18958
rect 4336 11096 4524 11398
rect 401 5016 581 5196
<< metal4 >>
rect 10515 30465 10607 30474
rect 11283 30465 11375 30474
rect 12051 30465 12143 30474
rect 12819 30465 12911 30474
rect 13587 30465 13679 30474
rect 14355 30465 14447 30474
rect 15123 30465 15215 30474
rect 15891 30465 15983 30474
rect 16659 30465 16751 30474
rect 17427 30465 17519 30474
rect 18195 30465 18287 30474
rect 18963 30465 19055 30474
rect 19731 30465 19823 30474
rect 20499 30465 20591 30474
rect 21267 30465 21359 30474
rect 22035 30465 22127 30474
rect 22803 30465 22895 30474
rect 23571 30465 23663 30474
rect 10508 30375 10515 30462
rect 10607 30375 10613 30462
rect 11276 30375 11283 30462
rect 11375 30375 11381 30462
rect 12044 30375 12051 30462
rect 12143 30375 12149 30462
rect 12812 30375 12819 30462
rect 12911 30375 12917 30462
rect 13580 30375 13587 30462
rect 13679 30375 13685 30462
rect 14348 30375 14355 30462
rect 14447 30375 14453 30462
rect 15116 30375 15123 30462
rect 15215 30375 15221 30462
rect 15884 30375 15891 30462
rect 15983 30375 15989 30462
rect 16652 30375 16659 30462
rect 16751 30375 16757 30462
rect 17420 30375 17427 30462
rect 17519 30375 17525 30462
rect 18188 30375 18195 30462
rect 18287 30375 18293 30462
rect 18956 30375 18963 30462
rect 19055 30375 19061 30462
rect 19724 30375 19731 30462
rect 19823 30375 19829 30462
rect 20492 30375 20499 30462
rect 20591 30375 20597 30462
rect 21260 30375 21267 30462
rect 21359 30375 21365 30462
rect 22028 30375 22035 30462
rect 22127 30375 22133 30462
rect 22796 30375 22803 30462
rect 22895 30375 22901 30462
rect 23564 30375 23571 30462
rect 23663 30375 23669 30462
rect 30480 30458 30576 30467
rect 31248 30458 31344 30467
rect 32016 30458 32112 30467
rect 32784 30458 32880 30467
rect 33552 30458 33648 30467
rect 34320 30458 34416 30467
rect 35088 30458 35184 30467
rect 35856 30458 35952 30467
rect 36624 30458 36720 30467
rect 37392 30458 37488 30467
rect 38160 30458 38256 30467
rect 10515 30364 10607 30373
rect 11283 30364 11375 30373
rect 12051 30364 12143 30373
rect 12819 30364 12911 30373
rect 13587 30364 13679 30373
rect 14355 30364 14447 30373
rect 15123 30364 15215 30373
rect 15891 30364 15983 30373
rect 16659 30364 16751 30373
rect 17427 30364 17519 30373
rect 18195 30364 18287 30373
rect 18963 30364 19055 30373
rect 19731 30364 19823 30373
rect 20499 30364 20591 30373
rect 21267 30364 21359 30373
rect 22035 30364 22127 30373
rect 22803 30364 22895 30373
rect 23571 30364 23663 30373
rect 30471 30362 30480 30458
rect 30576 30362 30585 30458
rect 31239 30362 31248 30458
rect 31344 30362 31353 30458
rect 32007 30362 32016 30458
rect 32112 30362 32121 30458
rect 32775 30362 32784 30458
rect 32880 30362 32889 30458
rect 33543 30362 33552 30458
rect 33648 30362 33657 30458
rect 34311 30362 34320 30458
rect 34416 30362 34425 30458
rect 35079 30362 35088 30458
rect 35184 30362 35193 30458
rect 35847 30362 35856 30458
rect 35952 30362 35961 30458
rect 36615 30362 36624 30458
rect 36720 30362 36729 30458
rect 37383 30362 37392 30458
rect 37488 30362 37497 30458
rect 38151 30362 38160 30458
rect 38256 30362 38265 30458
rect 30480 30353 30576 30362
rect 31248 30353 31344 30362
rect 32016 30353 32112 30362
rect 32784 30353 32880 30362
rect 33552 30353 33648 30362
rect 34320 30353 34416 30362
rect 35088 30353 35184 30362
rect 35856 30353 35952 30362
rect 36624 30353 36720 30362
rect 37392 30353 37488 30362
rect 38160 30353 38256 30362
rect 2026 30244 3192 30322
rect 2026 30118 2268 30244
rect 2936 30118 3192 30244
rect 2026 29124 2148 30118
rect 3040 30040 3192 30118
rect 4340 30118 4950 30256
rect 4340 30040 4496 30118
rect 2420 29730 2768 30014
rect 3040 29910 4496 30040
rect 3040 29750 3276 29910
rect 3484 29834 3630 29910
rect 3944 29882 4496 29910
rect 4768 30040 4950 30118
rect 4768 29916 7132 30040
rect 4768 29882 6184 29916
rect 3944 29750 4314 29882
rect 2420 29124 2768 29500
rect 3040 29124 3262 29750
rect 3652 29596 3846 29680
rect 3534 29124 3846 29596
rect 4118 29652 4314 29750
rect 4982 29876 6184 29882
rect 4982 29756 5250 29876
rect 5918 29756 6184 29876
rect 6392 29840 6538 29916
rect 6852 29756 7132 29916
rect 4982 29652 5174 29756
rect 4118 29124 4496 29652
rect 4768 29262 5174 29652
rect 5446 29354 5724 29646
rect 5996 29262 6170 29756
rect 6560 29602 6754 29686
rect 4768 29124 5258 29262
rect 5926 29130 6170 29262
rect 6442 29130 6754 29602
rect 7026 29130 7132 29756
rect 5926 29124 7132 29130
rect 2026 29012 7132 29124
rect 7314 29884 39350 29894
rect 7314 29817 38902 29884
rect 7314 29512 10528 29817
rect 10841 29512 18296 29817
rect 18609 29512 26055 29817
rect 26368 29512 33840 29817
rect 34153 29512 38902 29817
rect 7314 28856 7690 29512
rect 10528 29503 10841 29512
rect 18296 29503 18609 29512
rect 26055 29503 26368 29512
rect 33840 29503 34153 29512
rect 38644 29444 38902 29512
rect 39342 29444 39350 29884
rect 38644 29434 39350 29444
rect 3870 28480 7690 28856
rect 3870 28013 4246 28480
rect 3870 27708 3898 28013
rect 4203 27708 4246 28013
rect 3870 27680 4246 27708
rect 4316 26518 4544 26538
rect 4316 26216 4336 26518
rect 4524 26216 4544 26518
rect 4316 26196 4544 26216
rect 416 24596 425 24776
rect 605 24596 614 24776
rect 425 21976 605 24596
rect 416 21796 425 21976
rect 605 21796 614 21976
rect 427 21576 607 21585
rect 427 18808 607 21396
rect 4316 18958 4544 18978
rect 4316 18656 4336 18958
rect 4524 18656 4544 18958
rect 4316 18636 4544 18656
rect 427 18619 607 18628
rect 392 18196 401 18376
rect 581 18196 590 18376
rect 401 5196 581 18196
rect 4316 11398 4544 11418
rect 4316 11096 4336 11398
rect 4524 11096 4544 11398
rect 4316 11076 4544 11096
rect 392 5016 401 5196
rect 581 5016 590 5196
rect 3894 1628 35572 1706
rect 3894 1610 6140 1628
rect 3894 1100 3940 1610
rect 4550 1100 6140 1610
rect 6668 1584 35572 1628
rect 6668 1144 11718 1584
rect 12158 1144 19492 1584
rect 19932 1578 35572 1584
rect 19932 1144 27266 1578
rect 6668 1138 27266 1144
rect 27706 1570 35572 1578
rect 27706 1138 35040 1570
rect 6668 1130 35040 1138
rect 35480 1130 35572 1570
rect 6668 1100 35572 1130
rect 3894 1030 35572 1100
<< via4 >>
rect 10517 30375 10604 30462
rect 11285 30375 11372 30462
rect 12053 30375 12140 30462
rect 12821 30375 12908 30462
rect 13589 30375 13676 30462
rect 14357 30375 14444 30462
rect 15125 30375 15212 30462
rect 15893 30375 15980 30462
rect 16661 30375 16748 30462
rect 17429 30375 17516 30462
rect 18197 30375 18284 30462
rect 18965 30375 19052 30462
rect 19733 30375 19820 30462
rect 20501 30375 20588 30462
rect 21269 30375 21356 30462
rect 22037 30375 22124 30462
rect 22805 30375 22892 30462
rect 23573 30375 23660 30462
rect 30480 30362 30576 30458
rect 31248 30362 31344 30458
rect 32016 30362 32112 30458
rect 32784 30362 32880 30458
rect 33552 30362 33648 30458
rect 34320 30362 34416 30458
rect 35088 30362 35184 30458
rect 35856 30362 35952 30458
rect 36624 30362 36720 30458
rect 37392 30362 37488 30458
rect 38160 30362 38256 30458
rect 10528 29512 10841 29817
rect 18296 29512 18609 29817
rect 26055 29512 26368 29817
rect 33840 29512 34153 29817
rect 38902 29444 39342 29884
rect 3898 27708 4203 28013
rect 4336 26216 4524 26518
rect 425 24596 605 24776
rect 427 21396 607 21576
rect 4336 18656 4524 18958
rect 401 18196 581 18376
rect 4336 11096 4524 11398
rect 3940 1100 4550 1610
rect 6140 1100 6668 1628
rect 11718 1144 12158 1584
rect 19492 1144 19932 1584
rect 27266 1138 27706 1578
rect 35040 1130 35480 1570
<< metal5 >>
rect 958 30596 1732 30678
rect 791 30592 1732 30596
rect 5922 30592 5982 30996
rect 6690 30592 6750 30996
rect 7458 30592 7518 30996
rect 8226 30592 8286 30996
rect 8994 30592 9054 30996
rect 9762 30592 9822 30996
rect 791 30532 9822 30592
rect 791 30456 1732 30532
rect 10530 30522 10590 30996
rect 11298 30522 11358 30996
rect 12066 30522 12126 30996
rect 12834 30522 12894 30996
rect 13602 30522 13662 30996
rect 14370 30522 14430 30996
rect 15138 30522 15198 30996
rect 15906 30522 15966 30996
rect 16674 30522 16734 30996
rect 17442 30522 17502 30996
rect 18210 30522 18270 30996
rect 18978 30522 19038 30996
rect 19746 30522 19806 30996
rect 20514 30522 20574 30996
rect 21282 30522 21342 30996
rect 22050 30522 22110 30996
rect 22818 30522 22878 30996
rect 23586 30522 23646 30996
rect 24354 30796 24414 30996
rect 25122 30796 25182 30996
rect 25890 30796 25950 30996
rect 26658 30796 26718 30996
rect 27426 30796 27486 30996
rect 28194 30796 28254 30996
rect 28962 30796 29022 30996
rect 29730 30796 29790 30996
rect 30498 30522 30558 30996
rect 31266 30522 31326 30996
rect 32034 30522 32094 30996
rect 32802 30522 32862 30996
rect 33570 30522 33630 30996
rect 34338 30522 34398 30996
rect 35106 30522 35166 30996
rect 35874 30522 35934 30996
rect 36642 30522 36702 30996
rect 37410 30522 37470 30996
rect 38178 30522 38238 30996
rect 800 30446 1732 30456
rect 10517 30462 10604 30522
rect 800 28722 1600 30446
rect 10517 30366 10604 30375
rect 11285 30462 11372 30522
rect 11285 30366 11372 30375
rect 12053 30462 12140 30522
rect 12053 30366 12140 30375
rect 12821 30462 12908 30522
rect 12821 30366 12908 30375
rect 13589 30462 13676 30522
rect 13589 30366 13676 30375
rect 14357 30462 14444 30522
rect 14357 30366 14444 30375
rect 15125 30462 15212 30522
rect 15125 30366 15212 30375
rect 15893 30462 15980 30522
rect 15893 30366 15980 30375
rect 16661 30462 16748 30522
rect 16661 30366 16748 30375
rect 17429 30462 17516 30522
rect 17429 30366 17516 30375
rect 18197 30462 18284 30522
rect 18197 30366 18284 30375
rect 18965 30462 19052 30522
rect 18965 30366 19052 30375
rect 19733 30462 19820 30522
rect 19733 30366 19820 30375
rect 20501 30462 20588 30522
rect 20501 30366 20588 30375
rect 21269 30462 21356 30522
rect 21269 30366 21356 30375
rect 22037 30462 22124 30522
rect 22037 30366 22124 30375
rect 22805 30462 22892 30522
rect 22805 30366 22892 30375
rect 23573 30462 23660 30522
rect 23573 30366 23660 30375
rect 30480 30458 30576 30522
rect 1660 30320 1860 30360
rect 30480 30353 30576 30362
rect 31248 30458 31344 30522
rect 31248 30353 31344 30362
rect 32016 30458 32112 30522
rect 32016 30353 32112 30362
rect 32784 30458 32880 30522
rect 32784 30353 32880 30362
rect 33552 30458 33648 30522
rect 33552 30353 33648 30362
rect 34320 30458 34416 30522
rect 34320 30353 34416 30362
rect 35088 30458 35184 30522
rect 35088 30353 35184 30362
rect 35856 30458 35952 30522
rect 35856 30353 35952 30362
rect 36624 30458 36720 30522
rect 36624 30353 36720 30362
rect 37392 30458 37488 30522
rect 37392 30353 37488 30362
rect 38160 30458 38256 30522
rect 38160 30353 38256 30362
rect 1660 30300 1880 30320
rect 1820 30260 1900 30300
rect 1820 30240 1880 30260
rect 1800 30200 1860 30240
rect 1780 30180 1860 30200
rect 1660 30120 1900 30180
rect 2268 30118 2936 30244
rect 1700 30020 1860 30060
rect 1660 30000 1900 30020
rect 1660 29940 1740 30000
rect 1820 29940 1900 30000
rect 1660 29920 1900 29940
rect 2148 30014 3040 30118
rect 1700 29880 1860 29920
rect 1840 29760 1900 29820
rect 1660 29700 1980 29760
rect 2148 29730 2420 30014
rect 2768 29730 3040 30014
rect 3276 29834 3484 29910
rect 3630 29834 3944 29910
rect 4496 29882 4768 30118
rect 7482 30000 38626 30276
rect 3276 29750 3944 29834
rect 1840 29640 1900 29700
rect 1660 29540 1860 29580
rect 1660 29520 1880 29540
rect 1820 29480 1900 29520
rect 2148 29500 3040 29730
rect 1820 29460 1880 29480
rect 1800 29420 1860 29460
rect 1780 29400 1860 29420
rect 1660 29340 1900 29400
rect 1660 29240 1940 29280
rect 1660 29200 1980 29240
rect 1740 29120 1820 29200
rect 1900 29120 1980 29200
rect 2148 29124 2420 29500
rect 2768 29124 3040 29500
rect 3262 29680 4118 29750
rect 3262 29596 3652 29680
rect 3262 29124 3534 29596
rect 3846 29124 4118 29680
rect 4314 29652 4982 29882
rect 5250 29756 5918 29876
rect 6184 29840 6392 29916
rect 6538 29840 6852 29916
rect 6184 29756 6852 29840
rect 4496 29124 4768 29652
rect 5174 29646 5996 29756
rect 5174 29354 5446 29646
rect 5724 29354 5996 29646
rect 5174 29262 5996 29354
rect 6170 29686 7026 29756
rect 6170 29602 6560 29686
rect 5258 29124 5926 29262
rect 6170 29130 6442 29602
rect 6754 29130 7026 29686
rect 1660 29080 1980 29120
rect 1660 29040 1940 29080
rect 7482 28722 7758 30000
rect 10519 29512 10528 29817
rect 10841 29512 10850 29817
rect 10532 28760 10837 29512
rect 11792 28740 12068 30000
rect 18287 29512 18296 29817
rect 18609 29512 18618 29817
rect 18300 28812 18605 29512
rect 19562 28740 19838 30000
rect 26046 29512 26055 29817
rect 26368 29512 26377 29817
rect 26059 28838 26364 29512
rect 27348 28844 27624 30000
rect 33831 29512 33840 29817
rect 34153 29512 34162 29817
rect 33844 28812 34149 29512
rect 35100 28810 35376 30000
rect 39440 29884 40240 30596
rect 38893 29444 38902 29884
rect 39342 29444 40240 29884
rect 800 28446 7758 28722
rect 800 26538 1600 28446
rect 3881 28013 5333 28030
rect 2120 27886 2668 27992
rect 3300 27960 3500 28000
rect 2120 27858 2760 27886
rect 1740 27620 1800 27680
rect 1660 27560 1960 27620
rect 1740 27500 1800 27560
rect 2120 27514 2300 27858
rect 2462 27758 2760 27858
rect 3180 27840 3500 27960
rect 2562 27514 2760 27758
rect 3080 27720 3500 27840
rect 1740 27460 1920 27500
rect 2120 27460 2760 27514
rect 2920 27640 3500 27720
rect 3881 27708 3898 28013
rect 4203 27708 5333 28013
rect 3881 27691 5333 27708
rect 1740 27440 1900 27460
rect 1660 27360 1760 27380
rect 1660 27340 1780 27360
rect 2120 27346 2610 27460
rect 2920 27440 3120 27640
rect 3300 27440 3500 27640
rect 6240 27602 6516 28446
rect 1660 27320 1800 27340
rect 1720 27300 1940 27320
rect 1740 27280 1940 27300
rect 1760 27260 1960 27280
rect 1780 27200 1840 27260
rect 1900 27200 1960 27260
rect 1660 27120 1960 27200
rect 2120 27270 2760 27346
rect 2920 27300 3660 27440
rect 2120 26862 2294 27270
rect 2458 27208 2760 27270
rect 2562 26862 2760 27208
rect 3300 26860 3500 27300
rect 800 26518 4544 26538
rect 800 26216 4336 26518
rect 4524 26216 4544 26518
rect 800 26196 4544 26216
rect 425 24776 605 24785
rect 0 24596 425 24776
rect 425 24587 605 24596
rect 0 21396 427 21576
rect 607 21396 616 21576
rect 800 18978 1600 26196
rect 800 18958 4544 18978
rect 800 18656 4336 18958
rect 4524 18656 4544 18958
rect 800 18636 4544 18656
rect 401 18376 581 18385
rect 0 18196 401 18376
rect 401 18187 581 18196
rect 0 14996 200 15176
rect 800 11418 1600 18636
rect 800 11398 4544 11418
rect 800 11096 4336 11398
rect 4524 11096 4544 11398
rect 800 11076 4544 11096
rect 800 1840 1600 11076
rect 800 1610 4600 1840
rect 800 1100 3940 1610
rect 4550 1100 4600 1610
rect 800 1030 4600 1100
rect 800 0 1600 1030
rect 4890 796 5406 3116
rect 6102 1628 6707 3082
rect 6102 1100 6140 1628
rect 6668 1100 6707 1628
rect 6102 1040 6707 1100
rect 10448 796 10968 2534
rect 11718 1584 12158 2488
rect 11718 1135 12158 1144
rect 18214 796 18734 2540
rect 19492 1584 19932 2372
rect 19492 1135 19932 1144
rect 25998 796 26518 2556
rect 27266 1578 27706 2372
rect 27266 1129 27706 1138
rect 33750 796 34270 2482
rect 35040 1570 35480 2372
rect 35040 1121 35480 1130
rect 39440 796 40240 29444
rect 4890 34 40240 796
rect 39440 0 40240 34
use r2r_dac  blue_dac
timestamp 1747574105
transform 0 -1 3596 -1 0 8292
box -2862 -1084 3942 844
use controller  controller_0
timestamp 1747539407
transform 1 0 7402 0 1 1156
box 0 652 31452 29000
use r2r_dac  green_dac
timestamp 1747574105
transform 0 -1 3596 -1 0 15852
box -2862 -1084 3942 844
use r2r_dac  red_dac
timestamp 1747574105
transform 0 -1 3596 -1 0 23412
box -2862 -1084 3942 844
use rgb_buffers  rgb_buffers_0
timestamp 1747539407
transform 1 0 4652 0 1 2416
box 0 -56 2600 25760
<< labels >>
flabel metal5 s 37410 30796 37470 30996 4 FreeSans 320 0 0 0 clk
port 2 nsew
flabel metal5 s 38178 30796 38238 30996 4 FreeSans 320 0 0 0 ena
port 3 nsew
flabel metal5 s 36642 30796 36702 30996 4 FreeSans 320 0 0 0 rst_n
port 4 nsew
flabel metal5 s 35874 30796 35934 30996 4 FreeSans 320 0 0 0 ui_in[0]
port 5 nsew
flabel metal5 s 35106 30796 35166 30996 4 FreeSans 320 0 0 0 ui_in[1]
port 6 nsew
flabel metal5 s 34338 30796 34398 30996 4 FreeSans 320 0 0 0 ui_in[2]
port 7 nsew
flabel metal5 s 33570 30796 33630 30996 4 FreeSans 320 0 0 0 ui_in[3]
port 8 nsew
flabel metal5 s 32802 30796 32862 30996 4 FreeSans 320 0 0 0 ui_in[4]
port 9 nsew
flabel metal5 s 32034 30796 32094 30996 4 FreeSans 320 0 0 0 ui_in[5]
port 10 nsew
flabel metal5 s 31266 30796 31326 30996 4 FreeSans 320 0 0 0 ui_in[6]
port 11 nsew
flabel metal5 s 30498 30796 30558 30996 4 FreeSans 320 0 0 0 ui_in[7]
port 12 nsew
flabel metal5 s 29730 30796 29790 30996 4 FreeSans 320 0 0 0 uio_in[0]
port 13 nsew
flabel metal5 s 28962 30796 29022 30996 4 FreeSans 320 0 0 0 uio_in[1]
port 14 nsew
flabel metal5 s 28194 30796 28254 30996 4 FreeSans 320 0 0 0 uio_in[2]
port 15 nsew
flabel metal5 s 27426 30796 27486 30996 4 FreeSans 320 0 0 0 uio_in[3]
port 16 nsew
flabel metal5 s 26658 30796 26718 30996 4 FreeSans 320 0 0 0 uio_in[4]
port 17 nsew
flabel metal5 s 25890 30796 25950 30996 4 FreeSans 320 0 0 0 uio_in[5]
port 18 nsew
flabel metal5 s 25122 30796 25182 30996 4 FreeSans 320 0 0 0 uio_in[6]
port 19 nsew
flabel metal5 s 24354 30796 24414 30996 4 FreeSans 320 0 0 0 uio_in[7]
port 20 nsew
flabel metal5 s 11298 30796 11358 30996 4 FreeSans 320 0 0 0 uio_oe[0]
port 21 nsew
flabel metal5 s 10530 30796 10590 30996 4 FreeSans 320 0 0 0 uio_oe[1]
port 22 nsew
flabel metal5 s 9762 30796 9822 30996 4 FreeSans 320 0 0 0 uio_oe[2]
port 23 nsew
flabel metal5 s 8994 30796 9054 30996 4 FreeSans 320 0 0 0 uio_oe[3]
port 24 nsew
flabel metal5 s 8226 30796 8286 30996 4 FreeSans 320 0 0 0 uio_oe[4]
port 25 nsew
flabel metal5 s 7458 30796 7518 30996 4 FreeSans 320 0 0 0 uio_oe[5]
port 26 nsew
flabel metal5 s 6690 30796 6750 30996 4 FreeSans 320 0 0 0 uio_oe[6]
port 27 nsew
flabel metal5 s 5922 30796 5982 30996 4 FreeSans 320 0 0 0 uio_oe[7]
port 28 nsew
flabel metal5 s 17442 30796 17502 30996 4 FreeSans 320 0 0 0 uio_out[0]
port 29 nsew
flabel metal5 s 16674 30796 16734 30996 4 FreeSans 320 0 0 0 uio_out[1]
port 30 nsew
flabel metal5 s 15906 30796 15966 30996 4 FreeSans 320 0 0 0 uio_out[2]
port 31 nsew
flabel metal5 s 15138 30796 15198 30996 4 FreeSans 320 0 0 0 uio_out[3]
port 32 nsew
flabel metal5 s 14370 30796 14430 30996 4 FreeSans 320 0 0 0 uio_out[4]
port 33 nsew
flabel metal5 s 13602 30796 13662 30996 4 FreeSans 320 0 0 0 uio_out[5]
port 34 nsew
flabel metal5 s 12834 30796 12894 30996 4 FreeSans 320 0 0 0 uio_out[6]
port 35 nsew
flabel metal5 s 12066 30796 12126 30996 4 FreeSans 320 0 0 0 uio_out[7]
port 36 nsew
flabel metal5 s 23586 30796 23646 30996 4 FreeSans 320 0 0 0 uo_out[0]
port 37 nsew
flabel metal5 s 22818 30796 22878 30996 4 FreeSans 320 0 0 0 uo_out[1]
port 38 nsew
flabel metal5 s 22050 30796 22110 30996 4 FreeSans 320 0 0 0 uo_out[2]
port 39 nsew
flabel metal5 s 21282 30796 21342 30996 4 FreeSans 320 0 0 0 uo_out[3]
port 40 nsew
flabel metal5 s 20514 30796 20574 30996 4 FreeSans 320 0 0 0 uo_out[4]
port 41 nsew
flabel metal5 s 19746 30796 19806 30996 4 FreeSans 320 0 0 0 uo_out[5]
port 42 nsew
flabel metal5 s 18978 30796 19038 30996 4 FreeSans 320 0 0 0 uo_out[6]
port 43 nsew
flabel metal5 s 18210 30796 18270 30996 4 FreeSans 320 0 0 0 uo_out[7]
port 44 nsew
flabel metal5 s 0 24596 200 24776 0 FreeSans 320 0 0 0 ua[0]
port 45 nsew
flabel metal5 s 0 21396 200 21576 0 FreeSans 320 0 0 0 ua[1]
port 46 nsew
flabel metal5 s 0 18196 200 18376 0 FreeSans 320 0 0 0 ua[2]
port 47 nsew
flabel metal5 s 0 14996 200 15176 0 FreeSans 320 0 0 0 ua[3]
port 48 nsew
flabel metal5 s 800 0 1600 30596 0 FreeSans 3200 90 0 0 VGND
port 49 nsew
flabel metal5 s 39440 0 40240 30596 0 FreeSans 3200 90 0 0 VPWR
port 51 nsew
<< properties >>
string FIXED_BBOX 0 0 40416 30996
<< end >>
